// Benchmark "top" written by ABC on Mon Sep 21 03:43:19 2020

module top ( 
    \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] , \a[24] ,
    \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] , \a[32] ,
    \a[33] , \a[34] , \a[35] , \a[36] , \a[37] , \a[38] , \a[39] , \a[40] ,
    \a[41] , \a[42] , \a[43] , \a[44] , \a[45] , \a[46] , \a[47] , \a[48] ,
    \a[49] , \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] , \a[56] ,
    \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] , \a[64] ,
    \a[65] , \a[66] , \a[67] , \a[68] , \a[69] , \a[70] , \a[71] , \a[72] ,
    \a[73] , \a[74] , \a[75] , \a[76] , \a[77] , \a[78] , \a[79] , \a[80] ,
    \a[81] , \a[82] , \a[83] , \a[84] , \a[85] , \a[86] , \a[87] , \a[88] ,
    \a[89] , \a[90] , \a[91] , \a[92] , \a[93] , \a[94] , \a[95] , \a[96] ,
    \a[97] , \a[98] , \a[99] , \a[100] , \a[101] , \a[102] , \a[103] ,
    \a[104] , \a[105] , \a[106] , \a[107] , \a[108] , \a[109] , \a[110] ,
    \a[111] , \a[112] , \a[113] , \a[114] , \a[115] , \a[116] , \a[117] ,
    \a[118] , \a[119] , \a[120] , \a[121] , \a[122] , \a[123] , \a[124] ,
    \a[125] , \a[126] , \a[127] ,
    \asqrt[0] , \asqrt[1] , \asqrt[2] , \asqrt[3] , \asqrt[4] , \asqrt[5] ,
    \asqrt[6] , \asqrt[7] , \asqrt[8] , \asqrt[9] , \asqrt[10] ,
    \asqrt[11] , \asqrt[12] , \asqrt[13] , \asqrt[14] , \asqrt[15] ,
    \asqrt[16] , \asqrt[17] , \asqrt[18] , \asqrt[19] , \asqrt[20] ,
    \asqrt[21] , \asqrt[22] , \asqrt[23] , \asqrt[24] , \asqrt[25] ,
    \asqrt[26] , \asqrt[27] , \asqrt[28] , \asqrt[29] , \asqrt[30] ,
    \asqrt[31] , \asqrt[32] , \asqrt[33] , \asqrt[34] , \asqrt[35] ,
    \asqrt[36] , \asqrt[37] , \asqrt[38] , \asqrt[39] , \asqrt[40] ,
    \asqrt[41] , \asqrt[42] , \asqrt[43] , \asqrt[44] , \asqrt[45] ,
    \asqrt[46] , \asqrt[47] , \asqrt[48] , \asqrt[49] , \asqrt[50] ,
    \asqrt[51] , \asqrt[52] , \asqrt[53] , \asqrt[54] , \asqrt[55] ,
    \asqrt[56] , \asqrt[57] , \asqrt[58] , \asqrt[59] , \asqrt[60] ,
    \asqrt[61] , \asqrt[62] , \asqrt[63]   );
  input  \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] ,
    \a[8] , \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] ,
    \a[32] , \a[33] , \a[34] , \a[35] , \a[36] , \a[37] , \a[38] , \a[39] ,
    \a[40] , \a[41] , \a[42] , \a[43] , \a[44] , \a[45] , \a[46] , \a[47] ,
    \a[48] , \a[49] , \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] ,
    \a[56] , \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] ,
    \a[64] , \a[65] , \a[66] , \a[67] , \a[68] , \a[69] , \a[70] , \a[71] ,
    \a[72] , \a[73] , \a[74] , \a[75] , \a[76] , \a[77] , \a[78] , \a[79] ,
    \a[80] , \a[81] , \a[82] , \a[83] , \a[84] , \a[85] , \a[86] , \a[87] ,
    \a[88] , \a[89] , \a[90] , \a[91] , \a[92] , \a[93] , \a[94] , \a[95] ,
    \a[96] , \a[97] , \a[98] , \a[99] , \a[100] , \a[101] , \a[102] ,
    \a[103] , \a[104] , \a[105] , \a[106] , \a[107] , \a[108] , \a[109] ,
    \a[110] , \a[111] , \a[112] , \a[113] , \a[114] , \a[115] , \a[116] ,
    \a[117] , \a[118] , \a[119] , \a[120] , \a[121] , \a[122] , \a[123] ,
    \a[124] , \a[125] , \a[126] , \a[127] ;
  output \asqrt[0] , \asqrt[1] , \asqrt[2] , \asqrt[3] , \asqrt[4] ,
    \asqrt[5] , \asqrt[6] , \asqrt[7] , \asqrt[8] , \asqrt[9] ,
    \asqrt[10] , \asqrt[11] , \asqrt[12] , \asqrt[13] , \asqrt[14] ,
    \asqrt[15] , \asqrt[16] , \asqrt[17] , \asqrt[18] , \asqrt[19] ,
    \asqrt[20] , \asqrt[21] , \asqrt[22] , \asqrt[23] , \asqrt[24] ,
    \asqrt[25] , \asqrt[26] , \asqrt[27] , \asqrt[28] , \asqrt[29] ,
    \asqrt[30] , \asqrt[31] , \asqrt[32] , \asqrt[33] , \asqrt[34] ,
    \asqrt[35] , \asqrt[36] , \asqrt[37] , \asqrt[38] , \asqrt[39] ,
    \asqrt[40] , \asqrt[41] , \asqrt[42] , \asqrt[43] , \asqrt[44] ,
    \asqrt[45] , \asqrt[46] , \asqrt[47] , \asqrt[48] , \asqrt[49] ,
    \asqrt[50] , \asqrt[51] , \asqrt[52] , \asqrt[53] , \asqrt[54] ,
    \asqrt[55] , \asqrt[56] , \asqrt[57] , \asqrt[58] , \asqrt[59] ,
    \asqrt[60] , \asqrt[61] , \asqrt[62] , \asqrt[63] ;
  wire new_n193_, new_n194_, new_n197_, new_n198_, new_n199_, new_n200_,
    new_n201_, new_n202_, new_n203_, new_n204_, new_n205_, new_n206_,
    new_n207_, new_n208_, new_n209_, new_n210_, new_n211_, new_n212_,
    new_n213_, new_n214_, new_n215_, new_n216_, new_n217_, new_n218_,
    new_n219_, new_n220_, new_n221_, new_n222_, new_n223_, new_n224_,
    new_n225_, new_n226_, new_n227_, new_n228_, new_n229_, new_n230_,
    new_n231_, new_n232_, new_n233_, new_n234_, new_n235_, new_n236_,
    new_n237_, new_n238_, new_n239_, new_n240_, new_n241_, new_n242_,
    new_n243_, new_n244_, new_n245_, new_n246_, new_n247_, new_n248_,
    new_n249_, new_n250_, new_n251_, new_n252_, new_n255_, new_n256_,
    new_n257_, new_n258_, new_n259_, new_n260_, new_n261_, new_n262_,
    new_n263_, new_n264_, new_n265_, new_n266_, new_n267_, new_n268_,
    new_n269_, new_n270_, new_n271_, new_n272_, new_n273_, new_n274_,
    new_n275_, new_n276_, new_n277_, new_n278_, new_n279_, new_n280_,
    new_n281_, new_n282_, new_n283_, new_n284_, new_n285_, new_n286_,
    new_n287_, new_n288_, new_n289_, new_n290_, new_n291_, new_n292_,
    new_n293_, new_n294_, new_n295_, new_n296_, new_n297_, new_n298_,
    new_n299_, new_n300_, new_n301_, new_n302_, new_n303_, new_n304_,
    new_n305_, new_n306_, new_n307_, new_n308_, new_n309_, new_n310_,
    new_n311_, new_n312_, new_n313_, new_n314_, new_n315_, new_n317_,
    new_n318_, new_n319_, new_n320_, new_n321_, new_n322_, new_n323_,
    new_n324_, new_n325_, new_n326_, new_n327_, new_n328_, new_n329_,
    new_n330_, new_n331_, new_n332_, new_n333_, new_n334_, new_n335_,
    new_n336_, new_n337_, new_n338_, new_n339_, new_n340_, new_n341_,
    new_n342_, new_n343_, new_n344_, new_n345_, new_n346_, new_n347_,
    new_n348_, new_n349_, new_n350_, new_n351_, new_n352_, new_n353_,
    new_n354_, new_n355_, new_n356_, new_n357_, new_n358_, new_n359_,
    new_n360_, new_n361_, new_n362_, new_n363_, new_n364_, new_n365_,
    new_n366_, new_n367_, new_n368_, new_n369_, new_n370_, new_n371_,
    new_n372_, new_n373_, new_n374_, new_n375_, new_n376_, new_n377_,
    new_n378_, new_n379_, new_n380_, new_n381_, new_n382_, new_n383_,
    new_n384_, new_n385_, new_n386_, new_n387_, new_n388_, new_n389_,
    new_n390_, new_n391_, new_n392_, new_n393_, new_n394_, new_n395_,
    new_n396_, new_n397_, new_n399_, new_n400_, new_n401_, new_n402_,
    new_n403_, new_n404_, new_n405_, new_n406_, new_n407_, new_n408_,
    new_n409_, new_n410_, new_n411_, new_n412_, new_n413_, new_n414_,
    new_n415_, new_n416_, new_n417_, new_n418_, new_n419_, new_n420_,
    new_n421_, new_n422_, new_n423_, new_n424_, new_n425_, new_n426_,
    new_n427_, new_n428_, new_n429_, new_n430_, new_n431_, new_n432_,
    new_n433_, new_n434_, new_n435_, new_n436_, new_n437_, new_n438_,
    new_n439_, new_n440_, new_n441_, new_n442_, new_n443_, new_n444_,
    new_n445_, new_n446_, new_n447_, new_n448_, new_n449_, new_n450_,
    new_n451_, new_n452_, new_n453_, new_n454_, new_n455_, new_n456_,
    new_n457_, new_n458_, new_n459_, new_n460_, new_n461_, new_n462_,
    new_n463_, new_n464_, new_n465_, new_n466_, new_n467_, new_n468_,
    new_n469_, new_n470_, new_n471_, new_n472_, new_n473_, new_n474_,
    new_n475_, new_n476_, new_n477_, new_n478_, new_n479_, new_n480_,
    new_n481_, new_n483_, new_n484_, new_n485_, new_n486_, new_n487_,
    new_n488_, new_n489_, new_n490_, new_n491_, new_n492_, new_n493_,
    new_n494_, new_n495_, new_n496_, new_n497_, new_n498_, new_n499_,
    new_n500_, new_n501_, new_n502_, new_n503_, new_n504_, new_n505_,
    new_n506_, new_n507_, new_n508_, new_n509_, new_n510_, new_n511_,
    new_n512_, new_n513_, new_n514_, new_n515_, new_n516_, new_n517_,
    new_n518_, new_n519_, new_n520_, new_n521_, new_n522_, new_n523_,
    new_n524_, new_n525_, new_n526_, new_n527_, new_n528_, new_n529_,
    new_n530_, new_n531_, new_n532_, new_n533_, new_n534_, new_n535_,
    new_n536_, new_n537_, new_n538_, new_n539_, new_n540_, new_n541_,
    new_n542_, new_n543_, new_n544_, new_n545_, new_n546_, new_n547_,
    new_n548_, new_n549_, new_n550_, new_n551_, new_n552_, new_n553_,
    new_n554_, new_n555_, new_n556_, new_n557_, new_n558_, new_n559_,
    new_n560_, new_n561_, new_n562_, new_n563_, new_n564_, new_n565_,
    new_n566_, new_n567_, new_n568_, new_n569_, new_n570_, new_n571_,
    new_n572_, new_n573_, new_n574_, new_n575_, new_n576_, new_n577_,
    new_n578_, new_n579_, new_n580_, new_n581_, new_n582_, new_n583_,
    new_n584_, new_n585_, new_n586_, new_n587_, new_n588_, new_n589_,
    new_n590_, new_n591_, new_n592_, new_n594_, new_n595_, new_n596_,
    new_n597_, new_n598_, new_n599_, new_n600_, new_n601_, new_n602_,
    new_n603_, new_n604_, new_n605_, new_n606_, new_n607_, new_n608_,
    new_n609_, new_n610_, new_n611_, new_n612_, new_n613_, new_n614_,
    new_n615_, new_n616_, new_n617_, new_n618_, new_n619_, new_n620_,
    new_n621_, new_n622_, new_n623_, new_n624_, new_n625_, new_n626_,
    new_n627_, new_n628_, new_n629_, new_n630_, new_n631_, new_n632_,
    new_n633_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_,
    new_n639_, new_n640_, new_n641_, new_n642_, new_n643_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n790_, new_n791_, new_n792_, new_n793_, new_n794_, new_n795_,
    new_n796_, new_n797_, new_n798_, new_n799_, new_n800_, new_n801_,
    new_n802_, new_n803_, new_n804_, new_n805_, new_n806_, new_n807_,
    new_n808_, new_n809_, new_n810_, new_n811_, new_n812_, new_n813_,
    new_n815_, new_n816_, new_n817_, new_n818_, new_n819_, new_n820_,
    new_n821_, new_n822_, new_n823_, new_n824_, new_n825_, new_n826_,
    new_n827_, new_n828_, new_n829_, new_n830_, new_n831_, new_n832_,
    new_n833_, new_n834_, new_n835_, new_n836_, new_n837_, new_n838_,
    new_n839_, new_n840_, new_n841_, new_n842_, new_n843_, new_n844_,
    new_n845_, new_n846_, new_n847_, new_n848_, new_n849_, new_n850_,
    new_n851_, new_n852_, new_n853_, new_n854_, new_n855_, new_n856_,
    new_n857_, new_n858_, new_n859_, new_n860_, new_n861_, new_n862_,
    new_n863_, new_n864_, new_n865_, new_n866_, new_n867_, new_n868_,
    new_n869_, new_n870_, new_n871_, new_n872_, new_n873_, new_n874_,
    new_n875_, new_n876_, new_n877_, new_n878_, new_n879_, new_n880_,
    new_n881_, new_n882_, new_n883_, new_n884_, new_n885_, new_n886_,
    new_n887_, new_n888_, new_n889_, new_n890_, new_n891_, new_n892_,
    new_n893_, new_n894_, new_n895_, new_n896_, new_n897_, new_n898_,
    new_n899_, new_n900_, new_n901_, new_n902_, new_n903_, new_n904_,
    new_n905_, new_n906_, new_n907_, new_n908_, new_n909_, new_n910_,
    new_n911_, new_n912_, new_n913_, new_n914_, new_n915_, new_n916_,
    new_n917_, new_n918_, new_n919_, new_n920_, new_n921_, new_n922_,
    new_n923_, new_n924_, new_n925_, new_n926_, new_n927_, new_n928_,
    new_n929_, new_n930_, new_n931_, new_n932_, new_n933_, new_n934_,
    new_n935_, new_n936_, new_n937_, new_n938_, new_n939_, new_n940_,
    new_n941_, new_n942_, new_n943_, new_n944_, new_n945_, new_n946_,
    new_n947_, new_n948_, new_n949_, new_n950_, new_n951_, new_n952_,
    new_n953_, new_n954_, new_n955_, new_n956_, new_n957_, new_n958_,
    new_n959_, new_n961_, new_n962_, new_n963_, new_n964_, new_n965_,
    new_n966_, new_n967_, new_n968_, new_n969_, new_n970_, new_n971_,
    new_n972_, new_n973_, new_n974_, new_n975_, new_n976_, new_n977_,
    new_n978_, new_n979_, new_n980_, new_n981_, new_n982_, new_n983_,
    new_n984_, new_n985_, new_n986_, new_n987_, new_n988_, new_n989_,
    new_n990_, new_n991_, new_n992_, new_n993_, new_n994_, new_n995_,
    new_n996_, new_n997_, new_n998_, new_n999_, new_n1000_, new_n1001_,
    new_n1002_, new_n1003_, new_n1004_, new_n1005_, new_n1006_, new_n1007_,
    new_n1008_, new_n1009_, new_n1010_, new_n1011_, new_n1012_, new_n1013_,
    new_n1014_, new_n1015_, new_n1016_, new_n1017_, new_n1018_, new_n1019_,
    new_n1020_, new_n1021_, new_n1022_, new_n1023_, new_n1024_, new_n1025_,
    new_n1026_, new_n1027_, new_n1028_, new_n1029_, new_n1030_, new_n1031_,
    new_n1032_, new_n1033_, new_n1034_, new_n1035_, new_n1036_, new_n1037_,
    new_n1038_, new_n1039_, new_n1040_, new_n1041_, new_n1042_, new_n1043_,
    new_n1044_, new_n1045_, new_n1046_, new_n1047_, new_n1048_, new_n1049_,
    new_n1050_, new_n1051_, new_n1052_, new_n1053_, new_n1054_, new_n1055_,
    new_n1056_, new_n1057_, new_n1058_, new_n1059_, new_n1060_, new_n1061_,
    new_n1062_, new_n1063_, new_n1064_, new_n1065_, new_n1066_, new_n1067_,
    new_n1068_, new_n1069_, new_n1070_, new_n1071_, new_n1072_, new_n1073_,
    new_n1074_, new_n1075_, new_n1076_, new_n1077_, new_n1078_, new_n1079_,
    new_n1080_, new_n1081_, new_n1082_, new_n1083_, new_n1084_, new_n1085_,
    new_n1086_, new_n1087_, new_n1088_, new_n1089_, new_n1090_, new_n1091_,
    new_n1092_, new_n1093_, new_n1094_, new_n1095_, new_n1096_, new_n1097_,
    new_n1098_, new_n1099_, new_n1100_, new_n1101_, new_n1102_, new_n1103_,
    new_n1104_, new_n1105_, new_n1106_, new_n1107_, new_n1108_, new_n1109_,
    new_n1110_, new_n1111_, new_n1112_, new_n1113_, new_n1114_, new_n1115_,
    new_n1116_, new_n1117_, new_n1118_, new_n1119_, new_n1120_, new_n1121_,
    new_n1122_, new_n1123_, new_n1124_, new_n1125_, new_n1126_, new_n1127_,
    new_n1128_, new_n1129_, new_n1130_, new_n1131_, new_n1132_, new_n1133_,
    new_n1134_, new_n1135_, new_n1136_, new_n1137_, new_n1138_, new_n1139_,
    new_n1140_, new_n1141_, new_n1142_, new_n1143_, new_n1144_, new_n1145_,
    new_n1146_, new_n1147_, new_n1148_, new_n1149_, new_n1150_, new_n1151_,
    new_n1152_, new_n1153_, new_n1154_, new_n1155_, new_n1156_, new_n1157_,
    new_n1158_, new_n1159_, new_n1160_, new_n1161_, new_n1162_, new_n1163_,
    new_n1164_, new_n1165_, new_n1166_, new_n1167_, new_n1168_, new_n1169_,
    new_n1170_, new_n1171_, new_n1172_, new_n1173_, new_n1174_, new_n1175_,
    new_n1176_, new_n1177_, new_n1178_, new_n1179_, new_n1180_, new_n1181_,
    new_n1182_, new_n1183_, new_n1184_, new_n1185_, new_n1186_, new_n1187_,
    new_n1188_, new_n1190_, new_n1191_, new_n1192_, new_n1193_, new_n1194_,
    new_n1195_, new_n1196_, new_n1197_, new_n1198_, new_n1199_, new_n1200_,
    new_n1201_, new_n1202_, new_n1203_, new_n1204_, new_n1205_, new_n1206_,
    new_n1207_, new_n1208_, new_n1209_, new_n1210_, new_n1211_, new_n1212_,
    new_n1213_, new_n1214_, new_n1215_, new_n1216_, new_n1217_, new_n1218_,
    new_n1219_, new_n1220_, new_n1221_, new_n1222_, new_n1223_, new_n1224_,
    new_n1225_, new_n1226_, new_n1227_, new_n1228_, new_n1229_, new_n1230_,
    new_n1231_, new_n1232_, new_n1233_, new_n1234_, new_n1235_, new_n1236_,
    new_n1237_, new_n1238_, new_n1239_, new_n1240_, new_n1241_, new_n1242_,
    new_n1243_, new_n1244_, new_n1245_, new_n1246_, new_n1247_, new_n1248_,
    new_n1249_, new_n1250_, new_n1251_, new_n1252_, new_n1253_, new_n1254_,
    new_n1255_, new_n1256_, new_n1257_, new_n1258_, new_n1259_, new_n1260_,
    new_n1261_, new_n1262_, new_n1263_, new_n1264_, new_n1265_, new_n1266_,
    new_n1267_, new_n1268_, new_n1269_, new_n1270_, new_n1271_, new_n1272_,
    new_n1273_, new_n1274_, new_n1275_, new_n1277_, new_n1278_, new_n1279_,
    new_n1280_, new_n1281_, new_n1282_, new_n1283_, new_n1284_, new_n1285_,
    new_n1286_, new_n1287_, new_n1288_, new_n1289_, new_n1290_, new_n1291_,
    new_n1292_, new_n1293_, new_n1294_, new_n1295_, new_n1296_, new_n1297_,
    new_n1298_, new_n1299_, new_n1300_, new_n1301_, new_n1302_, new_n1303_,
    new_n1304_, new_n1305_, new_n1306_, new_n1307_, new_n1308_, new_n1309_,
    new_n1310_, new_n1311_, new_n1312_, new_n1313_, new_n1314_, new_n1315_,
    new_n1316_, new_n1317_, new_n1318_, new_n1319_, new_n1320_, new_n1321_,
    new_n1322_, new_n1323_, new_n1324_, new_n1325_, new_n1326_, new_n1327_,
    new_n1328_, new_n1329_, new_n1330_, new_n1331_, new_n1332_, new_n1333_,
    new_n1334_, new_n1335_, new_n1336_, new_n1337_, new_n1338_, new_n1339_,
    new_n1340_, new_n1341_, new_n1342_, new_n1343_, new_n1344_, new_n1345_,
    new_n1346_, new_n1347_, new_n1348_, new_n1349_, new_n1350_, new_n1351_,
    new_n1352_, new_n1353_, new_n1354_, new_n1355_, new_n1356_, new_n1357_,
    new_n1358_, new_n1359_, new_n1360_, new_n1361_, new_n1362_, new_n1363_,
    new_n1364_, new_n1365_, new_n1366_, new_n1367_, new_n1368_, new_n1369_,
    new_n1370_, new_n1371_, new_n1372_, new_n1373_, new_n1374_, new_n1375_,
    new_n1376_, new_n1377_, new_n1378_, new_n1379_, new_n1380_, new_n1381_,
    new_n1382_, new_n1383_, new_n1384_, new_n1385_, new_n1386_, new_n1387_,
    new_n1388_, new_n1389_, new_n1390_, new_n1391_, new_n1392_, new_n1393_,
    new_n1394_, new_n1395_, new_n1396_, new_n1397_, new_n1398_, new_n1399_,
    new_n1400_, new_n1401_, new_n1402_, new_n1403_, new_n1404_, new_n1405_,
    new_n1406_, new_n1407_, new_n1408_, new_n1409_, new_n1410_, new_n1411_,
    new_n1412_, new_n1413_, new_n1414_, new_n1415_, new_n1416_, new_n1417_,
    new_n1418_, new_n1419_, new_n1420_, new_n1421_, new_n1422_, new_n1423_,
    new_n1424_, new_n1425_, new_n1426_, new_n1427_, new_n1428_, new_n1429_,
    new_n1430_, new_n1431_, new_n1432_, new_n1433_, new_n1434_, new_n1435_,
    new_n1436_, new_n1437_, new_n1438_, new_n1439_, new_n1440_, new_n1441_,
    new_n1442_, new_n1443_, new_n1444_, new_n1445_, new_n1446_, new_n1447_,
    new_n1449_, new_n1450_, new_n1451_, new_n1452_, new_n1453_, new_n1454_,
    new_n1455_, new_n1456_, new_n1457_, new_n1458_, new_n1459_, new_n1460_,
    new_n1461_, new_n1462_, new_n1463_, new_n1464_, new_n1465_, new_n1466_,
    new_n1467_, new_n1468_, new_n1469_, new_n1470_, new_n1471_, new_n1472_,
    new_n1473_, new_n1474_, new_n1475_, new_n1476_, new_n1477_, new_n1478_,
    new_n1479_, new_n1480_, new_n1481_, new_n1482_, new_n1483_, new_n1484_,
    new_n1485_, new_n1486_, new_n1487_, new_n1488_, new_n1489_, new_n1490_,
    new_n1491_, new_n1492_, new_n1493_, new_n1494_, new_n1495_, new_n1496_,
    new_n1497_, new_n1498_, new_n1499_, new_n1500_, new_n1501_, new_n1502_,
    new_n1503_, new_n1504_, new_n1505_, new_n1506_, new_n1507_, new_n1508_,
    new_n1509_, new_n1510_, new_n1511_, new_n1512_, new_n1513_, new_n1514_,
    new_n1515_, new_n1516_, new_n1517_, new_n1518_, new_n1519_, new_n1520_,
    new_n1521_, new_n1522_, new_n1523_, new_n1524_, new_n1525_, new_n1526_,
    new_n1527_, new_n1528_, new_n1529_, new_n1530_, new_n1531_, new_n1532_,
    new_n1533_, new_n1534_, new_n1535_, new_n1536_, new_n1537_, new_n1538_,
    new_n1539_, new_n1540_, new_n1541_, new_n1542_, new_n1543_, new_n1544_,
    new_n1545_, new_n1546_, new_n1547_, new_n1548_, new_n1549_, new_n1550_,
    new_n1551_, new_n1552_, new_n1553_, new_n1554_, new_n1555_, new_n1556_,
    new_n1557_, new_n1558_, new_n1559_, new_n1560_, new_n1561_, new_n1562_,
    new_n1563_, new_n1564_, new_n1565_, new_n1566_, new_n1567_, new_n1568_,
    new_n1569_, new_n1570_, new_n1571_, new_n1572_, new_n1573_, new_n1574_,
    new_n1575_, new_n1576_, new_n1577_, new_n1578_, new_n1579_, new_n1580_,
    new_n1581_, new_n1582_, new_n1583_, new_n1584_, new_n1585_, new_n1586_,
    new_n1587_, new_n1588_, new_n1589_, new_n1590_, new_n1591_, new_n1592_,
    new_n1593_, new_n1594_, new_n1595_, new_n1596_, new_n1597_, new_n1598_,
    new_n1599_, new_n1600_, new_n1601_, new_n1602_, new_n1603_, new_n1604_,
    new_n1605_, new_n1606_, new_n1607_, new_n1608_, new_n1609_, new_n1610_,
    new_n1611_, new_n1612_, new_n1613_, new_n1614_, new_n1615_, new_n1616_,
    new_n1617_, new_n1618_, new_n1619_, new_n1620_, new_n1621_, new_n1622_,
    new_n1623_, new_n1624_, new_n1625_, new_n1626_, new_n1627_, new_n1628_,
    new_n1629_, new_n1630_, new_n1631_, new_n1632_, new_n1633_, new_n1634_,
    new_n1635_, new_n1636_, new_n1637_, new_n1638_, new_n1639_, new_n1640_,
    new_n1641_, new_n1642_, new_n1643_, new_n1644_, new_n1645_, new_n1646_,
    new_n1647_, new_n1648_, new_n1649_, new_n1650_, new_n1651_, new_n1652_,
    new_n1653_, new_n1654_, new_n1655_, new_n1656_, new_n1657_, new_n1658_,
    new_n1659_, new_n1660_, new_n1661_, new_n1662_, new_n1663_, new_n1664_,
    new_n1665_, new_n1666_, new_n1667_, new_n1668_, new_n1669_, new_n1670_,
    new_n1671_, new_n1672_, new_n1673_, new_n1674_, new_n1675_, new_n1676_,
    new_n1677_, new_n1678_, new_n1679_, new_n1680_, new_n1681_, new_n1682_,
    new_n1683_, new_n1684_, new_n1685_, new_n1686_, new_n1687_, new_n1688_,
    new_n1689_, new_n1690_, new_n1691_, new_n1692_, new_n1693_, new_n1694_,
    new_n1695_, new_n1696_, new_n1697_, new_n1698_, new_n1699_, new_n1700_,
    new_n1701_, new_n1702_, new_n1703_, new_n1704_, new_n1705_, new_n1706_,
    new_n1707_, new_n1708_, new_n1709_, new_n1710_, new_n1711_, new_n1713_,
    new_n1714_, new_n1715_, new_n1716_, new_n1717_, new_n1718_, new_n1719_,
    new_n1720_, new_n1721_, new_n1722_, new_n1723_, new_n1724_, new_n1725_,
    new_n1726_, new_n1727_, new_n1728_, new_n1729_, new_n1730_, new_n1731_,
    new_n1732_, new_n1733_, new_n1734_, new_n1735_, new_n1736_, new_n1737_,
    new_n1738_, new_n1739_, new_n1740_, new_n1741_, new_n1742_, new_n1743_,
    new_n1744_, new_n1745_, new_n1746_, new_n1747_, new_n1748_, new_n1749_,
    new_n1750_, new_n1751_, new_n1752_, new_n1753_, new_n1754_, new_n1755_,
    new_n1756_, new_n1757_, new_n1758_, new_n1759_, new_n1760_, new_n1761_,
    new_n1762_, new_n1763_, new_n1764_, new_n1765_, new_n1766_, new_n1767_,
    new_n1768_, new_n1769_, new_n1770_, new_n1771_, new_n1772_, new_n1773_,
    new_n1774_, new_n1775_, new_n1776_, new_n1777_, new_n1778_, new_n1779_,
    new_n1780_, new_n1781_, new_n1782_, new_n1783_, new_n1784_, new_n1785_,
    new_n1786_, new_n1787_, new_n1788_, new_n1789_, new_n1790_, new_n1791_,
    new_n1792_, new_n1793_, new_n1794_, new_n1795_, new_n1796_, new_n1797_,
    new_n1798_, new_n1799_, new_n1800_, new_n1801_, new_n1802_, new_n1803_,
    new_n1804_, new_n1805_, new_n1806_, new_n1807_, new_n1808_, new_n1809_,
    new_n1810_, new_n1811_, new_n1812_, new_n1813_, new_n1814_, new_n1815_,
    new_n1816_, new_n1817_, new_n1818_, new_n1819_, new_n1820_, new_n1821_,
    new_n1822_, new_n1823_, new_n1824_, new_n1825_, new_n1826_, new_n1827_,
    new_n1828_, new_n1829_, new_n1830_, new_n1831_, new_n1832_, new_n1833_,
    new_n1834_, new_n1836_, new_n1837_, new_n1838_, new_n1839_, new_n1840_,
    new_n1841_, new_n1842_, new_n1843_, new_n1844_, new_n1845_, new_n1846_,
    new_n1847_, new_n1848_, new_n1849_, new_n1850_, new_n1851_, new_n1852_,
    new_n1853_, new_n1854_, new_n1855_, new_n1856_, new_n1857_, new_n1858_,
    new_n1859_, new_n1860_, new_n1861_, new_n1862_, new_n1863_, new_n1864_,
    new_n1865_, new_n1866_, new_n1867_, new_n1868_, new_n1869_, new_n1870_,
    new_n1871_, new_n1872_, new_n1873_, new_n1874_, new_n1875_, new_n1876_,
    new_n1877_, new_n1878_, new_n1879_, new_n1880_, new_n1881_, new_n1882_,
    new_n1883_, new_n1884_, new_n1885_, new_n1886_, new_n1887_, new_n1888_,
    new_n1889_, new_n1890_, new_n1891_, new_n1892_, new_n1893_, new_n1894_,
    new_n1895_, new_n1896_, new_n1897_, new_n1898_, new_n1899_, new_n1900_,
    new_n1901_, new_n1902_, new_n1903_, new_n1904_, new_n1905_, new_n1906_,
    new_n1907_, new_n1908_, new_n1909_, new_n1910_, new_n1911_, new_n1912_,
    new_n1913_, new_n1914_, new_n1915_, new_n1916_, new_n1917_, new_n1918_,
    new_n1919_, new_n1920_, new_n1921_, new_n1922_, new_n1923_, new_n1924_,
    new_n1925_, new_n1926_, new_n1927_, new_n1928_, new_n1929_, new_n1930_,
    new_n1931_, new_n1932_, new_n1933_, new_n1934_, new_n1935_, new_n1936_,
    new_n1937_, new_n1938_, new_n1939_, new_n1940_, new_n1941_, new_n1942_,
    new_n1943_, new_n1944_, new_n1945_, new_n1946_, new_n1947_, new_n1948_,
    new_n1949_, new_n1950_, new_n1951_, new_n1952_, new_n1953_, new_n1954_,
    new_n1955_, new_n1956_, new_n1957_, new_n1958_, new_n1959_, new_n1960_,
    new_n1961_, new_n1962_, new_n1963_, new_n1964_, new_n1965_, new_n1966_,
    new_n1967_, new_n1968_, new_n1969_, new_n1970_, new_n1971_, new_n1972_,
    new_n1973_, new_n1974_, new_n1975_, new_n1976_, new_n1977_, new_n1978_,
    new_n1979_, new_n1980_, new_n1981_, new_n1982_, new_n1983_, new_n1984_,
    new_n1985_, new_n1986_, new_n1987_, new_n1988_, new_n1989_, new_n1990_,
    new_n1991_, new_n1992_, new_n1993_, new_n1994_, new_n1995_, new_n1996_,
    new_n1997_, new_n1998_, new_n1999_, new_n2000_, new_n2001_, new_n2002_,
    new_n2003_, new_n2004_, new_n2005_, new_n2006_, new_n2007_, new_n2008_,
    new_n2009_, new_n2010_, new_n2011_, new_n2012_, new_n2013_, new_n2014_,
    new_n2015_, new_n2016_, new_n2017_, new_n2018_, new_n2019_, new_n2020_,
    new_n2021_, new_n2022_, new_n2023_, new_n2024_, new_n2025_, new_n2026_,
    new_n2027_, new_n2028_, new_n2029_, new_n2030_, new_n2031_, new_n2032_,
    new_n2033_, new_n2034_, new_n2035_, new_n2036_, new_n2037_, new_n2038_,
    new_n2039_, new_n2040_, new_n2041_, new_n2042_, new_n2043_, new_n2044_,
    new_n2045_, new_n2046_, new_n2047_, new_n2048_, new_n2049_, new_n2050_,
    new_n2051_, new_n2052_, new_n2053_, new_n2054_, new_n2055_, new_n2056_,
    new_n2057_, new_n2058_, new_n2059_, new_n2060_, new_n2061_, new_n2062_,
    new_n2063_, new_n2064_, new_n2065_, new_n2067_, new_n2068_, new_n2069_,
    new_n2070_, new_n2071_, new_n2072_, new_n2073_, new_n2074_, new_n2075_,
    new_n2076_, new_n2077_, new_n2078_, new_n2079_, new_n2080_, new_n2081_,
    new_n2082_, new_n2083_, new_n2084_, new_n2085_, new_n2086_, new_n2087_,
    new_n2088_, new_n2089_, new_n2090_, new_n2091_, new_n2092_, new_n2093_,
    new_n2094_, new_n2095_, new_n2096_, new_n2097_, new_n2098_, new_n2099_,
    new_n2100_, new_n2101_, new_n2102_, new_n2103_, new_n2104_, new_n2105_,
    new_n2106_, new_n2107_, new_n2108_, new_n2109_, new_n2110_, new_n2111_,
    new_n2112_, new_n2113_, new_n2114_, new_n2115_, new_n2116_, new_n2117_,
    new_n2118_, new_n2119_, new_n2120_, new_n2121_, new_n2122_, new_n2123_,
    new_n2124_, new_n2125_, new_n2126_, new_n2127_, new_n2128_, new_n2129_,
    new_n2130_, new_n2131_, new_n2132_, new_n2133_, new_n2134_, new_n2135_,
    new_n2136_, new_n2137_, new_n2138_, new_n2139_, new_n2140_, new_n2141_,
    new_n2142_, new_n2143_, new_n2144_, new_n2145_, new_n2146_, new_n2147_,
    new_n2148_, new_n2149_, new_n2150_, new_n2151_, new_n2152_, new_n2153_,
    new_n2154_, new_n2155_, new_n2156_, new_n2157_, new_n2158_, new_n2159_,
    new_n2160_, new_n2161_, new_n2162_, new_n2163_, new_n2164_, new_n2165_,
    new_n2166_, new_n2167_, new_n2168_, new_n2169_, new_n2170_, new_n2171_,
    new_n2172_, new_n2173_, new_n2174_, new_n2175_, new_n2176_, new_n2177_,
    new_n2178_, new_n2179_, new_n2180_, new_n2181_, new_n2182_, new_n2183_,
    new_n2184_, new_n2185_, new_n2186_, new_n2187_, new_n2188_, new_n2189_,
    new_n2190_, new_n2191_, new_n2192_, new_n2193_, new_n2194_, new_n2195_,
    new_n2196_, new_n2197_, new_n2198_, new_n2199_, new_n2200_, new_n2201_,
    new_n2202_, new_n2203_, new_n2204_, new_n2205_, new_n2206_, new_n2207_,
    new_n2208_, new_n2209_, new_n2210_, new_n2211_, new_n2212_, new_n2213_,
    new_n2214_, new_n2215_, new_n2216_, new_n2217_, new_n2218_, new_n2219_,
    new_n2220_, new_n2221_, new_n2222_, new_n2223_, new_n2224_, new_n2225_,
    new_n2226_, new_n2227_, new_n2228_, new_n2229_, new_n2230_, new_n2231_,
    new_n2232_, new_n2233_, new_n2234_, new_n2235_, new_n2236_, new_n2237_,
    new_n2238_, new_n2239_, new_n2240_, new_n2241_, new_n2242_, new_n2243_,
    new_n2244_, new_n2245_, new_n2246_, new_n2247_, new_n2248_, new_n2249_,
    new_n2250_, new_n2251_, new_n2252_, new_n2253_, new_n2254_, new_n2255_,
    new_n2256_, new_n2257_, new_n2258_, new_n2259_, new_n2260_, new_n2261_,
    new_n2262_, new_n2263_, new_n2265_, new_n2266_, new_n2267_, new_n2268_,
    new_n2269_, new_n2270_, new_n2271_, new_n2272_, new_n2273_, new_n2274_,
    new_n2275_, new_n2276_, new_n2277_, new_n2278_, new_n2279_, new_n2280_,
    new_n2281_, new_n2282_, new_n2283_, new_n2284_, new_n2285_, new_n2286_,
    new_n2287_, new_n2288_, new_n2289_, new_n2290_, new_n2291_, new_n2292_,
    new_n2293_, new_n2294_, new_n2295_, new_n2296_, new_n2297_, new_n2298_,
    new_n2299_, new_n2300_, new_n2301_, new_n2302_, new_n2303_, new_n2304_,
    new_n2305_, new_n2306_, new_n2307_, new_n2308_, new_n2309_, new_n2310_,
    new_n2311_, new_n2312_, new_n2313_, new_n2314_, new_n2315_, new_n2316_,
    new_n2317_, new_n2318_, new_n2319_, new_n2320_, new_n2321_, new_n2322_,
    new_n2323_, new_n2324_, new_n2325_, new_n2326_, new_n2327_, new_n2328_,
    new_n2329_, new_n2330_, new_n2331_, new_n2332_, new_n2333_, new_n2334_,
    new_n2335_, new_n2336_, new_n2337_, new_n2338_, new_n2339_, new_n2340_,
    new_n2341_, new_n2342_, new_n2343_, new_n2344_, new_n2345_, new_n2346_,
    new_n2347_, new_n2348_, new_n2349_, new_n2350_, new_n2351_, new_n2352_,
    new_n2353_, new_n2354_, new_n2355_, new_n2356_, new_n2357_, new_n2358_,
    new_n2359_, new_n2360_, new_n2361_, new_n2362_, new_n2363_, new_n2364_,
    new_n2365_, new_n2366_, new_n2367_, new_n2368_, new_n2369_, new_n2370_,
    new_n2371_, new_n2372_, new_n2373_, new_n2374_, new_n2375_, new_n2376_,
    new_n2377_, new_n2378_, new_n2379_, new_n2380_, new_n2381_, new_n2382_,
    new_n2383_, new_n2384_, new_n2385_, new_n2386_, new_n2387_, new_n2388_,
    new_n2389_, new_n2390_, new_n2391_, new_n2392_, new_n2393_, new_n2394_,
    new_n2395_, new_n2396_, new_n2397_, new_n2398_, new_n2399_, new_n2400_,
    new_n2401_, new_n2402_, new_n2403_, new_n2404_, new_n2405_, new_n2406_,
    new_n2407_, new_n2408_, new_n2409_, new_n2410_, new_n2411_, new_n2412_,
    new_n2413_, new_n2414_, new_n2415_, new_n2416_, new_n2417_, new_n2418_,
    new_n2419_, new_n2420_, new_n2421_, new_n2422_, new_n2423_, new_n2424_,
    new_n2425_, new_n2426_, new_n2427_, new_n2428_, new_n2429_, new_n2430_,
    new_n2431_, new_n2432_, new_n2433_, new_n2434_, new_n2435_, new_n2436_,
    new_n2437_, new_n2438_, new_n2439_, new_n2440_, new_n2441_, new_n2442_,
    new_n2443_, new_n2444_, new_n2445_, new_n2446_, new_n2447_, new_n2448_,
    new_n2449_, new_n2450_, new_n2451_, new_n2452_, new_n2453_, new_n2454_,
    new_n2455_, new_n2456_, new_n2457_, new_n2458_, new_n2459_, new_n2460_,
    new_n2461_, new_n2462_, new_n2463_, new_n2464_, new_n2465_, new_n2466_,
    new_n2467_, new_n2468_, new_n2469_, new_n2470_, new_n2471_, new_n2472_,
    new_n2473_, new_n2474_, new_n2475_, new_n2476_, new_n2477_, new_n2478_,
    new_n2479_, new_n2480_, new_n2481_, new_n2482_, new_n2483_, new_n2484_,
    new_n2485_, new_n2486_, new_n2487_, new_n2488_, new_n2489_, new_n2490_,
    new_n2491_, new_n2492_, new_n2493_, new_n2494_, new_n2495_, new_n2496_,
    new_n2497_, new_n2498_, new_n2499_, new_n2500_, new_n2501_, new_n2503_,
    new_n2504_, new_n2505_, new_n2506_, new_n2507_, new_n2508_, new_n2509_,
    new_n2510_, new_n2511_, new_n2512_, new_n2513_, new_n2514_, new_n2515_,
    new_n2516_, new_n2517_, new_n2518_, new_n2519_, new_n2520_, new_n2521_,
    new_n2522_, new_n2523_, new_n2524_, new_n2525_, new_n2526_, new_n2527_,
    new_n2528_, new_n2529_, new_n2530_, new_n2531_, new_n2532_, new_n2533_,
    new_n2534_, new_n2535_, new_n2536_, new_n2537_, new_n2538_, new_n2539_,
    new_n2540_, new_n2541_, new_n2542_, new_n2543_, new_n2544_, new_n2545_,
    new_n2546_, new_n2547_, new_n2548_, new_n2549_, new_n2550_, new_n2551_,
    new_n2552_, new_n2553_, new_n2554_, new_n2555_, new_n2556_, new_n2557_,
    new_n2558_, new_n2559_, new_n2560_, new_n2561_, new_n2562_, new_n2563_,
    new_n2564_, new_n2565_, new_n2566_, new_n2567_, new_n2568_, new_n2569_,
    new_n2570_, new_n2571_, new_n2572_, new_n2573_, new_n2574_, new_n2575_,
    new_n2576_, new_n2577_, new_n2578_, new_n2579_, new_n2580_, new_n2581_,
    new_n2582_, new_n2583_, new_n2584_, new_n2585_, new_n2586_, new_n2587_,
    new_n2588_, new_n2589_, new_n2590_, new_n2591_, new_n2592_, new_n2593_,
    new_n2594_, new_n2595_, new_n2596_, new_n2597_, new_n2598_, new_n2599_,
    new_n2600_, new_n2601_, new_n2602_, new_n2603_, new_n2604_, new_n2605_,
    new_n2606_, new_n2607_, new_n2608_, new_n2609_, new_n2610_, new_n2611_,
    new_n2612_, new_n2613_, new_n2614_, new_n2615_, new_n2616_, new_n2617_,
    new_n2618_, new_n2619_, new_n2620_, new_n2621_, new_n2622_, new_n2623_,
    new_n2624_, new_n2625_, new_n2626_, new_n2627_, new_n2628_, new_n2629_,
    new_n2630_, new_n2631_, new_n2632_, new_n2633_, new_n2634_, new_n2635_,
    new_n2636_, new_n2637_, new_n2638_, new_n2639_, new_n2640_, new_n2641_,
    new_n2642_, new_n2643_, new_n2644_, new_n2645_, new_n2646_, new_n2647_,
    new_n2648_, new_n2649_, new_n2650_, new_n2651_, new_n2652_, new_n2653_,
    new_n2654_, new_n2655_, new_n2656_, new_n2657_, new_n2658_, new_n2659_,
    new_n2660_, new_n2661_, new_n2662_, new_n2663_, new_n2664_, new_n2665_,
    new_n2666_, new_n2667_, new_n2668_, new_n2669_, new_n2670_, new_n2671_,
    new_n2672_, new_n2673_, new_n2674_, new_n2675_, new_n2676_, new_n2677_,
    new_n2678_, new_n2679_, new_n2680_, new_n2681_, new_n2682_, new_n2683_,
    new_n2684_, new_n2685_, new_n2686_, new_n2687_, new_n2688_, new_n2689_,
    new_n2690_, new_n2691_, new_n2692_, new_n2693_, new_n2694_, new_n2695_,
    new_n2696_, new_n2697_, new_n2698_, new_n2699_, new_n2700_, new_n2701_,
    new_n2702_, new_n2703_, new_n2704_, new_n2705_, new_n2706_, new_n2707_,
    new_n2708_, new_n2709_, new_n2710_, new_n2711_, new_n2712_, new_n2713_,
    new_n2714_, new_n2715_, new_n2716_, new_n2717_, new_n2718_, new_n2719_,
    new_n2720_, new_n2721_, new_n2722_, new_n2723_, new_n2724_, new_n2725_,
    new_n2726_, new_n2727_, new_n2728_, new_n2729_, new_n2730_, new_n2731_,
    new_n2732_, new_n2733_, new_n2734_, new_n2735_, new_n2736_, new_n2737_,
    new_n2738_, new_n2739_, new_n2740_, new_n2741_, new_n2742_, new_n2743_,
    new_n2744_, new_n2745_, new_n2746_, new_n2747_, new_n2749_, new_n2750_,
    new_n2751_, new_n2752_, new_n2753_, new_n2754_, new_n2755_, new_n2756_,
    new_n2757_, new_n2758_, new_n2759_, new_n2760_, new_n2761_, new_n2762_,
    new_n2763_, new_n2764_, new_n2765_, new_n2766_, new_n2767_, new_n2768_,
    new_n2769_, new_n2770_, new_n2771_, new_n2772_, new_n2773_, new_n2774_,
    new_n2775_, new_n2776_, new_n2777_, new_n2778_, new_n2779_, new_n2780_,
    new_n2781_, new_n2782_, new_n2783_, new_n2784_, new_n2785_, new_n2786_,
    new_n2787_, new_n2788_, new_n2789_, new_n2790_, new_n2791_, new_n2792_,
    new_n2793_, new_n2794_, new_n2795_, new_n2796_, new_n2797_, new_n2798_,
    new_n2799_, new_n2800_, new_n2801_, new_n2802_, new_n2803_, new_n2804_,
    new_n2805_, new_n2806_, new_n2807_, new_n2808_, new_n2809_, new_n2810_,
    new_n2811_, new_n2812_, new_n2813_, new_n2814_, new_n2815_, new_n2816_,
    new_n2817_, new_n2818_, new_n2819_, new_n2820_, new_n2821_, new_n2822_,
    new_n2823_, new_n2824_, new_n2825_, new_n2826_, new_n2827_, new_n2828_,
    new_n2829_, new_n2830_, new_n2831_, new_n2832_, new_n2833_, new_n2834_,
    new_n2835_, new_n2836_, new_n2837_, new_n2838_, new_n2839_, new_n2840_,
    new_n2841_, new_n2842_, new_n2843_, new_n2844_, new_n2845_, new_n2846_,
    new_n2847_, new_n2848_, new_n2849_, new_n2850_, new_n2851_, new_n2852_,
    new_n2853_, new_n2854_, new_n2855_, new_n2856_, new_n2857_, new_n2858_,
    new_n2859_, new_n2860_, new_n2861_, new_n2862_, new_n2863_, new_n2864_,
    new_n2865_, new_n2866_, new_n2867_, new_n2868_, new_n2869_, new_n2870_,
    new_n2871_, new_n2872_, new_n2873_, new_n2874_, new_n2875_, new_n2876_,
    new_n2877_, new_n2878_, new_n2879_, new_n2880_, new_n2881_, new_n2882_,
    new_n2883_, new_n2884_, new_n2885_, new_n2886_, new_n2887_, new_n2888_,
    new_n2889_, new_n2890_, new_n2891_, new_n2892_, new_n2893_, new_n2894_,
    new_n2895_, new_n2896_, new_n2897_, new_n2898_, new_n2899_, new_n2900_,
    new_n2901_, new_n2902_, new_n2903_, new_n2904_, new_n2905_, new_n2906_,
    new_n2907_, new_n2908_, new_n2909_, new_n2910_, new_n2911_, new_n2912_,
    new_n2913_, new_n2914_, new_n2915_, new_n2916_, new_n2917_, new_n2918_,
    new_n2919_, new_n2920_, new_n2921_, new_n2922_, new_n2923_, new_n2924_,
    new_n2925_, new_n2926_, new_n2927_, new_n2928_, new_n2929_, new_n2930_,
    new_n2931_, new_n2932_, new_n2933_, new_n2934_, new_n2935_, new_n2936_,
    new_n2937_, new_n2938_, new_n2939_, new_n2940_, new_n2941_, new_n2942_,
    new_n2943_, new_n2944_, new_n2945_, new_n2946_, new_n2947_, new_n2948_,
    new_n2949_, new_n2950_, new_n2951_, new_n2952_, new_n2953_, new_n2954_,
    new_n2955_, new_n2956_, new_n2957_, new_n2958_, new_n2959_, new_n2960_,
    new_n2961_, new_n2962_, new_n2963_, new_n2964_, new_n2965_, new_n2966_,
    new_n2967_, new_n2968_, new_n2969_, new_n2970_, new_n2971_, new_n2972_,
    new_n2973_, new_n2974_, new_n2975_, new_n2976_, new_n2977_, new_n2978_,
    new_n2979_, new_n2980_, new_n2981_, new_n2982_, new_n2983_, new_n2984_,
    new_n2985_, new_n2986_, new_n2987_, new_n2988_, new_n2989_, new_n2990_,
    new_n2991_, new_n2992_, new_n2993_, new_n2994_, new_n2995_, new_n2996_,
    new_n2997_, new_n2998_, new_n2999_, new_n3000_, new_n3001_, new_n3002_,
    new_n3003_, new_n3004_, new_n3005_, new_n3006_, new_n3007_, new_n3008_,
    new_n3009_, new_n3010_, new_n3011_, new_n3012_, new_n3013_, new_n3014_,
    new_n3015_, new_n3016_, new_n3017_, new_n3018_, new_n3019_, new_n3020_,
    new_n3021_, new_n3022_, new_n3023_, new_n3024_, new_n3025_, new_n3026_,
    new_n3027_, new_n3028_, new_n3029_, new_n3030_, new_n3031_, new_n3032_,
    new_n3033_, new_n3034_, new_n3035_, new_n3036_, new_n3037_, new_n3038_,
    new_n3039_, new_n3040_, new_n3041_, new_n3042_, new_n3043_, new_n3044_,
    new_n3045_, new_n3046_, new_n3047_, new_n3048_, new_n3049_, new_n3050_,
    new_n3051_, new_n3052_, new_n3053_, new_n3054_, new_n3055_, new_n3056_,
    new_n3057_, new_n3058_, new_n3059_, new_n3060_, new_n3061_, new_n3062_,
    new_n3063_, new_n3064_, new_n3065_, new_n3066_, new_n3067_, new_n3068_,
    new_n3069_, new_n3070_, new_n3071_, new_n3072_, new_n3073_, new_n3074_,
    new_n3075_, new_n3076_, new_n3077_, new_n3078_, new_n3079_, new_n3080_,
    new_n3081_, new_n3082_, new_n3083_, new_n3084_, new_n3085_, new_n3087_,
    new_n3088_, new_n3089_, new_n3090_, new_n3091_, new_n3092_, new_n3093_,
    new_n3094_, new_n3095_, new_n3096_, new_n3097_, new_n3098_, new_n3099_,
    new_n3100_, new_n3101_, new_n3102_, new_n3103_, new_n3104_, new_n3105_,
    new_n3106_, new_n3107_, new_n3108_, new_n3109_, new_n3110_, new_n3111_,
    new_n3112_, new_n3113_, new_n3114_, new_n3115_, new_n3116_, new_n3117_,
    new_n3118_, new_n3119_, new_n3120_, new_n3121_, new_n3122_, new_n3123_,
    new_n3124_, new_n3125_, new_n3126_, new_n3127_, new_n3128_, new_n3129_,
    new_n3130_, new_n3131_, new_n3132_, new_n3133_, new_n3134_, new_n3135_,
    new_n3136_, new_n3137_, new_n3138_, new_n3139_, new_n3140_, new_n3141_,
    new_n3142_, new_n3143_, new_n3144_, new_n3145_, new_n3146_, new_n3147_,
    new_n3148_, new_n3149_, new_n3150_, new_n3151_, new_n3152_, new_n3153_,
    new_n3154_, new_n3155_, new_n3156_, new_n3157_, new_n3158_, new_n3159_,
    new_n3160_, new_n3161_, new_n3162_, new_n3163_, new_n3164_, new_n3165_,
    new_n3166_, new_n3167_, new_n3168_, new_n3169_, new_n3170_, new_n3171_,
    new_n3172_, new_n3173_, new_n3174_, new_n3175_, new_n3176_, new_n3177_,
    new_n3178_, new_n3179_, new_n3180_, new_n3181_, new_n3182_, new_n3183_,
    new_n3184_, new_n3185_, new_n3186_, new_n3187_, new_n3188_, new_n3189_,
    new_n3190_, new_n3191_, new_n3192_, new_n3193_, new_n3194_, new_n3195_,
    new_n3196_, new_n3197_, new_n3198_, new_n3199_, new_n3200_, new_n3201_,
    new_n3202_, new_n3203_, new_n3204_, new_n3205_, new_n3206_, new_n3207_,
    new_n3208_, new_n3209_, new_n3210_, new_n3211_, new_n3212_, new_n3213_,
    new_n3214_, new_n3215_, new_n3216_, new_n3217_, new_n3218_, new_n3219_,
    new_n3220_, new_n3221_, new_n3222_, new_n3223_, new_n3224_, new_n3225_,
    new_n3226_, new_n3227_, new_n3228_, new_n3229_, new_n3230_, new_n3231_,
    new_n3232_, new_n3233_, new_n3234_, new_n3235_, new_n3236_, new_n3237_,
    new_n3238_, new_n3239_, new_n3240_, new_n3241_, new_n3242_, new_n3243_,
    new_n3244_, new_n3245_, new_n3246_, new_n3247_, new_n3248_, new_n3249_,
    new_n3250_, new_n3251_, new_n3252_, new_n3253_, new_n3254_, new_n3255_,
    new_n3256_, new_n3257_, new_n3258_, new_n3259_, new_n3260_, new_n3261_,
    new_n3262_, new_n3263_, new_n3264_, new_n3265_, new_n3266_, new_n3267_,
    new_n3268_, new_n3269_, new_n3270_, new_n3271_, new_n3272_, new_n3273_,
    new_n3274_, new_n3275_, new_n3276_, new_n3277_, new_n3278_, new_n3279_,
    new_n3280_, new_n3281_, new_n3282_, new_n3283_, new_n3284_, new_n3285_,
    new_n3286_, new_n3287_, new_n3288_, new_n3289_, new_n3290_, new_n3291_,
    new_n3292_, new_n3293_, new_n3294_, new_n3295_, new_n3296_, new_n3297_,
    new_n3298_, new_n3299_, new_n3300_, new_n3301_, new_n3302_, new_n3303_,
    new_n3304_, new_n3305_, new_n3307_, new_n3308_, new_n3309_, new_n3310_,
    new_n3311_, new_n3312_, new_n3313_, new_n3314_, new_n3315_, new_n3316_,
    new_n3317_, new_n3318_, new_n3319_, new_n3320_, new_n3321_, new_n3322_,
    new_n3323_, new_n3324_, new_n3325_, new_n3326_, new_n3327_, new_n3328_,
    new_n3329_, new_n3330_, new_n3331_, new_n3332_, new_n3333_, new_n3334_,
    new_n3335_, new_n3336_, new_n3337_, new_n3338_, new_n3339_, new_n3340_,
    new_n3341_, new_n3342_, new_n3343_, new_n3344_, new_n3345_, new_n3346_,
    new_n3347_, new_n3348_, new_n3349_, new_n3350_, new_n3351_, new_n3352_,
    new_n3353_, new_n3354_, new_n3355_, new_n3356_, new_n3357_, new_n3358_,
    new_n3359_, new_n3360_, new_n3361_, new_n3362_, new_n3363_, new_n3364_,
    new_n3365_, new_n3366_, new_n3367_, new_n3368_, new_n3369_, new_n3370_,
    new_n3371_, new_n3372_, new_n3373_, new_n3374_, new_n3375_, new_n3376_,
    new_n3377_, new_n3378_, new_n3379_, new_n3380_, new_n3381_, new_n3382_,
    new_n3383_, new_n3384_, new_n3385_, new_n3386_, new_n3387_, new_n3388_,
    new_n3389_, new_n3390_, new_n3391_, new_n3392_, new_n3393_, new_n3394_,
    new_n3395_, new_n3396_, new_n3397_, new_n3398_, new_n3399_, new_n3400_,
    new_n3401_, new_n3402_, new_n3403_, new_n3404_, new_n3405_, new_n3406_,
    new_n3407_, new_n3408_, new_n3409_, new_n3410_, new_n3411_, new_n3412_,
    new_n3413_, new_n3414_, new_n3415_, new_n3416_, new_n3417_, new_n3418_,
    new_n3419_, new_n3420_, new_n3421_, new_n3422_, new_n3423_, new_n3424_,
    new_n3425_, new_n3426_, new_n3427_, new_n3428_, new_n3429_, new_n3430_,
    new_n3431_, new_n3432_, new_n3433_, new_n3434_, new_n3435_, new_n3436_,
    new_n3437_, new_n3438_, new_n3439_, new_n3440_, new_n3441_, new_n3442_,
    new_n3443_, new_n3444_, new_n3445_, new_n3446_, new_n3447_, new_n3448_,
    new_n3449_, new_n3450_, new_n3451_, new_n3452_, new_n3453_, new_n3454_,
    new_n3455_, new_n3456_, new_n3457_, new_n3458_, new_n3459_, new_n3460_,
    new_n3461_, new_n3462_, new_n3463_, new_n3464_, new_n3465_, new_n3466_,
    new_n3467_, new_n3468_, new_n3469_, new_n3470_, new_n3471_, new_n3472_,
    new_n3473_, new_n3474_, new_n3475_, new_n3476_, new_n3477_, new_n3478_,
    new_n3479_, new_n3480_, new_n3481_, new_n3482_, new_n3483_, new_n3484_,
    new_n3485_, new_n3486_, new_n3487_, new_n3488_, new_n3489_, new_n3490_,
    new_n3491_, new_n3492_, new_n3493_, new_n3494_, new_n3495_, new_n3496_,
    new_n3497_, new_n3498_, new_n3499_, new_n3500_, new_n3501_, new_n3502_,
    new_n3503_, new_n3504_, new_n3505_, new_n3506_, new_n3507_, new_n3508_,
    new_n3509_, new_n3510_, new_n3511_, new_n3512_, new_n3513_, new_n3514_,
    new_n3515_, new_n3516_, new_n3517_, new_n3518_, new_n3519_, new_n3520_,
    new_n3521_, new_n3522_, new_n3523_, new_n3524_, new_n3525_, new_n3526_,
    new_n3527_, new_n3528_, new_n3529_, new_n3530_, new_n3531_, new_n3532_,
    new_n3533_, new_n3534_, new_n3535_, new_n3536_, new_n3537_, new_n3538_,
    new_n3539_, new_n3540_, new_n3541_, new_n3542_, new_n3543_, new_n3544_,
    new_n3545_, new_n3546_, new_n3547_, new_n3548_, new_n3549_, new_n3550_,
    new_n3551_, new_n3552_, new_n3553_, new_n3554_, new_n3555_, new_n3556_,
    new_n3557_, new_n3558_, new_n3559_, new_n3560_, new_n3561_, new_n3562_,
    new_n3563_, new_n3564_, new_n3565_, new_n3566_, new_n3567_, new_n3568_,
    new_n3569_, new_n3570_, new_n3571_, new_n3572_, new_n3573_, new_n3574_,
    new_n3575_, new_n3576_, new_n3577_, new_n3578_, new_n3579_, new_n3580_,
    new_n3581_, new_n3582_, new_n3583_, new_n3584_, new_n3585_, new_n3586_,
    new_n3587_, new_n3588_, new_n3590_, new_n3591_, new_n3592_, new_n3593_,
    new_n3594_, new_n3595_, new_n3596_, new_n3597_, new_n3598_, new_n3599_,
    new_n3600_, new_n3601_, new_n3602_, new_n3603_, new_n3604_, new_n3605_,
    new_n3606_, new_n3607_, new_n3608_, new_n3609_, new_n3610_, new_n3611_,
    new_n3612_, new_n3613_, new_n3614_, new_n3615_, new_n3616_, new_n3617_,
    new_n3618_, new_n3619_, new_n3620_, new_n3621_, new_n3622_, new_n3623_,
    new_n3624_, new_n3625_, new_n3626_, new_n3627_, new_n3628_, new_n3629_,
    new_n3630_, new_n3631_, new_n3632_, new_n3633_, new_n3634_, new_n3635_,
    new_n3636_, new_n3637_, new_n3638_, new_n3639_, new_n3640_, new_n3641_,
    new_n3642_, new_n3643_, new_n3644_, new_n3645_, new_n3646_, new_n3647_,
    new_n3648_, new_n3649_, new_n3650_, new_n3651_, new_n3652_, new_n3653_,
    new_n3654_, new_n3655_, new_n3656_, new_n3657_, new_n3658_, new_n3659_,
    new_n3660_, new_n3661_, new_n3662_, new_n3663_, new_n3664_, new_n3665_,
    new_n3666_, new_n3667_, new_n3668_, new_n3669_, new_n3670_, new_n3671_,
    new_n3672_, new_n3673_, new_n3674_, new_n3675_, new_n3676_, new_n3677_,
    new_n3678_, new_n3679_, new_n3680_, new_n3681_, new_n3682_, new_n3683_,
    new_n3684_, new_n3685_, new_n3686_, new_n3687_, new_n3688_, new_n3689_,
    new_n3690_, new_n3691_, new_n3692_, new_n3693_, new_n3694_, new_n3695_,
    new_n3696_, new_n3697_, new_n3698_, new_n3699_, new_n3700_, new_n3701_,
    new_n3702_, new_n3703_, new_n3704_, new_n3705_, new_n3706_, new_n3707_,
    new_n3708_, new_n3709_, new_n3710_, new_n3711_, new_n3712_, new_n3713_,
    new_n3714_, new_n3715_, new_n3716_, new_n3717_, new_n3718_, new_n3719_,
    new_n3720_, new_n3721_, new_n3722_, new_n3723_, new_n3724_, new_n3725_,
    new_n3726_, new_n3727_, new_n3728_, new_n3729_, new_n3730_, new_n3731_,
    new_n3732_, new_n3733_, new_n3734_, new_n3735_, new_n3736_, new_n3737_,
    new_n3738_, new_n3739_, new_n3740_, new_n3741_, new_n3742_, new_n3743_,
    new_n3744_, new_n3745_, new_n3746_, new_n3747_, new_n3748_, new_n3749_,
    new_n3750_, new_n3751_, new_n3752_, new_n3753_, new_n3754_, new_n3755_,
    new_n3756_, new_n3757_, new_n3758_, new_n3759_, new_n3760_, new_n3761_,
    new_n3762_, new_n3763_, new_n3764_, new_n3765_, new_n3766_, new_n3767_,
    new_n3768_, new_n3769_, new_n3770_, new_n3771_, new_n3772_, new_n3773_,
    new_n3774_, new_n3775_, new_n3776_, new_n3777_, new_n3778_, new_n3779_,
    new_n3780_, new_n3781_, new_n3782_, new_n3783_, new_n3784_, new_n3785_,
    new_n3786_, new_n3787_, new_n3788_, new_n3789_, new_n3790_, new_n3791_,
    new_n3792_, new_n3793_, new_n3794_, new_n3795_, new_n3796_, new_n3797_,
    new_n3798_, new_n3799_, new_n3800_, new_n3801_, new_n3802_, new_n3803_,
    new_n3804_, new_n3805_, new_n3806_, new_n3807_, new_n3808_, new_n3809_,
    new_n3810_, new_n3811_, new_n3812_, new_n3813_, new_n3814_, new_n3815_,
    new_n3816_, new_n3817_, new_n3818_, new_n3819_, new_n3820_, new_n3821_,
    new_n3822_, new_n3823_, new_n3824_, new_n3825_, new_n3826_, new_n3827_,
    new_n3828_, new_n3829_, new_n3830_, new_n3831_, new_n3832_, new_n3833_,
    new_n3834_, new_n3835_, new_n3836_, new_n3837_, new_n3838_, new_n3839_,
    new_n3840_, new_n3841_, new_n3842_, new_n3843_, new_n3844_, new_n3845_,
    new_n3846_, new_n3847_, new_n3848_, new_n3849_, new_n3850_, new_n3851_,
    new_n3852_, new_n3853_, new_n3854_, new_n3855_, new_n3856_, new_n3857_,
    new_n3858_, new_n3859_, new_n3860_, new_n3861_, new_n3862_, new_n3863_,
    new_n3865_, new_n3866_, new_n3867_, new_n3868_, new_n3869_, new_n3870_,
    new_n3871_, new_n3872_, new_n3873_, new_n3874_, new_n3875_, new_n3876_,
    new_n3877_, new_n3878_, new_n3879_, new_n3880_, new_n3881_, new_n3882_,
    new_n3883_, new_n3884_, new_n3885_, new_n3886_, new_n3887_, new_n3888_,
    new_n3889_, new_n3890_, new_n3891_, new_n3892_, new_n3893_, new_n3894_,
    new_n3895_, new_n3896_, new_n3897_, new_n3898_, new_n3899_, new_n3900_,
    new_n3901_, new_n3902_, new_n3903_, new_n3904_, new_n3905_, new_n3906_,
    new_n3907_, new_n3908_, new_n3909_, new_n3910_, new_n3911_, new_n3912_,
    new_n3913_, new_n3914_, new_n3915_, new_n3916_, new_n3917_, new_n3918_,
    new_n3919_, new_n3920_, new_n3921_, new_n3922_, new_n3923_, new_n3924_,
    new_n3925_, new_n3926_, new_n3927_, new_n3928_, new_n3929_, new_n3930_,
    new_n3931_, new_n3932_, new_n3933_, new_n3934_, new_n3935_, new_n3936_,
    new_n3937_, new_n3938_, new_n3939_, new_n3940_, new_n3941_, new_n3942_,
    new_n3943_, new_n3944_, new_n3945_, new_n3946_, new_n3947_, new_n3948_,
    new_n3949_, new_n3950_, new_n3951_, new_n3952_, new_n3953_, new_n3954_,
    new_n3955_, new_n3956_, new_n3957_, new_n3958_, new_n3959_, new_n3960_,
    new_n3961_, new_n3962_, new_n3963_, new_n3964_, new_n3965_, new_n3966_,
    new_n3967_, new_n3968_, new_n3969_, new_n3970_, new_n3971_, new_n3972_,
    new_n3973_, new_n3974_, new_n3975_, new_n3976_, new_n3977_, new_n3978_,
    new_n3979_, new_n3980_, new_n3981_, new_n3982_, new_n3983_, new_n3984_,
    new_n3985_, new_n3986_, new_n3987_, new_n3988_, new_n3989_, new_n3990_,
    new_n3991_, new_n3992_, new_n3993_, new_n3994_, new_n3995_, new_n3996_,
    new_n3997_, new_n3998_, new_n3999_, new_n4000_, new_n4001_, new_n4002_,
    new_n4003_, new_n4004_, new_n4005_, new_n4006_, new_n4007_, new_n4008_,
    new_n4009_, new_n4010_, new_n4011_, new_n4012_, new_n4013_, new_n4014_,
    new_n4015_, new_n4016_, new_n4017_, new_n4018_, new_n4019_, new_n4020_,
    new_n4021_, new_n4022_, new_n4023_, new_n4024_, new_n4025_, new_n4026_,
    new_n4027_, new_n4028_, new_n4029_, new_n4030_, new_n4031_, new_n4032_,
    new_n4033_, new_n4034_, new_n4035_, new_n4036_, new_n4037_, new_n4038_,
    new_n4039_, new_n4040_, new_n4041_, new_n4042_, new_n4043_, new_n4044_,
    new_n4045_, new_n4046_, new_n4047_, new_n4048_, new_n4049_, new_n4050_,
    new_n4051_, new_n4052_, new_n4053_, new_n4054_, new_n4055_, new_n4056_,
    new_n4057_, new_n4058_, new_n4059_, new_n4060_, new_n4061_, new_n4062_,
    new_n4063_, new_n4064_, new_n4065_, new_n4066_, new_n4067_, new_n4068_,
    new_n4069_, new_n4070_, new_n4071_, new_n4072_, new_n4073_, new_n4074_,
    new_n4075_, new_n4076_, new_n4077_, new_n4078_, new_n4079_, new_n4080_,
    new_n4081_, new_n4082_, new_n4083_, new_n4084_, new_n4085_, new_n4086_,
    new_n4087_, new_n4088_, new_n4089_, new_n4090_, new_n4091_, new_n4092_,
    new_n4093_, new_n4094_, new_n4095_, new_n4096_, new_n4097_, new_n4098_,
    new_n4099_, new_n4100_, new_n4101_, new_n4102_, new_n4103_, new_n4104_,
    new_n4105_, new_n4106_, new_n4107_, new_n4108_, new_n4109_, new_n4110_,
    new_n4111_, new_n4112_, new_n4113_, new_n4114_, new_n4115_, new_n4116_,
    new_n4117_, new_n4118_, new_n4119_, new_n4120_, new_n4121_, new_n4122_,
    new_n4123_, new_n4124_, new_n4125_, new_n4126_, new_n4127_, new_n4128_,
    new_n4129_, new_n4130_, new_n4131_, new_n4132_, new_n4133_, new_n4134_,
    new_n4135_, new_n4136_, new_n4137_, new_n4138_, new_n4139_, new_n4140_,
    new_n4141_, new_n4142_, new_n4143_, new_n4144_, new_n4145_, new_n4146_,
    new_n4147_, new_n4148_, new_n4149_, new_n4150_, new_n4151_, new_n4152_,
    new_n4153_, new_n4154_, new_n4155_, new_n4156_, new_n4157_, new_n4158_,
    new_n4159_, new_n4160_, new_n4161_, new_n4162_, new_n4163_, new_n4164_,
    new_n4165_, new_n4167_, new_n4168_, new_n4169_, new_n4170_, new_n4171_,
    new_n4172_, new_n4173_, new_n4174_, new_n4175_, new_n4176_, new_n4177_,
    new_n4178_, new_n4179_, new_n4180_, new_n4181_, new_n4182_, new_n4183_,
    new_n4184_, new_n4185_, new_n4186_, new_n4187_, new_n4188_, new_n4189_,
    new_n4190_, new_n4191_, new_n4192_, new_n4193_, new_n4194_, new_n4195_,
    new_n4196_, new_n4197_, new_n4198_, new_n4199_, new_n4200_, new_n4201_,
    new_n4202_, new_n4203_, new_n4204_, new_n4205_, new_n4206_, new_n4207_,
    new_n4208_, new_n4209_, new_n4210_, new_n4211_, new_n4212_, new_n4213_,
    new_n4214_, new_n4215_, new_n4216_, new_n4217_, new_n4218_, new_n4219_,
    new_n4220_, new_n4221_, new_n4222_, new_n4223_, new_n4224_, new_n4225_,
    new_n4226_, new_n4227_, new_n4228_, new_n4229_, new_n4230_, new_n4231_,
    new_n4232_, new_n4233_, new_n4234_, new_n4235_, new_n4236_, new_n4237_,
    new_n4238_, new_n4239_, new_n4240_, new_n4241_, new_n4242_, new_n4243_,
    new_n4244_, new_n4245_, new_n4246_, new_n4247_, new_n4248_, new_n4249_,
    new_n4250_, new_n4251_, new_n4252_, new_n4253_, new_n4254_, new_n4255_,
    new_n4256_, new_n4257_, new_n4258_, new_n4259_, new_n4260_, new_n4261_,
    new_n4262_, new_n4263_, new_n4264_, new_n4265_, new_n4266_, new_n4267_,
    new_n4268_, new_n4269_, new_n4270_, new_n4271_, new_n4272_, new_n4273_,
    new_n4274_, new_n4275_, new_n4276_, new_n4277_, new_n4278_, new_n4279_,
    new_n4280_, new_n4281_, new_n4282_, new_n4283_, new_n4284_, new_n4285_,
    new_n4286_, new_n4287_, new_n4288_, new_n4289_, new_n4290_, new_n4291_,
    new_n4292_, new_n4293_, new_n4294_, new_n4295_, new_n4296_, new_n4297_,
    new_n4298_, new_n4299_, new_n4300_, new_n4301_, new_n4302_, new_n4303_,
    new_n4304_, new_n4305_, new_n4306_, new_n4307_, new_n4308_, new_n4309_,
    new_n4310_, new_n4311_, new_n4312_, new_n4313_, new_n4314_, new_n4315_,
    new_n4316_, new_n4317_, new_n4318_, new_n4319_, new_n4320_, new_n4321_,
    new_n4322_, new_n4323_, new_n4324_, new_n4325_, new_n4326_, new_n4327_,
    new_n4328_, new_n4329_, new_n4330_, new_n4331_, new_n4332_, new_n4333_,
    new_n4334_, new_n4335_, new_n4336_, new_n4337_, new_n4338_, new_n4339_,
    new_n4340_, new_n4341_, new_n4342_, new_n4343_, new_n4344_, new_n4345_,
    new_n4346_, new_n4347_, new_n4348_, new_n4349_, new_n4350_, new_n4351_,
    new_n4352_, new_n4353_, new_n4354_, new_n4355_, new_n4356_, new_n4357_,
    new_n4358_, new_n4359_, new_n4360_, new_n4361_, new_n4362_, new_n4363_,
    new_n4364_, new_n4365_, new_n4366_, new_n4367_, new_n4368_, new_n4369_,
    new_n4370_, new_n4371_, new_n4372_, new_n4373_, new_n4374_, new_n4375_,
    new_n4376_, new_n4377_, new_n4378_, new_n4379_, new_n4380_, new_n4381_,
    new_n4382_, new_n4383_, new_n4384_, new_n4385_, new_n4386_, new_n4387_,
    new_n4388_, new_n4389_, new_n4390_, new_n4391_, new_n4392_, new_n4393_,
    new_n4394_, new_n4395_, new_n4396_, new_n4397_, new_n4398_, new_n4399_,
    new_n4400_, new_n4401_, new_n4402_, new_n4403_, new_n4404_, new_n4405_,
    new_n4406_, new_n4407_, new_n4408_, new_n4409_, new_n4410_, new_n4411_,
    new_n4412_, new_n4413_, new_n4414_, new_n4415_, new_n4416_, new_n4417_,
    new_n4418_, new_n4419_, new_n4420_, new_n4421_, new_n4422_, new_n4423_,
    new_n4424_, new_n4425_, new_n4426_, new_n4427_, new_n4428_, new_n4429_,
    new_n4430_, new_n4431_, new_n4432_, new_n4433_, new_n4434_, new_n4435_,
    new_n4436_, new_n4437_, new_n4438_, new_n4439_, new_n4440_, new_n4441_,
    new_n4442_, new_n4443_, new_n4444_, new_n4445_, new_n4446_, new_n4447_,
    new_n4448_, new_n4449_, new_n4450_, new_n4451_, new_n4452_, new_n4453_,
    new_n4454_, new_n4455_, new_n4456_, new_n4457_, new_n4458_, new_n4459_,
    new_n4460_, new_n4461_, new_n4462_, new_n4463_, new_n4464_, new_n4465_,
    new_n4466_, new_n4467_, new_n4468_, new_n4469_, new_n4470_, new_n4471_,
    new_n4472_, new_n4473_, new_n4474_, new_n4475_, new_n4476_, new_n4477_,
    new_n4478_, new_n4479_, new_n4480_, new_n4481_, new_n4482_, new_n4483_,
    new_n4484_, new_n4485_, new_n4486_, new_n4487_, new_n4488_, new_n4489_,
    new_n4490_, new_n4491_, new_n4492_, new_n4493_, new_n4494_, new_n4495_,
    new_n4496_, new_n4497_, new_n4498_, new_n4499_, new_n4500_, new_n4501_,
    new_n4502_, new_n4503_, new_n4505_, new_n4506_, new_n4507_, new_n4508_,
    new_n4509_, new_n4510_, new_n4511_, new_n4512_, new_n4513_, new_n4514_,
    new_n4515_, new_n4516_, new_n4517_, new_n4518_, new_n4519_, new_n4520_,
    new_n4521_, new_n4522_, new_n4523_, new_n4524_, new_n4525_, new_n4526_,
    new_n4527_, new_n4528_, new_n4529_, new_n4530_, new_n4531_, new_n4532_,
    new_n4533_, new_n4534_, new_n4535_, new_n4536_, new_n4537_, new_n4538_,
    new_n4539_, new_n4540_, new_n4541_, new_n4542_, new_n4543_, new_n4544_,
    new_n4545_, new_n4546_, new_n4547_, new_n4548_, new_n4549_, new_n4550_,
    new_n4551_, new_n4552_, new_n4553_, new_n4554_, new_n4555_, new_n4556_,
    new_n4557_, new_n4558_, new_n4559_, new_n4560_, new_n4561_, new_n4562_,
    new_n4563_, new_n4564_, new_n4565_, new_n4566_, new_n4567_, new_n4568_,
    new_n4569_, new_n4570_, new_n4571_, new_n4572_, new_n4573_, new_n4574_,
    new_n4575_, new_n4576_, new_n4577_, new_n4578_, new_n4579_, new_n4580_,
    new_n4581_, new_n4582_, new_n4583_, new_n4584_, new_n4585_, new_n4586_,
    new_n4587_, new_n4588_, new_n4589_, new_n4590_, new_n4591_, new_n4592_,
    new_n4593_, new_n4594_, new_n4595_, new_n4596_, new_n4597_, new_n4598_,
    new_n4599_, new_n4600_, new_n4601_, new_n4602_, new_n4603_, new_n4604_,
    new_n4605_, new_n4606_, new_n4607_, new_n4608_, new_n4609_, new_n4610_,
    new_n4611_, new_n4612_, new_n4613_, new_n4614_, new_n4615_, new_n4616_,
    new_n4617_, new_n4618_, new_n4619_, new_n4620_, new_n4621_, new_n4622_,
    new_n4623_, new_n4624_, new_n4625_, new_n4626_, new_n4627_, new_n4628_,
    new_n4629_, new_n4630_, new_n4631_, new_n4632_, new_n4633_, new_n4634_,
    new_n4635_, new_n4636_, new_n4637_, new_n4638_, new_n4639_, new_n4640_,
    new_n4641_, new_n4642_, new_n4643_, new_n4644_, new_n4645_, new_n4646_,
    new_n4647_, new_n4648_, new_n4649_, new_n4650_, new_n4651_, new_n4652_,
    new_n4653_, new_n4654_, new_n4655_, new_n4656_, new_n4657_, new_n4658_,
    new_n4659_, new_n4660_, new_n4661_, new_n4662_, new_n4663_, new_n4664_,
    new_n4665_, new_n4666_, new_n4667_, new_n4668_, new_n4669_, new_n4670_,
    new_n4671_, new_n4672_, new_n4673_, new_n4674_, new_n4675_, new_n4676_,
    new_n4677_, new_n4678_, new_n4679_, new_n4680_, new_n4681_, new_n4682_,
    new_n4683_, new_n4684_, new_n4685_, new_n4686_, new_n4687_, new_n4688_,
    new_n4689_, new_n4690_, new_n4691_, new_n4692_, new_n4693_, new_n4694_,
    new_n4695_, new_n4696_, new_n4697_, new_n4698_, new_n4699_, new_n4700_,
    new_n4701_, new_n4702_, new_n4703_, new_n4704_, new_n4705_, new_n4706_,
    new_n4707_, new_n4708_, new_n4709_, new_n4710_, new_n4711_, new_n4712_,
    new_n4713_, new_n4714_, new_n4715_, new_n4716_, new_n4717_, new_n4718_,
    new_n4719_, new_n4720_, new_n4721_, new_n4722_, new_n4723_, new_n4724_,
    new_n4725_, new_n4726_, new_n4727_, new_n4728_, new_n4729_, new_n4730_,
    new_n4731_, new_n4732_, new_n4733_, new_n4734_, new_n4735_, new_n4736_,
    new_n4737_, new_n4738_, new_n4739_, new_n4740_, new_n4741_, new_n4742_,
    new_n4743_, new_n4744_, new_n4745_, new_n4746_, new_n4747_, new_n4748_,
    new_n4749_, new_n4750_, new_n4751_, new_n4752_, new_n4753_, new_n4754_,
    new_n4755_, new_n4756_, new_n4757_, new_n4758_, new_n4759_, new_n4760_,
    new_n4761_, new_n4762_, new_n4763_, new_n4764_, new_n4765_, new_n4766_,
    new_n4767_, new_n4768_, new_n4769_, new_n4770_, new_n4771_, new_n4772_,
    new_n4773_, new_n4774_, new_n4775_, new_n4776_, new_n4777_, new_n4778_,
    new_n4779_, new_n4780_, new_n4781_, new_n4782_, new_n4783_, new_n4784_,
    new_n4785_, new_n4786_, new_n4787_, new_n4788_, new_n4789_, new_n4790_,
    new_n4791_, new_n4792_, new_n4793_, new_n4794_, new_n4795_, new_n4796_,
    new_n4797_, new_n4798_, new_n4799_, new_n4800_, new_n4801_, new_n4802_,
    new_n4803_, new_n4804_, new_n4805_, new_n4806_, new_n4807_, new_n4808_,
    new_n4809_, new_n4810_, new_n4811_, new_n4812_, new_n4813_, new_n4814_,
    new_n4815_, new_n4816_, new_n4817_, new_n4818_, new_n4819_, new_n4820_,
    new_n4821_, new_n4822_, new_n4823_, new_n4824_, new_n4825_, new_n4826_,
    new_n4828_, new_n4829_, new_n4830_, new_n4831_, new_n4832_, new_n4833_,
    new_n4834_, new_n4835_, new_n4836_, new_n4837_, new_n4838_, new_n4839_,
    new_n4840_, new_n4841_, new_n4842_, new_n4843_, new_n4844_, new_n4845_,
    new_n4846_, new_n4847_, new_n4848_, new_n4849_, new_n4850_, new_n4851_,
    new_n4852_, new_n4853_, new_n4854_, new_n4855_, new_n4856_, new_n4857_,
    new_n4858_, new_n4859_, new_n4860_, new_n4861_, new_n4862_, new_n4863_,
    new_n4864_, new_n4865_, new_n4866_, new_n4867_, new_n4868_, new_n4869_,
    new_n4870_, new_n4871_, new_n4872_, new_n4873_, new_n4874_, new_n4875_,
    new_n4876_, new_n4877_, new_n4878_, new_n4879_, new_n4880_, new_n4881_,
    new_n4882_, new_n4883_, new_n4884_, new_n4885_, new_n4886_, new_n4887_,
    new_n4888_, new_n4889_, new_n4890_, new_n4891_, new_n4892_, new_n4893_,
    new_n4894_, new_n4895_, new_n4896_, new_n4897_, new_n4898_, new_n4899_,
    new_n4900_, new_n4901_, new_n4902_, new_n4903_, new_n4904_, new_n4905_,
    new_n4906_, new_n4907_, new_n4908_, new_n4909_, new_n4910_, new_n4911_,
    new_n4912_, new_n4913_, new_n4914_, new_n4915_, new_n4916_, new_n4917_,
    new_n4918_, new_n4919_, new_n4920_, new_n4921_, new_n4922_, new_n4923_,
    new_n4924_, new_n4925_, new_n4926_, new_n4927_, new_n4928_, new_n4929_,
    new_n4930_, new_n4931_, new_n4932_, new_n4933_, new_n4934_, new_n4935_,
    new_n4936_, new_n4937_, new_n4938_, new_n4939_, new_n4940_, new_n4941_,
    new_n4942_, new_n4943_, new_n4944_, new_n4945_, new_n4946_, new_n4947_,
    new_n4948_, new_n4949_, new_n4950_, new_n4951_, new_n4952_, new_n4953_,
    new_n4954_, new_n4955_, new_n4956_, new_n4957_, new_n4958_, new_n4959_,
    new_n4960_, new_n4961_, new_n4962_, new_n4963_, new_n4964_, new_n4965_,
    new_n4966_, new_n4967_, new_n4968_, new_n4969_, new_n4970_, new_n4971_,
    new_n4972_, new_n4973_, new_n4974_, new_n4975_, new_n4976_, new_n4977_,
    new_n4978_, new_n4979_, new_n4980_, new_n4981_, new_n4982_, new_n4983_,
    new_n4984_, new_n4985_, new_n4986_, new_n4987_, new_n4988_, new_n4989_,
    new_n4990_, new_n4991_, new_n4992_, new_n4993_, new_n4994_, new_n4995_,
    new_n4996_, new_n4997_, new_n4998_, new_n4999_, new_n5000_, new_n5001_,
    new_n5002_, new_n5003_, new_n5004_, new_n5005_, new_n5006_, new_n5007_,
    new_n5008_, new_n5009_, new_n5010_, new_n5011_, new_n5012_, new_n5013_,
    new_n5014_, new_n5015_, new_n5016_, new_n5017_, new_n5018_, new_n5019_,
    new_n5020_, new_n5021_, new_n5022_, new_n5023_, new_n5024_, new_n5025_,
    new_n5026_, new_n5027_, new_n5028_, new_n5029_, new_n5030_, new_n5031_,
    new_n5032_, new_n5033_, new_n5034_, new_n5035_, new_n5036_, new_n5037_,
    new_n5038_, new_n5039_, new_n5040_, new_n5041_, new_n5042_, new_n5043_,
    new_n5044_, new_n5045_, new_n5046_, new_n5047_, new_n5048_, new_n5049_,
    new_n5050_, new_n5051_, new_n5052_, new_n5053_, new_n5054_, new_n5055_,
    new_n5056_, new_n5057_, new_n5058_, new_n5059_, new_n5060_, new_n5061_,
    new_n5062_, new_n5063_, new_n5064_, new_n5065_, new_n5066_, new_n5067_,
    new_n5068_, new_n5069_, new_n5070_, new_n5071_, new_n5072_, new_n5073_,
    new_n5074_, new_n5075_, new_n5076_, new_n5077_, new_n5078_, new_n5079_,
    new_n5080_, new_n5081_, new_n5082_, new_n5083_, new_n5084_, new_n5085_,
    new_n5086_, new_n5087_, new_n5088_, new_n5089_, new_n5090_, new_n5091_,
    new_n5092_, new_n5093_, new_n5094_, new_n5095_, new_n5096_, new_n5097_,
    new_n5098_, new_n5099_, new_n5100_, new_n5101_, new_n5102_, new_n5103_,
    new_n5104_, new_n5105_, new_n5106_, new_n5107_, new_n5108_, new_n5109_,
    new_n5110_, new_n5111_, new_n5112_, new_n5113_, new_n5114_, new_n5115_,
    new_n5116_, new_n5117_, new_n5118_, new_n5119_, new_n5120_, new_n5121_,
    new_n5122_, new_n5123_, new_n5124_, new_n5125_, new_n5126_, new_n5127_,
    new_n5128_, new_n5129_, new_n5130_, new_n5131_, new_n5132_, new_n5133_,
    new_n5134_, new_n5135_, new_n5136_, new_n5137_, new_n5138_, new_n5139_,
    new_n5140_, new_n5141_, new_n5142_, new_n5143_, new_n5144_, new_n5145_,
    new_n5146_, new_n5147_, new_n5148_, new_n5149_, new_n5150_, new_n5151_,
    new_n5152_, new_n5153_, new_n5154_, new_n5155_, new_n5156_, new_n5157_,
    new_n5158_, new_n5159_, new_n5160_, new_n5161_, new_n5162_, new_n5163_,
    new_n5164_, new_n5165_, new_n5166_, new_n5167_, new_n5168_, new_n5169_,
    new_n5170_, new_n5171_, new_n5172_, new_n5173_, new_n5174_, new_n5175_,
    new_n5176_, new_n5177_, new_n5178_, new_n5179_, new_n5180_, new_n5181_,
    new_n5182_, new_n5183_, new_n5184_, new_n5185_, new_n5186_, new_n5187_,
    new_n5188_, new_n5189_, new_n5190_, new_n5191_, new_n5192_, new_n5193_,
    new_n5194_, new_n5195_, new_n5196_, new_n5197_, new_n5198_, new_n5199_,
    new_n5200_, new_n5201_, new_n5202_, new_n5203_, new_n5204_, new_n5205_,
    new_n5206_, new_n5207_, new_n5208_, new_n5210_, new_n5211_, new_n5212_,
    new_n5213_, new_n5214_, new_n5215_, new_n5216_, new_n5217_, new_n5218_,
    new_n5219_, new_n5220_, new_n5221_, new_n5222_, new_n5223_, new_n5224_,
    new_n5225_, new_n5226_, new_n5227_, new_n5228_, new_n5229_, new_n5230_,
    new_n5231_, new_n5232_, new_n5233_, new_n5234_, new_n5235_, new_n5236_,
    new_n5237_, new_n5238_, new_n5239_, new_n5240_, new_n5241_, new_n5242_,
    new_n5243_, new_n5244_, new_n5245_, new_n5246_, new_n5247_, new_n5248_,
    new_n5249_, new_n5250_, new_n5251_, new_n5252_, new_n5253_, new_n5254_,
    new_n5255_, new_n5256_, new_n5257_, new_n5258_, new_n5259_, new_n5260_,
    new_n5261_, new_n5262_, new_n5263_, new_n5264_, new_n5265_, new_n5266_,
    new_n5267_, new_n5268_, new_n5269_, new_n5270_, new_n5271_, new_n5272_,
    new_n5273_, new_n5274_, new_n5275_, new_n5276_, new_n5277_, new_n5278_,
    new_n5279_, new_n5280_, new_n5281_, new_n5282_, new_n5283_, new_n5284_,
    new_n5285_, new_n5286_, new_n5287_, new_n5288_, new_n5289_, new_n5290_,
    new_n5291_, new_n5292_, new_n5293_, new_n5294_, new_n5295_, new_n5296_,
    new_n5297_, new_n5298_, new_n5299_, new_n5300_, new_n5301_, new_n5302_,
    new_n5303_, new_n5304_, new_n5305_, new_n5306_, new_n5307_, new_n5308_,
    new_n5309_, new_n5310_, new_n5311_, new_n5312_, new_n5313_, new_n5314_,
    new_n5315_, new_n5316_, new_n5317_, new_n5318_, new_n5319_, new_n5320_,
    new_n5321_, new_n5322_, new_n5323_, new_n5324_, new_n5325_, new_n5326_,
    new_n5327_, new_n5328_, new_n5329_, new_n5330_, new_n5331_, new_n5332_,
    new_n5333_, new_n5334_, new_n5335_, new_n5336_, new_n5337_, new_n5338_,
    new_n5339_, new_n5340_, new_n5341_, new_n5342_, new_n5343_, new_n5344_,
    new_n5345_, new_n5346_, new_n5347_, new_n5348_, new_n5349_, new_n5350_,
    new_n5351_, new_n5352_, new_n5353_, new_n5354_, new_n5355_, new_n5356_,
    new_n5357_, new_n5358_, new_n5359_, new_n5360_, new_n5361_, new_n5362_,
    new_n5363_, new_n5364_, new_n5365_, new_n5366_, new_n5367_, new_n5368_,
    new_n5369_, new_n5370_, new_n5371_, new_n5372_, new_n5373_, new_n5374_,
    new_n5375_, new_n5376_, new_n5377_, new_n5378_, new_n5379_, new_n5380_,
    new_n5381_, new_n5382_, new_n5383_, new_n5384_, new_n5385_, new_n5386_,
    new_n5387_, new_n5388_, new_n5389_, new_n5390_, new_n5391_, new_n5392_,
    new_n5393_, new_n5394_, new_n5395_, new_n5396_, new_n5397_, new_n5398_,
    new_n5399_, new_n5400_, new_n5401_, new_n5402_, new_n5403_, new_n5404_,
    new_n5405_, new_n5406_, new_n5407_, new_n5408_, new_n5409_, new_n5410_,
    new_n5411_, new_n5412_, new_n5413_, new_n5414_, new_n5415_, new_n5416_,
    new_n5417_, new_n5418_, new_n5419_, new_n5420_, new_n5421_, new_n5422_,
    new_n5423_, new_n5424_, new_n5425_, new_n5426_, new_n5427_, new_n5428_,
    new_n5429_, new_n5430_, new_n5431_, new_n5432_, new_n5433_, new_n5434_,
    new_n5435_, new_n5436_, new_n5437_, new_n5438_, new_n5439_, new_n5440_,
    new_n5441_, new_n5442_, new_n5443_, new_n5444_, new_n5445_, new_n5446_,
    new_n5447_, new_n5448_, new_n5449_, new_n5450_, new_n5451_, new_n5452_,
    new_n5453_, new_n5454_, new_n5455_, new_n5456_, new_n5457_, new_n5458_,
    new_n5459_, new_n5460_, new_n5461_, new_n5462_, new_n5463_, new_n5464_,
    new_n5465_, new_n5466_, new_n5467_, new_n5468_, new_n5469_, new_n5470_,
    new_n5471_, new_n5472_, new_n5473_, new_n5474_, new_n5475_, new_n5476_,
    new_n5477_, new_n5478_, new_n5479_, new_n5480_, new_n5481_, new_n5482_,
    new_n5483_, new_n5484_, new_n5485_, new_n5486_, new_n5487_, new_n5488_,
    new_n5489_, new_n5490_, new_n5491_, new_n5492_, new_n5493_, new_n5494_,
    new_n5495_, new_n5496_, new_n5497_, new_n5498_, new_n5499_, new_n5500_,
    new_n5501_, new_n5502_, new_n5503_, new_n5504_, new_n5505_, new_n5506_,
    new_n5507_, new_n5508_, new_n5509_, new_n5510_, new_n5511_, new_n5512_,
    new_n5513_, new_n5514_, new_n5515_, new_n5516_, new_n5517_, new_n5518_,
    new_n5519_, new_n5520_, new_n5521_, new_n5522_, new_n5523_, new_n5524_,
    new_n5525_, new_n5526_, new_n5527_, new_n5528_, new_n5529_, new_n5530_,
    new_n5531_, new_n5532_, new_n5533_, new_n5534_, new_n5535_, new_n5536_,
    new_n5537_, new_n5538_, new_n5539_, new_n5540_, new_n5541_, new_n5542_,
    new_n5543_, new_n5544_, new_n5545_, new_n5546_, new_n5547_, new_n5548_,
    new_n5549_, new_n5550_, new_n5551_, new_n5552_, new_n5553_, new_n5554_,
    new_n5555_, new_n5556_, new_n5557_, new_n5558_, new_n5559_, new_n5560_,
    new_n5561_, new_n5562_, new_n5563_, new_n5564_, new_n5565_, new_n5567_,
    new_n5568_, new_n5569_, new_n5570_, new_n5571_, new_n5572_, new_n5573_,
    new_n5574_, new_n5575_, new_n5576_, new_n5577_, new_n5578_, new_n5579_,
    new_n5580_, new_n5581_, new_n5582_, new_n5583_, new_n5584_, new_n5585_,
    new_n5586_, new_n5587_, new_n5588_, new_n5589_, new_n5590_, new_n5591_,
    new_n5592_, new_n5593_, new_n5594_, new_n5595_, new_n5596_, new_n5597_,
    new_n5598_, new_n5599_, new_n5600_, new_n5601_, new_n5602_, new_n5603_,
    new_n5604_, new_n5605_, new_n5606_, new_n5607_, new_n5608_, new_n5609_,
    new_n5610_, new_n5611_, new_n5612_, new_n5613_, new_n5614_, new_n5615_,
    new_n5616_, new_n5617_, new_n5618_, new_n5619_, new_n5620_, new_n5621_,
    new_n5622_, new_n5623_, new_n5624_, new_n5625_, new_n5626_, new_n5627_,
    new_n5628_, new_n5629_, new_n5630_, new_n5631_, new_n5632_, new_n5633_,
    new_n5634_, new_n5635_, new_n5636_, new_n5637_, new_n5638_, new_n5639_,
    new_n5640_, new_n5641_, new_n5642_, new_n5643_, new_n5644_, new_n5645_,
    new_n5646_, new_n5647_, new_n5648_, new_n5649_, new_n5650_, new_n5651_,
    new_n5652_, new_n5653_, new_n5654_, new_n5655_, new_n5656_, new_n5657_,
    new_n5658_, new_n5659_, new_n5660_, new_n5661_, new_n5662_, new_n5663_,
    new_n5664_, new_n5665_, new_n5666_, new_n5667_, new_n5668_, new_n5669_,
    new_n5670_, new_n5671_, new_n5672_, new_n5673_, new_n5674_, new_n5675_,
    new_n5676_, new_n5677_, new_n5678_, new_n5679_, new_n5680_, new_n5681_,
    new_n5682_, new_n5683_, new_n5684_, new_n5685_, new_n5686_, new_n5687_,
    new_n5688_, new_n5689_, new_n5690_, new_n5691_, new_n5692_, new_n5693_,
    new_n5694_, new_n5695_, new_n5696_, new_n5697_, new_n5698_, new_n5699_,
    new_n5700_, new_n5701_, new_n5702_, new_n5703_, new_n5704_, new_n5705_,
    new_n5706_, new_n5707_, new_n5708_, new_n5709_, new_n5710_, new_n5711_,
    new_n5712_, new_n5713_, new_n5714_, new_n5715_, new_n5716_, new_n5717_,
    new_n5718_, new_n5719_, new_n5720_, new_n5721_, new_n5722_, new_n5723_,
    new_n5724_, new_n5725_, new_n5726_, new_n5727_, new_n5728_, new_n5729_,
    new_n5730_, new_n5731_, new_n5732_, new_n5733_, new_n5734_, new_n5735_,
    new_n5736_, new_n5737_, new_n5738_, new_n5739_, new_n5740_, new_n5741_,
    new_n5742_, new_n5743_, new_n5744_, new_n5745_, new_n5746_, new_n5747_,
    new_n5748_, new_n5749_, new_n5750_, new_n5751_, new_n5752_, new_n5753_,
    new_n5754_, new_n5755_, new_n5756_, new_n5757_, new_n5758_, new_n5759_,
    new_n5760_, new_n5761_, new_n5762_, new_n5763_, new_n5764_, new_n5765_,
    new_n5766_, new_n5767_, new_n5768_, new_n5769_, new_n5770_, new_n5771_,
    new_n5772_, new_n5773_, new_n5774_, new_n5775_, new_n5776_, new_n5777_,
    new_n5778_, new_n5779_, new_n5780_, new_n5781_, new_n5782_, new_n5783_,
    new_n5784_, new_n5785_, new_n5786_, new_n5787_, new_n5788_, new_n5789_,
    new_n5790_, new_n5791_, new_n5792_, new_n5793_, new_n5794_, new_n5795_,
    new_n5796_, new_n5797_, new_n5798_, new_n5799_, new_n5800_, new_n5801_,
    new_n5802_, new_n5803_, new_n5804_, new_n5805_, new_n5806_, new_n5807_,
    new_n5808_, new_n5809_, new_n5810_, new_n5811_, new_n5812_, new_n5813_,
    new_n5814_, new_n5815_, new_n5816_, new_n5817_, new_n5818_, new_n5819_,
    new_n5820_, new_n5821_, new_n5822_, new_n5823_, new_n5824_, new_n5825_,
    new_n5826_, new_n5827_, new_n5828_, new_n5829_, new_n5830_, new_n5831_,
    new_n5832_, new_n5833_, new_n5834_, new_n5835_, new_n5836_, new_n5837_,
    new_n5838_, new_n5839_, new_n5840_, new_n5841_, new_n5842_, new_n5843_,
    new_n5844_, new_n5845_, new_n5846_, new_n5847_, new_n5848_, new_n5849_,
    new_n5850_, new_n5851_, new_n5852_, new_n5853_, new_n5854_, new_n5855_,
    new_n5856_, new_n5857_, new_n5858_, new_n5859_, new_n5860_, new_n5861_,
    new_n5862_, new_n5863_, new_n5864_, new_n5865_, new_n5866_, new_n5867_,
    new_n5868_, new_n5869_, new_n5870_, new_n5871_, new_n5872_, new_n5873_,
    new_n5874_, new_n5875_, new_n5876_, new_n5877_, new_n5878_, new_n5879_,
    new_n5880_, new_n5881_, new_n5882_, new_n5883_, new_n5884_, new_n5885_,
    new_n5886_, new_n5887_, new_n5888_, new_n5889_, new_n5890_, new_n5891_,
    new_n5892_, new_n5893_, new_n5894_, new_n5895_, new_n5896_, new_n5897_,
    new_n5898_, new_n5899_, new_n5900_, new_n5901_, new_n5902_, new_n5903_,
    new_n5904_, new_n5905_, new_n5906_, new_n5907_, new_n5908_, new_n5910_,
    new_n5911_, new_n5912_, new_n5913_, new_n5914_, new_n5915_, new_n5916_,
    new_n5917_, new_n5918_, new_n5919_, new_n5920_, new_n5921_, new_n5922_,
    new_n5923_, new_n5924_, new_n5925_, new_n5926_, new_n5927_, new_n5928_,
    new_n5929_, new_n5930_, new_n5931_, new_n5932_, new_n5933_, new_n5934_,
    new_n5935_, new_n5936_, new_n5937_, new_n5938_, new_n5939_, new_n5940_,
    new_n5941_, new_n5942_, new_n5943_, new_n5944_, new_n5945_, new_n5946_,
    new_n5947_, new_n5948_, new_n5949_, new_n5950_, new_n5951_, new_n5952_,
    new_n5953_, new_n5954_, new_n5955_, new_n5956_, new_n5957_, new_n5958_,
    new_n5959_, new_n5960_, new_n5961_, new_n5962_, new_n5963_, new_n5964_,
    new_n5965_, new_n5966_, new_n5967_, new_n5968_, new_n5969_, new_n5970_,
    new_n5971_, new_n5972_, new_n5973_, new_n5974_, new_n5975_, new_n5976_,
    new_n5977_, new_n5978_, new_n5979_, new_n5980_, new_n5981_, new_n5982_,
    new_n5983_, new_n5984_, new_n5985_, new_n5986_, new_n5987_, new_n5988_,
    new_n5989_, new_n5990_, new_n5991_, new_n5992_, new_n5993_, new_n5994_,
    new_n5995_, new_n5996_, new_n5997_, new_n5998_, new_n5999_, new_n6000_,
    new_n6001_, new_n6002_, new_n6003_, new_n6004_, new_n6005_, new_n6006_,
    new_n6007_, new_n6008_, new_n6009_, new_n6010_, new_n6011_, new_n6012_,
    new_n6013_, new_n6014_, new_n6015_, new_n6016_, new_n6017_, new_n6018_,
    new_n6019_, new_n6020_, new_n6021_, new_n6022_, new_n6023_, new_n6024_,
    new_n6025_, new_n6026_, new_n6027_, new_n6028_, new_n6029_, new_n6030_,
    new_n6031_, new_n6032_, new_n6033_, new_n6034_, new_n6035_, new_n6036_,
    new_n6037_, new_n6038_, new_n6039_, new_n6040_, new_n6041_, new_n6042_,
    new_n6043_, new_n6044_, new_n6045_, new_n6046_, new_n6047_, new_n6048_,
    new_n6049_, new_n6050_, new_n6051_, new_n6052_, new_n6053_, new_n6054_,
    new_n6055_, new_n6056_, new_n6057_, new_n6058_, new_n6059_, new_n6060_,
    new_n6061_, new_n6062_, new_n6063_, new_n6064_, new_n6065_, new_n6066_,
    new_n6067_, new_n6068_, new_n6069_, new_n6070_, new_n6071_, new_n6072_,
    new_n6073_, new_n6074_, new_n6075_, new_n6076_, new_n6077_, new_n6078_,
    new_n6079_, new_n6080_, new_n6081_, new_n6082_, new_n6083_, new_n6084_,
    new_n6085_, new_n6086_, new_n6087_, new_n6088_, new_n6089_, new_n6090_,
    new_n6091_, new_n6092_, new_n6093_, new_n6094_, new_n6095_, new_n6096_,
    new_n6097_, new_n6098_, new_n6099_, new_n6100_, new_n6101_, new_n6102_,
    new_n6103_, new_n6104_, new_n6105_, new_n6106_, new_n6107_, new_n6108_,
    new_n6109_, new_n6110_, new_n6111_, new_n6112_, new_n6113_, new_n6114_,
    new_n6115_, new_n6116_, new_n6117_, new_n6118_, new_n6119_, new_n6120_,
    new_n6121_, new_n6122_, new_n6123_, new_n6124_, new_n6125_, new_n6126_,
    new_n6127_, new_n6128_, new_n6129_, new_n6130_, new_n6131_, new_n6132_,
    new_n6133_, new_n6134_, new_n6135_, new_n6136_, new_n6137_, new_n6138_,
    new_n6139_, new_n6140_, new_n6141_, new_n6142_, new_n6143_, new_n6144_,
    new_n6145_, new_n6146_, new_n6147_, new_n6148_, new_n6149_, new_n6150_,
    new_n6151_, new_n6152_, new_n6153_, new_n6154_, new_n6155_, new_n6156_,
    new_n6157_, new_n6158_, new_n6159_, new_n6160_, new_n6161_, new_n6162_,
    new_n6163_, new_n6164_, new_n6165_, new_n6166_, new_n6167_, new_n6168_,
    new_n6169_, new_n6170_, new_n6171_, new_n6172_, new_n6173_, new_n6174_,
    new_n6175_, new_n6176_, new_n6177_, new_n6178_, new_n6179_, new_n6180_,
    new_n6181_, new_n6182_, new_n6183_, new_n6184_, new_n6185_, new_n6186_,
    new_n6187_, new_n6188_, new_n6189_, new_n6190_, new_n6191_, new_n6192_,
    new_n6193_, new_n6194_, new_n6195_, new_n6196_, new_n6197_, new_n6198_,
    new_n6199_, new_n6200_, new_n6201_, new_n6202_, new_n6203_, new_n6204_,
    new_n6205_, new_n6206_, new_n6207_, new_n6208_, new_n6209_, new_n6210_,
    new_n6211_, new_n6212_, new_n6213_, new_n6214_, new_n6215_, new_n6216_,
    new_n6217_, new_n6218_, new_n6219_, new_n6220_, new_n6221_, new_n6222_,
    new_n6223_, new_n6224_, new_n6225_, new_n6226_, new_n6227_, new_n6228_,
    new_n6229_, new_n6230_, new_n6231_, new_n6232_, new_n6233_, new_n6234_,
    new_n6235_, new_n6236_, new_n6237_, new_n6238_, new_n6239_, new_n6240_,
    new_n6241_, new_n6242_, new_n6243_, new_n6244_, new_n6245_, new_n6246_,
    new_n6247_, new_n6248_, new_n6249_, new_n6250_, new_n6251_, new_n6252_,
    new_n6253_, new_n6254_, new_n6255_, new_n6256_, new_n6257_, new_n6258_,
    new_n6259_, new_n6260_, new_n6261_, new_n6262_, new_n6263_, new_n6264_,
    new_n6265_, new_n6266_, new_n6267_, new_n6268_, new_n6269_, new_n6270_,
    new_n6271_, new_n6272_, new_n6273_, new_n6274_, new_n6275_, new_n6276_,
    new_n6277_, new_n6278_, new_n6279_, new_n6280_, new_n6281_, new_n6282_,
    new_n6283_, new_n6284_, new_n6285_, new_n6286_, new_n6287_, new_n6288_,
    new_n6289_, new_n6290_, new_n6291_, new_n6292_, new_n6293_, new_n6294_,
    new_n6295_, new_n6296_, new_n6297_, new_n6298_, new_n6299_, new_n6300_,
    new_n6301_, new_n6302_, new_n6303_, new_n6304_, new_n6305_, new_n6306_,
    new_n6307_, new_n6308_, new_n6309_, new_n6310_, new_n6311_, new_n6312_,
    new_n6313_, new_n6314_, new_n6315_, new_n6316_, new_n6317_, new_n6318_,
    new_n6319_, new_n6320_, new_n6321_, new_n6322_, new_n6323_, new_n6324_,
    new_n6325_, new_n6326_, new_n6327_, new_n6328_, new_n6329_, new_n6330_,
    new_n6331_, new_n6332_, new_n6333_, new_n6334_, new_n6335_, new_n6336_,
    new_n6337_, new_n6338_, new_n6339_, new_n6340_, new_n6341_, new_n6342_,
    new_n6343_, new_n6344_, new_n6345_, new_n6346_, new_n6347_, new_n6348_,
    new_n6349_, new_n6350_, new_n6351_, new_n6352_, new_n6353_, new_n6354_,
    new_n6355_, new_n6356_, new_n6357_, new_n6358_, new_n6359_, new_n6360_,
    new_n6361_, new_n6362_, new_n6363_, new_n6364_, new_n6366_, new_n6367_,
    new_n6368_, new_n6369_, new_n6370_, new_n6371_, new_n6372_, new_n6373_,
    new_n6374_, new_n6375_, new_n6376_, new_n6377_, new_n6378_, new_n6379_,
    new_n6380_, new_n6381_, new_n6382_, new_n6383_, new_n6384_, new_n6385_,
    new_n6386_, new_n6387_, new_n6388_, new_n6389_, new_n6390_, new_n6391_,
    new_n6392_, new_n6393_, new_n6394_, new_n6395_, new_n6396_, new_n6397_,
    new_n6398_, new_n6399_, new_n6400_, new_n6401_, new_n6402_, new_n6403_,
    new_n6404_, new_n6405_, new_n6406_, new_n6407_, new_n6408_, new_n6409_,
    new_n6410_, new_n6411_, new_n6412_, new_n6413_, new_n6414_, new_n6415_,
    new_n6416_, new_n6417_, new_n6418_, new_n6419_, new_n6420_, new_n6421_,
    new_n6422_, new_n6423_, new_n6424_, new_n6425_, new_n6426_, new_n6427_,
    new_n6428_, new_n6429_, new_n6430_, new_n6431_, new_n6432_, new_n6433_,
    new_n6434_, new_n6435_, new_n6436_, new_n6437_, new_n6438_, new_n6439_,
    new_n6440_, new_n6441_, new_n6442_, new_n6443_, new_n6444_, new_n6445_,
    new_n6446_, new_n6447_, new_n6448_, new_n6449_, new_n6450_, new_n6451_,
    new_n6452_, new_n6453_, new_n6454_, new_n6455_, new_n6456_, new_n6457_,
    new_n6458_, new_n6459_, new_n6460_, new_n6461_, new_n6462_, new_n6463_,
    new_n6464_, new_n6465_, new_n6466_, new_n6467_, new_n6468_, new_n6469_,
    new_n6470_, new_n6471_, new_n6472_, new_n6473_, new_n6474_, new_n6475_,
    new_n6476_, new_n6477_, new_n6478_, new_n6479_, new_n6480_, new_n6481_,
    new_n6482_, new_n6483_, new_n6484_, new_n6485_, new_n6486_, new_n6487_,
    new_n6488_, new_n6489_, new_n6490_, new_n6491_, new_n6492_, new_n6493_,
    new_n6494_, new_n6495_, new_n6496_, new_n6497_, new_n6498_, new_n6499_,
    new_n6500_, new_n6501_, new_n6502_, new_n6503_, new_n6504_, new_n6505_,
    new_n6506_, new_n6507_, new_n6508_, new_n6509_, new_n6510_, new_n6511_,
    new_n6512_, new_n6513_, new_n6514_, new_n6515_, new_n6516_, new_n6517_,
    new_n6518_, new_n6519_, new_n6520_, new_n6521_, new_n6522_, new_n6523_,
    new_n6524_, new_n6525_, new_n6526_, new_n6527_, new_n6528_, new_n6529_,
    new_n6530_, new_n6531_, new_n6532_, new_n6533_, new_n6534_, new_n6535_,
    new_n6536_, new_n6537_, new_n6538_, new_n6539_, new_n6540_, new_n6541_,
    new_n6542_, new_n6543_, new_n6544_, new_n6545_, new_n6546_, new_n6547_,
    new_n6548_, new_n6549_, new_n6550_, new_n6551_, new_n6552_, new_n6553_,
    new_n6554_, new_n6555_, new_n6556_, new_n6557_, new_n6558_, new_n6559_,
    new_n6560_, new_n6561_, new_n6562_, new_n6563_, new_n6564_, new_n6565_,
    new_n6566_, new_n6567_, new_n6568_, new_n6569_, new_n6570_, new_n6571_,
    new_n6572_, new_n6573_, new_n6574_, new_n6575_, new_n6576_, new_n6577_,
    new_n6578_, new_n6579_, new_n6580_, new_n6581_, new_n6582_, new_n6583_,
    new_n6584_, new_n6585_, new_n6586_, new_n6587_, new_n6588_, new_n6589_,
    new_n6590_, new_n6591_, new_n6592_, new_n6593_, new_n6594_, new_n6595_,
    new_n6596_, new_n6597_, new_n6598_, new_n6599_, new_n6600_, new_n6601_,
    new_n6602_, new_n6603_, new_n6604_, new_n6605_, new_n6606_, new_n6607_,
    new_n6608_, new_n6609_, new_n6610_, new_n6611_, new_n6612_, new_n6613_,
    new_n6614_, new_n6615_, new_n6616_, new_n6617_, new_n6618_, new_n6619_,
    new_n6620_, new_n6621_, new_n6622_, new_n6623_, new_n6624_, new_n6625_,
    new_n6626_, new_n6627_, new_n6628_, new_n6629_, new_n6630_, new_n6631_,
    new_n6632_, new_n6633_, new_n6634_, new_n6635_, new_n6636_, new_n6637_,
    new_n6638_, new_n6639_, new_n6640_, new_n6641_, new_n6642_, new_n6643_,
    new_n6644_, new_n6645_, new_n6646_, new_n6647_, new_n6648_, new_n6649_,
    new_n6650_, new_n6651_, new_n6652_, new_n6653_, new_n6654_, new_n6655_,
    new_n6656_, new_n6657_, new_n6658_, new_n6659_, new_n6660_, new_n6661_,
    new_n6662_, new_n6663_, new_n6664_, new_n6665_, new_n6666_, new_n6667_,
    new_n6668_, new_n6669_, new_n6670_, new_n6671_, new_n6672_, new_n6673_,
    new_n6674_, new_n6675_, new_n6676_, new_n6677_, new_n6678_, new_n6679_,
    new_n6680_, new_n6681_, new_n6682_, new_n6683_, new_n6684_, new_n6685_,
    new_n6686_, new_n6687_, new_n6688_, new_n6689_, new_n6690_, new_n6691_,
    new_n6692_, new_n6693_, new_n6694_, new_n6695_, new_n6696_, new_n6697_,
    new_n6698_, new_n6699_, new_n6700_, new_n6701_, new_n6702_, new_n6703_,
    new_n6704_, new_n6705_, new_n6706_, new_n6707_, new_n6708_, new_n6709_,
    new_n6711_, new_n6712_, new_n6713_, new_n6714_, new_n6715_, new_n6716_,
    new_n6717_, new_n6718_, new_n6719_, new_n6720_, new_n6721_, new_n6722_,
    new_n6723_, new_n6724_, new_n6725_, new_n6726_, new_n6727_, new_n6728_,
    new_n6729_, new_n6730_, new_n6731_, new_n6732_, new_n6733_, new_n6734_,
    new_n6735_, new_n6736_, new_n6737_, new_n6738_, new_n6739_, new_n6740_,
    new_n6741_, new_n6742_, new_n6743_, new_n6744_, new_n6745_, new_n6746_,
    new_n6747_, new_n6748_, new_n6749_, new_n6750_, new_n6751_, new_n6752_,
    new_n6753_, new_n6754_, new_n6755_, new_n6756_, new_n6757_, new_n6758_,
    new_n6759_, new_n6760_, new_n6761_, new_n6762_, new_n6763_, new_n6764_,
    new_n6765_, new_n6766_, new_n6767_, new_n6768_, new_n6769_, new_n6770_,
    new_n6771_, new_n6772_, new_n6773_, new_n6774_, new_n6775_, new_n6776_,
    new_n6777_, new_n6778_, new_n6779_, new_n6780_, new_n6781_, new_n6782_,
    new_n6783_, new_n6784_, new_n6785_, new_n6786_, new_n6787_, new_n6788_,
    new_n6789_, new_n6790_, new_n6791_, new_n6792_, new_n6793_, new_n6794_,
    new_n6795_, new_n6796_, new_n6797_, new_n6798_, new_n6799_, new_n6800_,
    new_n6801_, new_n6802_, new_n6803_, new_n6804_, new_n6805_, new_n6806_,
    new_n6807_, new_n6808_, new_n6809_, new_n6810_, new_n6811_, new_n6812_,
    new_n6813_, new_n6814_, new_n6815_, new_n6816_, new_n6817_, new_n6818_,
    new_n6819_, new_n6820_, new_n6821_, new_n6822_, new_n6823_, new_n6824_,
    new_n6825_, new_n6826_, new_n6827_, new_n6828_, new_n6829_, new_n6830_,
    new_n6831_, new_n6832_, new_n6833_, new_n6834_, new_n6835_, new_n6836_,
    new_n6837_, new_n6838_, new_n6839_, new_n6840_, new_n6841_, new_n6842_,
    new_n6843_, new_n6844_, new_n6845_, new_n6846_, new_n6847_, new_n6848_,
    new_n6849_, new_n6850_, new_n6851_, new_n6852_, new_n6853_, new_n6854_,
    new_n6855_, new_n6856_, new_n6857_, new_n6858_, new_n6859_, new_n6860_,
    new_n6861_, new_n6862_, new_n6863_, new_n6864_, new_n6865_, new_n6866_,
    new_n6867_, new_n6868_, new_n6869_, new_n6870_, new_n6871_, new_n6872_,
    new_n6873_, new_n6874_, new_n6875_, new_n6876_, new_n6877_, new_n6878_,
    new_n6879_, new_n6880_, new_n6881_, new_n6882_, new_n6883_, new_n6884_,
    new_n6885_, new_n6886_, new_n6887_, new_n6888_, new_n6889_, new_n6890_,
    new_n6891_, new_n6892_, new_n6893_, new_n6894_, new_n6895_, new_n6896_,
    new_n6897_, new_n6898_, new_n6899_, new_n6900_, new_n6901_, new_n6902_,
    new_n6903_, new_n6904_, new_n6905_, new_n6906_, new_n6907_, new_n6908_,
    new_n6909_, new_n6910_, new_n6911_, new_n6912_, new_n6913_, new_n6914_,
    new_n6915_, new_n6916_, new_n6917_, new_n6918_, new_n6919_, new_n6920_,
    new_n6921_, new_n6922_, new_n6923_, new_n6924_, new_n6925_, new_n6926_,
    new_n6927_, new_n6928_, new_n6929_, new_n6930_, new_n6931_, new_n6932_,
    new_n6933_, new_n6934_, new_n6935_, new_n6936_, new_n6937_, new_n6938_,
    new_n6939_, new_n6940_, new_n6941_, new_n6942_, new_n6943_, new_n6944_,
    new_n6945_, new_n6946_, new_n6947_, new_n6948_, new_n6949_, new_n6950_,
    new_n6951_, new_n6952_, new_n6953_, new_n6954_, new_n6955_, new_n6956_,
    new_n6957_, new_n6958_, new_n6959_, new_n6960_, new_n6961_, new_n6962_,
    new_n6963_, new_n6964_, new_n6965_, new_n6966_, new_n6967_, new_n6968_,
    new_n6969_, new_n6970_, new_n6971_, new_n6972_, new_n6973_, new_n6974_,
    new_n6975_, new_n6976_, new_n6977_, new_n6978_, new_n6979_, new_n6980_,
    new_n6981_, new_n6982_, new_n6983_, new_n6984_, new_n6985_, new_n6986_,
    new_n6987_, new_n6988_, new_n6989_, new_n6990_, new_n6991_, new_n6992_,
    new_n6993_, new_n6994_, new_n6995_, new_n6996_, new_n6997_, new_n6998_,
    new_n6999_, new_n7000_, new_n7001_, new_n7002_, new_n7003_, new_n7004_,
    new_n7005_, new_n7006_, new_n7007_, new_n7008_, new_n7009_, new_n7010_,
    new_n7011_, new_n7012_, new_n7013_, new_n7014_, new_n7015_, new_n7016_,
    new_n7017_, new_n7018_, new_n7019_, new_n7020_, new_n7021_, new_n7022_,
    new_n7023_, new_n7024_, new_n7025_, new_n7026_, new_n7027_, new_n7028_,
    new_n7029_, new_n7030_, new_n7031_, new_n7032_, new_n7033_, new_n7034_,
    new_n7035_, new_n7036_, new_n7037_, new_n7038_, new_n7039_, new_n7040_,
    new_n7041_, new_n7042_, new_n7043_, new_n7044_, new_n7045_, new_n7046_,
    new_n7047_, new_n7048_, new_n7049_, new_n7050_, new_n7051_, new_n7052_,
    new_n7053_, new_n7054_, new_n7055_, new_n7056_, new_n7057_, new_n7058_,
    new_n7059_, new_n7060_, new_n7061_, new_n7062_, new_n7063_, new_n7064_,
    new_n7065_, new_n7066_, new_n7067_, new_n7068_, new_n7069_, new_n7070_,
    new_n7071_, new_n7072_, new_n7073_, new_n7074_, new_n7075_, new_n7076_,
    new_n7077_, new_n7078_, new_n7079_, new_n7080_, new_n7081_, new_n7082_,
    new_n7083_, new_n7084_, new_n7085_, new_n7086_, new_n7087_, new_n7088_,
    new_n7089_, new_n7090_, new_n7091_, new_n7092_, new_n7093_, new_n7094_,
    new_n7095_, new_n7096_, new_n7097_, new_n7098_, new_n7099_, new_n7100_,
    new_n7101_, new_n7102_, new_n7103_, new_n7105_, new_n7106_, new_n7107_,
    new_n7108_, new_n7109_, new_n7110_, new_n7111_, new_n7112_, new_n7113_,
    new_n7114_, new_n7115_, new_n7116_, new_n7117_, new_n7118_, new_n7119_,
    new_n7120_, new_n7121_, new_n7122_, new_n7123_, new_n7124_, new_n7125_,
    new_n7126_, new_n7127_, new_n7128_, new_n7129_, new_n7130_, new_n7131_,
    new_n7132_, new_n7133_, new_n7134_, new_n7135_, new_n7136_, new_n7137_,
    new_n7138_, new_n7139_, new_n7140_, new_n7141_, new_n7142_, new_n7143_,
    new_n7144_, new_n7145_, new_n7146_, new_n7147_, new_n7148_, new_n7149_,
    new_n7150_, new_n7151_, new_n7152_, new_n7153_, new_n7154_, new_n7155_,
    new_n7156_, new_n7157_, new_n7158_, new_n7159_, new_n7160_, new_n7161_,
    new_n7162_, new_n7163_, new_n7164_, new_n7165_, new_n7166_, new_n7167_,
    new_n7168_, new_n7169_, new_n7170_, new_n7171_, new_n7172_, new_n7173_,
    new_n7174_, new_n7175_, new_n7176_, new_n7177_, new_n7178_, new_n7179_,
    new_n7180_, new_n7181_, new_n7182_, new_n7183_, new_n7184_, new_n7185_,
    new_n7186_, new_n7187_, new_n7188_, new_n7189_, new_n7190_, new_n7191_,
    new_n7192_, new_n7193_, new_n7194_, new_n7195_, new_n7196_, new_n7197_,
    new_n7198_, new_n7199_, new_n7200_, new_n7201_, new_n7202_, new_n7203_,
    new_n7204_, new_n7205_, new_n7206_, new_n7207_, new_n7208_, new_n7209_,
    new_n7210_, new_n7211_, new_n7212_, new_n7213_, new_n7214_, new_n7215_,
    new_n7216_, new_n7217_, new_n7218_, new_n7219_, new_n7220_, new_n7221_,
    new_n7222_, new_n7223_, new_n7224_, new_n7225_, new_n7226_, new_n7227_,
    new_n7228_, new_n7229_, new_n7230_, new_n7231_, new_n7232_, new_n7233_,
    new_n7234_, new_n7235_, new_n7236_, new_n7237_, new_n7238_, new_n7239_,
    new_n7240_, new_n7241_, new_n7242_, new_n7243_, new_n7244_, new_n7245_,
    new_n7246_, new_n7247_, new_n7248_, new_n7249_, new_n7250_, new_n7251_,
    new_n7252_, new_n7253_, new_n7254_, new_n7255_, new_n7256_, new_n7257_,
    new_n7258_, new_n7259_, new_n7260_, new_n7261_, new_n7262_, new_n7263_,
    new_n7264_, new_n7265_, new_n7266_, new_n7267_, new_n7268_, new_n7269_,
    new_n7270_, new_n7271_, new_n7272_, new_n7273_, new_n7274_, new_n7275_,
    new_n7276_, new_n7277_, new_n7278_, new_n7279_, new_n7280_, new_n7281_,
    new_n7282_, new_n7283_, new_n7284_, new_n7285_, new_n7286_, new_n7287_,
    new_n7288_, new_n7289_, new_n7290_, new_n7291_, new_n7292_, new_n7293_,
    new_n7294_, new_n7295_, new_n7296_, new_n7297_, new_n7298_, new_n7299_,
    new_n7300_, new_n7301_, new_n7302_, new_n7303_, new_n7304_, new_n7305_,
    new_n7306_, new_n7307_, new_n7308_, new_n7309_, new_n7310_, new_n7311_,
    new_n7312_, new_n7313_, new_n7314_, new_n7315_, new_n7316_, new_n7317_,
    new_n7318_, new_n7319_, new_n7320_, new_n7321_, new_n7322_, new_n7323_,
    new_n7324_, new_n7325_, new_n7326_, new_n7327_, new_n7328_, new_n7329_,
    new_n7330_, new_n7331_, new_n7332_, new_n7333_, new_n7334_, new_n7335_,
    new_n7336_, new_n7337_, new_n7338_, new_n7339_, new_n7340_, new_n7341_,
    new_n7342_, new_n7343_, new_n7344_, new_n7345_, new_n7346_, new_n7347_,
    new_n7348_, new_n7349_, new_n7350_, new_n7351_, new_n7352_, new_n7353_,
    new_n7354_, new_n7355_, new_n7356_, new_n7357_, new_n7358_, new_n7359_,
    new_n7360_, new_n7361_, new_n7362_, new_n7363_, new_n7364_, new_n7365_,
    new_n7366_, new_n7367_, new_n7368_, new_n7369_, new_n7370_, new_n7371_,
    new_n7372_, new_n7373_, new_n7374_, new_n7375_, new_n7376_, new_n7377_,
    new_n7378_, new_n7379_, new_n7380_, new_n7381_, new_n7382_, new_n7383_,
    new_n7384_, new_n7385_, new_n7386_, new_n7387_, new_n7388_, new_n7389_,
    new_n7390_, new_n7391_, new_n7392_, new_n7393_, new_n7394_, new_n7395_,
    new_n7396_, new_n7397_, new_n7398_, new_n7399_, new_n7400_, new_n7401_,
    new_n7402_, new_n7403_, new_n7404_, new_n7405_, new_n7406_, new_n7407_,
    new_n7408_, new_n7409_, new_n7410_, new_n7411_, new_n7412_, new_n7413_,
    new_n7414_, new_n7415_, new_n7416_, new_n7417_, new_n7418_, new_n7419_,
    new_n7420_, new_n7421_, new_n7422_, new_n7423_, new_n7424_, new_n7425_,
    new_n7426_, new_n7427_, new_n7428_, new_n7429_, new_n7430_, new_n7431_,
    new_n7432_, new_n7433_, new_n7434_, new_n7435_, new_n7436_, new_n7437_,
    new_n7438_, new_n7439_, new_n7440_, new_n7441_, new_n7442_, new_n7443_,
    new_n7444_, new_n7445_, new_n7446_, new_n7447_, new_n7448_, new_n7449_,
    new_n7450_, new_n7451_, new_n7452_, new_n7453_, new_n7454_, new_n7455_,
    new_n7456_, new_n7457_, new_n7458_, new_n7459_, new_n7460_, new_n7461_,
    new_n7462_, new_n7463_, new_n7464_, new_n7465_, new_n7466_, new_n7467_,
    new_n7468_, new_n7469_, new_n7470_, new_n7471_, new_n7472_, new_n7473_,
    new_n7474_, new_n7475_, new_n7476_, new_n7477_, new_n7478_, new_n7479_,
    new_n7480_, new_n7481_, new_n7482_, new_n7483_, new_n7484_, new_n7485_,
    new_n7486_, new_n7487_, new_n7488_, new_n7489_, new_n7490_, new_n7491_,
    new_n7492_, new_n7493_, new_n7494_, new_n7495_, new_n7496_, new_n7497_,
    new_n7498_, new_n7499_, new_n7500_, new_n7501_, new_n7502_, new_n7503_,
    new_n7504_, new_n7505_, new_n7506_, new_n7507_, new_n7508_, new_n7509_,
    new_n7510_, new_n7511_, new_n7512_, new_n7513_, new_n7514_, new_n7515_,
    new_n7516_, new_n7517_, new_n7518_, new_n7519_, new_n7520_, new_n7521_,
    new_n7522_, new_n7523_, new_n7524_, new_n7525_, new_n7526_, new_n7527_,
    new_n7528_, new_n7529_, new_n7530_, new_n7531_, new_n7532_, new_n7533_,
    new_n7534_, new_n7535_, new_n7536_, new_n7537_, new_n7538_, new_n7539_,
    new_n7540_, new_n7541_, new_n7542_, new_n7543_, new_n7544_, new_n7545_,
    new_n7546_, new_n7547_, new_n7548_, new_n7549_, new_n7550_, new_n7551_,
    new_n7552_, new_n7553_, new_n7554_, new_n7555_, new_n7556_, new_n7557_,
    new_n7558_, new_n7559_, new_n7560_, new_n7561_, new_n7562_, new_n7563_,
    new_n7564_, new_n7565_, new_n7566_, new_n7567_, new_n7568_, new_n7569_,
    new_n7570_, new_n7571_, new_n7572_, new_n7573_, new_n7574_, new_n7575_,
    new_n7576_, new_n7577_, new_n7578_, new_n7579_, new_n7580_, new_n7581_,
    new_n7582_, new_n7583_, new_n7584_, new_n7585_, new_n7586_, new_n7587_,
    new_n7588_, new_n7589_, new_n7590_, new_n7591_, new_n7592_, new_n7593_,
    new_n7594_, new_n7595_, new_n7596_, new_n7597_, new_n7598_, new_n7599_,
    new_n7600_, new_n7601_, new_n7602_, new_n7603_, new_n7604_, new_n7605_,
    new_n7606_, new_n7607_, new_n7608_, new_n7609_, new_n7610_, new_n7611_,
    new_n7613_, new_n7614_, new_n7615_, new_n7616_, new_n7617_, new_n7618_,
    new_n7619_, new_n7620_, new_n7621_, new_n7622_, new_n7623_, new_n7624_,
    new_n7625_, new_n7626_, new_n7627_, new_n7628_, new_n7629_, new_n7630_,
    new_n7631_, new_n7632_, new_n7633_, new_n7634_, new_n7635_, new_n7636_,
    new_n7637_, new_n7638_, new_n7639_, new_n7640_, new_n7641_, new_n7642_,
    new_n7643_, new_n7644_, new_n7645_, new_n7646_, new_n7647_, new_n7648_,
    new_n7649_, new_n7650_, new_n7651_, new_n7652_, new_n7653_, new_n7654_,
    new_n7655_, new_n7656_, new_n7657_, new_n7658_, new_n7659_, new_n7660_,
    new_n7661_, new_n7662_, new_n7663_, new_n7664_, new_n7665_, new_n7666_,
    new_n7667_, new_n7668_, new_n7669_, new_n7670_, new_n7671_, new_n7672_,
    new_n7673_, new_n7674_, new_n7675_, new_n7676_, new_n7677_, new_n7678_,
    new_n7679_, new_n7680_, new_n7681_, new_n7682_, new_n7683_, new_n7684_,
    new_n7685_, new_n7686_, new_n7687_, new_n7688_, new_n7689_, new_n7690_,
    new_n7691_, new_n7692_, new_n7693_, new_n7694_, new_n7695_, new_n7696_,
    new_n7697_, new_n7698_, new_n7699_, new_n7700_, new_n7701_, new_n7702_,
    new_n7703_, new_n7704_, new_n7705_, new_n7706_, new_n7707_, new_n7708_,
    new_n7709_, new_n7710_, new_n7711_, new_n7712_, new_n7713_, new_n7714_,
    new_n7715_, new_n7716_, new_n7717_, new_n7718_, new_n7719_, new_n7720_,
    new_n7721_, new_n7722_, new_n7723_, new_n7724_, new_n7725_, new_n7726_,
    new_n7727_, new_n7728_, new_n7729_, new_n7730_, new_n7731_, new_n7732_,
    new_n7733_, new_n7734_, new_n7735_, new_n7736_, new_n7737_, new_n7738_,
    new_n7739_, new_n7740_, new_n7741_, new_n7742_, new_n7743_, new_n7744_,
    new_n7745_, new_n7746_, new_n7747_, new_n7748_, new_n7749_, new_n7750_,
    new_n7751_, new_n7752_, new_n7753_, new_n7754_, new_n7755_, new_n7756_,
    new_n7757_, new_n7758_, new_n7759_, new_n7760_, new_n7761_, new_n7762_,
    new_n7763_, new_n7764_, new_n7765_, new_n7766_, new_n7767_, new_n7768_,
    new_n7769_, new_n7770_, new_n7771_, new_n7772_, new_n7773_, new_n7774_,
    new_n7775_, new_n7776_, new_n7777_, new_n7778_, new_n7779_, new_n7780_,
    new_n7781_, new_n7782_, new_n7783_, new_n7784_, new_n7785_, new_n7786_,
    new_n7787_, new_n7788_, new_n7789_, new_n7790_, new_n7791_, new_n7792_,
    new_n7793_, new_n7794_, new_n7795_, new_n7796_, new_n7797_, new_n7798_,
    new_n7799_, new_n7800_, new_n7801_, new_n7802_, new_n7803_, new_n7804_,
    new_n7805_, new_n7806_, new_n7807_, new_n7808_, new_n7809_, new_n7810_,
    new_n7811_, new_n7812_, new_n7813_, new_n7814_, new_n7815_, new_n7816_,
    new_n7817_, new_n7818_, new_n7819_, new_n7820_, new_n7821_, new_n7822_,
    new_n7823_, new_n7824_, new_n7825_, new_n7826_, new_n7827_, new_n7828_,
    new_n7829_, new_n7830_, new_n7831_, new_n7832_, new_n7833_, new_n7834_,
    new_n7835_, new_n7836_, new_n7837_, new_n7838_, new_n7839_, new_n7840_,
    new_n7841_, new_n7842_, new_n7843_, new_n7844_, new_n7845_, new_n7846_,
    new_n7847_, new_n7848_, new_n7849_, new_n7850_, new_n7851_, new_n7852_,
    new_n7853_, new_n7854_, new_n7855_, new_n7856_, new_n7857_, new_n7858_,
    new_n7859_, new_n7860_, new_n7861_, new_n7862_, new_n7863_, new_n7864_,
    new_n7865_, new_n7866_, new_n7867_, new_n7868_, new_n7869_, new_n7870_,
    new_n7871_, new_n7872_, new_n7873_, new_n7874_, new_n7875_, new_n7876_,
    new_n7877_, new_n7878_, new_n7879_, new_n7880_, new_n7881_, new_n7882_,
    new_n7883_, new_n7884_, new_n7885_, new_n7886_, new_n7887_, new_n7888_,
    new_n7889_, new_n7890_, new_n7891_, new_n7892_, new_n7893_, new_n7894_,
    new_n7895_, new_n7896_, new_n7897_, new_n7898_, new_n7899_, new_n7900_,
    new_n7901_, new_n7902_, new_n7903_, new_n7904_, new_n7905_, new_n7906_,
    new_n7907_, new_n7908_, new_n7909_, new_n7910_, new_n7911_, new_n7912_,
    new_n7913_, new_n7914_, new_n7915_, new_n7916_, new_n7917_, new_n7918_,
    new_n7919_, new_n7920_, new_n7921_, new_n7922_, new_n7923_, new_n7924_,
    new_n7925_, new_n7926_, new_n7927_, new_n7928_, new_n7929_, new_n7930_,
    new_n7931_, new_n7932_, new_n7933_, new_n7934_, new_n7935_, new_n7936_,
    new_n7937_, new_n7938_, new_n7939_, new_n7940_, new_n7941_, new_n7942_,
    new_n7943_, new_n7944_, new_n7945_, new_n7946_, new_n7947_, new_n7948_,
    new_n7949_, new_n7950_, new_n7951_, new_n7952_, new_n7953_, new_n7954_,
    new_n7955_, new_n7956_, new_n7957_, new_n7958_, new_n7959_, new_n7960_,
    new_n7961_, new_n7962_, new_n7963_, new_n7964_, new_n7965_, new_n7966_,
    new_n7967_, new_n7968_, new_n7969_, new_n7970_, new_n7971_, new_n7972_,
    new_n7973_, new_n7974_, new_n7975_, new_n7976_, new_n7977_, new_n7978_,
    new_n7979_, new_n7980_, new_n7981_, new_n7982_, new_n7983_, new_n7984_,
    new_n7985_, new_n7986_, new_n7987_, new_n7988_, new_n7989_, new_n7990_,
    new_n7991_, new_n7992_, new_n7993_, new_n7994_, new_n7995_, new_n7996_,
    new_n7998_, new_n7999_, new_n8000_, new_n8001_, new_n8002_, new_n8003_,
    new_n8004_, new_n8005_, new_n8006_, new_n8007_, new_n8008_, new_n8009_,
    new_n8010_, new_n8011_, new_n8012_, new_n8013_, new_n8014_, new_n8015_,
    new_n8016_, new_n8017_, new_n8018_, new_n8019_, new_n8020_, new_n8021_,
    new_n8022_, new_n8023_, new_n8024_, new_n8025_, new_n8026_, new_n8027_,
    new_n8028_, new_n8029_, new_n8030_, new_n8031_, new_n8032_, new_n8033_,
    new_n8034_, new_n8035_, new_n8036_, new_n8037_, new_n8038_, new_n8039_,
    new_n8040_, new_n8041_, new_n8042_, new_n8043_, new_n8044_, new_n8045_,
    new_n8046_, new_n8047_, new_n8048_, new_n8049_, new_n8050_, new_n8051_,
    new_n8052_, new_n8053_, new_n8054_, new_n8055_, new_n8056_, new_n8057_,
    new_n8058_, new_n8059_, new_n8060_, new_n8061_, new_n8062_, new_n8063_,
    new_n8064_, new_n8065_, new_n8066_, new_n8067_, new_n8068_, new_n8069_,
    new_n8070_, new_n8071_, new_n8072_, new_n8073_, new_n8074_, new_n8075_,
    new_n8076_, new_n8077_, new_n8078_, new_n8079_, new_n8080_, new_n8081_,
    new_n8082_, new_n8083_, new_n8084_, new_n8085_, new_n8086_, new_n8087_,
    new_n8088_, new_n8089_, new_n8090_, new_n8091_, new_n8092_, new_n8093_,
    new_n8094_, new_n8095_, new_n8096_, new_n8097_, new_n8098_, new_n8099_,
    new_n8100_, new_n8101_, new_n8102_, new_n8103_, new_n8104_, new_n8105_,
    new_n8106_, new_n8107_, new_n8108_, new_n8109_, new_n8110_, new_n8111_,
    new_n8112_, new_n8113_, new_n8114_, new_n8115_, new_n8116_, new_n8117_,
    new_n8118_, new_n8119_, new_n8120_, new_n8121_, new_n8122_, new_n8123_,
    new_n8124_, new_n8125_, new_n8126_, new_n8127_, new_n8128_, new_n8129_,
    new_n8130_, new_n8131_, new_n8132_, new_n8133_, new_n8134_, new_n8135_,
    new_n8136_, new_n8137_, new_n8138_, new_n8139_, new_n8140_, new_n8141_,
    new_n8142_, new_n8143_, new_n8144_, new_n8145_, new_n8146_, new_n8147_,
    new_n8148_, new_n8149_, new_n8150_, new_n8151_, new_n8152_, new_n8153_,
    new_n8154_, new_n8155_, new_n8156_, new_n8157_, new_n8158_, new_n8159_,
    new_n8160_, new_n8161_, new_n8162_, new_n8163_, new_n8164_, new_n8165_,
    new_n8166_, new_n8167_, new_n8168_, new_n8169_, new_n8170_, new_n8171_,
    new_n8172_, new_n8173_, new_n8174_, new_n8175_, new_n8176_, new_n8177_,
    new_n8178_, new_n8179_, new_n8180_, new_n8181_, new_n8182_, new_n8183_,
    new_n8184_, new_n8185_, new_n8186_, new_n8187_, new_n8188_, new_n8189_,
    new_n8190_, new_n8191_, new_n8192_, new_n8193_, new_n8194_, new_n8195_,
    new_n8196_, new_n8197_, new_n8198_, new_n8199_, new_n8200_, new_n8201_,
    new_n8202_, new_n8203_, new_n8204_, new_n8205_, new_n8206_, new_n8207_,
    new_n8208_, new_n8209_, new_n8210_, new_n8211_, new_n8212_, new_n8213_,
    new_n8214_, new_n8215_, new_n8216_, new_n8217_, new_n8218_, new_n8219_,
    new_n8220_, new_n8221_, new_n8222_, new_n8223_, new_n8224_, new_n8225_,
    new_n8226_, new_n8227_, new_n8228_, new_n8229_, new_n8230_, new_n8231_,
    new_n8232_, new_n8233_, new_n8234_, new_n8235_, new_n8236_, new_n8237_,
    new_n8238_, new_n8239_, new_n8240_, new_n8241_, new_n8242_, new_n8243_,
    new_n8244_, new_n8245_, new_n8246_, new_n8247_, new_n8248_, new_n8249_,
    new_n8250_, new_n8251_, new_n8252_, new_n8253_, new_n8254_, new_n8255_,
    new_n8256_, new_n8257_, new_n8258_, new_n8259_, new_n8260_, new_n8261_,
    new_n8262_, new_n8263_, new_n8264_, new_n8265_, new_n8266_, new_n8267_,
    new_n8268_, new_n8269_, new_n8270_, new_n8271_, new_n8272_, new_n8273_,
    new_n8274_, new_n8275_, new_n8276_, new_n8277_, new_n8278_, new_n8279_,
    new_n8280_, new_n8281_, new_n8282_, new_n8283_, new_n8284_, new_n8285_,
    new_n8286_, new_n8287_, new_n8288_, new_n8289_, new_n8290_, new_n8291_,
    new_n8292_, new_n8293_, new_n8294_, new_n8295_, new_n8296_, new_n8297_,
    new_n8298_, new_n8299_, new_n8300_, new_n8301_, new_n8302_, new_n8303_,
    new_n8304_, new_n8305_, new_n8306_, new_n8307_, new_n8308_, new_n8309_,
    new_n8310_, new_n8311_, new_n8312_, new_n8313_, new_n8314_, new_n8315_,
    new_n8316_, new_n8317_, new_n8318_, new_n8319_, new_n8320_, new_n8321_,
    new_n8322_, new_n8323_, new_n8324_, new_n8325_, new_n8326_, new_n8327_,
    new_n8328_, new_n8329_, new_n8330_, new_n8331_, new_n8332_, new_n8333_,
    new_n8334_, new_n8335_, new_n8336_, new_n8337_, new_n8338_, new_n8339_,
    new_n8340_, new_n8341_, new_n8342_, new_n8343_, new_n8344_, new_n8345_,
    new_n8346_, new_n8347_, new_n8348_, new_n8349_, new_n8350_, new_n8351_,
    new_n8352_, new_n8353_, new_n8354_, new_n8355_, new_n8356_, new_n8357_,
    new_n8358_, new_n8359_, new_n8360_, new_n8361_, new_n8362_, new_n8363_,
    new_n8364_, new_n8365_, new_n8366_, new_n8367_, new_n8368_, new_n8369_,
    new_n8370_, new_n8371_, new_n8372_, new_n8373_, new_n8374_, new_n8375_,
    new_n8376_, new_n8377_, new_n8378_, new_n8379_, new_n8380_, new_n8381_,
    new_n8382_, new_n8383_, new_n8384_, new_n8385_, new_n8386_, new_n8387_,
    new_n8388_, new_n8389_, new_n8390_, new_n8391_, new_n8392_, new_n8393_,
    new_n8394_, new_n8395_, new_n8396_, new_n8397_, new_n8398_, new_n8399_,
    new_n8400_, new_n8401_, new_n8402_, new_n8403_, new_n8404_, new_n8405_,
    new_n8406_, new_n8407_, new_n8408_, new_n8409_, new_n8410_, new_n8411_,
    new_n8412_, new_n8414_, new_n8415_, new_n8416_, new_n8417_, new_n8418_,
    new_n8419_, new_n8420_, new_n8421_, new_n8422_, new_n8423_, new_n8424_,
    new_n8425_, new_n8426_, new_n8427_, new_n8428_, new_n8429_, new_n8430_,
    new_n8431_, new_n8432_, new_n8433_, new_n8434_, new_n8435_, new_n8436_,
    new_n8437_, new_n8438_, new_n8439_, new_n8440_, new_n8441_, new_n8442_,
    new_n8443_, new_n8444_, new_n8445_, new_n8446_, new_n8447_, new_n8448_,
    new_n8449_, new_n8450_, new_n8451_, new_n8452_, new_n8453_, new_n8454_,
    new_n8455_, new_n8456_, new_n8457_, new_n8458_, new_n8459_, new_n8460_,
    new_n8461_, new_n8462_, new_n8463_, new_n8464_, new_n8465_, new_n8466_,
    new_n8467_, new_n8468_, new_n8469_, new_n8470_, new_n8471_, new_n8472_,
    new_n8473_, new_n8474_, new_n8475_, new_n8476_, new_n8477_, new_n8478_,
    new_n8479_, new_n8480_, new_n8481_, new_n8482_, new_n8483_, new_n8484_,
    new_n8485_, new_n8486_, new_n8487_, new_n8488_, new_n8489_, new_n8490_,
    new_n8491_, new_n8492_, new_n8493_, new_n8494_, new_n8495_, new_n8496_,
    new_n8497_, new_n8498_, new_n8499_, new_n8500_, new_n8501_, new_n8502_,
    new_n8503_, new_n8504_, new_n8505_, new_n8506_, new_n8507_, new_n8508_,
    new_n8509_, new_n8510_, new_n8511_, new_n8512_, new_n8513_, new_n8514_,
    new_n8515_, new_n8516_, new_n8517_, new_n8518_, new_n8519_, new_n8520_,
    new_n8521_, new_n8522_, new_n8523_, new_n8524_, new_n8525_, new_n8526_,
    new_n8527_, new_n8528_, new_n8529_, new_n8530_, new_n8531_, new_n8532_,
    new_n8533_, new_n8534_, new_n8535_, new_n8536_, new_n8537_, new_n8538_,
    new_n8539_, new_n8540_, new_n8541_, new_n8542_, new_n8543_, new_n8544_,
    new_n8545_, new_n8546_, new_n8547_, new_n8548_, new_n8549_, new_n8550_,
    new_n8551_, new_n8552_, new_n8553_, new_n8554_, new_n8555_, new_n8556_,
    new_n8557_, new_n8558_, new_n8559_, new_n8560_, new_n8561_, new_n8562_,
    new_n8563_, new_n8564_, new_n8565_, new_n8566_, new_n8567_, new_n8568_,
    new_n8569_, new_n8570_, new_n8571_, new_n8572_, new_n8573_, new_n8574_,
    new_n8575_, new_n8576_, new_n8577_, new_n8578_, new_n8579_, new_n8580_,
    new_n8581_, new_n8582_, new_n8583_, new_n8584_, new_n8585_, new_n8586_,
    new_n8587_, new_n8588_, new_n8589_, new_n8590_, new_n8591_, new_n8592_,
    new_n8593_, new_n8594_, new_n8595_, new_n8596_, new_n8597_, new_n8598_,
    new_n8599_, new_n8600_, new_n8601_, new_n8602_, new_n8603_, new_n8604_,
    new_n8605_, new_n8606_, new_n8607_, new_n8608_, new_n8609_, new_n8610_,
    new_n8611_, new_n8612_, new_n8613_, new_n8614_, new_n8615_, new_n8616_,
    new_n8617_, new_n8618_, new_n8619_, new_n8620_, new_n8621_, new_n8622_,
    new_n8623_, new_n8624_, new_n8625_, new_n8626_, new_n8627_, new_n8628_,
    new_n8629_, new_n8630_, new_n8631_, new_n8632_, new_n8633_, new_n8634_,
    new_n8635_, new_n8636_, new_n8637_, new_n8638_, new_n8639_, new_n8640_,
    new_n8641_, new_n8642_, new_n8643_, new_n8644_, new_n8645_, new_n8646_,
    new_n8647_, new_n8648_, new_n8649_, new_n8650_, new_n8651_, new_n8652_,
    new_n8653_, new_n8654_, new_n8655_, new_n8656_, new_n8657_, new_n8658_,
    new_n8659_, new_n8660_, new_n8661_, new_n8662_, new_n8663_, new_n8664_,
    new_n8665_, new_n8666_, new_n8667_, new_n8668_, new_n8669_, new_n8670_,
    new_n8671_, new_n8672_, new_n8673_, new_n8674_, new_n8675_, new_n8676_,
    new_n8677_, new_n8678_, new_n8679_, new_n8680_, new_n8681_, new_n8682_,
    new_n8683_, new_n8684_, new_n8685_, new_n8686_, new_n8687_, new_n8688_,
    new_n8689_, new_n8690_, new_n8691_, new_n8692_, new_n8693_, new_n8694_,
    new_n8695_, new_n8696_, new_n8697_, new_n8698_, new_n8699_, new_n8700_,
    new_n8701_, new_n8702_, new_n8703_, new_n8704_, new_n8705_, new_n8706_,
    new_n8707_, new_n8708_, new_n8709_, new_n8710_, new_n8711_, new_n8712_,
    new_n8713_, new_n8714_, new_n8715_, new_n8716_, new_n8717_, new_n8718_,
    new_n8719_, new_n8720_, new_n8721_, new_n8722_, new_n8723_, new_n8724_,
    new_n8725_, new_n8726_, new_n8727_, new_n8728_, new_n8729_, new_n8730_,
    new_n8731_, new_n8732_, new_n8733_, new_n8734_, new_n8735_, new_n8736_,
    new_n8737_, new_n8738_, new_n8739_, new_n8740_, new_n8741_, new_n8742_,
    new_n8743_, new_n8744_, new_n8745_, new_n8746_, new_n8747_, new_n8748_,
    new_n8749_, new_n8750_, new_n8751_, new_n8752_, new_n8753_, new_n8754_,
    new_n8755_, new_n8756_, new_n8757_, new_n8758_, new_n8759_, new_n8760_,
    new_n8761_, new_n8762_, new_n8763_, new_n8764_, new_n8765_, new_n8766_,
    new_n8767_, new_n8768_, new_n8769_, new_n8770_, new_n8771_, new_n8772_,
    new_n8773_, new_n8774_, new_n8775_, new_n8776_, new_n8777_, new_n8778_,
    new_n8779_, new_n8780_, new_n8781_, new_n8782_, new_n8783_, new_n8784_,
    new_n8785_, new_n8786_, new_n8787_, new_n8788_, new_n8789_, new_n8790_,
    new_n8791_, new_n8792_, new_n8793_, new_n8794_, new_n8795_, new_n8796_,
    new_n8797_, new_n8798_, new_n8799_, new_n8800_, new_n8801_, new_n8802_,
    new_n8803_, new_n8804_, new_n8805_, new_n8806_, new_n8807_, new_n8808_,
    new_n8809_, new_n8810_, new_n8811_, new_n8812_, new_n8813_, new_n8814_,
    new_n8815_, new_n8816_, new_n8817_, new_n8818_, new_n8819_, new_n8820_,
    new_n8821_, new_n8822_, new_n8823_, new_n8824_, new_n8825_, new_n8826_,
    new_n8827_, new_n8828_, new_n8829_, new_n8830_, new_n8831_, new_n8832_,
    new_n8833_, new_n8834_, new_n8835_, new_n8836_, new_n8837_, new_n8838_,
    new_n8839_, new_n8840_, new_n8841_, new_n8842_, new_n8843_, new_n8844_,
    new_n8845_, new_n8846_, new_n8847_, new_n8848_, new_n8849_, new_n8850_,
    new_n8851_, new_n8852_, new_n8853_, new_n8854_, new_n8855_, new_n8856_,
    new_n8857_, new_n8858_, new_n8859_, new_n8860_, new_n8861_, new_n8862_,
    new_n8863_, new_n8864_, new_n8865_, new_n8866_, new_n8867_, new_n8868_,
    new_n8869_, new_n8870_, new_n8871_, new_n8872_, new_n8873_, new_n8874_,
    new_n8875_, new_n8876_, new_n8877_, new_n8878_, new_n8879_, new_n8880_,
    new_n8881_, new_n8882_, new_n8883_, new_n8884_, new_n8885_, new_n8886_,
    new_n8887_, new_n8888_, new_n8889_, new_n8890_, new_n8891_, new_n8892_,
    new_n8893_, new_n8894_, new_n8895_, new_n8896_, new_n8897_, new_n8898_,
    new_n8899_, new_n8900_, new_n8901_, new_n8902_, new_n8903_, new_n8904_,
    new_n8905_, new_n8906_, new_n8907_, new_n8908_, new_n8909_, new_n8910_,
    new_n8911_, new_n8912_, new_n8913_, new_n8914_, new_n8915_, new_n8916_,
    new_n8917_, new_n8918_, new_n8919_, new_n8920_, new_n8921_, new_n8922_,
    new_n8923_, new_n8924_, new_n8925_, new_n8926_, new_n8927_, new_n8928_,
    new_n8929_, new_n8930_, new_n8931_, new_n8932_, new_n8933_, new_n8934_,
    new_n8935_, new_n8936_, new_n8937_, new_n8938_, new_n8939_, new_n8940_,
    new_n8941_, new_n8942_, new_n8943_, new_n8944_, new_n8945_, new_n8947_,
    new_n8948_, new_n8949_, new_n8950_, new_n8951_, new_n8952_, new_n8953_,
    new_n8954_, new_n8955_, new_n8956_, new_n8957_, new_n8958_, new_n8959_,
    new_n8960_, new_n8961_, new_n8962_, new_n8963_, new_n8964_, new_n8965_,
    new_n8966_, new_n8967_, new_n8968_, new_n8969_, new_n8970_, new_n8971_,
    new_n8972_, new_n8973_, new_n8974_, new_n8975_, new_n8976_, new_n8977_,
    new_n8978_, new_n8979_, new_n8980_, new_n8981_, new_n8982_, new_n8983_,
    new_n8984_, new_n8985_, new_n8986_, new_n8987_, new_n8988_, new_n8989_,
    new_n8990_, new_n8991_, new_n8992_, new_n8993_, new_n8994_, new_n8995_,
    new_n8996_, new_n8997_, new_n8998_, new_n8999_, new_n9000_, new_n9001_,
    new_n9002_, new_n9003_, new_n9004_, new_n9005_, new_n9006_, new_n9007_,
    new_n9008_, new_n9009_, new_n9010_, new_n9011_, new_n9012_, new_n9013_,
    new_n9014_, new_n9015_, new_n9016_, new_n9017_, new_n9018_, new_n9019_,
    new_n9020_, new_n9021_, new_n9022_, new_n9023_, new_n9024_, new_n9025_,
    new_n9026_, new_n9027_, new_n9028_, new_n9029_, new_n9030_, new_n9031_,
    new_n9032_, new_n9033_, new_n9034_, new_n9035_, new_n9036_, new_n9037_,
    new_n9038_, new_n9039_, new_n9040_, new_n9041_, new_n9042_, new_n9043_,
    new_n9044_, new_n9045_, new_n9046_, new_n9047_, new_n9048_, new_n9049_,
    new_n9050_, new_n9051_, new_n9052_, new_n9053_, new_n9054_, new_n9055_,
    new_n9056_, new_n9057_, new_n9058_, new_n9059_, new_n9060_, new_n9061_,
    new_n9062_, new_n9063_, new_n9064_, new_n9065_, new_n9066_, new_n9067_,
    new_n9068_, new_n9069_, new_n9070_, new_n9071_, new_n9072_, new_n9073_,
    new_n9074_, new_n9075_, new_n9076_, new_n9077_, new_n9078_, new_n9079_,
    new_n9080_, new_n9081_, new_n9082_, new_n9083_, new_n9084_, new_n9085_,
    new_n9086_, new_n9087_, new_n9088_, new_n9089_, new_n9090_, new_n9091_,
    new_n9092_, new_n9093_, new_n9094_, new_n9095_, new_n9096_, new_n9097_,
    new_n9098_, new_n9099_, new_n9100_, new_n9101_, new_n9102_, new_n9103_,
    new_n9104_, new_n9105_, new_n9106_, new_n9107_, new_n9108_, new_n9109_,
    new_n9110_, new_n9111_, new_n9112_, new_n9113_, new_n9114_, new_n9115_,
    new_n9116_, new_n9117_, new_n9118_, new_n9119_, new_n9120_, new_n9121_,
    new_n9122_, new_n9123_, new_n9124_, new_n9125_, new_n9126_, new_n9127_,
    new_n9128_, new_n9129_, new_n9130_, new_n9131_, new_n9132_, new_n9133_,
    new_n9134_, new_n9135_, new_n9136_, new_n9137_, new_n9138_, new_n9139_,
    new_n9140_, new_n9141_, new_n9142_, new_n9143_, new_n9144_, new_n9145_,
    new_n9146_, new_n9147_, new_n9148_, new_n9149_, new_n9150_, new_n9151_,
    new_n9152_, new_n9153_, new_n9154_, new_n9155_, new_n9156_, new_n9157_,
    new_n9158_, new_n9159_, new_n9160_, new_n9161_, new_n9162_, new_n9163_,
    new_n9164_, new_n9165_, new_n9166_, new_n9167_, new_n9168_, new_n9169_,
    new_n9170_, new_n9171_, new_n9172_, new_n9173_, new_n9174_, new_n9175_,
    new_n9176_, new_n9177_, new_n9178_, new_n9179_, new_n9180_, new_n9181_,
    new_n9182_, new_n9183_, new_n9184_, new_n9185_, new_n9186_, new_n9187_,
    new_n9188_, new_n9189_, new_n9190_, new_n9191_, new_n9192_, new_n9193_,
    new_n9194_, new_n9195_, new_n9196_, new_n9197_, new_n9198_, new_n9199_,
    new_n9200_, new_n9201_, new_n9202_, new_n9203_, new_n9204_, new_n9205_,
    new_n9206_, new_n9207_, new_n9208_, new_n9209_, new_n9210_, new_n9211_,
    new_n9212_, new_n9213_, new_n9214_, new_n9215_, new_n9216_, new_n9217_,
    new_n9218_, new_n9219_, new_n9220_, new_n9221_, new_n9222_, new_n9223_,
    new_n9224_, new_n9225_, new_n9226_, new_n9227_, new_n9228_, new_n9229_,
    new_n9230_, new_n9231_, new_n9232_, new_n9233_, new_n9234_, new_n9235_,
    new_n9236_, new_n9237_, new_n9238_, new_n9239_, new_n9240_, new_n9241_,
    new_n9242_, new_n9243_, new_n9244_, new_n9245_, new_n9246_, new_n9247_,
    new_n9248_, new_n9249_, new_n9250_, new_n9251_, new_n9252_, new_n9253_,
    new_n9254_, new_n9255_, new_n9256_, new_n9257_, new_n9258_, new_n9259_,
    new_n9260_, new_n9261_, new_n9262_, new_n9263_, new_n9264_, new_n9265_,
    new_n9266_, new_n9267_, new_n9268_, new_n9269_, new_n9270_, new_n9271_,
    new_n9272_, new_n9273_, new_n9274_, new_n9275_, new_n9276_, new_n9277_,
    new_n9278_, new_n9279_, new_n9280_, new_n9281_, new_n9282_, new_n9283_,
    new_n9284_, new_n9285_, new_n9286_, new_n9287_, new_n9288_, new_n9289_,
    new_n9290_, new_n9291_, new_n9292_, new_n9293_, new_n9294_, new_n9295_,
    new_n9296_, new_n9297_, new_n9298_, new_n9299_, new_n9300_, new_n9301_,
    new_n9302_, new_n9303_, new_n9304_, new_n9305_, new_n9306_, new_n9307_,
    new_n9308_, new_n9309_, new_n9310_, new_n9311_, new_n9312_, new_n9313_,
    new_n9314_, new_n9315_, new_n9316_, new_n9317_, new_n9318_, new_n9319_,
    new_n9320_, new_n9321_, new_n9322_, new_n9323_, new_n9324_, new_n9325_,
    new_n9326_, new_n9327_, new_n9328_, new_n9329_, new_n9330_, new_n9331_,
    new_n9332_, new_n9333_, new_n9334_, new_n9335_, new_n9336_, new_n9337_,
    new_n9338_, new_n9339_, new_n9340_, new_n9341_, new_n9342_, new_n9343_,
    new_n9344_, new_n9345_, new_n9346_, new_n9347_, new_n9348_, new_n9349_,
    new_n9350_, new_n9351_, new_n9352_, new_n9353_, new_n9354_, new_n9355_,
    new_n9356_, new_n9357_, new_n9358_, new_n9359_, new_n9360_, new_n9361_,
    new_n9362_, new_n9363_, new_n9365_, new_n9366_, new_n9367_, new_n9368_,
    new_n9369_, new_n9370_, new_n9371_, new_n9372_, new_n9373_, new_n9374_,
    new_n9375_, new_n9376_, new_n9377_, new_n9378_, new_n9379_, new_n9380_,
    new_n9381_, new_n9382_, new_n9383_, new_n9384_, new_n9385_, new_n9386_,
    new_n9387_, new_n9388_, new_n9389_, new_n9390_, new_n9391_, new_n9392_,
    new_n9393_, new_n9394_, new_n9395_, new_n9396_, new_n9397_, new_n9398_,
    new_n9399_, new_n9400_, new_n9401_, new_n9402_, new_n9403_, new_n9404_,
    new_n9405_, new_n9406_, new_n9407_, new_n9408_, new_n9409_, new_n9410_,
    new_n9411_, new_n9412_, new_n9413_, new_n9414_, new_n9415_, new_n9416_,
    new_n9417_, new_n9418_, new_n9419_, new_n9420_, new_n9421_, new_n9422_,
    new_n9423_, new_n9424_, new_n9425_, new_n9426_, new_n9427_, new_n9428_,
    new_n9429_, new_n9430_, new_n9431_, new_n9432_, new_n9433_, new_n9434_,
    new_n9435_, new_n9436_, new_n9437_, new_n9438_, new_n9439_, new_n9440_,
    new_n9441_, new_n9442_, new_n9443_, new_n9444_, new_n9445_, new_n9446_,
    new_n9447_, new_n9448_, new_n9449_, new_n9450_, new_n9451_, new_n9452_,
    new_n9453_, new_n9454_, new_n9455_, new_n9456_, new_n9457_, new_n9458_,
    new_n9459_, new_n9460_, new_n9461_, new_n9462_, new_n9463_, new_n9464_,
    new_n9465_, new_n9466_, new_n9467_, new_n9468_, new_n9469_, new_n9470_,
    new_n9471_, new_n9472_, new_n9473_, new_n9474_, new_n9475_, new_n9476_,
    new_n9477_, new_n9478_, new_n9479_, new_n9480_, new_n9481_, new_n9482_,
    new_n9483_, new_n9484_, new_n9485_, new_n9486_, new_n9487_, new_n9488_,
    new_n9489_, new_n9490_, new_n9491_, new_n9492_, new_n9493_, new_n9494_,
    new_n9495_, new_n9496_, new_n9497_, new_n9498_, new_n9499_, new_n9500_,
    new_n9501_, new_n9502_, new_n9503_, new_n9504_, new_n9505_, new_n9506_,
    new_n9507_, new_n9508_, new_n9509_, new_n9510_, new_n9511_, new_n9512_,
    new_n9513_, new_n9514_, new_n9515_, new_n9516_, new_n9517_, new_n9518_,
    new_n9519_, new_n9520_, new_n9521_, new_n9522_, new_n9523_, new_n9524_,
    new_n9525_, new_n9526_, new_n9527_, new_n9528_, new_n9529_, new_n9530_,
    new_n9531_, new_n9532_, new_n9533_, new_n9534_, new_n9535_, new_n9536_,
    new_n9537_, new_n9538_, new_n9539_, new_n9540_, new_n9541_, new_n9542_,
    new_n9543_, new_n9544_, new_n9545_, new_n9546_, new_n9547_, new_n9548_,
    new_n9549_, new_n9550_, new_n9551_, new_n9552_, new_n9553_, new_n9554_,
    new_n9555_, new_n9556_, new_n9557_, new_n9558_, new_n9559_, new_n9560_,
    new_n9561_, new_n9562_, new_n9563_, new_n9564_, new_n9565_, new_n9566_,
    new_n9567_, new_n9568_, new_n9569_, new_n9570_, new_n9571_, new_n9572_,
    new_n9573_, new_n9574_, new_n9575_, new_n9576_, new_n9577_, new_n9578_,
    new_n9579_, new_n9580_, new_n9581_, new_n9582_, new_n9583_, new_n9584_,
    new_n9585_, new_n9586_, new_n9587_, new_n9588_, new_n9589_, new_n9590_,
    new_n9591_, new_n9592_, new_n9593_, new_n9594_, new_n9595_, new_n9596_,
    new_n9597_, new_n9598_, new_n9599_, new_n9600_, new_n9601_, new_n9602_,
    new_n9603_, new_n9604_, new_n9605_, new_n9606_, new_n9607_, new_n9608_,
    new_n9609_, new_n9610_, new_n9611_, new_n9612_, new_n9613_, new_n9614_,
    new_n9615_, new_n9616_, new_n9617_, new_n9618_, new_n9619_, new_n9620_,
    new_n9621_, new_n9622_, new_n9623_, new_n9624_, new_n9625_, new_n9626_,
    new_n9627_, new_n9628_, new_n9629_, new_n9630_, new_n9631_, new_n9632_,
    new_n9633_, new_n9634_, new_n9635_, new_n9636_, new_n9637_, new_n9638_,
    new_n9639_, new_n9640_, new_n9641_, new_n9642_, new_n9643_, new_n9644_,
    new_n9645_, new_n9646_, new_n9647_, new_n9648_, new_n9649_, new_n9650_,
    new_n9651_, new_n9652_, new_n9653_, new_n9654_, new_n9655_, new_n9656_,
    new_n9657_, new_n9658_, new_n9659_, new_n9660_, new_n9661_, new_n9662_,
    new_n9663_, new_n9664_, new_n9665_, new_n9666_, new_n9667_, new_n9668_,
    new_n9669_, new_n9670_, new_n9671_, new_n9672_, new_n9673_, new_n9674_,
    new_n9675_, new_n9676_, new_n9677_, new_n9678_, new_n9679_, new_n9680_,
    new_n9681_, new_n9682_, new_n9683_, new_n9684_, new_n9685_, new_n9686_,
    new_n9687_, new_n9688_, new_n9689_, new_n9690_, new_n9691_, new_n9692_,
    new_n9693_, new_n9694_, new_n9695_, new_n9696_, new_n9697_, new_n9698_,
    new_n9699_, new_n9700_, new_n9701_, new_n9702_, new_n9703_, new_n9704_,
    new_n9705_, new_n9706_, new_n9707_, new_n9708_, new_n9709_, new_n9710_,
    new_n9711_, new_n9712_, new_n9713_, new_n9714_, new_n9715_, new_n9716_,
    new_n9717_, new_n9718_, new_n9719_, new_n9720_, new_n9721_, new_n9722_,
    new_n9723_, new_n9724_, new_n9725_, new_n9726_, new_n9727_, new_n9728_,
    new_n9729_, new_n9730_, new_n9731_, new_n9732_, new_n9733_, new_n9734_,
    new_n9735_, new_n9736_, new_n9737_, new_n9738_, new_n9739_, new_n9740_,
    new_n9741_, new_n9742_, new_n9743_, new_n9744_, new_n9745_, new_n9746_,
    new_n9747_, new_n9748_, new_n9749_, new_n9750_, new_n9751_, new_n9752_,
    new_n9753_, new_n9754_, new_n9755_, new_n9756_, new_n9757_, new_n9758_,
    new_n9759_, new_n9760_, new_n9761_, new_n9762_, new_n9763_, new_n9764_,
    new_n9765_, new_n9766_, new_n9767_, new_n9768_, new_n9769_, new_n9770_,
    new_n9771_, new_n9772_, new_n9773_, new_n9774_, new_n9775_, new_n9776_,
    new_n9777_, new_n9778_, new_n9779_, new_n9780_, new_n9781_, new_n9782_,
    new_n9783_, new_n9784_, new_n9785_, new_n9786_, new_n9787_, new_n9788_,
    new_n9789_, new_n9790_, new_n9791_, new_n9792_, new_n9793_, new_n9794_,
    new_n9795_, new_n9796_, new_n9797_, new_n9798_, new_n9799_, new_n9800_,
    new_n9801_, new_n9802_, new_n9803_, new_n9804_, new_n9805_, new_n9806_,
    new_n9807_, new_n9808_, new_n9809_, new_n9810_, new_n9811_, new_n9812_,
    new_n9813_, new_n9814_, new_n9815_, new_n9816_, new_n9817_, new_n9818_,
    new_n9819_, new_n9820_, new_n9821_, new_n9822_, new_n9823_, new_n9824_,
    new_n9825_, new_n9826_, new_n9827_, new_n9828_, new_n9829_, new_n9830_,
    new_n9831_, new_n9832_, new_n9833_, new_n9835_, new_n9836_, new_n9837_,
    new_n9838_, new_n9839_, new_n9840_, new_n9841_, new_n9842_, new_n9843_,
    new_n9844_, new_n9845_, new_n9846_, new_n9847_, new_n9848_, new_n9849_,
    new_n9850_, new_n9851_, new_n9852_, new_n9853_, new_n9854_, new_n9855_,
    new_n9856_, new_n9857_, new_n9858_, new_n9859_, new_n9860_, new_n9861_,
    new_n9862_, new_n9863_, new_n9864_, new_n9865_, new_n9866_, new_n9867_,
    new_n9868_, new_n9869_, new_n9870_, new_n9871_, new_n9872_, new_n9873_,
    new_n9874_, new_n9875_, new_n9876_, new_n9877_, new_n9878_, new_n9879_,
    new_n9880_, new_n9881_, new_n9882_, new_n9883_, new_n9884_, new_n9885_,
    new_n9886_, new_n9887_, new_n9888_, new_n9889_, new_n9890_, new_n9891_,
    new_n9892_, new_n9893_, new_n9894_, new_n9895_, new_n9896_, new_n9897_,
    new_n9898_, new_n9899_, new_n9900_, new_n9901_, new_n9902_, new_n9903_,
    new_n9904_, new_n9905_, new_n9906_, new_n9907_, new_n9908_, new_n9909_,
    new_n9910_, new_n9911_, new_n9912_, new_n9913_, new_n9914_, new_n9915_,
    new_n9916_, new_n9917_, new_n9918_, new_n9919_, new_n9920_, new_n9921_,
    new_n9922_, new_n9923_, new_n9924_, new_n9925_, new_n9926_, new_n9927_,
    new_n9928_, new_n9929_, new_n9930_, new_n9931_, new_n9932_, new_n9933_,
    new_n9934_, new_n9935_, new_n9936_, new_n9937_, new_n9938_, new_n9939_,
    new_n9940_, new_n9941_, new_n9942_, new_n9943_, new_n9944_, new_n9945_,
    new_n9946_, new_n9947_, new_n9948_, new_n9949_, new_n9950_, new_n9951_,
    new_n9952_, new_n9953_, new_n9954_, new_n9955_, new_n9956_, new_n9957_,
    new_n9958_, new_n9959_, new_n9960_, new_n9961_, new_n9962_, new_n9963_,
    new_n9964_, new_n9965_, new_n9966_, new_n9967_, new_n9968_, new_n9969_,
    new_n9970_, new_n9971_, new_n9972_, new_n9973_, new_n9974_, new_n9975_,
    new_n9976_, new_n9977_, new_n9978_, new_n9979_, new_n9980_, new_n9981_,
    new_n9982_, new_n9983_, new_n9984_, new_n9985_, new_n9986_, new_n9987_,
    new_n9988_, new_n9989_, new_n9990_, new_n9991_, new_n9992_, new_n9993_,
    new_n9994_, new_n9995_, new_n9996_, new_n9997_, new_n9998_, new_n9999_,
    new_n10000_, new_n10001_, new_n10002_, new_n10003_, new_n10004_,
    new_n10005_, new_n10006_, new_n10007_, new_n10008_, new_n10009_,
    new_n10010_, new_n10011_, new_n10012_, new_n10013_, new_n10014_,
    new_n10015_, new_n10016_, new_n10017_, new_n10018_, new_n10019_,
    new_n10020_, new_n10021_, new_n10022_, new_n10023_, new_n10024_,
    new_n10025_, new_n10026_, new_n10027_, new_n10028_, new_n10029_,
    new_n10030_, new_n10031_, new_n10032_, new_n10033_, new_n10034_,
    new_n10035_, new_n10036_, new_n10037_, new_n10038_, new_n10039_,
    new_n10040_, new_n10041_, new_n10042_, new_n10043_, new_n10044_,
    new_n10045_, new_n10046_, new_n10047_, new_n10048_, new_n10049_,
    new_n10050_, new_n10051_, new_n10052_, new_n10053_, new_n10054_,
    new_n10055_, new_n10056_, new_n10057_, new_n10058_, new_n10059_,
    new_n10060_, new_n10061_, new_n10062_, new_n10063_, new_n10064_,
    new_n10065_, new_n10066_, new_n10067_, new_n10068_, new_n10069_,
    new_n10070_, new_n10071_, new_n10072_, new_n10073_, new_n10074_,
    new_n10075_, new_n10076_, new_n10077_, new_n10078_, new_n10079_,
    new_n10080_, new_n10081_, new_n10082_, new_n10083_, new_n10084_,
    new_n10085_, new_n10086_, new_n10087_, new_n10088_, new_n10089_,
    new_n10090_, new_n10091_, new_n10092_, new_n10093_, new_n10094_,
    new_n10095_, new_n10096_, new_n10097_, new_n10098_, new_n10099_,
    new_n10100_, new_n10101_, new_n10102_, new_n10103_, new_n10104_,
    new_n10105_, new_n10106_, new_n10107_, new_n10108_, new_n10109_,
    new_n10110_, new_n10111_, new_n10112_, new_n10113_, new_n10114_,
    new_n10115_, new_n10116_, new_n10117_, new_n10118_, new_n10119_,
    new_n10120_, new_n10121_, new_n10122_, new_n10123_, new_n10124_,
    new_n10125_, new_n10126_, new_n10127_, new_n10128_, new_n10129_,
    new_n10130_, new_n10131_, new_n10132_, new_n10133_, new_n10134_,
    new_n10135_, new_n10136_, new_n10137_, new_n10138_, new_n10139_,
    new_n10140_, new_n10141_, new_n10142_, new_n10143_, new_n10144_,
    new_n10145_, new_n10146_, new_n10147_, new_n10148_, new_n10149_,
    new_n10150_, new_n10151_, new_n10152_, new_n10153_, new_n10154_,
    new_n10155_, new_n10156_, new_n10157_, new_n10158_, new_n10159_,
    new_n10160_, new_n10161_, new_n10162_, new_n10163_, new_n10164_,
    new_n10165_, new_n10166_, new_n10167_, new_n10168_, new_n10169_,
    new_n10170_, new_n10171_, new_n10172_, new_n10173_, new_n10174_,
    new_n10175_, new_n10176_, new_n10177_, new_n10178_, new_n10179_,
    new_n10180_, new_n10181_, new_n10182_, new_n10183_, new_n10184_,
    new_n10185_, new_n10186_, new_n10187_, new_n10188_, new_n10189_,
    new_n10190_, new_n10191_, new_n10192_, new_n10193_, new_n10194_,
    new_n10195_, new_n10196_, new_n10197_, new_n10198_, new_n10199_,
    new_n10200_, new_n10201_, new_n10202_, new_n10203_, new_n10204_,
    new_n10205_, new_n10206_, new_n10207_, new_n10208_, new_n10209_,
    new_n10210_, new_n10211_, new_n10212_, new_n10213_, new_n10214_,
    new_n10215_, new_n10216_, new_n10217_, new_n10218_, new_n10219_,
    new_n10220_, new_n10221_, new_n10222_, new_n10223_, new_n10224_,
    new_n10225_, new_n10226_, new_n10227_, new_n10228_, new_n10229_,
    new_n10230_, new_n10231_, new_n10232_, new_n10233_, new_n10234_,
    new_n10235_, new_n10236_, new_n10237_, new_n10238_, new_n10239_,
    new_n10240_, new_n10241_, new_n10242_, new_n10243_, new_n10244_,
    new_n10245_, new_n10246_, new_n10247_, new_n10248_, new_n10249_,
    new_n10250_, new_n10251_, new_n10252_, new_n10253_, new_n10254_,
    new_n10255_, new_n10256_, new_n10257_, new_n10258_, new_n10259_,
    new_n10260_, new_n10261_, new_n10262_, new_n10263_, new_n10264_,
    new_n10265_, new_n10266_, new_n10267_, new_n10268_, new_n10269_,
    new_n10270_, new_n10271_, new_n10272_, new_n10273_, new_n10274_,
    new_n10275_, new_n10276_, new_n10277_, new_n10278_, new_n10279_,
    new_n10280_, new_n10281_, new_n10282_, new_n10283_, new_n10284_,
    new_n10285_, new_n10286_, new_n10287_, new_n10288_, new_n10289_,
    new_n10290_, new_n10291_, new_n10292_, new_n10293_, new_n10294_,
    new_n10295_, new_n10296_, new_n10297_, new_n10298_, new_n10299_,
    new_n10300_, new_n10301_, new_n10302_, new_n10303_, new_n10304_,
    new_n10305_, new_n10306_, new_n10307_, new_n10308_, new_n10309_,
    new_n10310_, new_n10311_, new_n10312_, new_n10313_, new_n10314_,
    new_n10315_, new_n10316_, new_n10317_, new_n10318_, new_n10319_,
    new_n10320_, new_n10321_, new_n10322_, new_n10323_, new_n10324_,
    new_n10325_, new_n10326_, new_n10327_, new_n10328_, new_n10329_,
    new_n10330_, new_n10331_, new_n10332_, new_n10333_, new_n10334_,
    new_n10335_, new_n10336_, new_n10337_, new_n10338_, new_n10339_,
    new_n10340_, new_n10341_, new_n10342_, new_n10343_, new_n10344_,
    new_n10345_, new_n10346_, new_n10347_, new_n10348_, new_n10349_,
    new_n10350_, new_n10351_, new_n10352_, new_n10353_, new_n10354_,
    new_n10355_, new_n10356_, new_n10357_, new_n10358_, new_n10359_,
    new_n10360_, new_n10361_, new_n10362_, new_n10363_, new_n10364_,
    new_n10365_, new_n10366_, new_n10367_, new_n10368_, new_n10369_,
    new_n10370_, new_n10371_, new_n10372_, new_n10373_, new_n10374_,
    new_n10375_, new_n10376_, new_n10377_, new_n10378_, new_n10379_,
    new_n10380_, new_n10381_, new_n10382_, new_n10383_, new_n10384_,
    new_n10385_, new_n10386_, new_n10387_, new_n10388_, new_n10389_,
    new_n10390_, new_n10391_, new_n10392_, new_n10393_, new_n10394_,
    new_n10395_, new_n10396_, new_n10397_, new_n10398_, new_n10399_,
    new_n10400_, new_n10401_, new_n10402_, new_n10403_, new_n10404_,
    new_n10405_, new_n10406_, new_n10407_, new_n10408_, new_n10409_,
    new_n10410_, new_n10411_, new_n10412_, new_n10413_, new_n10414_,
    new_n10415_, new_n10417_, new_n10418_, new_n10419_, new_n10420_,
    new_n10421_, new_n10422_, new_n10423_, new_n10424_, new_n10425_,
    new_n10426_, new_n10427_, new_n10428_, new_n10429_, new_n10430_,
    new_n10431_, new_n10432_, new_n10433_, new_n10434_, new_n10435_,
    new_n10436_, new_n10437_, new_n10438_, new_n10439_, new_n10440_,
    new_n10441_, new_n10442_, new_n10443_, new_n10444_, new_n10445_,
    new_n10446_, new_n10447_, new_n10448_, new_n10449_, new_n10450_,
    new_n10451_, new_n10452_, new_n10453_, new_n10454_, new_n10455_,
    new_n10456_, new_n10457_, new_n10458_, new_n10459_, new_n10460_,
    new_n10461_, new_n10462_, new_n10463_, new_n10464_, new_n10465_,
    new_n10466_, new_n10467_, new_n10468_, new_n10469_, new_n10470_,
    new_n10471_, new_n10472_, new_n10473_, new_n10474_, new_n10475_,
    new_n10476_, new_n10477_, new_n10478_, new_n10479_, new_n10480_,
    new_n10481_, new_n10482_, new_n10483_, new_n10484_, new_n10485_,
    new_n10486_, new_n10487_, new_n10488_, new_n10489_, new_n10490_,
    new_n10491_, new_n10492_, new_n10493_, new_n10494_, new_n10495_,
    new_n10496_, new_n10497_, new_n10498_, new_n10499_, new_n10500_,
    new_n10501_, new_n10502_, new_n10503_, new_n10504_, new_n10505_,
    new_n10506_, new_n10507_, new_n10508_, new_n10509_, new_n10510_,
    new_n10511_, new_n10512_, new_n10513_, new_n10514_, new_n10515_,
    new_n10516_, new_n10517_, new_n10518_, new_n10519_, new_n10520_,
    new_n10521_, new_n10522_, new_n10523_, new_n10524_, new_n10525_,
    new_n10526_, new_n10527_, new_n10528_, new_n10529_, new_n10530_,
    new_n10531_, new_n10532_, new_n10533_, new_n10534_, new_n10535_,
    new_n10536_, new_n10537_, new_n10538_, new_n10539_, new_n10540_,
    new_n10541_, new_n10542_, new_n10543_, new_n10544_, new_n10545_,
    new_n10546_, new_n10547_, new_n10548_, new_n10549_, new_n10550_,
    new_n10551_, new_n10552_, new_n10553_, new_n10554_, new_n10555_,
    new_n10556_, new_n10557_, new_n10558_, new_n10559_, new_n10560_,
    new_n10561_, new_n10562_, new_n10563_, new_n10564_, new_n10565_,
    new_n10566_, new_n10567_, new_n10568_, new_n10569_, new_n10570_,
    new_n10571_, new_n10572_, new_n10573_, new_n10574_, new_n10575_,
    new_n10576_, new_n10577_, new_n10578_, new_n10579_, new_n10580_,
    new_n10581_, new_n10582_, new_n10583_, new_n10584_, new_n10585_,
    new_n10586_, new_n10587_, new_n10588_, new_n10589_, new_n10590_,
    new_n10591_, new_n10592_, new_n10593_, new_n10594_, new_n10595_,
    new_n10596_, new_n10597_, new_n10598_, new_n10599_, new_n10600_,
    new_n10601_, new_n10602_, new_n10603_, new_n10604_, new_n10605_,
    new_n10606_, new_n10607_, new_n10608_, new_n10609_, new_n10610_,
    new_n10611_, new_n10612_, new_n10613_, new_n10614_, new_n10615_,
    new_n10616_, new_n10617_, new_n10618_, new_n10619_, new_n10620_,
    new_n10621_, new_n10622_, new_n10623_, new_n10624_, new_n10625_,
    new_n10626_, new_n10627_, new_n10628_, new_n10629_, new_n10630_,
    new_n10631_, new_n10632_, new_n10633_, new_n10634_, new_n10635_,
    new_n10636_, new_n10637_, new_n10638_, new_n10639_, new_n10640_,
    new_n10641_, new_n10642_, new_n10643_, new_n10644_, new_n10645_,
    new_n10646_, new_n10647_, new_n10648_, new_n10649_, new_n10650_,
    new_n10651_, new_n10652_, new_n10653_, new_n10654_, new_n10655_,
    new_n10656_, new_n10657_, new_n10658_, new_n10659_, new_n10660_,
    new_n10661_, new_n10662_, new_n10663_, new_n10664_, new_n10665_,
    new_n10666_, new_n10667_, new_n10668_, new_n10669_, new_n10670_,
    new_n10671_, new_n10672_, new_n10673_, new_n10674_, new_n10675_,
    new_n10676_, new_n10677_, new_n10678_, new_n10679_, new_n10680_,
    new_n10681_, new_n10682_, new_n10683_, new_n10684_, new_n10685_,
    new_n10686_, new_n10687_, new_n10688_, new_n10689_, new_n10690_,
    new_n10691_, new_n10692_, new_n10693_, new_n10694_, new_n10695_,
    new_n10696_, new_n10697_, new_n10698_, new_n10699_, new_n10700_,
    new_n10701_, new_n10702_, new_n10703_, new_n10704_, new_n10705_,
    new_n10706_, new_n10707_, new_n10708_, new_n10709_, new_n10710_,
    new_n10711_, new_n10712_, new_n10713_, new_n10714_, new_n10715_,
    new_n10716_, new_n10717_, new_n10718_, new_n10719_, new_n10720_,
    new_n10721_, new_n10722_, new_n10723_, new_n10724_, new_n10725_,
    new_n10726_, new_n10727_, new_n10728_, new_n10729_, new_n10730_,
    new_n10731_, new_n10732_, new_n10733_, new_n10734_, new_n10735_,
    new_n10736_, new_n10737_, new_n10738_, new_n10739_, new_n10740_,
    new_n10741_, new_n10742_, new_n10743_, new_n10744_, new_n10745_,
    new_n10746_, new_n10747_, new_n10748_, new_n10749_, new_n10750_,
    new_n10751_, new_n10752_, new_n10753_, new_n10754_, new_n10755_,
    new_n10756_, new_n10757_, new_n10758_, new_n10759_, new_n10760_,
    new_n10761_, new_n10762_, new_n10763_, new_n10764_, new_n10765_,
    new_n10766_, new_n10767_, new_n10768_, new_n10769_, new_n10770_,
    new_n10771_, new_n10772_, new_n10773_, new_n10774_, new_n10775_,
    new_n10776_, new_n10777_, new_n10778_, new_n10779_, new_n10780_,
    new_n10781_, new_n10782_, new_n10783_, new_n10784_, new_n10785_,
    new_n10786_, new_n10787_, new_n10788_, new_n10789_, new_n10790_,
    new_n10791_, new_n10792_, new_n10793_, new_n10794_, new_n10795_,
    new_n10796_, new_n10797_, new_n10798_, new_n10799_, new_n10800_,
    new_n10801_, new_n10802_, new_n10803_, new_n10804_, new_n10805_,
    new_n10806_, new_n10807_, new_n10808_, new_n10809_, new_n10810_,
    new_n10811_, new_n10812_, new_n10813_, new_n10814_, new_n10815_,
    new_n10816_, new_n10817_, new_n10818_, new_n10819_, new_n10820_,
    new_n10821_, new_n10822_, new_n10823_, new_n10824_, new_n10825_,
    new_n10826_, new_n10827_, new_n10828_, new_n10829_, new_n10830_,
    new_n10831_, new_n10832_, new_n10833_, new_n10834_, new_n10835_,
    new_n10836_, new_n10837_, new_n10838_, new_n10839_, new_n10840_,
    new_n10841_, new_n10842_, new_n10843_, new_n10844_, new_n10845_,
    new_n10846_, new_n10847_, new_n10848_, new_n10849_, new_n10850_,
    new_n10851_, new_n10852_, new_n10853_, new_n10854_, new_n10855_,
    new_n10856_, new_n10857_, new_n10858_, new_n10859_, new_n10860_,
    new_n10861_, new_n10862_, new_n10863_, new_n10864_, new_n10865_,
    new_n10866_, new_n10867_, new_n10868_, new_n10869_, new_n10870_,
    new_n10871_, new_n10872_, new_n10873_, new_n10874_, new_n10875_,
    new_n10877_, new_n10878_, new_n10879_, new_n10880_, new_n10881_,
    new_n10882_, new_n10883_, new_n10884_, new_n10885_, new_n10886_,
    new_n10887_, new_n10888_, new_n10889_, new_n10890_, new_n10891_,
    new_n10892_, new_n10893_, new_n10894_, new_n10895_, new_n10896_,
    new_n10897_, new_n10898_, new_n10899_, new_n10900_, new_n10901_,
    new_n10902_, new_n10903_, new_n10904_, new_n10905_, new_n10906_,
    new_n10907_, new_n10908_, new_n10909_, new_n10910_, new_n10911_,
    new_n10912_, new_n10913_, new_n10914_, new_n10915_, new_n10916_,
    new_n10917_, new_n10918_, new_n10919_, new_n10920_, new_n10921_,
    new_n10922_, new_n10923_, new_n10924_, new_n10925_, new_n10926_,
    new_n10927_, new_n10928_, new_n10929_, new_n10930_, new_n10931_,
    new_n10932_, new_n10933_, new_n10934_, new_n10935_, new_n10936_,
    new_n10937_, new_n10938_, new_n10939_, new_n10940_, new_n10941_,
    new_n10942_, new_n10943_, new_n10944_, new_n10945_, new_n10946_,
    new_n10947_, new_n10948_, new_n10949_, new_n10950_, new_n10951_,
    new_n10952_, new_n10953_, new_n10954_, new_n10955_, new_n10956_,
    new_n10957_, new_n10958_, new_n10959_, new_n10960_, new_n10961_,
    new_n10962_, new_n10963_, new_n10964_, new_n10965_, new_n10966_,
    new_n10967_, new_n10968_, new_n10969_, new_n10970_, new_n10971_,
    new_n10972_, new_n10973_, new_n10974_, new_n10975_, new_n10976_,
    new_n10977_, new_n10978_, new_n10979_, new_n10980_, new_n10981_,
    new_n10982_, new_n10983_, new_n10984_, new_n10985_, new_n10986_,
    new_n10987_, new_n10988_, new_n10989_, new_n10990_, new_n10991_,
    new_n10992_, new_n10993_, new_n10994_, new_n10995_, new_n10996_,
    new_n10997_, new_n10998_, new_n10999_, new_n11000_, new_n11001_,
    new_n11002_, new_n11003_, new_n11004_, new_n11005_, new_n11006_,
    new_n11007_, new_n11008_, new_n11009_, new_n11010_, new_n11011_,
    new_n11012_, new_n11013_, new_n11014_, new_n11015_, new_n11016_,
    new_n11017_, new_n11018_, new_n11019_, new_n11020_, new_n11021_,
    new_n11022_, new_n11023_, new_n11024_, new_n11025_, new_n11026_,
    new_n11027_, new_n11028_, new_n11029_, new_n11030_, new_n11031_,
    new_n11032_, new_n11033_, new_n11034_, new_n11035_, new_n11036_,
    new_n11037_, new_n11038_, new_n11039_, new_n11040_, new_n11041_,
    new_n11042_, new_n11043_, new_n11044_, new_n11045_, new_n11046_,
    new_n11047_, new_n11048_, new_n11049_, new_n11050_, new_n11051_,
    new_n11052_, new_n11053_, new_n11054_, new_n11055_, new_n11056_,
    new_n11057_, new_n11058_, new_n11059_, new_n11060_, new_n11061_,
    new_n11062_, new_n11063_, new_n11064_, new_n11065_, new_n11066_,
    new_n11067_, new_n11068_, new_n11069_, new_n11070_, new_n11071_,
    new_n11072_, new_n11073_, new_n11074_, new_n11075_, new_n11076_,
    new_n11077_, new_n11078_, new_n11079_, new_n11080_, new_n11081_,
    new_n11082_, new_n11083_, new_n11084_, new_n11085_, new_n11086_,
    new_n11087_, new_n11088_, new_n11089_, new_n11090_, new_n11091_,
    new_n11092_, new_n11093_, new_n11094_, new_n11095_, new_n11096_,
    new_n11097_, new_n11098_, new_n11099_, new_n11100_, new_n11101_,
    new_n11102_, new_n11103_, new_n11104_, new_n11105_, new_n11106_,
    new_n11107_, new_n11108_, new_n11109_, new_n11110_, new_n11111_,
    new_n11112_, new_n11113_, new_n11114_, new_n11115_, new_n11116_,
    new_n11117_, new_n11118_, new_n11119_, new_n11120_, new_n11121_,
    new_n11122_, new_n11123_, new_n11124_, new_n11125_, new_n11126_,
    new_n11127_, new_n11128_, new_n11129_, new_n11130_, new_n11131_,
    new_n11132_, new_n11133_, new_n11134_, new_n11135_, new_n11136_,
    new_n11137_, new_n11138_, new_n11139_, new_n11140_, new_n11141_,
    new_n11142_, new_n11143_, new_n11144_, new_n11145_, new_n11146_,
    new_n11147_, new_n11148_, new_n11149_, new_n11150_, new_n11151_,
    new_n11152_, new_n11153_, new_n11154_, new_n11155_, new_n11156_,
    new_n11157_, new_n11158_, new_n11159_, new_n11160_, new_n11161_,
    new_n11162_, new_n11163_, new_n11164_, new_n11165_, new_n11166_,
    new_n11167_, new_n11168_, new_n11169_, new_n11170_, new_n11171_,
    new_n11172_, new_n11173_, new_n11174_, new_n11175_, new_n11176_,
    new_n11177_, new_n11178_, new_n11179_, new_n11180_, new_n11181_,
    new_n11182_, new_n11183_, new_n11184_, new_n11185_, new_n11186_,
    new_n11187_, new_n11188_, new_n11189_, new_n11190_, new_n11191_,
    new_n11192_, new_n11193_, new_n11194_, new_n11195_, new_n11196_,
    new_n11197_, new_n11198_, new_n11199_, new_n11200_, new_n11201_,
    new_n11202_, new_n11203_, new_n11204_, new_n11205_, new_n11206_,
    new_n11207_, new_n11208_, new_n11209_, new_n11210_, new_n11211_,
    new_n11212_, new_n11213_, new_n11214_, new_n11215_, new_n11216_,
    new_n11217_, new_n11218_, new_n11219_, new_n11220_, new_n11221_,
    new_n11222_, new_n11223_, new_n11224_, new_n11225_, new_n11226_,
    new_n11227_, new_n11228_, new_n11229_, new_n11230_, new_n11231_,
    new_n11232_, new_n11233_, new_n11234_, new_n11235_, new_n11236_,
    new_n11237_, new_n11238_, new_n11239_, new_n11240_, new_n11241_,
    new_n11242_, new_n11243_, new_n11244_, new_n11245_, new_n11246_,
    new_n11247_, new_n11248_, new_n11249_, new_n11250_, new_n11251_,
    new_n11252_, new_n11253_, new_n11254_, new_n11255_, new_n11256_,
    new_n11257_, new_n11258_, new_n11259_, new_n11260_, new_n11261_,
    new_n11262_, new_n11263_, new_n11264_, new_n11265_, new_n11266_,
    new_n11267_, new_n11268_, new_n11269_, new_n11270_, new_n11271_,
    new_n11272_, new_n11273_, new_n11274_, new_n11275_, new_n11276_,
    new_n11277_, new_n11278_, new_n11279_, new_n11280_, new_n11281_,
    new_n11282_, new_n11283_, new_n11284_, new_n11285_, new_n11286_,
    new_n11287_, new_n11288_, new_n11289_, new_n11290_, new_n11291_,
    new_n11292_, new_n11293_, new_n11294_, new_n11295_, new_n11296_,
    new_n11297_, new_n11298_, new_n11299_, new_n11300_, new_n11301_,
    new_n11302_, new_n11303_, new_n11304_, new_n11305_, new_n11306_,
    new_n11307_, new_n11308_, new_n11309_, new_n11310_, new_n11311_,
    new_n11312_, new_n11313_, new_n11314_, new_n11315_, new_n11316_,
    new_n11317_, new_n11318_, new_n11319_, new_n11320_, new_n11321_,
    new_n11322_, new_n11323_, new_n11324_, new_n11325_, new_n11326_,
    new_n11327_, new_n11328_, new_n11329_, new_n11330_, new_n11331_,
    new_n11332_, new_n11333_, new_n11334_, new_n11335_, new_n11336_,
    new_n11337_, new_n11338_, new_n11339_, new_n11340_, new_n11341_,
    new_n11342_, new_n11343_, new_n11344_, new_n11345_, new_n11346_,
    new_n11347_, new_n11348_, new_n11349_, new_n11350_, new_n11351_,
    new_n11352_, new_n11353_, new_n11354_, new_n11355_, new_n11356_,
    new_n11357_, new_n11358_, new_n11359_, new_n11360_, new_n11361_,
    new_n11362_, new_n11364_, new_n11365_, new_n11366_, new_n11367_,
    new_n11368_, new_n11369_, new_n11370_, new_n11371_, new_n11372_,
    new_n11373_, new_n11374_, new_n11375_, new_n11376_, new_n11377_,
    new_n11378_, new_n11379_, new_n11380_, new_n11381_, new_n11382_,
    new_n11383_, new_n11384_, new_n11385_, new_n11386_, new_n11387_,
    new_n11388_, new_n11389_, new_n11390_, new_n11391_, new_n11392_,
    new_n11393_, new_n11394_, new_n11395_, new_n11396_, new_n11397_,
    new_n11398_, new_n11399_, new_n11400_, new_n11401_, new_n11402_,
    new_n11403_, new_n11404_, new_n11405_, new_n11406_, new_n11407_,
    new_n11408_, new_n11409_, new_n11410_, new_n11411_, new_n11412_,
    new_n11413_, new_n11414_, new_n11415_, new_n11416_, new_n11417_,
    new_n11418_, new_n11419_, new_n11420_, new_n11421_, new_n11422_,
    new_n11423_, new_n11424_, new_n11425_, new_n11426_, new_n11427_,
    new_n11428_, new_n11429_, new_n11430_, new_n11431_, new_n11432_,
    new_n11433_, new_n11434_, new_n11435_, new_n11436_, new_n11437_,
    new_n11438_, new_n11439_, new_n11440_, new_n11441_, new_n11442_,
    new_n11443_, new_n11444_, new_n11445_, new_n11446_, new_n11447_,
    new_n11448_, new_n11449_, new_n11450_, new_n11451_, new_n11452_,
    new_n11453_, new_n11454_, new_n11455_, new_n11456_, new_n11457_,
    new_n11458_, new_n11459_, new_n11460_, new_n11461_, new_n11462_,
    new_n11463_, new_n11464_, new_n11465_, new_n11466_, new_n11467_,
    new_n11468_, new_n11469_, new_n11470_, new_n11471_, new_n11472_,
    new_n11473_, new_n11474_, new_n11475_, new_n11476_, new_n11477_,
    new_n11478_, new_n11479_, new_n11480_, new_n11481_, new_n11482_,
    new_n11483_, new_n11484_, new_n11485_, new_n11486_, new_n11487_,
    new_n11488_, new_n11489_, new_n11490_, new_n11491_, new_n11492_,
    new_n11493_, new_n11494_, new_n11495_, new_n11496_, new_n11497_,
    new_n11498_, new_n11499_, new_n11500_, new_n11501_, new_n11502_,
    new_n11503_, new_n11504_, new_n11505_, new_n11506_, new_n11507_,
    new_n11508_, new_n11509_, new_n11510_, new_n11511_, new_n11512_,
    new_n11513_, new_n11514_, new_n11515_, new_n11516_, new_n11517_,
    new_n11518_, new_n11519_, new_n11520_, new_n11521_, new_n11522_,
    new_n11523_, new_n11524_, new_n11525_, new_n11526_, new_n11527_,
    new_n11528_, new_n11529_, new_n11530_, new_n11531_, new_n11532_,
    new_n11533_, new_n11534_, new_n11535_, new_n11536_, new_n11537_,
    new_n11538_, new_n11539_, new_n11540_, new_n11541_, new_n11542_,
    new_n11543_, new_n11544_, new_n11545_, new_n11546_, new_n11547_,
    new_n11548_, new_n11549_, new_n11550_, new_n11551_, new_n11552_,
    new_n11553_, new_n11554_, new_n11555_, new_n11556_, new_n11557_,
    new_n11558_, new_n11559_, new_n11560_, new_n11561_, new_n11562_,
    new_n11563_, new_n11564_, new_n11565_, new_n11566_, new_n11567_,
    new_n11568_, new_n11569_, new_n11570_, new_n11571_, new_n11572_,
    new_n11573_, new_n11574_, new_n11575_, new_n11576_, new_n11577_,
    new_n11578_, new_n11579_, new_n11580_, new_n11581_, new_n11582_,
    new_n11583_, new_n11584_, new_n11585_, new_n11586_, new_n11587_,
    new_n11588_, new_n11589_, new_n11590_, new_n11591_, new_n11592_,
    new_n11593_, new_n11594_, new_n11595_, new_n11596_, new_n11597_,
    new_n11598_, new_n11599_, new_n11600_, new_n11601_, new_n11602_,
    new_n11603_, new_n11604_, new_n11605_, new_n11606_, new_n11607_,
    new_n11608_, new_n11609_, new_n11610_, new_n11611_, new_n11612_,
    new_n11613_, new_n11614_, new_n11615_, new_n11616_, new_n11617_,
    new_n11618_, new_n11619_, new_n11620_, new_n11621_, new_n11622_,
    new_n11623_, new_n11624_, new_n11625_, new_n11626_, new_n11627_,
    new_n11628_, new_n11629_, new_n11630_, new_n11631_, new_n11632_,
    new_n11633_, new_n11634_, new_n11635_, new_n11636_, new_n11637_,
    new_n11638_, new_n11639_, new_n11640_, new_n11641_, new_n11642_,
    new_n11643_, new_n11644_, new_n11645_, new_n11646_, new_n11647_,
    new_n11648_, new_n11649_, new_n11650_, new_n11651_, new_n11652_,
    new_n11653_, new_n11654_, new_n11655_, new_n11656_, new_n11657_,
    new_n11658_, new_n11659_, new_n11660_, new_n11661_, new_n11662_,
    new_n11663_, new_n11664_, new_n11665_, new_n11666_, new_n11667_,
    new_n11668_, new_n11669_, new_n11670_, new_n11671_, new_n11672_,
    new_n11673_, new_n11674_, new_n11675_, new_n11676_, new_n11677_,
    new_n11678_, new_n11679_, new_n11680_, new_n11681_, new_n11682_,
    new_n11683_, new_n11684_, new_n11685_, new_n11686_, new_n11687_,
    new_n11688_, new_n11689_, new_n11690_, new_n11691_, new_n11692_,
    new_n11693_, new_n11694_, new_n11695_, new_n11696_, new_n11697_,
    new_n11698_, new_n11699_, new_n11700_, new_n11701_, new_n11702_,
    new_n11703_, new_n11704_, new_n11705_, new_n11706_, new_n11707_,
    new_n11708_, new_n11709_, new_n11710_, new_n11711_, new_n11712_,
    new_n11713_, new_n11714_, new_n11715_, new_n11716_, new_n11717_,
    new_n11718_, new_n11719_, new_n11720_, new_n11721_, new_n11722_,
    new_n11723_, new_n11724_, new_n11725_, new_n11726_, new_n11727_,
    new_n11728_, new_n11729_, new_n11730_, new_n11731_, new_n11732_,
    new_n11733_, new_n11734_, new_n11735_, new_n11736_, new_n11737_,
    new_n11738_, new_n11739_, new_n11740_, new_n11741_, new_n11742_,
    new_n11743_, new_n11744_, new_n11745_, new_n11746_, new_n11747_,
    new_n11748_, new_n11749_, new_n11750_, new_n11751_, new_n11752_,
    new_n11753_, new_n11754_, new_n11755_, new_n11756_, new_n11757_,
    new_n11758_, new_n11759_, new_n11760_, new_n11761_, new_n11762_,
    new_n11763_, new_n11764_, new_n11765_, new_n11766_, new_n11767_,
    new_n11768_, new_n11769_, new_n11770_, new_n11771_, new_n11772_,
    new_n11773_, new_n11774_, new_n11775_, new_n11776_, new_n11777_,
    new_n11778_, new_n11779_, new_n11780_, new_n11781_, new_n11782_,
    new_n11783_, new_n11784_, new_n11785_, new_n11786_, new_n11787_,
    new_n11788_, new_n11789_, new_n11790_, new_n11791_, new_n11792_,
    new_n11793_, new_n11794_, new_n11795_, new_n11796_, new_n11797_,
    new_n11798_, new_n11799_, new_n11800_, new_n11801_, new_n11802_,
    new_n11803_, new_n11804_, new_n11805_, new_n11806_, new_n11807_,
    new_n11808_, new_n11809_, new_n11810_, new_n11811_, new_n11812_,
    new_n11813_, new_n11814_, new_n11815_, new_n11816_, new_n11817_,
    new_n11818_, new_n11819_, new_n11820_, new_n11821_, new_n11822_,
    new_n11823_, new_n11824_, new_n11825_, new_n11826_, new_n11827_,
    new_n11828_, new_n11829_, new_n11830_, new_n11831_, new_n11832_,
    new_n11833_, new_n11834_, new_n11835_, new_n11836_, new_n11837_,
    new_n11838_, new_n11839_, new_n11840_, new_n11841_, new_n11842_,
    new_n11843_, new_n11844_, new_n11845_, new_n11846_, new_n11847_,
    new_n11848_, new_n11849_, new_n11850_, new_n11851_, new_n11852_,
    new_n11853_, new_n11854_, new_n11855_, new_n11856_, new_n11857_,
    new_n11858_, new_n11859_, new_n11860_, new_n11861_, new_n11862_,
    new_n11863_, new_n11864_, new_n11865_, new_n11866_, new_n11867_,
    new_n11868_, new_n11869_, new_n11870_, new_n11871_, new_n11872_,
    new_n11873_, new_n11874_, new_n11875_, new_n11876_, new_n11877_,
    new_n11878_, new_n11879_, new_n11880_, new_n11881_, new_n11882_,
    new_n11883_, new_n11884_, new_n11885_, new_n11886_, new_n11887_,
    new_n11888_, new_n11889_, new_n11890_, new_n11891_, new_n11892_,
    new_n11893_, new_n11894_, new_n11895_, new_n11896_, new_n11897_,
    new_n11898_, new_n11899_, new_n11900_, new_n11901_, new_n11902_,
    new_n11903_, new_n11904_, new_n11905_, new_n11906_, new_n11907_,
    new_n11908_, new_n11909_, new_n11910_, new_n11911_, new_n11912_,
    new_n11913_, new_n11914_, new_n11915_, new_n11916_, new_n11917_,
    new_n11918_, new_n11919_, new_n11920_, new_n11921_, new_n11922_,
    new_n11923_, new_n11924_, new_n11925_, new_n11926_, new_n11927_,
    new_n11928_, new_n11929_, new_n11930_, new_n11931_, new_n11932_,
    new_n11933_, new_n11934_, new_n11935_, new_n11936_, new_n11937_,
    new_n11938_, new_n11939_, new_n11940_, new_n11941_, new_n11942_,
    new_n11943_, new_n11944_, new_n11945_, new_n11946_, new_n11947_,
    new_n11948_, new_n11949_, new_n11950_, new_n11951_, new_n11952_,
    new_n11953_, new_n11954_, new_n11955_, new_n11956_, new_n11957_,
    new_n11958_, new_n11959_, new_n11960_, new_n11961_, new_n11962_,
    new_n11963_, new_n11964_, new_n11965_, new_n11967_, new_n11968_,
    new_n11969_, new_n11970_, new_n11971_, new_n11972_, new_n11973_,
    new_n11974_, new_n11975_, new_n11976_, new_n11977_, new_n11978_,
    new_n11979_, new_n11980_, new_n11981_, new_n11982_, new_n11983_,
    new_n11984_, new_n11985_, new_n11986_, new_n11987_, new_n11988_,
    new_n11989_, new_n11990_, new_n11991_, new_n11992_, new_n11993_,
    new_n11994_, new_n11995_, new_n11996_, new_n11997_, new_n11998_,
    new_n11999_, new_n12000_, new_n12001_, new_n12002_, new_n12003_,
    new_n12004_, new_n12005_, new_n12006_, new_n12007_, new_n12008_,
    new_n12009_, new_n12010_, new_n12011_, new_n12012_, new_n12013_,
    new_n12014_, new_n12015_, new_n12016_, new_n12017_, new_n12018_,
    new_n12019_, new_n12020_, new_n12021_, new_n12022_, new_n12023_,
    new_n12024_, new_n12025_, new_n12026_, new_n12027_, new_n12028_,
    new_n12029_, new_n12030_, new_n12031_, new_n12032_, new_n12033_,
    new_n12034_, new_n12035_, new_n12036_, new_n12037_, new_n12038_,
    new_n12039_, new_n12040_, new_n12041_, new_n12042_, new_n12043_,
    new_n12044_, new_n12045_, new_n12046_, new_n12047_, new_n12048_,
    new_n12049_, new_n12050_, new_n12051_, new_n12052_, new_n12053_,
    new_n12054_, new_n12055_, new_n12056_, new_n12057_, new_n12058_,
    new_n12059_, new_n12060_, new_n12061_, new_n12062_, new_n12063_,
    new_n12064_, new_n12065_, new_n12066_, new_n12067_, new_n12068_,
    new_n12069_, new_n12070_, new_n12071_, new_n12072_, new_n12073_,
    new_n12074_, new_n12075_, new_n12076_, new_n12077_, new_n12078_,
    new_n12079_, new_n12080_, new_n12081_, new_n12082_, new_n12083_,
    new_n12084_, new_n12085_, new_n12086_, new_n12087_, new_n12088_,
    new_n12089_, new_n12090_, new_n12091_, new_n12092_, new_n12093_,
    new_n12094_, new_n12095_, new_n12096_, new_n12097_, new_n12098_,
    new_n12099_, new_n12100_, new_n12101_, new_n12102_, new_n12103_,
    new_n12104_, new_n12105_, new_n12106_, new_n12107_, new_n12108_,
    new_n12109_, new_n12110_, new_n12111_, new_n12112_, new_n12113_,
    new_n12114_, new_n12115_, new_n12116_, new_n12117_, new_n12118_,
    new_n12119_, new_n12120_, new_n12121_, new_n12122_, new_n12123_,
    new_n12124_, new_n12125_, new_n12126_, new_n12127_, new_n12128_,
    new_n12129_, new_n12130_, new_n12131_, new_n12132_, new_n12133_,
    new_n12134_, new_n12135_, new_n12136_, new_n12137_, new_n12138_,
    new_n12139_, new_n12140_, new_n12141_, new_n12142_, new_n12143_,
    new_n12144_, new_n12145_, new_n12146_, new_n12147_, new_n12148_,
    new_n12149_, new_n12150_, new_n12151_, new_n12152_, new_n12153_,
    new_n12154_, new_n12155_, new_n12156_, new_n12157_, new_n12158_,
    new_n12159_, new_n12160_, new_n12161_, new_n12162_, new_n12163_,
    new_n12164_, new_n12165_, new_n12166_, new_n12167_, new_n12168_,
    new_n12169_, new_n12170_, new_n12171_, new_n12172_, new_n12173_,
    new_n12174_, new_n12175_, new_n12176_, new_n12177_, new_n12178_,
    new_n12179_, new_n12180_, new_n12181_, new_n12182_, new_n12183_,
    new_n12184_, new_n12185_, new_n12186_, new_n12187_, new_n12188_,
    new_n12189_, new_n12190_, new_n12191_, new_n12192_, new_n12193_,
    new_n12194_, new_n12195_, new_n12196_, new_n12197_, new_n12198_,
    new_n12199_, new_n12200_, new_n12201_, new_n12202_, new_n12203_,
    new_n12204_, new_n12205_, new_n12206_, new_n12207_, new_n12208_,
    new_n12209_, new_n12210_, new_n12211_, new_n12212_, new_n12213_,
    new_n12214_, new_n12215_, new_n12216_, new_n12217_, new_n12218_,
    new_n12219_, new_n12220_, new_n12221_, new_n12222_, new_n12223_,
    new_n12224_, new_n12225_, new_n12226_, new_n12227_, new_n12228_,
    new_n12229_, new_n12230_, new_n12231_, new_n12232_, new_n12233_,
    new_n12234_, new_n12235_, new_n12236_, new_n12237_, new_n12238_,
    new_n12239_, new_n12240_, new_n12241_, new_n12242_, new_n12243_,
    new_n12244_, new_n12245_, new_n12246_, new_n12247_, new_n12248_,
    new_n12249_, new_n12250_, new_n12251_, new_n12252_, new_n12253_,
    new_n12254_, new_n12255_, new_n12256_, new_n12257_, new_n12258_,
    new_n12259_, new_n12260_, new_n12261_, new_n12262_, new_n12263_,
    new_n12264_, new_n12265_, new_n12266_, new_n12267_, new_n12268_,
    new_n12269_, new_n12270_, new_n12271_, new_n12272_, new_n12273_,
    new_n12274_, new_n12275_, new_n12276_, new_n12277_, new_n12278_,
    new_n12279_, new_n12280_, new_n12281_, new_n12282_, new_n12283_,
    new_n12284_, new_n12285_, new_n12286_, new_n12287_, new_n12288_,
    new_n12289_, new_n12290_, new_n12291_, new_n12292_, new_n12293_,
    new_n12294_, new_n12295_, new_n12296_, new_n12297_, new_n12298_,
    new_n12299_, new_n12300_, new_n12301_, new_n12302_, new_n12303_,
    new_n12304_, new_n12305_, new_n12306_, new_n12307_, new_n12308_,
    new_n12309_, new_n12310_, new_n12311_, new_n12312_, new_n12313_,
    new_n12314_, new_n12315_, new_n12316_, new_n12317_, new_n12318_,
    new_n12319_, new_n12320_, new_n12321_, new_n12322_, new_n12323_,
    new_n12324_, new_n12325_, new_n12326_, new_n12327_, new_n12328_,
    new_n12329_, new_n12330_, new_n12331_, new_n12332_, new_n12333_,
    new_n12334_, new_n12335_, new_n12336_, new_n12337_, new_n12338_,
    new_n12339_, new_n12340_, new_n12341_, new_n12342_, new_n12343_,
    new_n12344_, new_n12345_, new_n12346_, new_n12347_, new_n12348_,
    new_n12349_, new_n12350_, new_n12351_, new_n12352_, new_n12353_,
    new_n12354_, new_n12355_, new_n12356_, new_n12357_, new_n12358_,
    new_n12359_, new_n12360_, new_n12361_, new_n12362_, new_n12363_,
    new_n12364_, new_n12365_, new_n12366_, new_n12367_, new_n12368_,
    new_n12369_, new_n12370_, new_n12371_, new_n12372_, new_n12373_,
    new_n12374_, new_n12375_, new_n12376_, new_n12377_, new_n12378_,
    new_n12379_, new_n12380_, new_n12381_, new_n12382_, new_n12383_,
    new_n12384_, new_n12385_, new_n12386_, new_n12387_, new_n12388_,
    new_n12389_, new_n12390_, new_n12391_, new_n12392_, new_n12393_,
    new_n12394_, new_n12395_, new_n12396_, new_n12397_, new_n12398_,
    new_n12399_, new_n12400_, new_n12401_, new_n12402_, new_n12403_,
    new_n12404_, new_n12405_, new_n12406_, new_n12407_, new_n12408_,
    new_n12409_, new_n12410_, new_n12411_, new_n12412_, new_n12413_,
    new_n12414_, new_n12415_, new_n12416_, new_n12417_, new_n12418_,
    new_n12419_, new_n12420_, new_n12421_, new_n12422_, new_n12423_,
    new_n12424_, new_n12425_, new_n12426_, new_n12427_, new_n12428_,
    new_n12429_, new_n12430_, new_n12431_, new_n12432_, new_n12433_,
    new_n12434_, new_n12435_, new_n12436_, new_n12437_, new_n12438_,
    new_n12439_, new_n12440_, new_n12441_, new_n12442_, new_n12443_,
    new_n12444_, new_n12445_, new_n12446_, new_n12447_, new_n12448_,
    new_n12449_, new_n12450_, new_n12451_, new_n12452_, new_n12453_,
    new_n12454_, new_n12455_, new_n12456_, new_n12457_, new_n12459_,
    new_n12460_, new_n12461_, new_n12462_, new_n12463_, new_n12464_,
    new_n12465_, new_n12466_, new_n12467_, new_n12468_, new_n12469_,
    new_n12470_, new_n12471_, new_n12472_, new_n12473_, new_n12474_,
    new_n12475_, new_n12476_, new_n12477_, new_n12478_, new_n12479_,
    new_n12480_, new_n12481_, new_n12482_, new_n12483_, new_n12484_,
    new_n12485_, new_n12486_, new_n12487_, new_n12488_, new_n12489_,
    new_n12490_, new_n12491_, new_n12492_, new_n12493_, new_n12494_,
    new_n12495_, new_n12496_, new_n12497_, new_n12498_, new_n12499_,
    new_n12500_, new_n12501_, new_n12502_, new_n12503_, new_n12504_,
    new_n12505_, new_n12506_, new_n12507_, new_n12508_, new_n12509_,
    new_n12510_, new_n12511_, new_n12512_, new_n12513_, new_n12514_,
    new_n12515_, new_n12516_, new_n12517_, new_n12518_, new_n12519_,
    new_n12520_, new_n12521_, new_n12522_, new_n12523_, new_n12524_,
    new_n12525_, new_n12526_, new_n12527_, new_n12528_, new_n12529_,
    new_n12530_, new_n12531_, new_n12532_, new_n12533_, new_n12534_,
    new_n12535_, new_n12536_, new_n12537_, new_n12538_, new_n12539_,
    new_n12540_, new_n12541_, new_n12542_, new_n12543_, new_n12544_,
    new_n12545_, new_n12546_, new_n12547_, new_n12548_, new_n12549_,
    new_n12550_, new_n12551_, new_n12552_, new_n12553_, new_n12554_,
    new_n12555_, new_n12556_, new_n12557_, new_n12558_, new_n12559_,
    new_n12560_, new_n12561_, new_n12562_, new_n12563_, new_n12564_,
    new_n12565_, new_n12566_, new_n12567_, new_n12568_, new_n12569_,
    new_n12570_, new_n12571_, new_n12572_, new_n12573_, new_n12574_,
    new_n12575_, new_n12576_, new_n12577_, new_n12578_, new_n12579_,
    new_n12580_, new_n12581_, new_n12582_, new_n12583_, new_n12584_,
    new_n12585_, new_n12586_, new_n12587_, new_n12588_, new_n12589_,
    new_n12590_, new_n12591_, new_n12592_, new_n12593_, new_n12594_,
    new_n12595_, new_n12596_, new_n12597_, new_n12598_, new_n12599_,
    new_n12600_, new_n12601_, new_n12602_, new_n12603_, new_n12604_,
    new_n12605_, new_n12606_, new_n12607_, new_n12608_, new_n12609_,
    new_n12610_, new_n12611_, new_n12612_, new_n12613_, new_n12614_,
    new_n12615_, new_n12616_, new_n12617_, new_n12618_, new_n12619_,
    new_n12620_, new_n12621_, new_n12622_, new_n12623_, new_n12624_,
    new_n12625_, new_n12626_, new_n12627_, new_n12628_, new_n12629_,
    new_n12630_, new_n12631_, new_n12632_, new_n12633_, new_n12634_,
    new_n12635_, new_n12636_, new_n12637_, new_n12638_, new_n12639_,
    new_n12640_, new_n12641_, new_n12642_, new_n12643_, new_n12644_,
    new_n12645_, new_n12646_, new_n12647_, new_n12648_, new_n12649_,
    new_n12650_, new_n12651_, new_n12652_, new_n12653_, new_n12654_,
    new_n12655_, new_n12656_, new_n12657_, new_n12658_, new_n12659_,
    new_n12660_, new_n12661_, new_n12662_, new_n12663_, new_n12664_,
    new_n12665_, new_n12666_, new_n12667_, new_n12668_, new_n12669_,
    new_n12670_, new_n12671_, new_n12672_, new_n12673_, new_n12674_,
    new_n12675_, new_n12676_, new_n12677_, new_n12678_, new_n12679_,
    new_n12680_, new_n12681_, new_n12682_, new_n12683_, new_n12684_,
    new_n12685_, new_n12686_, new_n12687_, new_n12688_, new_n12689_,
    new_n12690_, new_n12691_, new_n12692_, new_n12693_, new_n12694_,
    new_n12695_, new_n12696_, new_n12697_, new_n12698_, new_n12699_,
    new_n12700_, new_n12701_, new_n12702_, new_n12703_, new_n12704_,
    new_n12705_, new_n12706_, new_n12707_, new_n12708_, new_n12709_,
    new_n12710_, new_n12711_, new_n12712_, new_n12713_, new_n12714_,
    new_n12715_, new_n12716_, new_n12717_, new_n12718_, new_n12719_,
    new_n12720_, new_n12721_, new_n12722_, new_n12723_, new_n12724_,
    new_n12725_, new_n12726_, new_n12727_, new_n12728_, new_n12729_,
    new_n12730_, new_n12731_, new_n12732_, new_n12733_, new_n12734_,
    new_n12735_, new_n12736_, new_n12737_, new_n12738_, new_n12739_,
    new_n12740_, new_n12741_, new_n12742_, new_n12743_, new_n12744_,
    new_n12745_, new_n12746_, new_n12747_, new_n12748_, new_n12749_,
    new_n12750_, new_n12751_, new_n12752_, new_n12753_, new_n12754_,
    new_n12755_, new_n12756_, new_n12757_, new_n12758_, new_n12759_,
    new_n12760_, new_n12761_, new_n12762_, new_n12763_, new_n12764_,
    new_n12765_, new_n12766_, new_n12767_, new_n12768_, new_n12769_,
    new_n12770_, new_n12771_, new_n12772_, new_n12773_, new_n12774_,
    new_n12775_, new_n12776_, new_n12777_, new_n12778_, new_n12779_,
    new_n12780_, new_n12781_, new_n12782_, new_n12783_, new_n12784_,
    new_n12785_, new_n12786_, new_n12787_, new_n12788_, new_n12789_,
    new_n12790_, new_n12791_, new_n12792_, new_n12793_, new_n12794_,
    new_n12795_, new_n12796_, new_n12797_, new_n12798_, new_n12799_,
    new_n12800_, new_n12801_, new_n12802_, new_n12803_, new_n12804_,
    new_n12805_, new_n12806_, new_n12807_, new_n12808_, new_n12809_,
    new_n12810_, new_n12811_, new_n12812_, new_n12813_, new_n12814_,
    new_n12815_, new_n12816_, new_n12817_, new_n12818_, new_n12819_,
    new_n12820_, new_n12821_, new_n12822_, new_n12823_, new_n12824_,
    new_n12825_, new_n12826_, new_n12827_, new_n12828_, new_n12829_,
    new_n12830_, new_n12831_, new_n12832_, new_n12833_, new_n12834_,
    new_n12835_, new_n12836_, new_n12837_, new_n12838_, new_n12839_,
    new_n12840_, new_n12841_, new_n12842_, new_n12843_, new_n12844_,
    new_n12845_, new_n12846_, new_n12847_, new_n12848_, new_n12849_,
    new_n12850_, new_n12851_, new_n12852_, new_n12853_, new_n12854_,
    new_n12855_, new_n12856_, new_n12857_, new_n12858_, new_n12859_,
    new_n12860_, new_n12861_, new_n12862_, new_n12863_, new_n12864_,
    new_n12865_, new_n12866_, new_n12867_, new_n12868_, new_n12869_,
    new_n12870_, new_n12871_, new_n12872_, new_n12873_, new_n12874_,
    new_n12875_, new_n12876_, new_n12877_, new_n12878_, new_n12879_,
    new_n12880_, new_n12881_, new_n12882_, new_n12883_, new_n12884_,
    new_n12885_, new_n12886_, new_n12887_, new_n12888_, new_n12889_,
    new_n12890_, new_n12891_, new_n12892_, new_n12893_, new_n12894_,
    new_n12895_, new_n12896_, new_n12897_, new_n12898_, new_n12899_,
    new_n12900_, new_n12901_, new_n12902_, new_n12903_, new_n12904_,
    new_n12905_, new_n12906_, new_n12907_, new_n12908_, new_n12909_,
    new_n12910_, new_n12911_, new_n12912_, new_n12913_, new_n12914_,
    new_n12915_, new_n12916_, new_n12917_, new_n12918_, new_n12919_,
    new_n12920_, new_n12921_, new_n12922_, new_n12923_, new_n12924_,
    new_n12925_, new_n12926_, new_n12927_, new_n12928_, new_n12929_,
    new_n12930_, new_n12931_, new_n12932_, new_n12933_, new_n12934_,
    new_n12935_, new_n12936_, new_n12937_, new_n12938_, new_n12939_,
    new_n12940_, new_n12941_, new_n12942_, new_n12943_, new_n12944_,
    new_n12945_, new_n12946_, new_n12947_, new_n12948_, new_n12949_,
    new_n12950_, new_n12951_, new_n12952_, new_n12953_, new_n12954_,
    new_n12955_, new_n12956_, new_n12957_, new_n12958_, new_n12959_,
    new_n12960_, new_n12961_, new_n12962_, new_n12963_, new_n12964_,
    new_n12965_, new_n12966_, new_n12967_, new_n12968_, new_n12969_,
    new_n12970_, new_n12971_, new_n12972_, new_n12973_, new_n12974_,
    new_n12975_, new_n12976_, new_n12977_, new_n12978_, new_n12979_,
    new_n12980_, new_n12981_, new_n12982_, new_n12983_, new_n12984_,
    new_n12985_, new_n12986_, new_n12987_, new_n12988_, new_n12989_,
    new_n12990_, new_n12991_, new_n12992_, new_n12993_, new_n12994_,
    new_n12995_, new_n12996_, new_n12997_, new_n12998_, new_n12999_,
    new_n13000_, new_n13002_, new_n13003_, new_n13004_, new_n13005_,
    new_n13006_, new_n13007_, new_n13008_, new_n13009_, new_n13010_,
    new_n13011_, new_n13012_, new_n13013_, new_n13014_, new_n13015_,
    new_n13016_, new_n13017_, new_n13018_, new_n13019_, new_n13020_,
    new_n13021_, new_n13022_, new_n13023_, new_n13024_, new_n13025_,
    new_n13026_, new_n13027_, new_n13028_, new_n13029_, new_n13030_,
    new_n13031_, new_n13032_, new_n13033_, new_n13034_, new_n13035_,
    new_n13036_, new_n13037_, new_n13038_, new_n13039_, new_n13040_,
    new_n13041_, new_n13042_, new_n13043_, new_n13044_, new_n13045_,
    new_n13046_, new_n13047_, new_n13048_, new_n13049_, new_n13050_,
    new_n13051_, new_n13052_, new_n13053_, new_n13054_, new_n13055_,
    new_n13056_, new_n13057_, new_n13058_, new_n13059_, new_n13060_,
    new_n13061_, new_n13062_, new_n13063_, new_n13064_, new_n13065_,
    new_n13066_, new_n13067_, new_n13068_, new_n13069_, new_n13070_,
    new_n13071_, new_n13072_, new_n13073_, new_n13074_, new_n13075_,
    new_n13076_, new_n13077_, new_n13078_, new_n13079_, new_n13080_,
    new_n13081_, new_n13082_, new_n13083_, new_n13084_, new_n13085_,
    new_n13086_, new_n13087_, new_n13088_, new_n13089_, new_n13090_,
    new_n13091_, new_n13092_, new_n13093_, new_n13094_, new_n13095_,
    new_n13096_, new_n13097_, new_n13098_, new_n13099_, new_n13100_,
    new_n13101_, new_n13102_, new_n13103_, new_n13104_, new_n13105_,
    new_n13106_, new_n13107_, new_n13108_, new_n13109_, new_n13110_,
    new_n13111_, new_n13112_, new_n13113_, new_n13114_, new_n13115_,
    new_n13116_, new_n13117_, new_n13118_, new_n13119_, new_n13120_,
    new_n13121_, new_n13122_, new_n13123_, new_n13124_, new_n13125_,
    new_n13126_, new_n13127_, new_n13128_, new_n13129_, new_n13130_,
    new_n13131_, new_n13132_, new_n13133_, new_n13134_, new_n13135_,
    new_n13136_, new_n13137_, new_n13138_, new_n13139_, new_n13140_,
    new_n13141_, new_n13142_, new_n13143_, new_n13144_, new_n13145_,
    new_n13146_, new_n13147_, new_n13148_, new_n13149_, new_n13150_,
    new_n13151_, new_n13152_, new_n13153_, new_n13154_, new_n13155_,
    new_n13156_, new_n13157_, new_n13158_, new_n13159_, new_n13160_,
    new_n13161_, new_n13162_, new_n13163_, new_n13164_, new_n13165_,
    new_n13166_, new_n13167_, new_n13168_, new_n13169_, new_n13170_,
    new_n13171_, new_n13172_, new_n13173_, new_n13174_, new_n13175_,
    new_n13176_, new_n13177_, new_n13178_, new_n13179_, new_n13180_,
    new_n13181_, new_n13182_, new_n13183_, new_n13184_, new_n13185_,
    new_n13186_, new_n13187_, new_n13188_, new_n13189_, new_n13190_,
    new_n13191_, new_n13192_, new_n13193_, new_n13194_, new_n13195_,
    new_n13196_, new_n13197_, new_n13198_, new_n13199_, new_n13200_,
    new_n13201_, new_n13202_, new_n13203_, new_n13204_, new_n13205_,
    new_n13206_, new_n13207_, new_n13208_, new_n13209_, new_n13210_,
    new_n13211_, new_n13212_, new_n13213_, new_n13214_, new_n13215_,
    new_n13216_, new_n13217_, new_n13218_, new_n13219_, new_n13220_,
    new_n13221_, new_n13222_, new_n13223_, new_n13224_, new_n13225_,
    new_n13226_, new_n13227_, new_n13228_, new_n13229_, new_n13230_,
    new_n13231_, new_n13232_, new_n13233_, new_n13234_, new_n13235_,
    new_n13236_, new_n13237_, new_n13238_, new_n13239_, new_n13240_,
    new_n13241_, new_n13242_, new_n13243_, new_n13244_, new_n13245_,
    new_n13246_, new_n13247_, new_n13248_, new_n13249_, new_n13250_,
    new_n13251_, new_n13252_, new_n13253_, new_n13254_, new_n13255_,
    new_n13256_, new_n13257_, new_n13258_, new_n13259_, new_n13260_,
    new_n13261_, new_n13262_, new_n13263_, new_n13264_, new_n13265_,
    new_n13266_, new_n13267_, new_n13268_, new_n13269_, new_n13270_,
    new_n13271_, new_n13272_, new_n13273_, new_n13274_, new_n13275_,
    new_n13276_, new_n13277_, new_n13278_, new_n13279_, new_n13280_,
    new_n13281_, new_n13282_, new_n13283_, new_n13284_, new_n13285_,
    new_n13286_, new_n13287_, new_n13288_, new_n13289_, new_n13290_,
    new_n13291_, new_n13292_, new_n13293_, new_n13294_, new_n13295_,
    new_n13296_, new_n13297_, new_n13298_, new_n13299_, new_n13300_,
    new_n13301_, new_n13302_, new_n13303_, new_n13304_, new_n13305_,
    new_n13306_, new_n13307_, new_n13308_, new_n13309_, new_n13310_,
    new_n13311_, new_n13312_, new_n13313_, new_n13314_, new_n13315_,
    new_n13316_, new_n13317_, new_n13318_, new_n13319_, new_n13320_,
    new_n13321_, new_n13322_, new_n13323_, new_n13324_, new_n13325_,
    new_n13326_, new_n13327_, new_n13328_, new_n13329_, new_n13330_,
    new_n13331_, new_n13332_, new_n13333_, new_n13334_, new_n13335_,
    new_n13336_, new_n13337_, new_n13338_, new_n13339_, new_n13340_,
    new_n13341_, new_n13342_, new_n13343_, new_n13344_, new_n13345_,
    new_n13346_, new_n13347_, new_n13348_, new_n13349_, new_n13350_,
    new_n13351_, new_n13352_, new_n13353_, new_n13354_, new_n13355_,
    new_n13356_, new_n13357_, new_n13358_, new_n13359_, new_n13360_,
    new_n13361_, new_n13362_, new_n13363_, new_n13364_, new_n13365_,
    new_n13366_, new_n13367_, new_n13368_, new_n13369_, new_n13370_,
    new_n13371_, new_n13372_, new_n13373_, new_n13374_, new_n13375_,
    new_n13376_, new_n13377_, new_n13378_, new_n13379_, new_n13380_,
    new_n13381_, new_n13382_, new_n13383_, new_n13384_, new_n13385_,
    new_n13386_, new_n13387_, new_n13388_, new_n13389_, new_n13390_,
    new_n13391_, new_n13392_, new_n13393_, new_n13394_, new_n13395_,
    new_n13396_, new_n13397_, new_n13398_, new_n13399_, new_n13400_,
    new_n13401_, new_n13402_, new_n13403_, new_n13404_, new_n13405_,
    new_n13406_, new_n13407_, new_n13408_, new_n13409_, new_n13410_,
    new_n13411_, new_n13412_, new_n13413_, new_n13414_, new_n13415_,
    new_n13416_, new_n13417_, new_n13418_, new_n13419_, new_n13420_,
    new_n13421_, new_n13422_, new_n13423_, new_n13424_, new_n13425_,
    new_n13426_, new_n13427_, new_n13428_, new_n13429_, new_n13430_,
    new_n13431_, new_n13432_, new_n13433_, new_n13434_, new_n13435_,
    new_n13436_, new_n13437_, new_n13438_, new_n13439_, new_n13440_,
    new_n13441_, new_n13442_, new_n13443_, new_n13444_, new_n13445_,
    new_n13446_, new_n13447_, new_n13448_, new_n13449_, new_n13450_,
    new_n13451_, new_n13452_, new_n13453_, new_n13454_, new_n13455_,
    new_n13456_, new_n13457_, new_n13458_, new_n13459_, new_n13460_,
    new_n13461_, new_n13462_, new_n13463_, new_n13464_, new_n13465_,
    new_n13466_, new_n13467_, new_n13468_, new_n13469_, new_n13470_,
    new_n13471_, new_n13472_, new_n13473_, new_n13474_, new_n13475_,
    new_n13476_, new_n13477_, new_n13478_, new_n13479_, new_n13480_,
    new_n13481_, new_n13482_, new_n13483_, new_n13484_, new_n13485_,
    new_n13486_, new_n13487_, new_n13488_, new_n13489_, new_n13490_,
    new_n13491_, new_n13492_, new_n13493_, new_n13494_, new_n13495_,
    new_n13496_, new_n13497_, new_n13498_, new_n13499_, new_n13500_,
    new_n13501_, new_n13502_, new_n13503_, new_n13504_, new_n13505_,
    new_n13506_, new_n13507_, new_n13508_, new_n13509_, new_n13510_,
    new_n13511_, new_n13512_, new_n13513_, new_n13514_, new_n13515_,
    new_n13516_, new_n13517_, new_n13518_, new_n13519_, new_n13520_,
    new_n13521_, new_n13522_, new_n13523_, new_n13524_, new_n13525_,
    new_n13526_, new_n13527_, new_n13528_, new_n13529_, new_n13530_,
    new_n13531_, new_n13532_, new_n13533_, new_n13534_, new_n13535_,
    new_n13536_, new_n13537_, new_n13538_, new_n13539_, new_n13540_,
    new_n13541_, new_n13542_, new_n13543_, new_n13544_, new_n13545_,
    new_n13546_, new_n13547_, new_n13548_, new_n13549_, new_n13550_,
    new_n13551_, new_n13552_, new_n13553_, new_n13554_, new_n13555_,
    new_n13556_, new_n13557_, new_n13558_, new_n13559_, new_n13560_,
    new_n13561_, new_n13562_, new_n13563_, new_n13564_, new_n13565_,
    new_n13566_, new_n13567_, new_n13568_, new_n13569_, new_n13570_,
    new_n13571_, new_n13572_, new_n13573_, new_n13574_, new_n13575_,
    new_n13576_, new_n13577_, new_n13578_, new_n13579_, new_n13580_,
    new_n13581_, new_n13582_, new_n13583_, new_n13584_, new_n13585_,
    new_n13586_, new_n13587_, new_n13588_, new_n13589_, new_n13590_,
    new_n13591_, new_n13592_, new_n13593_, new_n13594_, new_n13595_,
    new_n13596_, new_n13597_, new_n13598_, new_n13599_, new_n13600_,
    new_n13601_, new_n13602_, new_n13603_, new_n13604_, new_n13605_,
    new_n13606_, new_n13607_, new_n13608_, new_n13609_, new_n13610_,
    new_n13611_, new_n13612_, new_n13613_, new_n13614_, new_n13615_,
    new_n13616_, new_n13617_, new_n13618_, new_n13619_, new_n13620_,
    new_n13621_, new_n13622_, new_n13623_, new_n13624_, new_n13625_,
    new_n13626_, new_n13627_, new_n13628_, new_n13629_, new_n13630_,
    new_n13631_, new_n13632_, new_n13633_, new_n13634_, new_n13635_,
    new_n13636_, new_n13637_, new_n13638_, new_n13639_, new_n13640_,
    new_n13641_, new_n13642_, new_n13643_, new_n13644_, new_n13645_,
    new_n13646_, new_n13647_, new_n13648_, new_n13649_, new_n13650_,
    new_n13651_, new_n13652_, new_n13653_, new_n13654_, new_n13656_,
    new_n13657_, new_n13658_, new_n13659_, new_n13660_, new_n13661_,
    new_n13662_, new_n13663_, new_n13664_, new_n13665_, new_n13666_,
    new_n13667_, new_n13668_, new_n13669_, new_n13670_, new_n13671_,
    new_n13672_, new_n13673_, new_n13674_, new_n13675_, new_n13676_,
    new_n13677_, new_n13678_, new_n13679_, new_n13680_, new_n13681_,
    new_n13682_, new_n13683_, new_n13684_, new_n13685_, new_n13686_,
    new_n13687_, new_n13688_, new_n13689_, new_n13690_, new_n13691_,
    new_n13692_, new_n13693_, new_n13694_, new_n13695_, new_n13696_,
    new_n13697_, new_n13698_, new_n13699_, new_n13700_, new_n13701_,
    new_n13702_, new_n13703_, new_n13704_, new_n13705_, new_n13706_,
    new_n13707_, new_n13708_, new_n13709_, new_n13710_, new_n13711_,
    new_n13712_, new_n13713_, new_n13714_, new_n13715_, new_n13716_,
    new_n13717_, new_n13718_, new_n13719_, new_n13720_, new_n13721_,
    new_n13722_, new_n13723_, new_n13724_, new_n13725_, new_n13726_,
    new_n13727_, new_n13728_, new_n13729_, new_n13730_, new_n13731_,
    new_n13732_, new_n13733_, new_n13734_, new_n13735_, new_n13736_,
    new_n13737_, new_n13738_, new_n13739_, new_n13740_, new_n13741_,
    new_n13742_, new_n13743_, new_n13744_, new_n13745_, new_n13746_,
    new_n13747_, new_n13748_, new_n13749_, new_n13750_, new_n13751_,
    new_n13752_, new_n13753_, new_n13754_, new_n13755_, new_n13756_,
    new_n13757_, new_n13758_, new_n13759_, new_n13760_, new_n13761_,
    new_n13762_, new_n13763_, new_n13764_, new_n13765_, new_n13766_,
    new_n13767_, new_n13768_, new_n13769_, new_n13770_, new_n13771_,
    new_n13772_, new_n13773_, new_n13774_, new_n13775_, new_n13776_,
    new_n13777_, new_n13778_, new_n13779_, new_n13780_, new_n13781_,
    new_n13782_, new_n13783_, new_n13784_, new_n13785_, new_n13786_,
    new_n13787_, new_n13788_, new_n13789_, new_n13790_, new_n13791_,
    new_n13792_, new_n13793_, new_n13794_, new_n13795_, new_n13796_,
    new_n13797_, new_n13798_, new_n13799_, new_n13800_, new_n13801_,
    new_n13802_, new_n13803_, new_n13804_, new_n13805_, new_n13806_,
    new_n13807_, new_n13808_, new_n13809_, new_n13810_, new_n13811_,
    new_n13812_, new_n13813_, new_n13814_, new_n13815_, new_n13816_,
    new_n13817_, new_n13818_, new_n13819_, new_n13820_, new_n13821_,
    new_n13822_, new_n13823_, new_n13824_, new_n13825_, new_n13826_,
    new_n13827_, new_n13828_, new_n13829_, new_n13830_, new_n13831_,
    new_n13832_, new_n13833_, new_n13834_, new_n13835_, new_n13836_,
    new_n13837_, new_n13838_, new_n13839_, new_n13840_, new_n13841_,
    new_n13842_, new_n13843_, new_n13844_, new_n13845_, new_n13846_,
    new_n13847_, new_n13848_, new_n13849_, new_n13850_, new_n13851_,
    new_n13852_, new_n13853_, new_n13854_, new_n13855_, new_n13856_,
    new_n13857_, new_n13858_, new_n13859_, new_n13860_, new_n13861_,
    new_n13862_, new_n13863_, new_n13864_, new_n13865_, new_n13866_,
    new_n13867_, new_n13868_, new_n13869_, new_n13870_, new_n13871_,
    new_n13872_, new_n13873_, new_n13874_, new_n13875_, new_n13876_,
    new_n13877_, new_n13878_, new_n13879_, new_n13880_, new_n13881_,
    new_n13882_, new_n13883_, new_n13884_, new_n13885_, new_n13886_,
    new_n13887_, new_n13888_, new_n13889_, new_n13890_, new_n13891_,
    new_n13892_, new_n13893_, new_n13894_, new_n13895_, new_n13896_,
    new_n13897_, new_n13898_, new_n13899_, new_n13900_, new_n13901_,
    new_n13902_, new_n13903_, new_n13904_, new_n13905_, new_n13906_,
    new_n13907_, new_n13908_, new_n13909_, new_n13910_, new_n13911_,
    new_n13912_, new_n13913_, new_n13914_, new_n13915_, new_n13916_,
    new_n13917_, new_n13918_, new_n13919_, new_n13920_, new_n13921_,
    new_n13922_, new_n13923_, new_n13924_, new_n13925_, new_n13926_,
    new_n13927_, new_n13928_, new_n13929_, new_n13930_, new_n13931_,
    new_n13932_, new_n13933_, new_n13934_, new_n13935_, new_n13936_,
    new_n13937_, new_n13938_, new_n13939_, new_n13940_, new_n13941_,
    new_n13942_, new_n13943_, new_n13944_, new_n13945_, new_n13946_,
    new_n13947_, new_n13948_, new_n13949_, new_n13950_, new_n13951_,
    new_n13952_, new_n13953_, new_n13954_, new_n13955_, new_n13956_,
    new_n13957_, new_n13958_, new_n13959_, new_n13960_, new_n13961_,
    new_n13962_, new_n13963_, new_n13964_, new_n13965_, new_n13966_,
    new_n13967_, new_n13968_, new_n13969_, new_n13970_, new_n13971_,
    new_n13972_, new_n13973_, new_n13974_, new_n13975_, new_n13976_,
    new_n13977_, new_n13978_, new_n13979_, new_n13980_, new_n13981_,
    new_n13982_, new_n13983_, new_n13984_, new_n13985_, new_n13986_,
    new_n13987_, new_n13988_, new_n13989_, new_n13990_, new_n13991_,
    new_n13992_, new_n13993_, new_n13994_, new_n13995_, new_n13996_,
    new_n13997_, new_n13998_, new_n13999_, new_n14000_, new_n14001_,
    new_n14002_, new_n14003_, new_n14004_, new_n14005_, new_n14006_,
    new_n14007_, new_n14008_, new_n14009_, new_n14010_, new_n14011_,
    new_n14012_, new_n14013_, new_n14014_, new_n14015_, new_n14016_,
    new_n14017_, new_n14018_, new_n14019_, new_n14020_, new_n14021_,
    new_n14022_, new_n14023_, new_n14024_, new_n14025_, new_n14026_,
    new_n14027_, new_n14028_, new_n14029_, new_n14030_, new_n14031_,
    new_n14032_, new_n14033_, new_n14034_, new_n14035_, new_n14036_,
    new_n14037_, new_n14038_, new_n14039_, new_n14040_, new_n14041_,
    new_n14042_, new_n14043_, new_n14044_, new_n14045_, new_n14046_,
    new_n14047_, new_n14048_, new_n14049_, new_n14050_, new_n14051_,
    new_n14052_, new_n14053_, new_n14054_, new_n14055_, new_n14056_,
    new_n14057_, new_n14058_, new_n14059_, new_n14060_, new_n14061_,
    new_n14062_, new_n14063_, new_n14064_, new_n14065_, new_n14066_,
    new_n14067_, new_n14068_, new_n14069_, new_n14070_, new_n14071_,
    new_n14072_, new_n14073_, new_n14074_, new_n14075_, new_n14076_,
    new_n14077_, new_n14078_, new_n14079_, new_n14080_, new_n14081_,
    new_n14082_, new_n14083_, new_n14084_, new_n14085_, new_n14086_,
    new_n14087_, new_n14088_, new_n14089_, new_n14090_, new_n14091_,
    new_n14092_, new_n14093_, new_n14094_, new_n14095_, new_n14096_,
    new_n14097_, new_n14098_, new_n14099_, new_n14100_, new_n14101_,
    new_n14102_, new_n14103_, new_n14104_, new_n14105_, new_n14106_,
    new_n14107_, new_n14108_, new_n14109_, new_n14110_, new_n14111_,
    new_n14112_, new_n14113_, new_n14114_, new_n14115_, new_n14116_,
    new_n14117_, new_n14118_, new_n14119_, new_n14120_, new_n14121_,
    new_n14122_, new_n14123_, new_n14124_, new_n14125_, new_n14126_,
    new_n14127_, new_n14128_, new_n14129_, new_n14130_, new_n14131_,
    new_n14132_, new_n14133_, new_n14134_, new_n14135_, new_n14136_,
    new_n14137_, new_n14138_, new_n14139_, new_n14140_, new_n14141_,
    new_n14142_, new_n14143_, new_n14144_, new_n14145_, new_n14146_,
    new_n14147_, new_n14148_, new_n14149_, new_n14150_, new_n14151_,
    new_n14152_, new_n14153_, new_n14154_, new_n14155_, new_n14156_,
    new_n14157_, new_n14158_, new_n14159_, new_n14160_, new_n14161_,
    new_n14162_, new_n14163_, new_n14164_, new_n14165_, new_n14166_,
    new_n14167_, new_n14168_, new_n14169_, new_n14170_, new_n14171_,
    new_n14172_, new_n14173_, new_n14174_, new_n14175_, new_n14176_,
    new_n14177_, new_n14178_, new_n14179_, new_n14180_, new_n14181_,
    new_n14182_, new_n14183_, new_n14184_, new_n14185_, new_n14186_,
    new_n14187_, new_n14188_, new_n14189_, new_n14190_, new_n14191_,
    new_n14193_, new_n14194_, new_n14195_, new_n14196_, new_n14197_,
    new_n14198_, new_n14199_, new_n14200_, new_n14201_, new_n14202_,
    new_n14203_, new_n14204_, new_n14205_, new_n14206_, new_n14207_,
    new_n14208_, new_n14209_, new_n14210_, new_n14211_, new_n14212_,
    new_n14213_, new_n14214_, new_n14215_, new_n14216_, new_n14217_,
    new_n14218_, new_n14219_, new_n14220_, new_n14221_, new_n14222_,
    new_n14223_, new_n14224_, new_n14225_, new_n14226_, new_n14227_,
    new_n14228_, new_n14229_, new_n14230_, new_n14231_, new_n14232_,
    new_n14233_, new_n14234_, new_n14235_, new_n14236_, new_n14237_,
    new_n14238_, new_n14239_, new_n14240_, new_n14241_, new_n14242_,
    new_n14243_, new_n14244_, new_n14245_, new_n14246_, new_n14247_,
    new_n14248_, new_n14249_, new_n14250_, new_n14251_, new_n14252_,
    new_n14253_, new_n14254_, new_n14255_, new_n14256_, new_n14257_,
    new_n14258_, new_n14259_, new_n14260_, new_n14261_, new_n14262_,
    new_n14263_, new_n14264_, new_n14265_, new_n14266_, new_n14267_,
    new_n14268_, new_n14269_, new_n14270_, new_n14271_, new_n14272_,
    new_n14273_, new_n14274_, new_n14275_, new_n14276_, new_n14277_,
    new_n14278_, new_n14279_, new_n14280_, new_n14281_, new_n14282_,
    new_n14283_, new_n14284_, new_n14285_, new_n14286_, new_n14287_,
    new_n14288_, new_n14289_, new_n14290_, new_n14291_, new_n14292_,
    new_n14293_, new_n14294_, new_n14295_, new_n14296_, new_n14297_,
    new_n14298_, new_n14299_, new_n14300_, new_n14301_, new_n14302_,
    new_n14303_, new_n14304_, new_n14305_, new_n14306_, new_n14307_,
    new_n14308_, new_n14309_, new_n14310_, new_n14311_, new_n14312_,
    new_n14313_, new_n14314_, new_n14315_, new_n14316_, new_n14317_,
    new_n14318_, new_n14319_, new_n14320_, new_n14321_, new_n14322_,
    new_n14323_, new_n14324_, new_n14325_, new_n14326_, new_n14327_,
    new_n14328_, new_n14329_, new_n14330_, new_n14331_, new_n14332_,
    new_n14333_, new_n14334_, new_n14335_, new_n14336_, new_n14337_,
    new_n14338_, new_n14339_, new_n14340_, new_n14341_, new_n14342_,
    new_n14343_, new_n14344_, new_n14345_, new_n14346_, new_n14347_,
    new_n14348_, new_n14349_, new_n14350_, new_n14351_, new_n14352_,
    new_n14353_, new_n14354_, new_n14355_, new_n14356_, new_n14357_,
    new_n14358_, new_n14359_, new_n14360_, new_n14361_, new_n14362_,
    new_n14363_, new_n14364_, new_n14365_, new_n14366_, new_n14367_,
    new_n14368_, new_n14369_, new_n14370_, new_n14371_, new_n14372_,
    new_n14373_, new_n14374_, new_n14375_, new_n14376_, new_n14377_,
    new_n14378_, new_n14379_, new_n14380_, new_n14381_, new_n14382_,
    new_n14383_, new_n14384_, new_n14385_, new_n14386_, new_n14387_,
    new_n14388_, new_n14389_, new_n14390_, new_n14391_, new_n14392_,
    new_n14393_, new_n14394_, new_n14395_, new_n14396_, new_n14397_,
    new_n14398_, new_n14399_, new_n14400_, new_n14401_, new_n14402_,
    new_n14403_, new_n14404_, new_n14405_, new_n14406_, new_n14407_,
    new_n14408_, new_n14409_, new_n14410_, new_n14411_, new_n14412_,
    new_n14413_, new_n14414_, new_n14415_, new_n14416_, new_n14417_,
    new_n14418_, new_n14419_, new_n14420_, new_n14421_, new_n14422_,
    new_n14423_, new_n14424_, new_n14425_, new_n14426_, new_n14427_,
    new_n14428_, new_n14429_, new_n14430_, new_n14431_, new_n14432_,
    new_n14433_, new_n14434_, new_n14435_, new_n14436_, new_n14437_,
    new_n14438_, new_n14439_, new_n14440_, new_n14441_, new_n14442_,
    new_n14443_, new_n14444_, new_n14445_, new_n14446_, new_n14447_,
    new_n14448_, new_n14449_, new_n14450_, new_n14451_, new_n14452_,
    new_n14453_, new_n14454_, new_n14455_, new_n14456_, new_n14457_,
    new_n14458_, new_n14459_, new_n14460_, new_n14461_, new_n14462_,
    new_n14463_, new_n14464_, new_n14465_, new_n14466_, new_n14467_,
    new_n14468_, new_n14469_, new_n14470_, new_n14471_, new_n14472_,
    new_n14473_, new_n14474_, new_n14475_, new_n14476_, new_n14477_,
    new_n14478_, new_n14479_, new_n14480_, new_n14481_, new_n14482_,
    new_n14483_, new_n14484_, new_n14485_, new_n14486_, new_n14487_,
    new_n14488_, new_n14489_, new_n14490_, new_n14491_, new_n14492_,
    new_n14493_, new_n14494_, new_n14495_, new_n14496_, new_n14497_,
    new_n14498_, new_n14499_, new_n14500_, new_n14501_, new_n14502_,
    new_n14503_, new_n14504_, new_n14505_, new_n14506_, new_n14507_,
    new_n14508_, new_n14509_, new_n14510_, new_n14511_, new_n14512_,
    new_n14513_, new_n14514_, new_n14515_, new_n14516_, new_n14517_,
    new_n14518_, new_n14519_, new_n14520_, new_n14521_, new_n14522_,
    new_n14523_, new_n14524_, new_n14525_, new_n14526_, new_n14527_,
    new_n14528_, new_n14529_, new_n14530_, new_n14531_, new_n14532_,
    new_n14533_, new_n14534_, new_n14535_, new_n14536_, new_n14537_,
    new_n14538_, new_n14539_, new_n14540_, new_n14541_, new_n14542_,
    new_n14543_, new_n14544_, new_n14545_, new_n14546_, new_n14547_,
    new_n14548_, new_n14549_, new_n14550_, new_n14551_, new_n14552_,
    new_n14553_, new_n14554_, new_n14555_, new_n14556_, new_n14557_,
    new_n14558_, new_n14559_, new_n14560_, new_n14561_, new_n14562_,
    new_n14563_, new_n14564_, new_n14565_, new_n14566_, new_n14567_,
    new_n14568_, new_n14569_, new_n14570_, new_n14571_, new_n14572_,
    new_n14573_, new_n14574_, new_n14575_, new_n14576_, new_n14577_,
    new_n14578_, new_n14579_, new_n14580_, new_n14581_, new_n14582_,
    new_n14583_, new_n14584_, new_n14585_, new_n14586_, new_n14587_,
    new_n14588_, new_n14589_, new_n14590_, new_n14591_, new_n14592_,
    new_n14593_, new_n14594_, new_n14595_, new_n14596_, new_n14597_,
    new_n14598_, new_n14599_, new_n14600_, new_n14601_, new_n14602_,
    new_n14603_, new_n14604_, new_n14605_, new_n14606_, new_n14607_,
    new_n14608_, new_n14609_, new_n14610_, new_n14611_, new_n14612_,
    new_n14613_, new_n14614_, new_n14615_, new_n14616_, new_n14617_,
    new_n14618_, new_n14619_, new_n14620_, new_n14621_, new_n14622_,
    new_n14623_, new_n14624_, new_n14625_, new_n14626_, new_n14627_,
    new_n14628_, new_n14629_, new_n14630_, new_n14631_, new_n14632_,
    new_n14633_, new_n14634_, new_n14635_, new_n14636_, new_n14637_,
    new_n14638_, new_n14639_, new_n14640_, new_n14641_, new_n14642_,
    new_n14643_, new_n14644_, new_n14645_, new_n14646_, new_n14647_,
    new_n14648_, new_n14649_, new_n14650_, new_n14651_, new_n14652_,
    new_n14653_, new_n14654_, new_n14655_, new_n14656_, new_n14657_,
    new_n14658_, new_n14659_, new_n14660_, new_n14661_, new_n14662_,
    new_n14663_, new_n14664_, new_n14665_, new_n14666_, new_n14667_,
    new_n14668_, new_n14669_, new_n14670_, new_n14671_, new_n14672_,
    new_n14673_, new_n14674_, new_n14675_, new_n14676_, new_n14677_,
    new_n14678_, new_n14679_, new_n14680_, new_n14681_, new_n14682_,
    new_n14683_, new_n14684_, new_n14685_, new_n14686_, new_n14687_,
    new_n14688_, new_n14689_, new_n14690_, new_n14691_, new_n14692_,
    new_n14693_, new_n14694_, new_n14695_, new_n14696_, new_n14697_,
    new_n14698_, new_n14699_, new_n14700_, new_n14701_, new_n14702_,
    new_n14703_, new_n14704_, new_n14705_, new_n14706_, new_n14707_,
    new_n14708_, new_n14709_, new_n14710_, new_n14711_, new_n14712_,
    new_n14713_, new_n14714_, new_n14715_, new_n14716_, new_n14717_,
    new_n14718_, new_n14719_, new_n14720_, new_n14721_, new_n14722_,
    new_n14723_, new_n14724_, new_n14725_, new_n14726_, new_n14727_,
    new_n14728_, new_n14729_, new_n14730_, new_n14731_, new_n14732_,
    new_n14733_, new_n14734_, new_n14735_, new_n14736_, new_n14737_,
    new_n14738_, new_n14739_, new_n14740_, new_n14741_, new_n14742_,
    new_n14743_, new_n14744_, new_n14745_, new_n14746_, new_n14747_,
    new_n14748_, new_n14749_, new_n14750_, new_n14751_, new_n14752_,
    new_n14753_, new_n14754_, new_n14756_, new_n14757_, new_n14758_,
    new_n14759_, new_n14760_, new_n14761_, new_n14762_, new_n14763_,
    new_n14764_, new_n14765_, new_n14766_, new_n14767_, new_n14768_,
    new_n14769_, new_n14770_, new_n14771_, new_n14772_, new_n14773_,
    new_n14774_, new_n14775_, new_n14776_, new_n14777_, new_n14778_,
    new_n14779_, new_n14780_, new_n14781_, new_n14782_, new_n14783_,
    new_n14784_, new_n14785_, new_n14786_, new_n14787_, new_n14788_,
    new_n14789_, new_n14790_, new_n14791_, new_n14792_, new_n14793_,
    new_n14794_, new_n14795_, new_n14796_, new_n14797_, new_n14798_,
    new_n14799_, new_n14800_, new_n14801_, new_n14802_, new_n14803_,
    new_n14804_, new_n14805_, new_n14806_, new_n14807_, new_n14808_,
    new_n14809_, new_n14810_, new_n14811_, new_n14812_, new_n14813_,
    new_n14814_, new_n14815_, new_n14816_, new_n14817_, new_n14818_,
    new_n14819_, new_n14820_, new_n14821_, new_n14822_, new_n14823_,
    new_n14824_, new_n14825_, new_n14826_, new_n14827_, new_n14828_,
    new_n14829_, new_n14830_, new_n14831_, new_n14832_, new_n14833_,
    new_n14834_, new_n14835_, new_n14836_, new_n14837_, new_n14838_,
    new_n14839_, new_n14840_, new_n14841_, new_n14842_, new_n14843_,
    new_n14844_, new_n14845_, new_n14846_, new_n14847_, new_n14848_,
    new_n14849_, new_n14850_, new_n14851_, new_n14852_, new_n14853_,
    new_n14854_, new_n14855_, new_n14856_, new_n14857_, new_n14858_,
    new_n14859_, new_n14860_, new_n14861_, new_n14862_, new_n14863_,
    new_n14864_, new_n14865_, new_n14866_, new_n14867_, new_n14868_,
    new_n14869_, new_n14870_, new_n14871_, new_n14872_, new_n14873_,
    new_n14874_, new_n14875_, new_n14876_, new_n14877_, new_n14878_,
    new_n14879_, new_n14880_, new_n14881_, new_n14882_, new_n14883_,
    new_n14884_, new_n14885_, new_n14886_, new_n14887_, new_n14888_,
    new_n14889_, new_n14890_, new_n14891_, new_n14892_, new_n14893_,
    new_n14894_, new_n14895_, new_n14896_, new_n14897_, new_n14898_,
    new_n14899_, new_n14900_, new_n14901_, new_n14902_, new_n14903_,
    new_n14904_, new_n14905_, new_n14906_, new_n14907_, new_n14908_,
    new_n14909_, new_n14910_, new_n14911_, new_n14912_, new_n14913_,
    new_n14914_, new_n14915_, new_n14916_, new_n14917_, new_n14918_,
    new_n14919_, new_n14920_, new_n14921_, new_n14922_, new_n14923_,
    new_n14924_, new_n14925_, new_n14926_, new_n14927_, new_n14928_,
    new_n14929_, new_n14930_, new_n14931_, new_n14932_, new_n14933_,
    new_n14934_, new_n14935_, new_n14936_, new_n14937_, new_n14938_,
    new_n14939_, new_n14940_, new_n14941_, new_n14942_, new_n14943_,
    new_n14944_, new_n14945_, new_n14946_, new_n14947_, new_n14948_,
    new_n14949_, new_n14950_, new_n14951_, new_n14952_, new_n14953_,
    new_n14954_, new_n14955_, new_n14956_, new_n14957_, new_n14958_,
    new_n14959_, new_n14960_, new_n14961_, new_n14962_, new_n14963_,
    new_n14964_, new_n14965_, new_n14966_, new_n14967_, new_n14968_,
    new_n14969_, new_n14970_, new_n14971_, new_n14972_, new_n14973_,
    new_n14974_, new_n14975_, new_n14976_, new_n14977_, new_n14978_,
    new_n14979_, new_n14980_, new_n14981_, new_n14982_, new_n14983_,
    new_n14984_, new_n14985_, new_n14986_, new_n14987_, new_n14988_,
    new_n14989_, new_n14990_, new_n14991_, new_n14992_, new_n14993_,
    new_n14994_, new_n14995_, new_n14996_, new_n14997_, new_n14998_,
    new_n14999_, new_n15000_, new_n15001_, new_n15002_, new_n15003_,
    new_n15004_, new_n15005_, new_n15006_, new_n15007_, new_n15008_,
    new_n15009_, new_n15010_, new_n15011_, new_n15012_, new_n15013_,
    new_n15014_, new_n15015_, new_n15016_, new_n15017_, new_n15018_,
    new_n15019_, new_n15020_, new_n15021_, new_n15022_, new_n15023_,
    new_n15024_, new_n15025_, new_n15026_, new_n15027_, new_n15028_,
    new_n15029_, new_n15030_, new_n15031_, new_n15032_, new_n15033_,
    new_n15034_, new_n15035_, new_n15036_, new_n15037_, new_n15038_,
    new_n15039_, new_n15040_, new_n15041_, new_n15042_, new_n15043_,
    new_n15044_, new_n15045_, new_n15046_, new_n15047_, new_n15048_,
    new_n15049_, new_n15050_, new_n15051_, new_n15052_, new_n15053_,
    new_n15054_, new_n15055_, new_n15056_, new_n15057_, new_n15058_,
    new_n15059_, new_n15060_, new_n15061_, new_n15062_, new_n15063_,
    new_n15064_, new_n15065_, new_n15066_, new_n15067_, new_n15068_,
    new_n15069_, new_n15070_, new_n15071_, new_n15072_, new_n15073_,
    new_n15074_, new_n15075_, new_n15076_, new_n15077_, new_n15078_,
    new_n15079_, new_n15080_, new_n15081_, new_n15082_, new_n15083_,
    new_n15084_, new_n15085_, new_n15086_, new_n15087_, new_n15088_,
    new_n15089_, new_n15090_, new_n15091_, new_n15092_, new_n15093_,
    new_n15094_, new_n15095_, new_n15096_, new_n15097_, new_n15098_,
    new_n15099_, new_n15100_, new_n15101_, new_n15102_, new_n15103_,
    new_n15104_, new_n15105_, new_n15106_, new_n15107_, new_n15108_,
    new_n15109_, new_n15110_, new_n15111_, new_n15112_, new_n15113_,
    new_n15114_, new_n15115_, new_n15116_, new_n15117_, new_n15118_,
    new_n15119_, new_n15120_, new_n15121_, new_n15122_, new_n15123_,
    new_n15124_, new_n15125_, new_n15126_, new_n15127_, new_n15128_,
    new_n15129_, new_n15130_, new_n15131_, new_n15132_, new_n15133_,
    new_n15134_, new_n15135_, new_n15136_, new_n15137_, new_n15138_,
    new_n15139_, new_n15140_, new_n15141_, new_n15142_, new_n15143_,
    new_n15144_, new_n15145_, new_n15146_, new_n15147_, new_n15148_,
    new_n15149_, new_n15150_, new_n15151_, new_n15152_, new_n15153_,
    new_n15154_, new_n15155_, new_n15156_, new_n15157_, new_n15158_,
    new_n15159_, new_n15160_, new_n15161_, new_n15162_, new_n15163_,
    new_n15164_, new_n15165_, new_n15166_, new_n15167_, new_n15168_,
    new_n15169_, new_n15170_, new_n15171_, new_n15172_, new_n15173_,
    new_n15174_, new_n15175_, new_n15176_, new_n15177_, new_n15178_,
    new_n15179_, new_n15180_, new_n15181_, new_n15182_, new_n15183_,
    new_n15184_, new_n15185_, new_n15186_, new_n15187_, new_n15188_,
    new_n15189_, new_n15190_, new_n15191_, new_n15192_, new_n15193_,
    new_n15194_, new_n15195_, new_n15196_, new_n15197_, new_n15198_,
    new_n15199_, new_n15200_, new_n15201_, new_n15202_, new_n15203_,
    new_n15204_, new_n15205_, new_n15206_, new_n15207_, new_n15208_,
    new_n15209_, new_n15210_, new_n15211_, new_n15212_, new_n15213_,
    new_n15214_, new_n15215_, new_n15216_, new_n15217_, new_n15218_,
    new_n15219_, new_n15220_, new_n15221_, new_n15222_, new_n15223_,
    new_n15224_, new_n15225_, new_n15226_, new_n15227_, new_n15228_,
    new_n15229_, new_n15230_, new_n15231_, new_n15232_, new_n15233_,
    new_n15234_, new_n15235_, new_n15236_, new_n15237_, new_n15238_,
    new_n15239_, new_n15240_, new_n15241_, new_n15242_, new_n15243_,
    new_n15244_, new_n15245_, new_n15246_, new_n15247_, new_n15248_,
    new_n15249_, new_n15250_, new_n15251_, new_n15252_, new_n15253_,
    new_n15254_, new_n15255_, new_n15256_, new_n15257_, new_n15258_,
    new_n15259_, new_n15260_, new_n15261_, new_n15262_, new_n15263_,
    new_n15264_, new_n15265_, new_n15266_, new_n15267_, new_n15268_,
    new_n15269_, new_n15270_, new_n15271_, new_n15272_, new_n15273_,
    new_n15274_, new_n15275_, new_n15276_, new_n15277_, new_n15278_,
    new_n15279_, new_n15280_, new_n15281_, new_n15282_, new_n15283_,
    new_n15284_, new_n15285_, new_n15286_, new_n15287_, new_n15288_,
    new_n15289_, new_n15290_, new_n15291_, new_n15292_, new_n15293_,
    new_n15294_, new_n15295_, new_n15296_, new_n15297_, new_n15298_,
    new_n15299_, new_n15300_, new_n15301_, new_n15302_, new_n15303_,
    new_n15304_, new_n15305_, new_n15306_, new_n15307_, new_n15308_,
    new_n15309_, new_n15310_, new_n15311_, new_n15312_, new_n15313_,
    new_n15314_, new_n15315_, new_n15316_, new_n15317_, new_n15318_,
    new_n15319_, new_n15320_, new_n15321_, new_n15322_, new_n15323_,
    new_n15324_, new_n15325_, new_n15326_, new_n15327_, new_n15328_,
    new_n15329_, new_n15330_, new_n15331_, new_n15332_, new_n15333_,
    new_n15334_, new_n15335_, new_n15336_, new_n15337_, new_n15338_,
    new_n15339_, new_n15340_, new_n15341_, new_n15342_, new_n15343_,
    new_n15344_, new_n15345_, new_n15346_, new_n15347_, new_n15348_,
    new_n15349_, new_n15350_, new_n15351_, new_n15352_, new_n15353_,
    new_n15354_, new_n15355_, new_n15356_, new_n15357_, new_n15358_,
    new_n15359_, new_n15360_, new_n15361_, new_n15362_, new_n15363_,
    new_n15364_, new_n15365_, new_n15366_, new_n15367_, new_n15368_,
    new_n15369_, new_n15370_, new_n15371_, new_n15372_, new_n15373_,
    new_n15374_, new_n15375_, new_n15376_, new_n15377_, new_n15378_,
    new_n15379_, new_n15380_, new_n15381_, new_n15382_, new_n15383_,
    new_n15384_, new_n15385_, new_n15386_, new_n15387_, new_n15388_,
    new_n15389_, new_n15390_, new_n15391_, new_n15392_, new_n15393_,
    new_n15394_, new_n15395_, new_n15396_, new_n15397_, new_n15398_,
    new_n15399_, new_n15400_, new_n15401_, new_n15402_, new_n15403_,
    new_n15404_, new_n15405_, new_n15406_, new_n15407_, new_n15408_,
    new_n15409_, new_n15410_, new_n15411_, new_n15412_, new_n15413_,
    new_n15414_, new_n15415_, new_n15416_, new_n15417_, new_n15418_,
    new_n15419_, new_n15420_, new_n15421_, new_n15422_, new_n15423_,
    new_n15424_, new_n15425_, new_n15426_, new_n15427_, new_n15428_,
    new_n15429_, new_n15430_, new_n15431_, new_n15432_, new_n15433_,
    new_n15434_, new_n15436_, new_n15437_, new_n15438_, new_n15439_,
    new_n15440_, new_n15441_, new_n15442_, new_n15443_, new_n15444_,
    new_n15445_, new_n15446_, new_n15447_, new_n15448_, new_n15449_,
    new_n15450_, new_n15451_, new_n15452_, new_n15453_, new_n15454_,
    new_n15455_, new_n15456_, new_n15457_, new_n15458_, new_n15459_,
    new_n15460_, new_n15461_, new_n15462_, new_n15463_, new_n15464_,
    new_n15465_, new_n15466_, new_n15467_, new_n15468_, new_n15469_,
    new_n15470_, new_n15471_, new_n15472_, new_n15473_, new_n15474_,
    new_n15475_, new_n15476_, new_n15477_, new_n15478_, new_n15479_,
    new_n15480_, new_n15481_, new_n15482_, new_n15483_, new_n15484_,
    new_n15485_, new_n15486_, new_n15487_, new_n15488_, new_n15489_,
    new_n15490_, new_n15491_, new_n15492_, new_n15493_, new_n15494_,
    new_n15495_, new_n15496_, new_n15497_, new_n15498_, new_n15499_,
    new_n15500_, new_n15501_, new_n15502_, new_n15503_, new_n15504_,
    new_n15505_, new_n15506_, new_n15507_, new_n15508_, new_n15509_,
    new_n15510_, new_n15511_, new_n15512_, new_n15513_, new_n15514_,
    new_n15515_, new_n15516_, new_n15517_, new_n15518_, new_n15519_,
    new_n15520_, new_n15521_, new_n15522_, new_n15523_, new_n15524_,
    new_n15525_, new_n15526_, new_n15527_, new_n15528_, new_n15529_,
    new_n15530_, new_n15531_, new_n15532_, new_n15533_, new_n15534_,
    new_n15535_, new_n15536_, new_n15537_, new_n15538_, new_n15539_,
    new_n15540_, new_n15541_, new_n15542_, new_n15543_, new_n15544_,
    new_n15545_, new_n15546_, new_n15547_, new_n15548_, new_n15549_,
    new_n15550_, new_n15551_, new_n15552_, new_n15553_, new_n15554_,
    new_n15555_, new_n15556_, new_n15557_, new_n15558_, new_n15559_,
    new_n15560_, new_n15561_, new_n15562_, new_n15563_, new_n15564_,
    new_n15565_, new_n15566_, new_n15567_, new_n15568_, new_n15569_,
    new_n15570_, new_n15571_, new_n15572_, new_n15573_, new_n15574_,
    new_n15575_, new_n15576_, new_n15577_, new_n15578_, new_n15579_,
    new_n15580_, new_n15581_, new_n15582_, new_n15583_, new_n15584_,
    new_n15585_, new_n15586_, new_n15587_, new_n15588_, new_n15589_,
    new_n15590_, new_n15591_, new_n15592_, new_n15593_, new_n15594_,
    new_n15595_, new_n15596_, new_n15597_, new_n15598_, new_n15599_,
    new_n15600_, new_n15601_, new_n15602_, new_n15603_, new_n15604_,
    new_n15605_, new_n15606_, new_n15607_, new_n15608_, new_n15609_,
    new_n15610_, new_n15611_, new_n15612_, new_n15613_, new_n15614_,
    new_n15615_, new_n15616_, new_n15617_, new_n15618_, new_n15619_,
    new_n15620_, new_n15621_, new_n15622_, new_n15623_, new_n15624_,
    new_n15625_, new_n15626_, new_n15627_, new_n15628_, new_n15629_,
    new_n15630_, new_n15631_, new_n15632_, new_n15633_, new_n15634_,
    new_n15635_, new_n15636_, new_n15637_, new_n15638_, new_n15639_,
    new_n15640_, new_n15641_, new_n15642_, new_n15643_, new_n15644_,
    new_n15645_, new_n15646_, new_n15647_, new_n15648_, new_n15649_,
    new_n15650_, new_n15651_, new_n15652_, new_n15653_, new_n15654_,
    new_n15655_, new_n15656_, new_n15657_, new_n15658_, new_n15659_,
    new_n15660_, new_n15661_, new_n15662_, new_n15663_, new_n15664_,
    new_n15665_, new_n15666_, new_n15667_, new_n15668_, new_n15669_,
    new_n15670_, new_n15671_, new_n15672_, new_n15673_, new_n15674_,
    new_n15675_, new_n15676_, new_n15677_, new_n15678_, new_n15679_,
    new_n15680_, new_n15681_, new_n15682_, new_n15683_, new_n15684_,
    new_n15685_, new_n15686_, new_n15687_, new_n15688_, new_n15689_,
    new_n15690_, new_n15691_, new_n15692_, new_n15693_, new_n15694_,
    new_n15695_, new_n15696_, new_n15697_, new_n15698_, new_n15699_,
    new_n15700_, new_n15701_, new_n15702_, new_n15703_, new_n15704_,
    new_n15705_, new_n15706_, new_n15707_, new_n15708_, new_n15709_,
    new_n15710_, new_n15711_, new_n15712_, new_n15713_, new_n15714_,
    new_n15715_, new_n15716_, new_n15717_, new_n15718_, new_n15719_,
    new_n15720_, new_n15721_, new_n15722_, new_n15723_, new_n15724_,
    new_n15725_, new_n15726_, new_n15727_, new_n15728_, new_n15729_,
    new_n15730_, new_n15731_, new_n15732_, new_n15733_, new_n15734_,
    new_n15735_, new_n15736_, new_n15737_, new_n15738_, new_n15739_,
    new_n15740_, new_n15741_, new_n15742_, new_n15743_, new_n15744_,
    new_n15745_, new_n15746_, new_n15747_, new_n15748_, new_n15749_,
    new_n15750_, new_n15751_, new_n15752_, new_n15753_, new_n15754_,
    new_n15755_, new_n15756_, new_n15757_, new_n15758_, new_n15759_,
    new_n15760_, new_n15761_, new_n15762_, new_n15763_, new_n15764_,
    new_n15765_, new_n15766_, new_n15767_, new_n15768_, new_n15769_,
    new_n15770_, new_n15771_, new_n15772_, new_n15773_, new_n15774_,
    new_n15775_, new_n15776_, new_n15777_, new_n15778_, new_n15779_,
    new_n15780_, new_n15781_, new_n15782_, new_n15783_, new_n15784_,
    new_n15785_, new_n15786_, new_n15787_, new_n15788_, new_n15789_,
    new_n15790_, new_n15791_, new_n15792_, new_n15793_, new_n15794_,
    new_n15795_, new_n15796_, new_n15797_, new_n15798_, new_n15799_,
    new_n15800_, new_n15801_, new_n15802_, new_n15803_, new_n15804_,
    new_n15805_, new_n15806_, new_n15807_, new_n15808_, new_n15809_,
    new_n15810_, new_n15811_, new_n15812_, new_n15813_, new_n15814_,
    new_n15815_, new_n15816_, new_n15817_, new_n15818_, new_n15819_,
    new_n15820_, new_n15821_, new_n15822_, new_n15823_, new_n15824_,
    new_n15825_, new_n15826_, new_n15827_, new_n15828_, new_n15829_,
    new_n15830_, new_n15831_, new_n15832_, new_n15833_, new_n15834_,
    new_n15835_, new_n15836_, new_n15837_, new_n15838_, new_n15839_,
    new_n15840_, new_n15841_, new_n15842_, new_n15843_, new_n15844_,
    new_n15845_, new_n15846_, new_n15847_, new_n15848_, new_n15849_,
    new_n15850_, new_n15851_, new_n15852_, new_n15853_, new_n15854_,
    new_n15855_, new_n15856_, new_n15857_, new_n15858_, new_n15859_,
    new_n15860_, new_n15861_, new_n15862_, new_n15863_, new_n15864_,
    new_n15865_, new_n15866_, new_n15867_, new_n15868_, new_n15869_,
    new_n15870_, new_n15871_, new_n15872_, new_n15873_, new_n15874_,
    new_n15875_, new_n15876_, new_n15877_, new_n15878_, new_n15879_,
    new_n15880_, new_n15881_, new_n15882_, new_n15883_, new_n15884_,
    new_n15885_, new_n15886_, new_n15887_, new_n15888_, new_n15889_,
    new_n15890_, new_n15891_, new_n15892_, new_n15893_, new_n15894_,
    new_n15895_, new_n15896_, new_n15897_, new_n15898_, new_n15899_,
    new_n15900_, new_n15901_, new_n15902_, new_n15903_, new_n15904_,
    new_n15905_, new_n15906_, new_n15907_, new_n15908_, new_n15909_,
    new_n15910_, new_n15911_, new_n15912_, new_n15913_, new_n15914_,
    new_n15915_, new_n15916_, new_n15917_, new_n15918_, new_n15919_,
    new_n15920_, new_n15921_, new_n15922_, new_n15923_, new_n15924_,
    new_n15925_, new_n15926_, new_n15927_, new_n15928_, new_n15929_,
    new_n15930_, new_n15931_, new_n15932_, new_n15933_, new_n15934_,
    new_n15935_, new_n15936_, new_n15937_, new_n15938_, new_n15939_,
    new_n15940_, new_n15941_, new_n15942_, new_n15943_, new_n15944_,
    new_n15945_, new_n15946_, new_n15947_, new_n15948_, new_n15949_,
    new_n15950_, new_n15951_, new_n15952_, new_n15953_, new_n15954_,
    new_n15955_, new_n15956_, new_n15957_, new_n15958_, new_n15959_,
    new_n15960_, new_n15961_, new_n15962_, new_n15963_, new_n15964_,
    new_n15965_, new_n15966_, new_n15967_, new_n15968_, new_n15969_,
    new_n15970_, new_n15971_, new_n15972_, new_n15973_, new_n15974_,
    new_n15975_, new_n15976_, new_n15977_, new_n15978_, new_n15979_,
    new_n15980_, new_n15981_, new_n15982_, new_n15983_, new_n15984_,
    new_n15985_, new_n15986_, new_n15987_, new_n15988_, new_n15989_,
    new_n15990_, new_n15991_, new_n15992_, new_n15993_, new_n15994_,
    new_n15995_, new_n15996_, new_n15997_, new_n15998_, new_n15999_,
    new_n16000_, new_n16002_, new_n16003_, new_n16004_, new_n16005_,
    new_n16006_, new_n16007_, new_n16008_, new_n16009_, new_n16010_,
    new_n16011_, new_n16012_, new_n16013_, new_n16014_, new_n16015_,
    new_n16016_, new_n16017_, new_n16018_, new_n16019_, new_n16020_,
    new_n16021_, new_n16022_, new_n16023_, new_n16024_, new_n16025_,
    new_n16026_, new_n16027_, new_n16028_, new_n16029_, new_n16030_,
    new_n16031_, new_n16032_, new_n16033_, new_n16034_, new_n16035_,
    new_n16036_, new_n16037_, new_n16038_, new_n16039_, new_n16040_,
    new_n16041_, new_n16042_, new_n16043_, new_n16044_, new_n16045_,
    new_n16046_, new_n16047_, new_n16048_, new_n16049_, new_n16050_,
    new_n16051_, new_n16052_, new_n16053_, new_n16054_, new_n16055_,
    new_n16056_, new_n16057_, new_n16058_, new_n16059_, new_n16060_,
    new_n16061_, new_n16062_, new_n16063_, new_n16064_, new_n16065_,
    new_n16066_, new_n16067_, new_n16068_, new_n16069_, new_n16070_,
    new_n16071_, new_n16072_, new_n16073_, new_n16074_, new_n16075_,
    new_n16076_, new_n16077_, new_n16078_, new_n16079_, new_n16080_,
    new_n16081_, new_n16082_, new_n16083_, new_n16084_, new_n16085_,
    new_n16086_, new_n16087_, new_n16088_, new_n16089_, new_n16090_,
    new_n16091_, new_n16092_, new_n16093_, new_n16094_, new_n16095_,
    new_n16096_, new_n16097_, new_n16098_, new_n16099_, new_n16100_,
    new_n16101_, new_n16102_, new_n16103_, new_n16104_, new_n16105_,
    new_n16106_, new_n16107_, new_n16108_, new_n16109_, new_n16110_,
    new_n16111_, new_n16112_, new_n16113_, new_n16114_, new_n16115_,
    new_n16116_, new_n16117_, new_n16118_, new_n16119_, new_n16120_,
    new_n16121_, new_n16122_, new_n16123_, new_n16124_, new_n16125_,
    new_n16126_, new_n16127_, new_n16128_, new_n16129_, new_n16130_,
    new_n16131_, new_n16132_, new_n16133_, new_n16134_, new_n16135_,
    new_n16136_, new_n16137_, new_n16138_, new_n16139_, new_n16140_,
    new_n16141_, new_n16142_, new_n16143_, new_n16144_, new_n16145_,
    new_n16146_, new_n16147_, new_n16148_, new_n16149_, new_n16150_,
    new_n16151_, new_n16152_, new_n16153_, new_n16154_, new_n16155_,
    new_n16156_, new_n16157_, new_n16158_, new_n16159_, new_n16160_,
    new_n16161_, new_n16162_, new_n16163_, new_n16164_, new_n16165_,
    new_n16166_, new_n16167_, new_n16168_, new_n16169_, new_n16170_,
    new_n16171_, new_n16172_, new_n16173_, new_n16174_, new_n16175_,
    new_n16176_, new_n16177_, new_n16178_, new_n16179_, new_n16180_,
    new_n16181_, new_n16182_, new_n16183_, new_n16184_, new_n16185_,
    new_n16186_, new_n16187_, new_n16188_, new_n16189_, new_n16190_,
    new_n16191_, new_n16192_, new_n16193_, new_n16194_, new_n16195_,
    new_n16196_, new_n16197_, new_n16198_, new_n16199_, new_n16200_,
    new_n16201_, new_n16202_, new_n16203_, new_n16204_, new_n16205_,
    new_n16206_, new_n16207_, new_n16208_, new_n16209_, new_n16210_,
    new_n16211_, new_n16212_, new_n16213_, new_n16214_, new_n16215_,
    new_n16216_, new_n16217_, new_n16218_, new_n16219_, new_n16220_,
    new_n16221_, new_n16222_, new_n16223_, new_n16224_, new_n16225_,
    new_n16226_, new_n16227_, new_n16228_, new_n16229_, new_n16230_,
    new_n16231_, new_n16232_, new_n16233_, new_n16234_, new_n16235_,
    new_n16236_, new_n16237_, new_n16238_, new_n16239_, new_n16240_,
    new_n16241_, new_n16242_, new_n16243_, new_n16244_, new_n16245_,
    new_n16246_, new_n16247_, new_n16248_, new_n16249_, new_n16250_,
    new_n16251_, new_n16252_, new_n16253_, new_n16254_, new_n16255_,
    new_n16256_, new_n16257_, new_n16258_, new_n16259_, new_n16260_,
    new_n16261_, new_n16262_, new_n16263_, new_n16264_, new_n16265_,
    new_n16266_, new_n16267_, new_n16268_, new_n16269_, new_n16270_,
    new_n16271_, new_n16272_, new_n16273_, new_n16274_, new_n16275_,
    new_n16276_, new_n16277_, new_n16278_, new_n16279_, new_n16280_,
    new_n16281_, new_n16282_, new_n16283_, new_n16284_, new_n16285_,
    new_n16286_, new_n16287_, new_n16288_, new_n16289_, new_n16290_,
    new_n16291_, new_n16292_, new_n16293_, new_n16294_, new_n16295_,
    new_n16296_, new_n16297_, new_n16298_, new_n16299_, new_n16300_,
    new_n16301_, new_n16302_, new_n16303_, new_n16304_, new_n16305_,
    new_n16306_, new_n16307_, new_n16308_, new_n16309_, new_n16310_,
    new_n16311_, new_n16312_, new_n16313_, new_n16314_, new_n16315_,
    new_n16316_, new_n16317_, new_n16318_, new_n16319_, new_n16320_,
    new_n16321_, new_n16322_, new_n16323_, new_n16324_, new_n16325_,
    new_n16326_, new_n16327_, new_n16328_, new_n16329_, new_n16330_,
    new_n16331_, new_n16332_, new_n16333_, new_n16334_, new_n16335_,
    new_n16336_, new_n16337_, new_n16338_, new_n16339_, new_n16340_,
    new_n16341_, new_n16342_, new_n16343_, new_n16344_, new_n16345_,
    new_n16346_, new_n16347_, new_n16348_, new_n16349_, new_n16350_,
    new_n16351_, new_n16352_, new_n16353_, new_n16354_, new_n16355_,
    new_n16356_, new_n16357_, new_n16358_, new_n16359_, new_n16360_,
    new_n16361_, new_n16362_, new_n16363_, new_n16364_, new_n16365_,
    new_n16366_, new_n16367_, new_n16368_, new_n16369_, new_n16370_,
    new_n16371_, new_n16372_, new_n16373_, new_n16374_, new_n16375_,
    new_n16376_, new_n16377_, new_n16378_, new_n16379_, new_n16380_,
    new_n16381_, new_n16382_, new_n16383_, new_n16384_, new_n16385_,
    new_n16386_, new_n16387_, new_n16388_, new_n16389_, new_n16390_,
    new_n16391_, new_n16392_, new_n16393_, new_n16394_, new_n16395_,
    new_n16396_, new_n16397_, new_n16398_, new_n16399_, new_n16400_,
    new_n16401_, new_n16402_, new_n16403_, new_n16404_, new_n16405_,
    new_n16406_, new_n16407_, new_n16408_, new_n16409_, new_n16410_,
    new_n16411_, new_n16412_, new_n16413_, new_n16414_, new_n16415_,
    new_n16416_, new_n16417_, new_n16418_, new_n16419_, new_n16420_,
    new_n16421_, new_n16422_, new_n16423_, new_n16424_, new_n16425_,
    new_n16426_, new_n16427_, new_n16428_, new_n16429_, new_n16430_,
    new_n16431_, new_n16432_, new_n16433_, new_n16434_, new_n16435_,
    new_n16436_, new_n16437_, new_n16438_, new_n16439_, new_n16440_,
    new_n16441_, new_n16442_, new_n16443_, new_n16444_, new_n16445_,
    new_n16446_, new_n16447_, new_n16448_, new_n16449_, new_n16450_,
    new_n16451_, new_n16452_, new_n16453_, new_n16454_, new_n16455_,
    new_n16456_, new_n16457_, new_n16458_, new_n16459_, new_n16460_,
    new_n16461_, new_n16462_, new_n16463_, new_n16464_, new_n16465_,
    new_n16466_, new_n16467_, new_n16468_, new_n16469_, new_n16470_,
    new_n16471_, new_n16472_, new_n16473_, new_n16474_, new_n16475_,
    new_n16476_, new_n16477_, new_n16478_, new_n16479_, new_n16480_,
    new_n16481_, new_n16482_, new_n16483_, new_n16484_, new_n16485_,
    new_n16486_, new_n16487_, new_n16488_, new_n16489_, new_n16490_,
    new_n16491_, new_n16492_, new_n16493_, new_n16494_, new_n16495_,
    new_n16496_, new_n16497_, new_n16498_, new_n16499_, new_n16500_,
    new_n16501_, new_n16502_, new_n16503_, new_n16504_, new_n16505_,
    new_n16506_, new_n16507_, new_n16508_, new_n16509_, new_n16510_,
    new_n16511_, new_n16512_, new_n16513_, new_n16514_, new_n16515_,
    new_n16516_, new_n16517_, new_n16518_, new_n16519_, new_n16520_,
    new_n16521_, new_n16522_, new_n16523_, new_n16524_, new_n16525_,
    new_n16526_, new_n16527_, new_n16528_, new_n16529_, new_n16530_,
    new_n16531_, new_n16532_, new_n16533_, new_n16534_, new_n16535_,
    new_n16536_, new_n16537_, new_n16538_, new_n16539_, new_n16540_,
    new_n16541_, new_n16542_, new_n16543_, new_n16544_, new_n16545_,
    new_n16546_, new_n16547_, new_n16548_, new_n16549_, new_n16550_,
    new_n16551_, new_n16552_, new_n16553_, new_n16554_, new_n16555_,
    new_n16556_, new_n16557_, new_n16558_, new_n16559_, new_n16560_,
    new_n16561_, new_n16562_, new_n16563_, new_n16564_, new_n16565_,
    new_n16566_, new_n16567_, new_n16568_, new_n16569_, new_n16570_,
    new_n16571_, new_n16572_, new_n16573_, new_n16574_, new_n16575_,
    new_n16576_, new_n16577_, new_n16578_, new_n16579_, new_n16580_,
    new_n16581_, new_n16582_, new_n16583_, new_n16584_, new_n16585_,
    new_n16586_, new_n16587_, new_n16588_, new_n16589_, new_n16590_,
    new_n16591_, new_n16592_, new_n16593_, new_n16594_, new_n16595_,
    new_n16596_, new_n16597_, new_n16598_, new_n16599_, new_n16600_,
    new_n16601_, new_n16602_, new_n16603_, new_n16604_, new_n16605_,
    new_n16606_, new_n16607_, new_n16608_, new_n16609_, new_n16610_,
    new_n16611_, new_n16612_, new_n16613_, new_n16614_, new_n16615_,
    new_n16616_, new_n16617_, new_n16619_, new_n16620_, new_n16621_,
    new_n16622_, new_n16623_, new_n16624_, new_n16625_, new_n16626_,
    new_n16627_, new_n16628_, new_n16629_, new_n16630_, new_n16631_,
    new_n16632_, new_n16633_, new_n16634_, new_n16635_, new_n16636_,
    new_n16637_, new_n16638_, new_n16639_, new_n16640_, new_n16641_,
    new_n16642_, new_n16643_, new_n16644_, new_n16645_, new_n16646_,
    new_n16647_, new_n16648_, new_n16649_, new_n16650_, new_n16651_,
    new_n16652_, new_n16653_, new_n16654_, new_n16655_, new_n16656_,
    new_n16657_, new_n16658_, new_n16659_, new_n16660_, new_n16661_,
    new_n16662_, new_n16663_, new_n16664_, new_n16665_, new_n16666_,
    new_n16667_, new_n16668_, new_n16669_, new_n16670_, new_n16671_,
    new_n16672_, new_n16673_, new_n16674_, new_n16675_, new_n16676_,
    new_n16677_, new_n16678_, new_n16679_, new_n16680_, new_n16681_,
    new_n16682_, new_n16683_, new_n16684_, new_n16685_, new_n16686_,
    new_n16687_, new_n16688_, new_n16689_, new_n16690_, new_n16691_,
    new_n16692_, new_n16693_, new_n16694_, new_n16695_, new_n16696_,
    new_n16697_, new_n16698_, new_n16699_, new_n16700_, new_n16701_,
    new_n16702_, new_n16703_, new_n16704_, new_n16705_, new_n16706_,
    new_n16707_, new_n16708_, new_n16709_, new_n16710_, new_n16711_,
    new_n16712_, new_n16713_, new_n16714_, new_n16715_, new_n16716_,
    new_n16717_, new_n16718_, new_n16719_, new_n16720_, new_n16721_,
    new_n16722_, new_n16723_, new_n16724_, new_n16725_, new_n16726_,
    new_n16727_, new_n16728_, new_n16729_, new_n16730_, new_n16731_,
    new_n16732_, new_n16733_, new_n16734_, new_n16735_, new_n16736_,
    new_n16737_, new_n16738_, new_n16739_, new_n16740_, new_n16741_,
    new_n16742_, new_n16743_, new_n16744_, new_n16745_, new_n16746_,
    new_n16747_, new_n16748_, new_n16749_, new_n16750_, new_n16751_,
    new_n16752_, new_n16753_, new_n16754_, new_n16755_, new_n16756_,
    new_n16757_, new_n16758_, new_n16759_, new_n16760_, new_n16761_,
    new_n16762_, new_n16763_, new_n16764_, new_n16765_, new_n16766_,
    new_n16767_, new_n16768_, new_n16769_, new_n16770_, new_n16771_,
    new_n16772_, new_n16773_, new_n16774_, new_n16775_, new_n16776_,
    new_n16777_, new_n16778_, new_n16779_, new_n16780_, new_n16781_,
    new_n16782_, new_n16783_, new_n16784_, new_n16785_, new_n16786_,
    new_n16787_, new_n16788_, new_n16789_, new_n16790_, new_n16791_,
    new_n16792_, new_n16793_, new_n16794_, new_n16795_, new_n16796_,
    new_n16797_, new_n16798_, new_n16799_, new_n16800_, new_n16801_,
    new_n16802_, new_n16803_, new_n16804_, new_n16805_, new_n16806_,
    new_n16807_, new_n16808_, new_n16809_, new_n16810_, new_n16811_,
    new_n16812_, new_n16813_, new_n16814_, new_n16815_, new_n16816_,
    new_n16817_, new_n16818_, new_n16819_, new_n16820_, new_n16821_,
    new_n16822_, new_n16823_, new_n16824_, new_n16825_, new_n16826_,
    new_n16827_, new_n16828_, new_n16829_, new_n16830_, new_n16831_,
    new_n16832_, new_n16833_, new_n16834_, new_n16835_, new_n16836_,
    new_n16837_, new_n16838_, new_n16839_, new_n16840_, new_n16841_,
    new_n16842_, new_n16843_, new_n16844_, new_n16845_, new_n16846_,
    new_n16847_, new_n16848_, new_n16849_, new_n16850_, new_n16851_,
    new_n16852_, new_n16853_, new_n16854_, new_n16855_, new_n16856_,
    new_n16857_, new_n16858_, new_n16859_, new_n16860_, new_n16861_,
    new_n16862_, new_n16863_, new_n16864_, new_n16865_, new_n16866_,
    new_n16867_, new_n16868_, new_n16869_, new_n16870_, new_n16871_,
    new_n16872_, new_n16873_, new_n16874_, new_n16875_, new_n16876_,
    new_n16877_, new_n16878_, new_n16879_, new_n16880_, new_n16881_,
    new_n16882_, new_n16883_, new_n16884_, new_n16885_, new_n16886_,
    new_n16887_, new_n16888_, new_n16889_, new_n16890_, new_n16891_,
    new_n16892_, new_n16893_, new_n16894_, new_n16895_, new_n16896_,
    new_n16897_, new_n16898_, new_n16899_, new_n16900_, new_n16901_,
    new_n16902_, new_n16903_, new_n16904_, new_n16905_, new_n16906_,
    new_n16907_, new_n16908_, new_n16909_, new_n16910_, new_n16911_,
    new_n16912_, new_n16913_, new_n16914_, new_n16915_, new_n16916_,
    new_n16917_, new_n16918_, new_n16919_, new_n16920_, new_n16921_,
    new_n16922_, new_n16923_, new_n16924_, new_n16925_, new_n16926_,
    new_n16927_, new_n16928_, new_n16929_, new_n16930_, new_n16931_,
    new_n16932_, new_n16933_, new_n16934_, new_n16935_, new_n16936_,
    new_n16937_, new_n16938_, new_n16939_, new_n16940_, new_n16941_,
    new_n16942_, new_n16943_, new_n16944_, new_n16945_, new_n16946_,
    new_n16947_, new_n16948_, new_n16949_, new_n16950_, new_n16951_,
    new_n16952_, new_n16953_, new_n16954_, new_n16955_, new_n16956_,
    new_n16957_, new_n16958_, new_n16959_, new_n16960_, new_n16961_,
    new_n16962_, new_n16963_, new_n16964_, new_n16965_, new_n16966_,
    new_n16967_, new_n16968_, new_n16969_, new_n16970_, new_n16971_,
    new_n16972_, new_n16973_, new_n16974_, new_n16975_, new_n16976_,
    new_n16977_, new_n16978_, new_n16979_, new_n16980_, new_n16981_,
    new_n16982_, new_n16983_, new_n16984_, new_n16985_, new_n16986_,
    new_n16987_, new_n16988_, new_n16989_, new_n16990_, new_n16991_,
    new_n16992_, new_n16993_, new_n16994_, new_n16995_, new_n16996_,
    new_n16997_, new_n16998_, new_n16999_, new_n17000_, new_n17001_,
    new_n17002_, new_n17003_, new_n17004_, new_n17005_, new_n17006_,
    new_n17007_, new_n17008_, new_n17009_, new_n17010_, new_n17011_,
    new_n17012_, new_n17013_, new_n17014_, new_n17015_, new_n17016_,
    new_n17017_, new_n17018_, new_n17019_, new_n17020_, new_n17021_,
    new_n17022_, new_n17023_, new_n17024_, new_n17025_, new_n17026_,
    new_n17027_, new_n17028_, new_n17029_, new_n17030_, new_n17031_,
    new_n17032_, new_n17033_, new_n17034_, new_n17035_, new_n17036_,
    new_n17037_, new_n17038_, new_n17039_, new_n17040_, new_n17041_,
    new_n17042_, new_n17043_, new_n17044_, new_n17045_, new_n17046_,
    new_n17047_, new_n17048_, new_n17049_, new_n17050_, new_n17051_,
    new_n17052_, new_n17053_, new_n17054_, new_n17055_, new_n17056_,
    new_n17057_, new_n17058_, new_n17059_, new_n17060_, new_n17061_,
    new_n17062_, new_n17063_, new_n17064_, new_n17065_, new_n17066_,
    new_n17067_, new_n17068_, new_n17069_, new_n17070_, new_n17071_,
    new_n17072_, new_n17073_, new_n17074_, new_n17075_, new_n17076_,
    new_n17077_, new_n17078_, new_n17079_, new_n17080_, new_n17081_,
    new_n17082_, new_n17083_, new_n17084_, new_n17085_, new_n17086_,
    new_n17087_, new_n17088_, new_n17089_, new_n17090_, new_n17091_,
    new_n17092_, new_n17093_, new_n17094_, new_n17095_, new_n17096_,
    new_n17097_, new_n17098_, new_n17099_, new_n17100_, new_n17101_,
    new_n17102_, new_n17103_, new_n17104_, new_n17105_, new_n17106_,
    new_n17107_, new_n17108_, new_n17109_, new_n17110_, new_n17111_,
    new_n17112_, new_n17113_, new_n17114_, new_n17115_, new_n17116_,
    new_n17117_, new_n17118_, new_n17119_, new_n17120_, new_n17121_,
    new_n17122_, new_n17123_, new_n17124_, new_n17125_, new_n17126_,
    new_n17127_, new_n17128_, new_n17129_, new_n17130_, new_n17131_,
    new_n17132_, new_n17133_, new_n17134_, new_n17135_, new_n17136_,
    new_n17137_, new_n17138_, new_n17139_, new_n17140_, new_n17141_,
    new_n17142_, new_n17143_, new_n17144_, new_n17145_, new_n17146_,
    new_n17147_, new_n17148_, new_n17149_, new_n17150_, new_n17151_,
    new_n17152_, new_n17153_, new_n17154_, new_n17155_, new_n17156_,
    new_n17157_, new_n17158_, new_n17159_, new_n17160_, new_n17161_,
    new_n17162_, new_n17163_, new_n17164_, new_n17165_, new_n17166_,
    new_n17167_, new_n17168_, new_n17169_, new_n17170_, new_n17171_,
    new_n17172_, new_n17173_, new_n17174_, new_n17175_, new_n17176_,
    new_n17177_, new_n17178_, new_n17179_, new_n17180_, new_n17181_,
    new_n17182_, new_n17183_, new_n17184_, new_n17185_, new_n17186_,
    new_n17187_, new_n17188_, new_n17189_, new_n17190_, new_n17191_,
    new_n17192_, new_n17193_, new_n17194_, new_n17195_, new_n17196_,
    new_n17197_, new_n17198_, new_n17199_, new_n17200_, new_n17201_,
    new_n17202_, new_n17203_, new_n17204_, new_n17205_, new_n17206_,
    new_n17207_, new_n17208_, new_n17209_, new_n17210_, new_n17211_,
    new_n17212_, new_n17213_, new_n17214_, new_n17215_, new_n17216_,
    new_n17217_, new_n17218_, new_n17219_, new_n17220_, new_n17221_,
    new_n17222_, new_n17223_, new_n17224_, new_n17225_, new_n17226_,
    new_n17227_, new_n17228_, new_n17229_, new_n17230_, new_n17231_,
    new_n17232_, new_n17233_, new_n17234_, new_n17235_, new_n17236_,
    new_n17237_, new_n17238_, new_n17239_, new_n17240_, new_n17241_,
    new_n17242_, new_n17243_, new_n17244_, new_n17245_, new_n17246_,
    new_n17247_, new_n17248_, new_n17249_, new_n17250_, new_n17251_,
    new_n17252_, new_n17253_, new_n17254_, new_n17255_, new_n17256_,
    new_n17257_, new_n17258_, new_n17259_, new_n17260_, new_n17261_,
    new_n17262_, new_n17263_, new_n17264_, new_n17265_, new_n17266_,
    new_n17267_, new_n17268_, new_n17269_, new_n17270_, new_n17271_,
    new_n17272_, new_n17273_, new_n17274_, new_n17275_, new_n17276_,
    new_n17277_, new_n17278_, new_n17279_, new_n17280_, new_n17281_,
    new_n17282_, new_n17283_, new_n17284_, new_n17285_, new_n17286_,
    new_n17287_, new_n17288_, new_n17289_, new_n17290_, new_n17291_,
    new_n17292_, new_n17293_, new_n17294_, new_n17295_, new_n17296_,
    new_n17297_, new_n17298_, new_n17299_, new_n17300_, new_n17301_,
    new_n17302_, new_n17303_, new_n17304_, new_n17305_, new_n17306_,
    new_n17307_, new_n17308_, new_n17309_, new_n17310_, new_n17311_,
    new_n17312_, new_n17313_, new_n17314_, new_n17315_, new_n17316_,
    new_n17317_, new_n17318_, new_n17319_, new_n17320_, new_n17321_,
    new_n17322_, new_n17323_, new_n17324_, new_n17325_, new_n17326_,
    new_n17327_, new_n17328_, new_n17329_, new_n17330_, new_n17331_,
    new_n17332_, new_n17333_, new_n17334_, new_n17335_, new_n17336_,
    new_n17337_, new_n17338_, new_n17339_, new_n17340_, new_n17341_,
    new_n17342_, new_n17344_, new_n17345_, new_n17346_, new_n17347_,
    new_n17348_, new_n17349_, new_n17350_, new_n17351_, new_n17352_,
    new_n17353_, new_n17354_, new_n17355_, new_n17356_, new_n17357_,
    new_n17358_, new_n17359_, new_n17360_, new_n17361_, new_n17362_,
    new_n17363_, new_n17364_, new_n17365_, new_n17366_, new_n17367_,
    new_n17368_, new_n17369_, new_n17370_, new_n17371_, new_n17372_,
    new_n17373_, new_n17374_, new_n17375_, new_n17376_, new_n17377_,
    new_n17378_, new_n17379_, new_n17380_, new_n17381_, new_n17382_,
    new_n17383_, new_n17384_, new_n17385_, new_n17386_, new_n17387_,
    new_n17388_, new_n17389_, new_n17390_, new_n17391_, new_n17392_,
    new_n17393_, new_n17394_, new_n17395_, new_n17396_, new_n17397_,
    new_n17398_, new_n17399_, new_n17400_, new_n17401_, new_n17402_,
    new_n17403_, new_n17404_, new_n17405_, new_n17406_, new_n17407_,
    new_n17408_, new_n17409_, new_n17410_, new_n17411_, new_n17412_,
    new_n17413_, new_n17414_, new_n17415_, new_n17416_, new_n17417_,
    new_n17418_, new_n17419_, new_n17420_, new_n17421_, new_n17422_,
    new_n17423_, new_n17424_, new_n17425_, new_n17426_, new_n17427_,
    new_n17428_, new_n17429_, new_n17430_, new_n17431_, new_n17432_,
    new_n17433_, new_n17434_, new_n17435_, new_n17436_, new_n17437_,
    new_n17438_, new_n17439_, new_n17440_, new_n17441_, new_n17442_,
    new_n17443_, new_n17444_, new_n17445_, new_n17446_, new_n17447_,
    new_n17448_, new_n17449_, new_n17450_, new_n17451_, new_n17452_,
    new_n17453_, new_n17454_, new_n17455_, new_n17456_, new_n17457_,
    new_n17458_, new_n17459_, new_n17460_, new_n17461_, new_n17462_,
    new_n17463_, new_n17464_, new_n17465_, new_n17466_, new_n17467_,
    new_n17468_, new_n17469_, new_n17470_, new_n17471_, new_n17472_,
    new_n17473_, new_n17474_, new_n17475_, new_n17476_, new_n17477_,
    new_n17478_, new_n17479_, new_n17480_, new_n17481_, new_n17482_,
    new_n17483_, new_n17484_, new_n17485_, new_n17486_, new_n17487_,
    new_n17488_, new_n17489_, new_n17490_, new_n17491_, new_n17492_,
    new_n17493_, new_n17494_, new_n17495_, new_n17496_, new_n17497_,
    new_n17498_, new_n17499_, new_n17500_, new_n17501_, new_n17502_,
    new_n17503_, new_n17504_, new_n17505_, new_n17506_, new_n17507_,
    new_n17508_, new_n17509_, new_n17510_, new_n17511_, new_n17512_,
    new_n17513_, new_n17514_, new_n17515_, new_n17516_, new_n17517_,
    new_n17518_, new_n17519_, new_n17520_, new_n17521_, new_n17522_,
    new_n17523_, new_n17524_, new_n17525_, new_n17526_, new_n17527_,
    new_n17528_, new_n17529_, new_n17530_, new_n17531_, new_n17532_,
    new_n17533_, new_n17534_, new_n17535_, new_n17536_, new_n17537_,
    new_n17538_, new_n17539_, new_n17540_, new_n17541_, new_n17542_,
    new_n17543_, new_n17544_, new_n17545_, new_n17546_, new_n17547_,
    new_n17548_, new_n17549_, new_n17550_, new_n17551_, new_n17552_,
    new_n17553_, new_n17554_, new_n17555_, new_n17556_, new_n17557_,
    new_n17558_, new_n17559_, new_n17560_, new_n17561_, new_n17562_,
    new_n17563_, new_n17564_, new_n17565_, new_n17566_, new_n17567_,
    new_n17568_, new_n17569_, new_n17570_, new_n17571_, new_n17572_,
    new_n17573_, new_n17574_, new_n17575_, new_n17576_, new_n17577_,
    new_n17578_, new_n17579_, new_n17580_, new_n17581_, new_n17582_,
    new_n17583_, new_n17584_, new_n17585_, new_n17586_, new_n17587_,
    new_n17588_, new_n17589_, new_n17590_, new_n17591_, new_n17592_,
    new_n17593_, new_n17594_, new_n17595_, new_n17596_, new_n17597_,
    new_n17598_, new_n17599_, new_n17600_, new_n17601_, new_n17602_,
    new_n17603_, new_n17604_, new_n17605_, new_n17606_, new_n17607_,
    new_n17608_, new_n17609_, new_n17610_, new_n17611_, new_n17612_,
    new_n17613_, new_n17614_, new_n17615_, new_n17616_, new_n17617_,
    new_n17618_, new_n17619_, new_n17620_, new_n17621_, new_n17622_,
    new_n17623_, new_n17624_, new_n17625_, new_n17626_, new_n17627_,
    new_n17628_, new_n17629_, new_n17630_, new_n17631_, new_n17632_,
    new_n17633_, new_n17634_, new_n17635_, new_n17636_, new_n17637_,
    new_n17638_, new_n17639_, new_n17640_, new_n17641_, new_n17642_,
    new_n17643_, new_n17644_, new_n17645_, new_n17646_, new_n17647_,
    new_n17648_, new_n17649_, new_n17650_, new_n17651_, new_n17652_,
    new_n17653_, new_n17654_, new_n17655_, new_n17656_, new_n17657_,
    new_n17658_, new_n17659_, new_n17660_, new_n17661_, new_n17662_,
    new_n17663_, new_n17664_, new_n17665_, new_n17666_, new_n17667_,
    new_n17668_, new_n17669_, new_n17670_, new_n17671_, new_n17672_,
    new_n17673_, new_n17674_, new_n17675_, new_n17676_, new_n17677_,
    new_n17678_, new_n17679_, new_n17680_, new_n17681_, new_n17682_,
    new_n17683_, new_n17684_, new_n17685_, new_n17686_, new_n17687_,
    new_n17688_, new_n17689_, new_n17690_, new_n17691_, new_n17692_,
    new_n17693_, new_n17694_, new_n17695_, new_n17696_, new_n17697_,
    new_n17698_, new_n17699_, new_n17700_, new_n17701_, new_n17702_,
    new_n17703_, new_n17704_, new_n17705_, new_n17706_, new_n17707_,
    new_n17708_, new_n17709_, new_n17710_, new_n17711_, new_n17712_,
    new_n17713_, new_n17714_, new_n17715_, new_n17716_, new_n17717_,
    new_n17718_, new_n17719_, new_n17720_, new_n17721_, new_n17722_,
    new_n17723_, new_n17724_, new_n17725_, new_n17726_, new_n17727_,
    new_n17728_, new_n17729_, new_n17730_, new_n17731_, new_n17732_,
    new_n17733_, new_n17734_, new_n17735_, new_n17736_, new_n17737_,
    new_n17738_, new_n17739_, new_n17740_, new_n17741_, new_n17742_,
    new_n17743_, new_n17744_, new_n17745_, new_n17746_, new_n17747_,
    new_n17748_, new_n17749_, new_n17750_, new_n17751_, new_n17752_,
    new_n17753_, new_n17754_, new_n17755_, new_n17756_, new_n17757_,
    new_n17758_, new_n17759_, new_n17760_, new_n17761_, new_n17762_,
    new_n17763_, new_n17764_, new_n17765_, new_n17766_, new_n17767_,
    new_n17768_, new_n17769_, new_n17770_, new_n17771_, new_n17772_,
    new_n17773_, new_n17774_, new_n17775_, new_n17776_, new_n17777_,
    new_n17778_, new_n17779_, new_n17780_, new_n17781_, new_n17782_,
    new_n17783_, new_n17784_, new_n17785_, new_n17786_, new_n17787_,
    new_n17788_, new_n17789_, new_n17790_, new_n17791_, new_n17792_,
    new_n17793_, new_n17794_, new_n17795_, new_n17796_, new_n17797_,
    new_n17798_, new_n17799_, new_n17800_, new_n17801_, new_n17802_,
    new_n17803_, new_n17804_, new_n17805_, new_n17806_, new_n17807_,
    new_n17808_, new_n17809_, new_n17810_, new_n17811_, new_n17812_,
    new_n17813_, new_n17814_, new_n17815_, new_n17816_, new_n17817_,
    new_n17818_, new_n17819_, new_n17820_, new_n17821_, new_n17822_,
    new_n17823_, new_n17824_, new_n17825_, new_n17826_, new_n17827_,
    new_n17828_, new_n17829_, new_n17830_, new_n17831_, new_n17832_,
    new_n17833_, new_n17834_, new_n17835_, new_n17836_, new_n17837_,
    new_n17838_, new_n17839_, new_n17840_, new_n17841_, new_n17842_,
    new_n17843_, new_n17844_, new_n17845_, new_n17846_, new_n17847_,
    new_n17848_, new_n17849_, new_n17850_, new_n17851_, new_n17852_,
    new_n17853_, new_n17854_, new_n17855_, new_n17856_, new_n17857_,
    new_n17858_, new_n17859_, new_n17860_, new_n17861_, new_n17862_,
    new_n17863_, new_n17864_, new_n17865_, new_n17866_, new_n17867_,
    new_n17868_, new_n17869_, new_n17870_, new_n17871_, new_n17872_,
    new_n17873_, new_n17874_, new_n17875_, new_n17876_, new_n17877_,
    new_n17878_, new_n17879_, new_n17880_, new_n17881_, new_n17882_,
    new_n17883_, new_n17884_, new_n17885_, new_n17886_, new_n17887_,
    new_n17888_, new_n17889_, new_n17890_, new_n17891_, new_n17892_,
    new_n17893_, new_n17894_, new_n17895_, new_n17896_, new_n17897_,
    new_n17898_, new_n17899_, new_n17900_, new_n17901_, new_n17902_,
    new_n17903_, new_n17904_, new_n17905_, new_n17906_, new_n17907_,
    new_n17908_, new_n17909_, new_n17910_, new_n17911_, new_n17912_,
    new_n17913_, new_n17914_, new_n17915_, new_n17916_, new_n17917_,
    new_n17918_, new_n17919_, new_n17920_, new_n17921_, new_n17922_,
    new_n17923_, new_n17924_, new_n17925_, new_n17926_, new_n17927_,
    new_n17928_, new_n17929_, new_n17930_, new_n17931_, new_n17932_,
    new_n17933_, new_n17934_, new_n17935_, new_n17936_, new_n17937_,
    new_n17938_, new_n17939_, new_n17940_, new_n17941_, new_n17942_,
    new_n17943_, new_n17944_, new_n17945_, new_n17946_, new_n17947_,
    new_n17948_, new_n17949_, new_n17950_, new_n17951_, new_n17952_,
    new_n17953_, new_n17955_, new_n17956_, new_n17957_, new_n17958_,
    new_n17959_, new_n17960_, new_n17961_, new_n17962_, new_n17963_,
    new_n17964_, new_n17965_, new_n17966_, new_n17967_, new_n17968_,
    new_n17969_, new_n17970_, new_n17971_, new_n17972_, new_n17973_,
    new_n17974_, new_n17975_, new_n17976_, new_n17977_, new_n17978_,
    new_n17979_, new_n17980_, new_n17981_, new_n17982_, new_n17983_,
    new_n17984_, new_n17985_, new_n17986_, new_n17987_, new_n17988_,
    new_n17989_, new_n17990_, new_n17991_, new_n17992_, new_n17993_,
    new_n17994_, new_n17995_, new_n17996_, new_n17997_, new_n17998_,
    new_n17999_, new_n18000_, new_n18001_, new_n18002_, new_n18003_,
    new_n18004_, new_n18005_, new_n18006_, new_n18007_, new_n18008_,
    new_n18009_, new_n18010_, new_n18011_, new_n18012_, new_n18013_,
    new_n18014_, new_n18015_, new_n18016_, new_n18017_, new_n18018_,
    new_n18019_, new_n18020_, new_n18021_, new_n18022_, new_n18023_,
    new_n18024_, new_n18025_, new_n18026_, new_n18027_, new_n18028_,
    new_n18029_, new_n18030_, new_n18031_, new_n18032_, new_n18033_,
    new_n18034_, new_n18035_, new_n18036_, new_n18037_, new_n18038_,
    new_n18039_, new_n18040_, new_n18041_, new_n18042_, new_n18043_,
    new_n18044_, new_n18045_, new_n18046_, new_n18047_, new_n18048_,
    new_n18049_, new_n18050_, new_n18051_, new_n18052_, new_n18053_,
    new_n18054_, new_n18055_, new_n18056_, new_n18057_, new_n18058_,
    new_n18059_, new_n18060_, new_n18061_, new_n18062_, new_n18063_,
    new_n18064_, new_n18065_, new_n18066_, new_n18067_, new_n18068_,
    new_n18069_, new_n18070_, new_n18071_, new_n18072_, new_n18073_,
    new_n18074_, new_n18075_, new_n18076_, new_n18077_, new_n18078_,
    new_n18079_, new_n18080_, new_n18081_, new_n18082_, new_n18083_,
    new_n18084_, new_n18085_, new_n18086_, new_n18087_, new_n18088_,
    new_n18089_, new_n18090_, new_n18091_, new_n18092_, new_n18093_,
    new_n18094_, new_n18095_, new_n18096_, new_n18097_, new_n18098_,
    new_n18099_, new_n18100_, new_n18101_, new_n18102_, new_n18103_,
    new_n18104_, new_n18105_, new_n18106_, new_n18107_, new_n18108_,
    new_n18109_, new_n18110_, new_n18111_, new_n18112_, new_n18113_,
    new_n18114_, new_n18115_, new_n18116_, new_n18117_, new_n18118_,
    new_n18119_, new_n18120_, new_n18121_, new_n18122_, new_n18123_,
    new_n18124_, new_n18125_, new_n18126_, new_n18127_, new_n18128_,
    new_n18129_, new_n18130_, new_n18131_, new_n18132_, new_n18133_,
    new_n18134_, new_n18135_, new_n18136_, new_n18137_, new_n18138_,
    new_n18139_, new_n18140_, new_n18141_, new_n18142_, new_n18143_,
    new_n18144_, new_n18145_, new_n18146_, new_n18147_, new_n18148_,
    new_n18149_, new_n18150_, new_n18151_, new_n18152_, new_n18153_,
    new_n18154_, new_n18155_, new_n18156_, new_n18157_, new_n18158_,
    new_n18159_, new_n18160_, new_n18161_, new_n18162_, new_n18163_,
    new_n18164_, new_n18165_, new_n18166_, new_n18167_, new_n18168_,
    new_n18169_, new_n18170_, new_n18171_, new_n18172_, new_n18173_,
    new_n18174_, new_n18175_, new_n18176_, new_n18177_, new_n18178_,
    new_n18179_, new_n18180_, new_n18181_, new_n18182_, new_n18183_,
    new_n18184_, new_n18185_, new_n18186_, new_n18187_, new_n18188_,
    new_n18189_, new_n18190_, new_n18191_, new_n18192_, new_n18193_,
    new_n18194_, new_n18195_, new_n18196_, new_n18197_, new_n18198_,
    new_n18199_, new_n18200_, new_n18201_, new_n18202_, new_n18203_,
    new_n18204_, new_n18205_, new_n18206_, new_n18207_, new_n18208_,
    new_n18209_, new_n18210_, new_n18211_, new_n18212_, new_n18213_,
    new_n18214_, new_n18215_, new_n18216_, new_n18217_, new_n18218_,
    new_n18219_, new_n18220_, new_n18221_, new_n18222_, new_n18223_,
    new_n18224_, new_n18225_, new_n18226_, new_n18227_, new_n18228_,
    new_n18229_, new_n18230_, new_n18231_, new_n18232_, new_n18233_,
    new_n18234_, new_n18235_, new_n18236_, new_n18237_, new_n18238_,
    new_n18239_, new_n18240_, new_n18241_, new_n18242_, new_n18243_,
    new_n18244_, new_n18245_, new_n18246_, new_n18247_, new_n18248_,
    new_n18249_, new_n18250_, new_n18251_, new_n18252_, new_n18253_,
    new_n18254_, new_n18255_, new_n18256_, new_n18257_, new_n18258_,
    new_n18259_, new_n18260_, new_n18261_, new_n18262_, new_n18263_,
    new_n18264_, new_n18265_, new_n18266_, new_n18267_, new_n18268_,
    new_n18269_, new_n18270_, new_n18271_, new_n18272_, new_n18273_,
    new_n18274_, new_n18275_, new_n18276_, new_n18277_, new_n18278_,
    new_n18279_, new_n18280_, new_n18281_, new_n18282_, new_n18283_,
    new_n18284_, new_n18285_, new_n18286_, new_n18287_, new_n18288_,
    new_n18289_, new_n18290_, new_n18291_, new_n18292_, new_n18293_,
    new_n18294_, new_n18295_, new_n18296_, new_n18297_, new_n18298_,
    new_n18299_, new_n18300_, new_n18301_, new_n18302_, new_n18303_,
    new_n18304_, new_n18305_, new_n18306_, new_n18307_, new_n18308_,
    new_n18309_, new_n18310_, new_n18311_, new_n18312_, new_n18313_,
    new_n18314_, new_n18315_, new_n18316_, new_n18317_, new_n18318_,
    new_n18319_, new_n18320_, new_n18321_, new_n18322_, new_n18323_,
    new_n18324_, new_n18325_, new_n18326_, new_n18327_, new_n18328_,
    new_n18329_, new_n18330_, new_n18331_, new_n18332_, new_n18333_,
    new_n18334_, new_n18335_, new_n18336_, new_n18337_, new_n18338_,
    new_n18339_, new_n18340_, new_n18341_, new_n18342_, new_n18343_,
    new_n18344_, new_n18345_, new_n18346_, new_n18347_, new_n18348_,
    new_n18349_, new_n18350_, new_n18351_, new_n18352_, new_n18353_,
    new_n18354_, new_n18355_, new_n18356_, new_n18357_, new_n18358_,
    new_n18359_, new_n18360_, new_n18361_, new_n18362_, new_n18363_,
    new_n18364_, new_n18365_, new_n18366_, new_n18367_, new_n18368_,
    new_n18369_, new_n18370_, new_n18371_, new_n18372_, new_n18373_,
    new_n18374_, new_n18375_, new_n18376_, new_n18377_, new_n18378_,
    new_n18379_, new_n18380_, new_n18381_, new_n18382_, new_n18383_,
    new_n18384_, new_n18385_, new_n18386_, new_n18387_, new_n18388_,
    new_n18389_, new_n18390_, new_n18391_, new_n18392_, new_n18393_,
    new_n18394_, new_n18395_, new_n18396_, new_n18397_, new_n18398_,
    new_n18399_, new_n18400_, new_n18401_, new_n18402_, new_n18403_,
    new_n18404_, new_n18405_, new_n18406_, new_n18407_, new_n18408_,
    new_n18409_, new_n18410_, new_n18411_, new_n18412_, new_n18413_,
    new_n18414_, new_n18415_, new_n18416_, new_n18417_, new_n18418_,
    new_n18419_, new_n18420_, new_n18421_, new_n18422_, new_n18423_,
    new_n18424_, new_n18425_, new_n18426_, new_n18427_, new_n18428_,
    new_n18429_, new_n18430_, new_n18431_, new_n18432_, new_n18433_,
    new_n18434_, new_n18435_, new_n18436_, new_n18437_, new_n18438_,
    new_n18439_, new_n18440_, new_n18441_, new_n18442_, new_n18443_,
    new_n18444_, new_n18445_, new_n18446_, new_n18447_, new_n18448_,
    new_n18449_, new_n18450_, new_n18451_, new_n18452_, new_n18453_,
    new_n18454_, new_n18455_, new_n18456_, new_n18457_, new_n18458_,
    new_n18459_, new_n18460_, new_n18461_, new_n18462_, new_n18463_,
    new_n18464_, new_n18465_, new_n18466_, new_n18467_, new_n18468_,
    new_n18469_, new_n18470_, new_n18471_, new_n18472_, new_n18473_,
    new_n18474_, new_n18475_, new_n18476_, new_n18477_, new_n18478_,
    new_n18479_, new_n18480_, new_n18481_, new_n18482_, new_n18483_,
    new_n18484_, new_n18485_, new_n18486_, new_n18487_, new_n18488_,
    new_n18489_, new_n18490_, new_n18491_, new_n18492_, new_n18493_,
    new_n18494_, new_n18495_, new_n18496_, new_n18497_, new_n18498_,
    new_n18499_, new_n18500_, new_n18501_, new_n18502_, new_n18503_,
    new_n18504_, new_n18505_, new_n18506_, new_n18507_, new_n18508_,
    new_n18509_, new_n18510_, new_n18511_, new_n18512_, new_n18513_,
    new_n18514_, new_n18515_, new_n18516_, new_n18517_, new_n18518_,
    new_n18519_, new_n18520_, new_n18521_, new_n18522_, new_n18523_,
    new_n18524_, new_n18525_, new_n18526_, new_n18527_, new_n18528_,
    new_n18529_, new_n18530_, new_n18531_, new_n18532_, new_n18533_,
    new_n18534_, new_n18535_, new_n18536_, new_n18537_, new_n18538_,
    new_n18539_, new_n18540_, new_n18541_, new_n18542_, new_n18543_,
    new_n18544_, new_n18545_, new_n18546_, new_n18547_, new_n18548_,
    new_n18549_, new_n18550_, new_n18551_, new_n18552_, new_n18553_,
    new_n18554_, new_n18555_, new_n18556_, new_n18557_, new_n18558_,
    new_n18559_, new_n18560_, new_n18561_, new_n18562_, new_n18563_,
    new_n18564_, new_n18565_, new_n18566_, new_n18567_, new_n18568_,
    new_n18569_, new_n18570_, new_n18571_, new_n18572_, new_n18573_,
    new_n18574_, new_n18575_, new_n18576_, new_n18577_, new_n18578_,
    new_n18579_, new_n18580_, new_n18581_, new_n18582_, new_n18583_,
    new_n18584_, new_n18585_, new_n18586_, new_n18587_, new_n18588_,
    new_n18589_, new_n18590_, new_n18591_, new_n18593_, new_n18594_,
    new_n18595_, new_n18596_, new_n18597_, new_n18598_, new_n18599_,
    new_n18600_, new_n18601_, new_n18602_, new_n18603_, new_n18604_,
    new_n18605_, new_n18606_, new_n18607_, new_n18608_, new_n18609_,
    new_n18610_, new_n18611_, new_n18612_, new_n18613_, new_n18614_,
    new_n18615_, new_n18616_, new_n18617_, new_n18618_, new_n18619_,
    new_n18620_, new_n18621_, new_n18622_, new_n18623_, new_n18624_,
    new_n18625_, new_n18626_, new_n18627_, new_n18628_, new_n18629_,
    new_n18630_, new_n18631_, new_n18632_, new_n18633_, new_n18634_,
    new_n18635_, new_n18636_, new_n18637_, new_n18638_, new_n18639_,
    new_n18640_, new_n18641_, new_n18642_, new_n18643_, new_n18644_,
    new_n18645_, new_n18646_, new_n18647_, new_n18648_, new_n18649_,
    new_n18650_, new_n18651_, new_n18652_, new_n18653_, new_n18654_,
    new_n18655_, new_n18656_, new_n18657_, new_n18658_, new_n18659_,
    new_n18660_, new_n18661_, new_n18662_, new_n18663_, new_n18664_,
    new_n18665_, new_n18666_, new_n18667_, new_n18668_, new_n18669_,
    new_n18670_, new_n18671_, new_n18672_, new_n18673_, new_n18674_,
    new_n18675_, new_n18676_, new_n18677_, new_n18678_, new_n18679_,
    new_n18680_, new_n18681_, new_n18682_, new_n18683_, new_n18684_,
    new_n18685_, new_n18686_, new_n18687_, new_n18688_, new_n18689_,
    new_n18690_, new_n18691_, new_n18692_, new_n18693_, new_n18694_,
    new_n18695_, new_n18696_, new_n18697_, new_n18698_, new_n18699_,
    new_n18700_, new_n18701_, new_n18702_, new_n18703_, new_n18704_,
    new_n18705_, new_n18706_, new_n18707_, new_n18708_, new_n18709_,
    new_n18710_, new_n18711_, new_n18712_, new_n18713_, new_n18714_,
    new_n18715_, new_n18716_, new_n18717_, new_n18718_, new_n18719_,
    new_n18720_, new_n18721_, new_n18722_, new_n18723_, new_n18724_,
    new_n18725_, new_n18726_, new_n18727_, new_n18728_, new_n18729_,
    new_n18730_, new_n18731_, new_n18732_, new_n18733_, new_n18734_,
    new_n18735_, new_n18736_, new_n18737_, new_n18738_, new_n18739_,
    new_n18740_, new_n18741_, new_n18742_, new_n18743_, new_n18744_,
    new_n18745_, new_n18746_, new_n18747_, new_n18748_, new_n18749_,
    new_n18750_, new_n18751_, new_n18752_, new_n18753_, new_n18754_,
    new_n18755_, new_n18756_, new_n18757_, new_n18758_, new_n18759_,
    new_n18760_, new_n18761_, new_n18762_, new_n18763_, new_n18764_,
    new_n18765_, new_n18766_, new_n18767_, new_n18768_, new_n18769_,
    new_n18770_, new_n18771_, new_n18772_, new_n18773_, new_n18774_,
    new_n18775_, new_n18776_, new_n18777_, new_n18778_, new_n18779_,
    new_n18780_, new_n18781_, new_n18782_, new_n18783_, new_n18784_,
    new_n18785_, new_n18786_, new_n18787_, new_n18788_, new_n18789_,
    new_n18790_, new_n18791_, new_n18792_, new_n18793_, new_n18794_,
    new_n18795_, new_n18796_, new_n18797_, new_n18798_, new_n18799_,
    new_n18800_, new_n18801_, new_n18802_, new_n18803_, new_n18804_,
    new_n18805_, new_n18806_, new_n18807_, new_n18808_, new_n18809_,
    new_n18810_, new_n18811_, new_n18812_, new_n18813_, new_n18814_,
    new_n18815_, new_n18816_, new_n18817_, new_n18818_, new_n18819_,
    new_n18820_, new_n18821_, new_n18822_, new_n18823_, new_n18824_,
    new_n18825_, new_n18826_, new_n18827_, new_n18828_, new_n18829_,
    new_n18830_, new_n18831_, new_n18832_, new_n18833_, new_n18834_,
    new_n18835_, new_n18836_, new_n18837_, new_n18838_, new_n18839_,
    new_n18840_, new_n18841_, new_n18842_, new_n18843_, new_n18844_,
    new_n18845_, new_n18846_, new_n18847_, new_n18848_, new_n18849_,
    new_n18850_, new_n18851_, new_n18852_, new_n18853_, new_n18854_,
    new_n18855_, new_n18856_, new_n18857_, new_n18858_, new_n18859_,
    new_n18860_, new_n18861_, new_n18862_, new_n18863_, new_n18864_,
    new_n18865_, new_n18866_, new_n18867_, new_n18868_, new_n18869_,
    new_n18870_, new_n18871_, new_n18872_, new_n18873_, new_n18874_,
    new_n18875_, new_n18876_, new_n18877_, new_n18878_, new_n18879_,
    new_n18880_, new_n18881_, new_n18882_, new_n18883_, new_n18884_,
    new_n18885_, new_n18886_, new_n18887_, new_n18888_, new_n18889_,
    new_n18890_, new_n18891_, new_n18892_, new_n18893_, new_n18894_,
    new_n18895_, new_n18896_, new_n18897_, new_n18898_, new_n18899_,
    new_n18900_, new_n18901_, new_n18902_, new_n18903_, new_n18904_,
    new_n18905_, new_n18906_, new_n18907_, new_n18908_, new_n18909_,
    new_n18910_, new_n18911_, new_n18912_, new_n18913_, new_n18914_,
    new_n18915_, new_n18916_, new_n18917_, new_n18918_, new_n18919_,
    new_n18920_, new_n18921_, new_n18922_, new_n18923_, new_n18924_,
    new_n18925_, new_n18926_, new_n18927_, new_n18928_, new_n18929_,
    new_n18930_, new_n18931_, new_n18932_, new_n18933_, new_n18934_,
    new_n18935_, new_n18936_, new_n18937_, new_n18938_, new_n18939_,
    new_n18940_, new_n18941_, new_n18942_, new_n18943_, new_n18944_,
    new_n18945_, new_n18946_, new_n18947_, new_n18948_, new_n18949_,
    new_n18950_, new_n18951_, new_n18952_, new_n18953_, new_n18954_,
    new_n18955_, new_n18956_, new_n18957_, new_n18958_, new_n18959_,
    new_n18960_, new_n18961_, new_n18962_, new_n18963_, new_n18964_,
    new_n18965_, new_n18966_, new_n18967_, new_n18968_, new_n18969_,
    new_n18970_, new_n18971_, new_n18972_, new_n18973_, new_n18974_,
    new_n18975_, new_n18976_, new_n18977_, new_n18978_, new_n18979_,
    new_n18980_, new_n18981_, new_n18982_, new_n18983_, new_n18984_,
    new_n18985_, new_n18986_, new_n18987_, new_n18988_, new_n18989_,
    new_n18990_, new_n18991_, new_n18992_, new_n18993_, new_n18994_,
    new_n18995_, new_n18996_, new_n18997_, new_n18998_, new_n18999_,
    new_n19000_, new_n19001_, new_n19002_, new_n19003_, new_n19004_,
    new_n19005_, new_n19006_, new_n19007_, new_n19008_, new_n19009_,
    new_n19010_, new_n19011_, new_n19012_, new_n19013_, new_n19014_,
    new_n19015_, new_n19016_, new_n19017_, new_n19018_, new_n19019_,
    new_n19020_, new_n19021_, new_n19022_, new_n19023_, new_n19024_,
    new_n19025_, new_n19026_, new_n19027_, new_n19028_, new_n19029_,
    new_n19030_, new_n19031_, new_n19032_, new_n19033_, new_n19034_,
    new_n19035_, new_n19036_, new_n19037_, new_n19038_, new_n19039_,
    new_n19040_, new_n19041_, new_n19042_, new_n19043_, new_n19044_,
    new_n19045_, new_n19046_, new_n19047_, new_n19048_, new_n19049_,
    new_n19050_, new_n19051_, new_n19052_, new_n19053_, new_n19054_,
    new_n19055_, new_n19056_, new_n19057_, new_n19058_, new_n19059_,
    new_n19060_, new_n19061_, new_n19062_, new_n19063_, new_n19064_,
    new_n19065_, new_n19066_, new_n19067_, new_n19068_, new_n19069_,
    new_n19070_, new_n19071_, new_n19072_, new_n19073_, new_n19074_,
    new_n19075_, new_n19076_, new_n19077_, new_n19078_, new_n19079_,
    new_n19080_, new_n19081_, new_n19082_, new_n19083_, new_n19084_,
    new_n19085_, new_n19086_, new_n19087_, new_n19088_, new_n19089_,
    new_n19090_, new_n19091_, new_n19092_, new_n19093_, new_n19094_,
    new_n19095_, new_n19096_, new_n19097_, new_n19098_, new_n19099_,
    new_n19100_, new_n19101_, new_n19102_, new_n19103_, new_n19104_,
    new_n19105_, new_n19106_, new_n19107_, new_n19108_, new_n19109_,
    new_n19110_, new_n19111_, new_n19112_, new_n19113_, new_n19114_,
    new_n19115_, new_n19116_, new_n19117_, new_n19118_, new_n19119_,
    new_n19120_, new_n19121_, new_n19122_, new_n19123_, new_n19124_,
    new_n19125_, new_n19126_, new_n19127_, new_n19128_, new_n19129_,
    new_n19130_, new_n19131_, new_n19132_, new_n19133_, new_n19134_,
    new_n19135_, new_n19136_, new_n19137_, new_n19138_, new_n19139_,
    new_n19140_, new_n19141_, new_n19142_, new_n19143_, new_n19144_,
    new_n19145_, new_n19146_, new_n19147_, new_n19148_, new_n19149_,
    new_n19150_, new_n19151_, new_n19152_, new_n19153_, new_n19154_,
    new_n19155_, new_n19156_, new_n19157_, new_n19158_, new_n19159_,
    new_n19160_, new_n19161_, new_n19162_, new_n19163_, new_n19164_,
    new_n19165_, new_n19166_, new_n19167_, new_n19168_, new_n19169_,
    new_n19170_, new_n19171_, new_n19172_, new_n19173_, new_n19174_,
    new_n19175_, new_n19176_, new_n19177_, new_n19178_, new_n19179_,
    new_n19180_, new_n19181_, new_n19182_, new_n19183_, new_n19184_,
    new_n19185_, new_n19186_, new_n19187_, new_n19188_, new_n19189_,
    new_n19190_, new_n19191_, new_n19192_, new_n19193_, new_n19194_,
    new_n19195_, new_n19196_, new_n19197_, new_n19198_, new_n19199_,
    new_n19200_, new_n19201_, new_n19202_, new_n19203_, new_n19204_,
    new_n19205_, new_n19206_, new_n19207_, new_n19208_, new_n19209_,
    new_n19210_, new_n19211_, new_n19212_, new_n19213_, new_n19214_,
    new_n19215_, new_n19216_, new_n19217_, new_n19218_, new_n19219_,
    new_n19220_, new_n19221_, new_n19222_, new_n19223_, new_n19224_,
    new_n19225_, new_n19226_, new_n19227_, new_n19228_, new_n19229_,
    new_n19230_, new_n19231_, new_n19232_, new_n19233_, new_n19234_,
    new_n19235_, new_n19236_, new_n19237_, new_n19238_, new_n19239_,
    new_n19240_, new_n19241_, new_n19242_, new_n19243_, new_n19244_,
    new_n19245_, new_n19246_, new_n19247_, new_n19248_, new_n19249_,
    new_n19250_, new_n19251_, new_n19252_, new_n19253_, new_n19254_,
    new_n19255_, new_n19256_, new_n19257_, new_n19258_, new_n19259_,
    new_n19260_, new_n19261_, new_n19262_, new_n19263_, new_n19264_,
    new_n19265_, new_n19266_, new_n19267_, new_n19268_, new_n19269_,
    new_n19270_, new_n19271_, new_n19272_, new_n19273_, new_n19274_,
    new_n19275_, new_n19276_, new_n19277_, new_n19278_, new_n19279_,
    new_n19280_, new_n19281_, new_n19282_, new_n19283_, new_n19284_,
    new_n19285_, new_n19286_, new_n19287_, new_n19288_, new_n19289_,
    new_n19290_, new_n19291_, new_n19292_, new_n19293_, new_n19294_,
    new_n19295_, new_n19296_, new_n19297_, new_n19298_, new_n19299_,
    new_n19300_, new_n19301_, new_n19302_, new_n19303_, new_n19304_,
    new_n19305_, new_n19306_, new_n19307_, new_n19308_, new_n19309_,
    new_n19310_, new_n19311_, new_n19312_, new_n19313_, new_n19314_,
    new_n19315_, new_n19316_, new_n19317_, new_n19318_, new_n19319_,
    new_n19320_, new_n19321_, new_n19322_, new_n19323_, new_n19324_,
    new_n19325_, new_n19326_, new_n19327_, new_n19328_, new_n19329_,
    new_n19330_, new_n19331_, new_n19332_, new_n19333_, new_n19334_,
    new_n19335_, new_n19336_, new_n19337_, new_n19338_, new_n19339_,
    new_n19340_, new_n19341_, new_n19342_, new_n19343_, new_n19344_,
    new_n19345_, new_n19347_, new_n19348_, new_n19349_, new_n19350_,
    new_n19351_, new_n19352_, new_n19353_, new_n19354_, new_n19355_,
    new_n19356_, new_n19357_, new_n19358_, new_n19359_, new_n19360_,
    new_n19361_, new_n19362_, new_n19363_, new_n19364_, new_n19365_,
    new_n19366_, new_n19367_, new_n19368_, new_n19369_, new_n19370_,
    new_n19371_, new_n19372_, new_n19373_, new_n19374_, new_n19375_,
    new_n19376_, new_n19377_, new_n19378_, new_n19379_, new_n19380_,
    new_n19381_, new_n19382_, new_n19383_, new_n19384_, new_n19385_,
    new_n19386_, new_n19387_, new_n19388_, new_n19389_, new_n19390_,
    new_n19391_, new_n19392_, new_n19393_, new_n19394_, new_n19395_,
    new_n19396_, new_n19397_, new_n19398_, new_n19399_, new_n19400_,
    new_n19401_, new_n19402_, new_n19403_, new_n19404_, new_n19405_,
    new_n19406_, new_n19407_, new_n19408_, new_n19409_, new_n19410_,
    new_n19411_, new_n19412_, new_n19413_, new_n19414_, new_n19415_,
    new_n19416_, new_n19417_, new_n19418_, new_n19419_, new_n19420_,
    new_n19421_, new_n19422_, new_n19423_, new_n19424_, new_n19425_,
    new_n19426_, new_n19427_, new_n19428_, new_n19429_, new_n19430_,
    new_n19431_, new_n19432_, new_n19433_, new_n19434_, new_n19435_,
    new_n19436_, new_n19437_, new_n19438_, new_n19439_, new_n19440_,
    new_n19441_, new_n19442_, new_n19443_, new_n19444_, new_n19445_,
    new_n19446_, new_n19447_, new_n19448_, new_n19449_, new_n19450_,
    new_n19451_, new_n19452_, new_n19453_, new_n19454_, new_n19455_,
    new_n19456_, new_n19457_, new_n19458_, new_n19459_, new_n19460_,
    new_n19461_, new_n19462_, new_n19463_, new_n19464_, new_n19465_,
    new_n19466_, new_n19467_, new_n19468_, new_n19469_, new_n19470_,
    new_n19471_, new_n19472_, new_n19473_, new_n19474_, new_n19475_,
    new_n19476_, new_n19477_, new_n19478_, new_n19479_, new_n19480_,
    new_n19481_, new_n19482_, new_n19483_, new_n19484_, new_n19485_,
    new_n19486_, new_n19487_, new_n19488_, new_n19489_, new_n19490_,
    new_n19491_, new_n19492_, new_n19493_, new_n19494_, new_n19495_,
    new_n19496_, new_n19497_, new_n19498_, new_n19499_, new_n19500_,
    new_n19501_, new_n19502_, new_n19503_, new_n19504_, new_n19505_,
    new_n19506_, new_n19507_, new_n19508_, new_n19509_, new_n19510_,
    new_n19511_, new_n19512_, new_n19513_, new_n19514_, new_n19515_,
    new_n19516_, new_n19517_, new_n19518_, new_n19519_, new_n19520_,
    new_n19521_, new_n19522_, new_n19523_, new_n19524_, new_n19525_,
    new_n19526_, new_n19527_, new_n19528_, new_n19529_, new_n19530_,
    new_n19531_, new_n19532_, new_n19533_, new_n19534_, new_n19535_,
    new_n19536_, new_n19537_, new_n19538_, new_n19539_, new_n19540_,
    new_n19541_, new_n19542_, new_n19543_, new_n19544_, new_n19545_,
    new_n19546_, new_n19547_, new_n19548_, new_n19549_, new_n19550_,
    new_n19551_, new_n19552_, new_n19553_, new_n19554_, new_n19555_,
    new_n19556_, new_n19557_, new_n19558_, new_n19559_, new_n19560_,
    new_n19561_, new_n19562_, new_n19563_, new_n19564_, new_n19565_,
    new_n19566_, new_n19567_, new_n19568_, new_n19569_, new_n19570_,
    new_n19571_, new_n19572_, new_n19573_, new_n19574_, new_n19575_,
    new_n19576_, new_n19577_, new_n19578_, new_n19579_, new_n19580_,
    new_n19581_, new_n19582_, new_n19583_, new_n19584_, new_n19585_,
    new_n19586_, new_n19587_, new_n19588_, new_n19589_, new_n19590_,
    new_n19591_, new_n19592_, new_n19593_, new_n19594_, new_n19595_,
    new_n19596_, new_n19597_, new_n19598_, new_n19599_, new_n19600_,
    new_n19601_, new_n19602_, new_n19603_, new_n19604_, new_n19605_,
    new_n19606_, new_n19607_, new_n19608_, new_n19609_, new_n19610_,
    new_n19611_, new_n19612_, new_n19613_, new_n19614_, new_n19615_,
    new_n19616_, new_n19617_, new_n19618_, new_n19619_, new_n19620_,
    new_n19621_, new_n19622_, new_n19623_, new_n19624_, new_n19625_,
    new_n19626_, new_n19627_, new_n19628_, new_n19629_, new_n19630_,
    new_n19631_, new_n19632_, new_n19633_, new_n19634_, new_n19635_,
    new_n19636_, new_n19637_, new_n19638_, new_n19639_, new_n19640_,
    new_n19641_, new_n19642_, new_n19643_, new_n19644_, new_n19645_,
    new_n19646_, new_n19647_, new_n19648_, new_n19649_, new_n19650_,
    new_n19651_, new_n19652_, new_n19653_, new_n19654_, new_n19655_,
    new_n19656_, new_n19657_, new_n19658_, new_n19659_, new_n19660_,
    new_n19661_, new_n19662_, new_n19663_, new_n19664_, new_n19665_,
    new_n19666_, new_n19667_, new_n19668_, new_n19669_, new_n19670_,
    new_n19671_, new_n19672_, new_n19673_, new_n19674_, new_n19675_,
    new_n19676_, new_n19677_, new_n19678_, new_n19679_, new_n19680_,
    new_n19681_, new_n19682_, new_n19683_, new_n19684_, new_n19685_,
    new_n19686_, new_n19687_, new_n19688_, new_n19689_, new_n19690_,
    new_n19691_, new_n19692_, new_n19693_, new_n19694_, new_n19695_,
    new_n19696_, new_n19697_, new_n19698_, new_n19699_, new_n19700_,
    new_n19701_, new_n19702_, new_n19703_, new_n19704_, new_n19705_,
    new_n19706_, new_n19707_, new_n19708_, new_n19709_, new_n19710_,
    new_n19711_, new_n19712_, new_n19713_, new_n19714_, new_n19715_,
    new_n19716_, new_n19717_, new_n19718_, new_n19719_, new_n19720_,
    new_n19721_, new_n19722_, new_n19723_, new_n19724_, new_n19725_,
    new_n19726_, new_n19727_, new_n19728_, new_n19729_, new_n19730_,
    new_n19731_, new_n19732_, new_n19733_, new_n19734_, new_n19735_,
    new_n19736_, new_n19737_, new_n19738_, new_n19739_, new_n19740_,
    new_n19741_, new_n19742_, new_n19743_, new_n19744_, new_n19745_,
    new_n19746_, new_n19747_, new_n19748_, new_n19749_, new_n19750_,
    new_n19751_, new_n19752_, new_n19753_, new_n19754_, new_n19755_,
    new_n19756_, new_n19757_, new_n19758_, new_n19759_, new_n19760_,
    new_n19761_, new_n19762_, new_n19763_, new_n19764_, new_n19765_,
    new_n19766_, new_n19767_, new_n19768_, new_n19769_, new_n19770_,
    new_n19771_, new_n19772_, new_n19773_, new_n19774_, new_n19775_,
    new_n19776_, new_n19777_, new_n19778_, new_n19779_, new_n19780_,
    new_n19781_, new_n19782_, new_n19783_, new_n19784_, new_n19785_,
    new_n19786_, new_n19787_, new_n19788_, new_n19789_, new_n19790_,
    new_n19791_, new_n19792_, new_n19793_, new_n19794_, new_n19795_,
    new_n19796_, new_n19797_, new_n19798_, new_n19799_, new_n19800_,
    new_n19801_, new_n19802_, new_n19803_, new_n19804_, new_n19805_,
    new_n19806_, new_n19807_, new_n19808_, new_n19809_, new_n19810_,
    new_n19811_, new_n19812_, new_n19813_, new_n19814_, new_n19815_,
    new_n19816_, new_n19817_, new_n19818_, new_n19819_, new_n19820_,
    new_n19821_, new_n19822_, new_n19823_, new_n19824_, new_n19825_,
    new_n19826_, new_n19827_, new_n19828_, new_n19829_, new_n19830_,
    new_n19831_, new_n19832_, new_n19833_, new_n19834_, new_n19835_,
    new_n19836_, new_n19837_, new_n19838_, new_n19839_, new_n19840_,
    new_n19841_, new_n19842_, new_n19843_, new_n19844_, new_n19845_,
    new_n19846_, new_n19847_, new_n19848_, new_n19849_, new_n19850_,
    new_n19851_, new_n19852_, new_n19853_, new_n19854_, new_n19855_,
    new_n19856_, new_n19857_, new_n19858_, new_n19859_, new_n19860_,
    new_n19861_, new_n19862_, new_n19863_, new_n19864_, new_n19865_,
    new_n19866_, new_n19867_, new_n19868_, new_n19869_, new_n19870_,
    new_n19871_, new_n19872_, new_n19873_, new_n19874_, new_n19875_,
    new_n19876_, new_n19877_, new_n19878_, new_n19879_, new_n19880_,
    new_n19881_, new_n19882_, new_n19883_, new_n19884_, new_n19885_,
    new_n19886_, new_n19887_, new_n19888_, new_n19889_, new_n19890_,
    new_n19891_, new_n19892_, new_n19893_, new_n19894_, new_n19895_,
    new_n19896_, new_n19897_, new_n19898_, new_n19899_, new_n19900_,
    new_n19901_, new_n19902_, new_n19903_, new_n19904_, new_n19905_,
    new_n19906_, new_n19907_, new_n19908_, new_n19909_, new_n19910_,
    new_n19911_, new_n19912_, new_n19913_, new_n19914_, new_n19915_,
    new_n19916_, new_n19917_, new_n19918_, new_n19919_, new_n19920_,
    new_n19921_, new_n19922_, new_n19923_, new_n19924_, new_n19925_,
    new_n19926_, new_n19927_, new_n19928_, new_n19929_, new_n19930_,
    new_n19931_, new_n19932_, new_n19933_, new_n19934_, new_n19935_,
    new_n19936_, new_n19937_, new_n19938_, new_n19939_, new_n19940_,
    new_n19941_, new_n19942_, new_n19943_, new_n19944_, new_n19945_,
    new_n19946_, new_n19947_, new_n19948_, new_n19949_, new_n19950_,
    new_n19951_, new_n19952_, new_n19953_, new_n19954_, new_n19955_,
    new_n19956_, new_n19957_, new_n19958_, new_n19959_, new_n19960_,
    new_n19961_, new_n19962_, new_n19963_, new_n19964_, new_n19965_,
    new_n19966_, new_n19967_, new_n19968_, new_n19969_, new_n19970_,
    new_n19971_, new_n19972_, new_n19973_, new_n19974_, new_n19975_,
    new_n19976_, new_n19977_, new_n19978_, new_n19979_, new_n19980_,
    new_n19981_, new_n19982_, new_n19983_, new_n19984_, new_n19985_,
    new_n19986_, new_n19988_, new_n19989_, new_n19990_, new_n19991_,
    new_n19992_, new_n19993_, new_n19994_, new_n19995_, new_n19996_,
    new_n19997_, new_n19998_, new_n19999_, new_n20000_, new_n20001_,
    new_n20002_, new_n20003_, new_n20004_, new_n20005_, new_n20006_,
    new_n20007_, new_n20008_, new_n20009_, new_n20010_, new_n20011_,
    new_n20012_, new_n20013_, new_n20014_, new_n20015_, new_n20016_,
    new_n20017_, new_n20018_, new_n20019_, new_n20020_, new_n20021_,
    new_n20022_, new_n20023_, new_n20024_, new_n20025_, new_n20026_,
    new_n20027_, new_n20028_, new_n20029_, new_n20030_, new_n20031_,
    new_n20032_, new_n20033_, new_n20034_, new_n20035_, new_n20036_,
    new_n20037_, new_n20038_, new_n20039_, new_n20040_, new_n20041_,
    new_n20042_, new_n20043_, new_n20044_, new_n20045_, new_n20046_,
    new_n20047_, new_n20048_, new_n20049_, new_n20050_, new_n20051_,
    new_n20052_, new_n20053_, new_n20054_, new_n20055_, new_n20056_,
    new_n20057_, new_n20058_, new_n20059_, new_n20060_, new_n20061_,
    new_n20062_, new_n20063_, new_n20064_, new_n20065_, new_n20066_,
    new_n20067_, new_n20068_, new_n20069_, new_n20070_, new_n20071_,
    new_n20072_, new_n20073_, new_n20074_, new_n20075_, new_n20076_,
    new_n20077_, new_n20078_, new_n20079_, new_n20080_, new_n20081_,
    new_n20082_, new_n20083_, new_n20084_, new_n20085_, new_n20086_,
    new_n20087_, new_n20088_, new_n20089_, new_n20090_, new_n20091_,
    new_n20092_, new_n20093_, new_n20094_, new_n20095_, new_n20096_,
    new_n20097_, new_n20098_, new_n20099_, new_n20100_, new_n20101_,
    new_n20102_, new_n20103_, new_n20104_, new_n20105_, new_n20106_,
    new_n20107_, new_n20108_, new_n20109_, new_n20110_, new_n20111_,
    new_n20112_, new_n20113_, new_n20114_, new_n20115_, new_n20116_,
    new_n20117_, new_n20118_, new_n20119_, new_n20120_, new_n20121_,
    new_n20122_, new_n20123_, new_n20124_, new_n20125_, new_n20126_,
    new_n20127_, new_n20128_, new_n20129_, new_n20130_, new_n20131_,
    new_n20132_, new_n20133_, new_n20134_, new_n20135_, new_n20136_,
    new_n20137_, new_n20138_, new_n20139_, new_n20140_, new_n20141_,
    new_n20142_, new_n20143_, new_n20144_, new_n20145_, new_n20146_,
    new_n20147_, new_n20148_, new_n20149_, new_n20150_, new_n20151_,
    new_n20152_, new_n20153_, new_n20154_, new_n20155_, new_n20156_,
    new_n20157_, new_n20158_, new_n20159_, new_n20160_, new_n20161_,
    new_n20162_, new_n20163_, new_n20164_, new_n20165_, new_n20166_,
    new_n20167_, new_n20168_, new_n20169_, new_n20170_, new_n20171_,
    new_n20172_, new_n20173_, new_n20174_, new_n20175_, new_n20176_,
    new_n20177_, new_n20178_, new_n20179_, new_n20180_, new_n20181_,
    new_n20182_, new_n20183_, new_n20184_, new_n20185_, new_n20186_,
    new_n20187_, new_n20188_, new_n20189_, new_n20190_, new_n20191_,
    new_n20192_, new_n20193_, new_n20194_, new_n20195_, new_n20196_,
    new_n20197_, new_n20198_, new_n20199_, new_n20200_, new_n20201_,
    new_n20202_, new_n20203_, new_n20204_, new_n20205_, new_n20206_,
    new_n20207_, new_n20208_, new_n20209_, new_n20210_, new_n20211_,
    new_n20212_, new_n20213_, new_n20214_, new_n20215_, new_n20216_,
    new_n20217_, new_n20218_, new_n20219_, new_n20220_, new_n20221_,
    new_n20222_, new_n20223_, new_n20224_, new_n20225_, new_n20226_,
    new_n20227_, new_n20228_, new_n20229_, new_n20230_, new_n20231_,
    new_n20232_, new_n20233_, new_n20234_, new_n20235_, new_n20236_,
    new_n20237_, new_n20238_, new_n20239_, new_n20240_, new_n20241_,
    new_n20242_, new_n20243_, new_n20244_, new_n20245_, new_n20246_,
    new_n20247_, new_n20248_, new_n20249_, new_n20250_, new_n20251_,
    new_n20252_, new_n20253_, new_n20254_, new_n20255_, new_n20256_,
    new_n20257_, new_n20258_, new_n20259_, new_n20260_, new_n20261_,
    new_n20262_, new_n20263_, new_n20264_, new_n20265_, new_n20266_,
    new_n20267_, new_n20268_, new_n20269_, new_n20270_, new_n20271_,
    new_n20272_, new_n20273_, new_n20274_, new_n20275_, new_n20276_,
    new_n20277_, new_n20278_, new_n20279_, new_n20280_, new_n20281_,
    new_n20282_, new_n20283_, new_n20284_, new_n20285_, new_n20286_,
    new_n20287_, new_n20288_, new_n20289_, new_n20290_, new_n20291_,
    new_n20292_, new_n20293_, new_n20294_, new_n20295_, new_n20296_,
    new_n20297_, new_n20298_, new_n20299_, new_n20300_, new_n20301_,
    new_n20302_, new_n20303_, new_n20304_, new_n20305_, new_n20306_,
    new_n20307_, new_n20308_, new_n20309_, new_n20310_, new_n20311_,
    new_n20312_, new_n20313_, new_n20314_, new_n20315_, new_n20316_,
    new_n20317_, new_n20318_, new_n20319_, new_n20320_, new_n20321_,
    new_n20322_, new_n20323_, new_n20324_, new_n20325_, new_n20326_,
    new_n20327_, new_n20328_, new_n20329_, new_n20330_, new_n20331_,
    new_n20332_, new_n20333_, new_n20334_, new_n20335_, new_n20336_,
    new_n20337_, new_n20338_, new_n20339_, new_n20340_, new_n20341_,
    new_n20342_, new_n20343_, new_n20344_, new_n20345_, new_n20346_,
    new_n20347_, new_n20348_, new_n20349_, new_n20350_, new_n20351_,
    new_n20352_, new_n20353_, new_n20354_, new_n20355_, new_n20356_,
    new_n20357_, new_n20358_, new_n20359_, new_n20360_, new_n20361_,
    new_n20362_, new_n20363_, new_n20364_, new_n20365_, new_n20366_,
    new_n20367_, new_n20368_, new_n20369_, new_n20370_, new_n20371_,
    new_n20372_, new_n20373_, new_n20374_, new_n20375_, new_n20376_,
    new_n20377_, new_n20378_, new_n20379_, new_n20380_, new_n20381_,
    new_n20382_, new_n20383_, new_n20384_, new_n20385_, new_n20386_,
    new_n20387_, new_n20388_, new_n20389_, new_n20390_, new_n20391_,
    new_n20392_, new_n20393_, new_n20394_, new_n20395_, new_n20396_,
    new_n20397_, new_n20398_, new_n20399_, new_n20400_, new_n20401_,
    new_n20402_, new_n20403_, new_n20404_, new_n20405_, new_n20406_,
    new_n20407_, new_n20408_, new_n20409_, new_n20410_, new_n20411_,
    new_n20412_, new_n20413_, new_n20414_, new_n20415_, new_n20416_,
    new_n20417_, new_n20418_, new_n20419_, new_n20420_, new_n20421_,
    new_n20422_, new_n20423_, new_n20424_, new_n20425_, new_n20426_,
    new_n20427_, new_n20428_, new_n20429_, new_n20430_, new_n20431_,
    new_n20432_, new_n20433_, new_n20434_, new_n20435_, new_n20436_,
    new_n20437_, new_n20438_, new_n20439_, new_n20440_, new_n20441_,
    new_n20442_, new_n20443_, new_n20444_, new_n20445_, new_n20446_,
    new_n20447_, new_n20448_, new_n20449_, new_n20450_, new_n20451_,
    new_n20452_, new_n20453_, new_n20454_, new_n20455_, new_n20456_,
    new_n20457_, new_n20458_, new_n20459_, new_n20460_, new_n20461_,
    new_n20462_, new_n20463_, new_n20464_, new_n20465_, new_n20466_,
    new_n20467_, new_n20468_, new_n20469_, new_n20470_, new_n20471_,
    new_n20472_, new_n20473_, new_n20474_, new_n20475_, new_n20476_,
    new_n20477_, new_n20478_, new_n20479_, new_n20480_, new_n20481_,
    new_n20482_, new_n20483_, new_n20484_, new_n20485_, new_n20486_,
    new_n20487_, new_n20488_, new_n20489_, new_n20490_, new_n20491_,
    new_n20492_, new_n20493_, new_n20494_, new_n20495_, new_n20496_,
    new_n20497_, new_n20498_, new_n20499_, new_n20500_, new_n20501_,
    new_n20502_, new_n20503_, new_n20504_, new_n20505_, new_n20506_,
    new_n20507_, new_n20508_, new_n20509_, new_n20510_, new_n20511_,
    new_n20512_, new_n20513_, new_n20514_, new_n20515_, new_n20516_,
    new_n20517_, new_n20518_, new_n20519_, new_n20520_, new_n20521_,
    new_n20522_, new_n20523_, new_n20524_, new_n20525_, new_n20526_,
    new_n20527_, new_n20528_, new_n20529_, new_n20530_, new_n20531_,
    new_n20532_, new_n20533_, new_n20534_, new_n20535_, new_n20536_,
    new_n20537_, new_n20538_, new_n20539_, new_n20540_, new_n20541_,
    new_n20542_, new_n20543_, new_n20544_, new_n20545_, new_n20546_,
    new_n20547_, new_n20548_, new_n20549_, new_n20550_, new_n20551_,
    new_n20552_, new_n20553_, new_n20554_, new_n20555_, new_n20556_,
    new_n20557_, new_n20558_, new_n20559_, new_n20560_, new_n20561_,
    new_n20562_, new_n20563_, new_n20564_, new_n20565_, new_n20566_,
    new_n20567_, new_n20568_, new_n20569_, new_n20570_, new_n20571_,
    new_n20572_, new_n20573_, new_n20574_, new_n20575_, new_n20576_,
    new_n20577_, new_n20578_, new_n20579_, new_n20580_, new_n20581_,
    new_n20582_, new_n20583_, new_n20584_, new_n20585_, new_n20586_,
    new_n20587_, new_n20588_, new_n20589_, new_n20590_, new_n20591_,
    new_n20592_, new_n20593_, new_n20594_, new_n20595_, new_n20596_,
    new_n20597_, new_n20598_, new_n20599_, new_n20600_, new_n20601_,
    new_n20602_, new_n20603_, new_n20604_, new_n20605_, new_n20606_,
    new_n20607_, new_n20608_, new_n20609_, new_n20610_, new_n20611_,
    new_n20612_, new_n20613_, new_n20614_, new_n20615_, new_n20616_,
    new_n20617_, new_n20618_, new_n20619_, new_n20620_, new_n20621_,
    new_n20622_, new_n20623_, new_n20624_, new_n20625_, new_n20626_,
    new_n20627_, new_n20628_, new_n20629_, new_n20630_, new_n20631_,
    new_n20632_, new_n20633_, new_n20634_, new_n20635_, new_n20636_,
    new_n20637_, new_n20638_, new_n20639_, new_n20640_, new_n20641_,
    new_n20642_, new_n20643_, new_n20644_, new_n20645_, new_n20646_,
    new_n20647_, new_n20648_, new_n20649_, new_n20650_, new_n20651_,
    new_n20652_, new_n20653_, new_n20654_, new_n20655_, new_n20656_,
    new_n20657_, new_n20658_, new_n20659_, new_n20660_, new_n20661_,
    new_n20662_, new_n20663_, new_n20664_, new_n20665_, new_n20666_,
    new_n20667_, new_n20668_, new_n20669_, new_n20670_, new_n20671_,
    new_n20672_, new_n20673_, new_n20674_, new_n20675_, new_n20676_,
    new_n20678_, new_n20679_, new_n20680_, new_n20681_, new_n20682_,
    new_n20683_, new_n20684_, new_n20685_, new_n20686_, new_n20687_,
    new_n20688_, new_n20689_, new_n20690_, new_n20691_, new_n20692_,
    new_n20693_, new_n20694_, new_n20695_, new_n20696_, new_n20697_,
    new_n20698_, new_n20699_, new_n20700_, new_n20701_, new_n20702_,
    new_n20703_, new_n20704_, new_n20705_, new_n20706_, new_n20707_,
    new_n20708_, new_n20709_, new_n20710_, new_n20711_, new_n20712_,
    new_n20713_, new_n20714_, new_n20715_, new_n20716_, new_n20717_,
    new_n20718_, new_n20719_, new_n20720_, new_n20721_, new_n20722_,
    new_n20723_, new_n20724_, new_n20725_, new_n20726_, new_n20727_,
    new_n20728_, new_n20729_, new_n20730_, new_n20731_, new_n20732_,
    new_n20733_, new_n20734_, new_n20735_, new_n20736_, new_n20737_,
    new_n20738_, new_n20739_, new_n20740_, new_n20741_, new_n20742_,
    new_n20743_, new_n20744_, new_n20745_, new_n20746_, new_n20747_,
    new_n20748_, new_n20749_, new_n20750_, new_n20751_, new_n20752_,
    new_n20753_, new_n20754_, new_n20755_, new_n20756_, new_n20757_,
    new_n20758_, new_n20759_, new_n20760_, new_n20761_, new_n20762_,
    new_n20763_, new_n20764_, new_n20765_, new_n20766_, new_n20767_,
    new_n20768_, new_n20769_, new_n20770_, new_n20771_, new_n20772_,
    new_n20773_, new_n20774_, new_n20775_, new_n20776_, new_n20777_,
    new_n20778_, new_n20779_, new_n20780_, new_n20781_, new_n20782_,
    new_n20783_, new_n20784_, new_n20785_, new_n20786_, new_n20787_,
    new_n20788_, new_n20789_, new_n20790_, new_n20791_, new_n20792_,
    new_n20793_, new_n20794_, new_n20795_, new_n20796_, new_n20797_,
    new_n20798_, new_n20799_, new_n20800_, new_n20801_, new_n20802_,
    new_n20803_, new_n20804_, new_n20805_, new_n20806_, new_n20807_,
    new_n20808_, new_n20809_, new_n20810_, new_n20811_, new_n20812_,
    new_n20813_, new_n20814_, new_n20815_, new_n20816_, new_n20817_,
    new_n20818_, new_n20819_, new_n20820_, new_n20821_, new_n20822_,
    new_n20823_, new_n20824_, new_n20825_, new_n20826_, new_n20827_,
    new_n20828_, new_n20829_, new_n20830_, new_n20831_, new_n20832_,
    new_n20833_, new_n20834_, new_n20835_, new_n20836_, new_n20837_,
    new_n20838_, new_n20839_, new_n20840_, new_n20841_, new_n20842_,
    new_n20843_, new_n20844_, new_n20845_, new_n20846_, new_n20847_,
    new_n20848_, new_n20849_, new_n20850_, new_n20851_, new_n20852_,
    new_n20853_, new_n20854_, new_n20855_, new_n20856_, new_n20857_,
    new_n20858_, new_n20859_, new_n20860_, new_n20861_, new_n20862_,
    new_n20863_, new_n20864_, new_n20865_, new_n20866_, new_n20867_,
    new_n20868_, new_n20869_, new_n20870_, new_n20871_, new_n20872_,
    new_n20873_, new_n20874_, new_n20875_, new_n20876_, new_n20877_,
    new_n20878_, new_n20879_, new_n20880_, new_n20881_, new_n20882_,
    new_n20883_, new_n20884_, new_n20885_, new_n20886_, new_n20887_,
    new_n20888_, new_n20889_, new_n20890_, new_n20891_, new_n20892_,
    new_n20893_, new_n20894_, new_n20895_, new_n20896_, new_n20897_,
    new_n20898_, new_n20899_, new_n20900_, new_n20901_, new_n20902_,
    new_n20903_, new_n20904_, new_n20905_, new_n20906_, new_n20907_,
    new_n20908_, new_n20909_, new_n20910_, new_n20911_, new_n20912_,
    new_n20913_, new_n20914_, new_n20915_, new_n20916_, new_n20917_,
    new_n20918_, new_n20919_, new_n20920_, new_n20921_, new_n20922_,
    new_n20923_, new_n20924_, new_n20925_, new_n20926_, new_n20927_,
    new_n20928_, new_n20929_, new_n20930_, new_n20931_, new_n20932_,
    new_n20933_, new_n20934_, new_n20935_, new_n20936_, new_n20937_,
    new_n20938_, new_n20939_, new_n20940_, new_n20941_, new_n20942_,
    new_n20943_, new_n20944_, new_n20945_, new_n20946_, new_n20947_,
    new_n20948_, new_n20949_, new_n20950_, new_n20951_, new_n20952_,
    new_n20953_, new_n20954_, new_n20955_, new_n20956_, new_n20957_,
    new_n20958_, new_n20959_, new_n20960_, new_n20961_, new_n20962_,
    new_n20963_, new_n20964_, new_n20965_, new_n20966_, new_n20967_,
    new_n20968_, new_n20969_, new_n20970_, new_n20971_, new_n20972_,
    new_n20973_, new_n20974_, new_n20975_, new_n20976_, new_n20977_,
    new_n20978_, new_n20979_, new_n20980_, new_n20981_, new_n20982_,
    new_n20983_, new_n20984_, new_n20985_, new_n20986_, new_n20987_,
    new_n20988_, new_n20989_, new_n20990_, new_n20991_, new_n20992_,
    new_n20993_, new_n20994_, new_n20995_, new_n20996_, new_n20997_,
    new_n20998_, new_n20999_, new_n21000_, new_n21001_, new_n21002_,
    new_n21003_, new_n21004_, new_n21005_, new_n21006_, new_n21007_,
    new_n21008_, new_n21009_, new_n21010_, new_n21011_, new_n21012_,
    new_n21013_, new_n21014_, new_n21015_, new_n21016_, new_n21017_,
    new_n21018_, new_n21019_, new_n21020_, new_n21021_, new_n21022_,
    new_n21023_, new_n21024_, new_n21025_, new_n21026_, new_n21027_,
    new_n21028_, new_n21029_, new_n21030_, new_n21031_, new_n21032_,
    new_n21033_, new_n21034_, new_n21035_, new_n21036_, new_n21037_,
    new_n21038_, new_n21039_, new_n21040_, new_n21041_, new_n21042_,
    new_n21043_, new_n21044_, new_n21045_, new_n21046_, new_n21047_,
    new_n21048_, new_n21049_, new_n21050_, new_n21051_, new_n21052_,
    new_n21053_, new_n21054_, new_n21055_, new_n21056_, new_n21057_,
    new_n21058_, new_n21059_, new_n21060_, new_n21061_, new_n21062_,
    new_n21063_, new_n21064_, new_n21065_, new_n21066_, new_n21067_,
    new_n21068_, new_n21069_, new_n21070_, new_n21071_, new_n21072_,
    new_n21073_, new_n21074_, new_n21075_, new_n21076_, new_n21077_,
    new_n21078_, new_n21079_, new_n21080_, new_n21081_, new_n21082_,
    new_n21083_, new_n21084_, new_n21085_, new_n21086_, new_n21087_,
    new_n21088_, new_n21089_, new_n21090_, new_n21091_, new_n21092_,
    new_n21093_, new_n21094_, new_n21095_, new_n21096_, new_n21097_,
    new_n21098_, new_n21099_, new_n21100_, new_n21101_, new_n21102_,
    new_n21103_, new_n21104_, new_n21105_, new_n21106_, new_n21107_,
    new_n21108_, new_n21109_, new_n21110_, new_n21111_, new_n21112_,
    new_n21113_, new_n21114_, new_n21115_, new_n21116_, new_n21117_,
    new_n21118_, new_n21119_, new_n21120_, new_n21121_, new_n21122_,
    new_n21123_, new_n21124_, new_n21125_, new_n21126_, new_n21127_,
    new_n21128_, new_n21129_, new_n21130_, new_n21131_, new_n21132_,
    new_n21133_, new_n21134_, new_n21135_, new_n21136_, new_n21137_,
    new_n21138_, new_n21139_, new_n21140_, new_n21141_, new_n21142_,
    new_n21143_, new_n21144_, new_n21145_, new_n21146_, new_n21147_,
    new_n21148_, new_n21149_, new_n21150_, new_n21151_, new_n21152_,
    new_n21153_, new_n21154_, new_n21155_, new_n21156_, new_n21157_,
    new_n21158_, new_n21159_, new_n21160_, new_n21161_, new_n21162_,
    new_n21163_, new_n21164_, new_n21165_, new_n21166_, new_n21167_,
    new_n21168_, new_n21169_, new_n21170_, new_n21171_, new_n21172_,
    new_n21173_, new_n21174_, new_n21175_, new_n21176_, new_n21177_,
    new_n21178_, new_n21179_, new_n21180_, new_n21181_, new_n21182_,
    new_n21183_, new_n21184_, new_n21185_, new_n21186_, new_n21187_,
    new_n21188_, new_n21189_, new_n21190_, new_n21191_, new_n21192_,
    new_n21193_, new_n21194_, new_n21195_, new_n21196_, new_n21197_,
    new_n21198_, new_n21199_, new_n21200_, new_n21201_, new_n21202_,
    new_n21203_, new_n21204_, new_n21205_, new_n21206_, new_n21207_,
    new_n21208_, new_n21209_, new_n21210_, new_n21211_, new_n21212_,
    new_n21213_, new_n21214_, new_n21215_, new_n21216_, new_n21217_,
    new_n21218_, new_n21219_, new_n21220_, new_n21221_, new_n21222_,
    new_n21223_, new_n21224_, new_n21225_, new_n21226_, new_n21227_,
    new_n21228_, new_n21229_, new_n21230_, new_n21231_, new_n21232_,
    new_n21233_, new_n21234_, new_n21235_, new_n21236_, new_n21237_,
    new_n21238_, new_n21239_, new_n21240_, new_n21241_, new_n21242_,
    new_n21243_, new_n21244_, new_n21245_, new_n21246_, new_n21247_,
    new_n21248_, new_n21249_, new_n21250_, new_n21251_, new_n21252_,
    new_n21253_, new_n21254_, new_n21255_, new_n21256_, new_n21257_,
    new_n21258_, new_n21259_, new_n21260_, new_n21261_, new_n21262_,
    new_n21263_, new_n21264_, new_n21265_, new_n21266_, new_n21267_,
    new_n21268_, new_n21269_, new_n21270_, new_n21271_, new_n21272_,
    new_n21273_, new_n21274_, new_n21275_, new_n21276_, new_n21277_,
    new_n21278_, new_n21279_, new_n21280_, new_n21281_, new_n21282_,
    new_n21283_, new_n21284_, new_n21285_, new_n21286_, new_n21287_,
    new_n21288_, new_n21289_, new_n21290_, new_n21291_, new_n21292_,
    new_n21293_, new_n21294_, new_n21295_, new_n21296_, new_n21297_,
    new_n21298_, new_n21299_, new_n21300_, new_n21301_, new_n21302_,
    new_n21303_, new_n21304_, new_n21305_, new_n21306_, new_n21307_,
    new_n21308_, new_n21309_, new_n21310_, new_n21311_, new_n21312_,
    new_n21313_, new_n21314_, new_n21315_, new_n21316_, new_n21317_,
    new_n21318_, new_n21319_, new_n21320_, new_n21321_, new_n21322_,
    new_n21323_, new_n21324_, new_n21325_, new_n21326_, new_n21327_,
    new_n21328_, new_n21329_, new_n21330_, new_n21331_, new_n21332_,
    new_n21333_, new_n21334_, new_n21335_, new_n21336_, new_n21337_,
    new_n21338_, new_n21339_, new_n21340_, new_n21341_, new_n21342_,
    new_n21343_, new_n21344_, new_n21345_, new_n21346_, new_n21347_,
    new_n21348_, new_n21349_, new_n21350_, new_n21351_, new_n21352_,
    new_n21353_, new_n21354_, new_n21355_, new_n21356_, new_n21357_,
    new_n21358_, new_n21359_, new_n21360_, new_n21361_, new_n21362_,
    new_n21363_, new_n21364_, new_n21365_, new_n21366_, new_n21367_,
    new_n21368_, new_n21369_, new_n21370_, new_n21371_, new_n21372_,
    new_n21373_, new_n21374_, new_n21375_, new_n21376_, new_n21377_,
    new_n21378_, new_n21379_, new_n21380_, new_n21381_, new_n21382_,
    new_n21383_, new_n21384_, new_n21385_, new_n21386_, new_n21387_,
    new_n21388_, new_n21389_, new_n21390_, new_n21391_, new_n21392_,
    new_n21393_, new_n21394_, new_n21395_, new_n21396_, new_n21397_,
    new_n21398_, new_n21399_, new_n21400_, new_n21401_, new_n21402_,
    new_n21403_, new_n21404_, new_n21405_, new_n21406_, new_n21407_,
    new_n21408_, new_n21409_, new_n21410_, new_n21411_, new_n21412_,
    new_n21413_, new_n21414_, new_n21415_, new_n21416_, new_n21417_,
    new_n21418_, new_n21419_, new_n21420_, new_n21421_, new_n21422_,
    new_n21423_, new_n21424_, new_n21425_, new_n21426_, new_n21427_,
    new_n21428_, new_n21429_, new_n21430_, new_n21431_, new_n21432_,
    new_n21433_, new_n21434_, new_n21435_, new_n21436_, new_n21437_,
    new_n21438_, new_n21439_, new_n21440_, new_n21441_, new_n21442_,
    new_n21443_, new_n21444_, new_n21445_, new_n21446_, new_n21447_,
    new_n21448_, new_n21449_, new_n21450_, new_n21451_, new_n21452_,
    new_n21453_, new_n21454_, new_n21455_, new_n21456_, new_n21457_,
    new_n21458_, new_n21459_, new_n21460_, new_n21461_, new_n21462_,
    new_n21463_, new_n21464_, new_n21465_, new_n21466_, new_n21467_,
    new_n21468_, new_n21469_, new_n21470_, new_n21471_, new_n21472_,
    new_n21473_, new_n21474_, new_n21475_, new_n21477_, new_n21478_,
    new_n21479_, new_n21480_, new_n21481_, new_n21482_, new_n21483_,
    new_n21484_, new_n21485_, new_n21486_, new_n21487_, new_n21488_,
    new_n21489_, new_n21490_, new_n21491_, new_n21492_, new_n21493_,
    new_n21494_, new_n21495_, new_n21496_, new_n21497_, new_n21498_,
    new_n21499_, new_n21500_, new_n21501_, new_n21502_, new_n21503_,
    new_n21504_, new_n21505_, new_n21506_, new_n21507_, new_n21508_,
    new_n21509_, new_n21510_, new_n21511_, new_n21512_, new_n21513_,
    new_n21514_, new_n21515_, new_n21516_, new_n21517_, new_n21518_,
    new_n21519_, new_n21520_, new_n21521_, new_n21522_, new_n21523_,
    new_n21524_, new_n21525_, new_n21526_, new_n21527_, new_n21528_,
    new_n21529_, new_n21530_, new_n21531_, new_n21532_, new_n21533_,
    new_n21534_, new_n21535_, new_n21536_, new_n21537_, new_n21538_,
    new_n21539_, new_n21540_, new_n21541_, new_n21542_, new_n21543_,
    new_n21544_, new_n21545_, new_n21546_, new_n21547_, new_n21548_,
    new_n21549_, new_n21550_, new_n21551_, new_n21552_, new_n21553_,
    new_n21554_, new_n21555_, new_n21556_, new_n21557_, new_n21558_,
    new_n21559_, new_n21560_, new_n21561_, new_n21562_, new_n21563_,
    new_n21564_, new_n21565_, new_n21566_, new_n21567_, new_n21568_,
    new_n21569_, new_n21570_, new_n21571_, new_n21572_, new_n21573_,
    new_n21574_, new_n21575_, new_n21576_, new_n21577_, new_n21578_,
    new_n21579_, new_n21580_, new_n21581_, new_n21582_, new_n21583_,
    new_n21584_, new_n21585_, new_n21586_, new_n21587_, new_n21588_,
    new_n21589_, new_n21590_, new_n21591_, new_n21592_, new_n21593_,
    new_n21594_, new_n21595_, new_n21596_, new_n21597_, new_n21598_,
    new_n21599_, new_n21600_, new_n21601_, new_n21602_, new_n21603_,
    new_n21604_, new_n21605_, new_n21606_, new_n21607_, new_n21608_,
    new_n21609_, new_n21610_, new_n21611_, new_n21612_, new_n21613_,
    new_n21614_, new_n21615_, new_n21616_, new_n21617_, new_n21618_,
    new_n21619_, new_n21620_, new_n21621_, new_n21622_, new_n21623_,
    new_n21624_, new_n21625_, new_n21626_, new_n21627_, new_n21628_,
    new_n21629_, new_n21630_, new_n21631_, new_n21632_, new_n21633_,
    new_n21634_, new_n21635_, new_n21636_, new_n21637_, new_n21638_,
    new_n21639_, new_n21640_, new_n21641_, new_n21642_, new_n21643_,
    new_n21644_, new_n21645_, new_n21646_, new_n21647_, new_n21648_,
    new_n21649_, new_n21650_, new_n21651_, new_n21652_, new_n21653_,
    new_n21654_, new_n21655_, new_n21656_, new_n21657_, new_n21658_,
    new_n21659_, new_n21660_, new_n21661_, new_n21662_, new_n21663_,
    new_n21664_, new_n21665_, new_n21666_, new_n21667_, new_n21668_,
    new_n21669_, new_n21670_, new_n21671_, new_n21672_, new_n21673_,
    new_n21674_, new_n21675_, new_n21676_, new_n21677_, new_n21678_,
    new_n21679_, new_n21680_, new_n21681_, new_n21682_, new_n21683_,
    new_n21684_, new_n21685_, new_n21686_, new_n21687_, new_n21688_,
    new_n21689_, new_n21690_, new_n21691_, new_n21692_, new_n21693_,
    new_n21694_, new_n21695_, new_n21696_, new_n21697_, new_n21698_,
    new_n21699_, new_n21700_, new_n21701_, new_n21702_, new_n21703_,
    new_n21704_, new_n21705_, new_n21706_, new_n21707_, new_n21708_,
    new_n21709_, new_n21710_, new_n21711_, new_n21712_, new_n21713_,
    new_n21714_, new_n21715_, new_n21716_, new_n21717_, new_n21718_,
    new_n21719_, new_n21720_, new_n21721_, new_n21722_, new_n21723_,
    new_n21724_, new_n21725_, new_n21726_, new_n21727_, new_n21728_,
    new_n21729_, new_n21730_, new_n21731_, new_n21732_, new_n21733_,
    new_n21734_, new_n21735_, new_n21736_, new_n21737_, new_n21738_,
    new_n21739_, new_n21740_, new_n21741_, new_n21742_, new_n21743_,
    new_n21744_, new_n21745_, new_n21746_, new_n21747_, new_n21748_,
    new_n21749_, new_n21750_, new_n21751_, new_n21752_, new_n21753_,
    new_n21754_, new_n21755_, new_n21756_, new_n21757_, new_n21758_,
    new_n21759_, new_n21760_, new_n21761_, new_n21762_, new_n21763_,
    new_n21764_, new_n21765_, new_n21766_, new_n21767_, new_n21768_,
    new_n21769_, new_n21770_, new_n21771_, new_n21772_, new_n21773_,
    new_n21774_, new_n21775_, new_n21776_, new_n21777_, new_n21778_,
    new_n21779_, new_n21780_, new_n21781_, new_n21782_, new_n21783_,
    new_n21784_, new_n21785_, new_n21786_, new_n21787_, new_n21788_,
    new_n21789_, new_n21790_, new_n21791_, new_n21792_, new_n21793_,
    new_n21794_, new_n21795_, new_n21796_, new_n21797_, new_n21798_,
    new_n21799_, new_n21800_, new_n21801_, new_n21802_, new_n21803_,
    new_n21804_, new_n21805_, new_n21806_, new_n21807_, new_n21808_,
    new_n21809_, new_n21810_, new_n21811_, new_n21812_, new_n21813_,
    new_n21814_, new_n21815_, new_n21816_, new_n21817_, new_n21818_,
    new_n21819_, new_n21820_, new_n21821_, new_n21822_, new_n21823_,
    new_n21824_, new_n21825_, new_n21826_, new_n21827_, new_n21828_,
    new_n21829_, new_n21830_, new_n21831_, new_n21832_, new_n21833_,
    new_n21834_, new_n21835_, new_n21836_, new_n21837_, new_n21838_,
    new_n21839_, new_n21840_, new_n21841_, new_n21842_, new_n21843_,
    new_n21844_, new_n21845_, new_n21846_, new_n21847_, new_n21848_,
    new_n21849_, new_n21850_, new_n21851_, new_n21852_, new_n21853_,
    new_n21854_, new_n21855_, new_n21856_, new_n21857_, new_n21858_,
    new_n21859_, new_n21860_, new_n21861_, new_n21862_, new_n21863_,
    new_n21864_, new_n21865_, new_n21866_, new_n21867_, new_n21868_,
    new_n21869_, new_n21870_, new_n21871_, new_n21872_, new_n21873_,
    new_n21874_, new_n21875_, new_n21876_, new_n21877_, new_n21878_,
    new_n21879_, new_n21880_, new_n21881_, new_n21882_, new_n21883_,
    new_n21884_, new_n21885_, new_n21886_, new_n21887_, new_n21888_,
    new_n21889_, new_n21890_, new_n21891_, new_n21892_, new_n21893_,
    new_n21894_, new_n21895_, new_n21896_, new_n21897_, new_n21898_,
    new_n21899_, new_n21900_, new_n21901_, new_n21902_, new_n21903_,
    new_n21904_, new_n21905_, new_n21906_, new_n21907_, new_n21908_,
    new_n21909_, new_n21910_, new_n21911_, new_n21912_, new_n21913_,
    new_n21914_, new_n21915_, new_n21916_, new_n21917_, new_n21918_,
    new_n21919_, new_n21920_, new_n21921_, new_n21922_, new_n21923_,
    new_n21924_, new_n21925_, new_n21926_, new_n21927_, new_n21928_,
    new_n21929_, new_n21930_, new_n21931_, new_n21932_, new_n21933_,
    new_n21934_, new_n21935_, new_n21936_, new_n21937_, new_n21938_,
    new_n21939_, new_n21940_, new_n21941_, new_n21942_, new_n21943_,
    new_n21944_, new_n21945_, new_n21946_, new_n21947_, new_n21948_,
    new_n21949_, new_n21950_, new_n21951_, new_n21952_, new_n21953_,
    new_n21954_, new_n21955_, new_n21956_, new_n21957_, new_n21958_,
    new_n21959_, new_n21960_, new_n21961_, new_n21962_, new_n21963_,
    new_n21964_, new_n21965_, new_n21966_, new_n21967_, new_n21968_,
    new_n21969_, new_n21970_, new_n21971_, new_n21972_, new_n21973_,
    new_n21974_, new_n21975_, new_n21976_, new_n21977_, new_n21978_,
    new_n21979_, new_n21980_, new_n21981_, new_n21982_, new_n21983_,
    new_n21984_, new_n21985_, new_n21986_, new_n21987_, new_n21988_,
    new_n21989_, new_n21990_, new_n21991_, new_n21992_, new_n21993_,
    new_n21994_, new_n21995_, new_n21996_, new_n21997_, new_n21998_,
    new_n21999_, new_n22000_, new_n22001_, new_n22002_, new_n22003_,
    new_n22004_, new_n22005_, new_n22006_, new_n22007_, new_n22008_,
    new_n22009_, new_n22010_, new_n22011_, new_n22012_, new_n22013_,
    new_n22014_, new_n22015_, new_n22016_, new_n22017_, new_n22018_,
    new_n22019_, new_n22020_, new_n22021_, new_n22022_, new_n22023_,
    new_n22024_, new_n22025_, new_n22026_, new_n22027_, new_n22028_,
    new_n22029_, new_n22030_, new_n22031_, new_n22032_, new_n22033_,
    new_n22034_, new_n22035_, new_n22036_, new_n22037_, new_n22038_,
    new_n22039_, new_n22040_, new_n22041_, new_n22042_, new_n22043_,
    new_n22044_, new_n22045_, new_n22046_, new_n22047_, new_n22048_,
    new_n22049_, new_n22050_, new_n22051_, new_n22052_, new_n22053_,
    new_n22054_, new_n22055_, new_n22056_, new_n22057_, new_n22058_,
    new_n22059_, new_n22060_, new_n22061_, new_n22062_, new_n22063_,
    new_n22064_, new_n22065_, new_n22066_, new_n22067_, new_n22068_,
    new_n22069_, new_n22070_, new_n22071_, new_n22072_, new_n22073_,
    new_n22074_, new_n22075_, new_n22076_, new_n22077_, new_n22078_,
    new_n22079_, new_n22080_, new_n22081_, new_n22082_, new_n22083_,
    new_n22084_, new_n22085_, new_n22086_, new_n22087_, new_n22088_,
    new_n22089_, new_n22090_, new_n22091_, new_n22092_, new_n22093_,
    new_n22094_, new_n22095_, new_n22096_, new_n22097_, new_n22098_,
    new_n22099_, new_n22100_, new_n22101_, new_n22102_, new_n22103_,
    new_n22104_, new_n22105_, new_n22106_, new_n22107_, new_n22108_,
    new_n22109_, new_n22110_, new_n22111_, new_n22112_, new_n22113_,
    new_n22114_, new_n22115_, new_n22116_, new_n22117_, new_n22118_,
    new_n22119_, new_n22120_, new_n22121_, new_n22122_, new_n22123_,
    new_n22124_, new_n22125_, new_n22126_, new_n22127_, new_n22128_,
    new_n22129_, new_n22130_, new_n22131_, new_n22132_, new_n22133_,
    new_n22134_, new_n22135_, new_n22136_, new_n22137_, new_n22138_,
    new_n22140_, new_n22141_, new_n22142_, new_n22143_, new_n22144_,
    new_n22145_, new_n22146_, new_n22147_, new_n22148_, new_n22149_,
    new_n22150_, new_n22151_, new_n22152_, new_n22153_, new_n22154_,
    new_n22155_, new_n22156_, new_n22157_, new_n22158_, new_n22159_,
    new_n22160_, new_n22161_, new_n22162_, new_n22163_, new_n22164_,
    new_n22165_, new_n22166_, new_n22167_, new_n22168_, new_n22169_,
    new_n22170_, new_n22171_, new_n22172_, new_n22173_, new_n22174_,
    new_n22175_, new_n22176_, new_n22177_, new_n22178_, new_n22179_,
    new_n22180_, new_n22181_, new_n22182_, new_n22183_, new_n22184_,
    new_n22185_, new_n22186_, new_n22187_, new_n22188_, new_n22189_,
    new_n22190_, new_n22191_, new_n22192_, new_n22193_, new_n22194_,
    new_n22195_, new_n22196_, new_n22197_, new_n22198_, new_n22199_,
    new_n22200_, new_n22201_, new_n22202_, new_n22203_, new_n22204_,
    new_n22205_, new_n22206_, new_n22207_, new_n22208_, new_n22209_,
    new_n22210_, new_n22211_, new_n22212_, new_n22213_, new_n22214_,
    new_n22215_, new_n22216_, new_n22217_, new_n22218_, new_n22219_,
    new_n22220_, new_n22221_, new_n22222_, new_n22223_, new_n22224_,
    new_n22225_, new_n22226_, new_n22227_, new_n22228_, new_n22229_,
    new_n22230_, new_n22231_, new_n22232_, new_n22233_, new_n22234_,
    new_n22235_, new_n22236_, new_n22237_, new_n22238_, new_n22239_,
    new_n22240_, new_n22241_, new_n22242_, new_n22243_, new_n22244_,
    new_n22245_, new_n22246_, new_n22247_, new_n22248_, new_n22249_,
    new_n22250_, new_n22251_, new_n22252_, new_n22253_, new_n22254_,
    new_n22255_, new_n22256_, new_n22257_, new_n22258_, new_n22259_,
    new_n22260_, new_n22261_, new_n22262_, new_n22263_, new_n22264_,
    new_n22265_, new_n22266_, new_n22267_, new_n22268_, new_n22269_,
    new_n22270_, new_n22271_, new_n22272_, new_n22273_, new_n22274_,
    new_n22275_, new_n22276_, new_n22277_, new_n22278_, new_n22279_,
    new_n22280_, new_n22281_, new_n22282_, new_n22283_, new_n22284_,
    new_n22285_, new_n22286_, new_n22287_, new_n22288_, new_n22289_,
    new_n22290_, new_n22291_, new_n22292_, new_n22293_, new_n22294_,
    new_n22295_, new_n22296_, new_n22297_, new_n22298_, new_n22299_,
    new_n22300_, new_n22301_, new_n22302_, new_n22303_, new_n22304_,
    new_n22305_, new_n22306_, new_n22307_, new_n22308_, new_n22309_,
    new_n22310_, new_n22311_, new_n22312_, new_n22313_, new_n22314_,
    new_n22315_, new_n22316_, new_n22317_, new_n22318_, new_n22319_,
    new_n22320_, new_n22321_, new_n22322_, new_n22323_, new_n22324_,
    new_n22325_, new_n22326_, new_n22327_, new_n22328_, new_n22329_,
    new_n22330_, new_n22331_, new_n22332_, new_n22333_, new_n22334_,
    new_n22335_, new_n22336_, new_n22337_, new_n22338_, new_n22339_,
    new_n22340_, new_n22341_, new_n22342_, new_n22343_, new_n22344_,
    new_n22345_, new_n22346_, new_n22347_, new_n22348_, new_n22349_,
    new_n22350_, new_n22351_, new_n22352_, new_n22353_, new_n22354_,
    new_n22355_, new_n22356_, new_n22357_, new_n22358_, new_n22359_,
    new_n22360_, new_n22361_, new_n22362_, new_n22363_, new_n22364_,
    new_n22365_, new_n22366_, new_n22367_, new_n22368_, new_n22369_,
    new_n22370_, new_n22371_, new_n22372_, new_n22373_, new_n22374_,
    new_n22375_, new_n22376_, new_n22377_, new_n22378_, new_n22379_,
    new_n22380_, new_n22381_, new_n22382_, new_n22383_, new_n22384_,
    new_n22385_, new_n22386_, new_n22387_, new_n22388_, new_n22389_,
    new_n22390_, new_n22391_, new_n22392_, new_n22393_, new_n22394_,
    new_n22395_, new_n22396_, new_n22397_, new_n22398_, new_n22399_,
    new_n22400_, new_n22401_, new_n22402_, new_n22403_, new_n22404_,
    new_n22405_, new_n22406_, new_n22407_, new_n22408_, new_n22409_,
    new_n22410_, new_n22411_, new_n22412_, new_n22413_, new_n22414_,
    new_n22415_, new_n22416_, new_n22417_, new_n22418_, new_n22419_,
    new_n22420_, new_n22421_, new_n22422_, new_n22423_, new_n22424_,
    new_n22425_, new_n22426_, new_n22427_, new_n22428_, new_n22429_,
    new_n22430_, new_n22431_, new_n22432_, new_n22433_, new_n22434_,
    new_n22435_, new_n22436_, new_n22437_, new_n22438_, new_n22439_,
    new_n22440_, new_n22441_, new_n22442_, new_n22443_, new_n22444_,
    new_n22445_, new_n22446_, new_n22447_, new_n22448_, new_n22449_,
    new_n22450_, new_n22451_, new_n22452_, new_n22453_, new_n22454_,
    new_n22455_, new_n22456_, new_n22457_, new_n22458_, new_n22459_,
    new_n22460_, new_n22461_, new_n22462_, new_n22463_, new_n22464_,
    new_n22465_, new_n22466_, new_n22467_, new_n22468_, new_n22469_,
    new_n22470_, new_n22471_, new_n22472_, new_n22473_, new_n22474_,
    new_n22475_, new_n22476_, new_n22477_, new_n22478_, new_n22479_,
    new_n22480_, new_n22481_, new_n22482_, new_n22483_, new_n22484_,
    new_n22485_, new_n22486_, new_n22487_, new_n22488_, new_n22489_,
    new_n22490_, new_n22491_, new_n22492_, new_n22493_, new_n22494_,
    new_n22495_, new_n22496_, new_n22497_, new_n22498_, new_n22499_,
    new_n22500_, new_n22501_, new_n22502_, new_n22503_, new_n22504_,
    new_n22505_, new_n22506_, new_n22507_, new_n22508_, new_n22509_,
    new_n22510_, new_n22511_, new_n22512_, new_n22513_, new_n22514_,
    new_n22515_, new_n22516_, new_n22517_, new_n22518_, new_n22519_,
    new_n22520_, new_n22521_, new_n22522_, new_n22523_, new_n22524_,
    new_n22525_, new_n22526_, new_n22527_, new_n22528_, new_n22529_,
    new_n22530_, new_n22531_, new_n22532_, new_n22533_, new_n22534_,
    new_n22535_, new_n22536_, new_n22537_, new_n22538_, new_n22539_,
    new_n22540_, new_n22541_, new_n22542_, new_n22543_, new_n22544_,
    new_n22545_, new_n22546_, new_n22547_, new_n22548_, new_n22549_,
    new_n22550_, new_n22551_, new_n22552_, new_n22553_, new_n22554_,
    new_n22555_, new_n22556_, new_n22557_, new_n22558_, new_n22559_,
    new_n22560_, new_n22561_, new_n22562_, new_n22563_, new_n22564_,
    new_n22565_, new_n22566_, new_n22567_, new_n22568_, new_n22569_,
    new_n22570_, new_n22571_, new_n22572_, new_n22573_, new_n22574_,
    new_n22575_, new_n22576_, new_n22577_, new_n22578_, new_n22579_,
    new_n22580_, new_n22581_, new_n22582_, new_n22583_, new_n22584_,
    new_n22585_, new_n22586_, new_n22587_, new_n22588_, new_n22589_,
    new_n22590_, new_n22591_, new_n22592_, new_n22593_, new_n22594_,
    new_n22595_, new_n22596_, new_n22597_, new_n22598_, new_n22599_,
    new_n22600_, new_n22601_, new_n22602_, new_n22603_, new_n22604_,
    new_n22605_, new_n22606_, new_n22607_, new_n22608_, new_n22609_,
    new_n22610_, new_n22611_, new_n22612_, new_n22613_, new_n22614_,
    new_n22615_, new_n22616_, new_n22617_, new_n22618_, new_n22619_,
    new_n22620_, new_n22621_, new_n22622_, new_n22623_, new_n22624_,
    new_n22625_, new_n22626_, new_n22627_, new_n22628_, new_n22629_,
    new_n22630_, new_n22631_, new_n22632_, new_n22633_, new_n22634_,
    new_n22635_, new_n22636_, new_n22637_, new_n22638_, new_n22639_,
    new_n22640_, new_n22641_, new_n22642_, new_n22643_, new_n22644_,
    new_n22645_, new_n22646_, new_n22647_, new_n22648_, new_n22649_,
    new_n22650_, new_n22651_, new_n22652_, new_n22653_, new_n22654_,
    new_n22655_, new_n22656_, new_n22657_, new_n22658_, new_n22659_,
    new_n22660_, new_n22661_, new_n22662_, new_n22663_, new_n22664_,
    new_n22665_, new_n22666_, new_n22667_, new_n22668_, new_n22669_,
    new_n22670_, new_n22671_, new_n22672_, new_n22673_, new_n22674_,
    new_n22675_, new_n22676_, new_n22677_, new_n22678_, new_n22679_,
    new_n22680_, new_n22681_, new_n22682_, new_n22683_, new_n22684_,
    new_n22685_, new_n22686_, new_n22687_, new_n22688_, new_n22689_,
    new_n22690_, new_n22691_, new_n22692_, new_n22693_, new_n22694_,
    new_n22695_, new_n22696_, new_n22697_, new_n22698_, new_n22699_,
    new_n22700_, new_n22701_, new_n22702_, new_n22703_, new_n22704_,
    new_n22705_, new_n22706_, new_n22707_, new_n22708_, new_n22709_,
    new_n22710_, new_n22711_, new_n22712_, new_n22713_, new_n22714_,
    new_n22715_, new_n22716_, new_n22717_, new_n22718_, new_n22719_,
    new_n22720_, new_n22721_, new_n22722_, new_n22723_, new_n22724_,
    new_n22725_, new_n22726_, new_n22727_, new_n22728_, new_n22729_,
    new_n22730_, new_n22731_, new_n22732_, new_n22733_, new_n22734_,
    new_n22735_, new_n22736_, new_n22737_, new_n22738_, new_n22739_,
    new_n22740_, new_n22741_, new_n22742_, new_n22743_, new_n22744_,
    new_n22745_, new_n22746_, new_n22747_, new_n22748_, new_n22749_,
    new_n22750_, new_n22751_, new_n22752_, new_n22753_, new_n22754_,
    new_n22755_, new_n22756_, new_n22757_, new_n22758_, new_n22759_,
    new_n22760_, new_n22761_, new_n22762_, new_n22763_, new_n22764_,
    new_n22765_, new_n22766_, new_n22767_, new_n22768_, new_n22769_,
    new_n22770_, new_n22771_, new_n22772_, new_n22773_, new_n22774_,
    new_n22775_, new_n22776_, new_n22777_, new_n22778_, new_n22779_,
    new_n22780_, new_n22781_, new_n22782_, new_n22783_, new_n22784_,
    new_n22785_, new_n22786_, new_n22787_, new_n22788_, new_n22789_,
    new_n22790_, new_n22791_, new_n22792_, new_n22793_, new_n22794_,
    new_n22795_, new_n22796_, new_n22797_, new_n22798_, new_n22799_,
    new_n22800_, new_n22801_, new_n22802_, new_n22803_, new_n22804_,
    new_n22805_, new_n22806_, new_n22807_, new_n22808_, new_n22809_,
    new_n22810_, new_n22811_, new_n22812_, new_n22813_, new_n22814_,
    new_n22815_, new_n22816_, new_n22817_, new_n22818_, new_n22819_,
    new_n22820_, new_n22821_, new_n22822_, new_n22823_, new_n22824_,
    new_n22825_, new_n22826_, new_n22827_, new_n22828_, new_n22829_,
    new_n22830_, new_n22831_, new_n22832_, new_n22833_, new_n22834_,
    new_n22835_, new_n22836_, new_n22837_, new_n22838_, new_n22839_,
    new_n22840_, new_n22841_, new_n22842_, new_n22843_, new_n22844_,
    new_n22845_, new_n22846_, new_n22847_, new_n22848_, new_n22849_,
    new_n22850_, new_n22851_, new_n22852_, new_n22853_, new_n22854_,
    new_n22855_, new_n22856_, new_n22857_, new_n22858_, new_n22859_,
    new_n22860_, new_n22861_, new_n22862_, new_n22863_, new_n22864_,
    new_n22865_, new_n22866_, new_n22867_, new_n22868_, new_n22869_,
    new_n22870_, new_n22871_, new_n22872_, new_n22873_, new_n22874_,
    new_n22876_, new_n22877_, new_n22878_, new_n22879_, new_n22880_,
    new_n22881_, new_n22882_, new_n22883_, new_n22884_, new_n22885_,
    new_n22886_, new_n22887_, new_n22888_, new_n22889_, new_n22890_,
    new_n22891_, new_n22892_, new_n22893_, new_n22894_, new_n22895_,
    new_n22896_, new_n22897_, new_n22898_, new_n22899_, new_n22900_,
    new_n22901_, new_n22902_, new_n22903_, new_n22904_, new_n22905_,
    new_n22906_, new_n22907_, new_n22908_, new_n22909_, new_n22910_,
    new_n22911_, new_n22912_, new_n22913_, new_n22914_, new_n22915_,
    new_n22916_, new_n22917_, new_n22918_, new_n22919_, new_n22920_,
    new_n22921_, new_n22922_, new_n22923_, new_n22924_, new_n22925_,
    new_n22926_, new_n22927_, new_n22928_, new_n22929_, new_n22930_,
    new_n22931_, new_n22932_, new_n22933_, new_n22934_, new_n22935_,
    new_n22936_, new_n22937_, new_n22938_, new_n22939_, new_n22940_,
    new_n22941_, new_n22942_, new_n22943_, new_n22944_, new_n22945_,
    new_n22946_, new_n22947_, new_n22948_, new_n22949_, new_n22950_,
    new_n22951_, new_n22952_, new_n22953_, new_n22954_, new_n22955_,
    new_n22956_, new_n22957_, new_n22958_, new_n22959_, new_n22960_,
    new_n22961_, new_n22962_, new_n22963_, new_n22964_, new_n22965_,
    new_n22966_, new_n22967_, new_n22968_, new_n22969_, new_n22970_,
    new_n22971_, new_n22972_, new_n22973_, new_n22974_, new_n22975_,
    new_n22976_, new_n22977_, new_n22978_, new_n22979_, new_n22980_,
    new_n22981_, new_n22982_, new_n22983_, new_n22984_, new_n22985_,
    new_n22986_, new_n22987_, new_n22988_, new_n22989_, new_n22990_,
    new_n22991_, new_n22992_, new_n22993_, new_n22994_, new_n22995_,
    new_n22996_, new_n22997_, new_n22998_, new_n22999_, new_n23000_,
    new_n23001_, new_n23002_, new_n23003_, new_n23004_, new_n23005_,
    new_n23006_, new_n23007_, new_n23008_, new_n23009_, new_n23010_,
    new_n23011_, new_n23012_, new_n23013_, new_n23014_, new_n23015_,
    new_n23016_, new_n23017_, new_n23018_, new_n23019_, new_n23020_,
    new_n23021_, new_n23022_, new_n23023_, new_n23024_, new_n23025_,
    new_n23026_, new_n23027_, new_n23028_, new_n23029_, new_n23030_,
    new_n23031_, new_n23032_, new_n23033_, new_n23034_, new_n23035_,
    new_n23036_, new_n23037_, new_n23038_, new_n23039_, new_n23040_,
    new_n23041_, new_n23042_, new_n23043_, new_n23044_, new_n23045_,
    new_n23046_, new_n23047_, new_n23048_, new_n23049_, new_n23050_,
    new_n23051_, new_n23052_, new_n23053_, new_n23054_, new_n23055_,
    new_n23056_, new_n23057_, new_n23058_, new_n23059_, new_n23060_,
    new_n23061_, new_n23062_, new_n23063_, new_n23064_, new_n23065_,
    new_n23066_, new_n23067_, new_n23068_, new_n23069_, new_n23070_,
    new_n23071_, new_n23072_, new_n23073_, new_n23074_, new_n23075_,
    new_n23076_, new_n23077_, new_n23078_, new_n23079_, new_n23080_,
    new_n23081_, new_n23082_, new_n23083_, new_n23084_, new_n23085_,
    new_n23086_, new_n23087_, new_n23088_, new_n23089_, new_n23090_,
    new_n23091_, new_n23092_, new_n23093_, new_n23094_, new_n23095_,
    new_n23096_, new_n23097_, new_n23098_, new_n23099_, new_n23100_,
    new_n23101_, new_n23102_, new_n23103_, new_n23104_, new_n23105_,
    new_n23106_, new_n23107_, new_n23108_, new_n23109_, new_n23110_,
    new_n23111_, new_n23112_, new_n23113_, new_n23114_, new_n23115_,
    new_n23116_, new_n23117_, new_n23118_, new_n23119_, new_n23120_,
    new_n23121_, new_n23122_, new_n23123_, new_n23124_, new_n23125_,
    new_n23126_, new_n23127_, new_n23128_, new_n23129_, new_n23130_,
    new_n23131_, new_n23132_, new_n23133_, new_n23134_, new_n23135_,
    new_n23136_, new_n23137_, new_n23138_, new_n23139_, new_n23140_,
    new_n23141_, new_n23142_, new_n23143_, new_n23144_, new_n23145_,
    new_n23146_, new_n23147_, new_n23148_, new_n23149_, new_n23150_,
    new_n23151_, new_n23152_, new_n23153_, new_n23154_, new_n23155_,
    new_n23156_, new_n23157_, new_n23158_, new_n23159_, new_n23160_,
    new_n23161_, new_n23162_, new_n23163_, new_n23164_, new_n23165_,
    new_n23166_, new_n23167_, new_n23168_, new_n23169_, new_n23170_,
    new_n23171_, new_n23172_, new_n23173_, new_n23174_, new_n23175_,
    new_n23176_, new_n23177_, new_n23178_, new_n23179_, new_n23180_,
    new_n23181_, new_n23182_, new_n23183_, new_n23184_, new_n23185_,
    new_n23186_, new_n23187_, new_n23188_, new_n23189_, new_n23190_,
    new_n23191_, new_n23192_, new_n23193_, new_n23194_, new_n23195_,
    new_n23196_, new_n23197_, new_n23198_, new_n23199_, new_n23200_,
    new_n23201_, new_n23202_, new_n23203_, new_n23204_, new_n23205_,
    new_n23206_, new_n23207_, new_n23208_, new_n23209_, new_n23210_,
    new_n23211_, new_n23212_, new_n23213_, new_n23214_, new_n23215_,
    new_n23216_, new_n23217_, new_n23218_, new_n23219_, new_n23220_,
    new_n23221_, new_n23222_, new_n23223_, new_n23224_, new_n23225_,
    new_n23226_, new_n23227_, new_n23228_, new_n23229_, new_n23230_,
    new_n23231_, new_n23232_, new_n23233_, new_n23234_, new_n23235_,
    new_n23236_, new_n23237_, new_n23238_, new_n23239_, new_n23240_,
    new_n23241_, new_n23242_, new_n23243_, new_n23244_, new_n23245_,
    new_n23246_, new_n23247_, new_n23248_, new_n23249_, new_n23250_,
    new_n23251_, new_n23252_, new_n23253_, new_n23254_, new_n23255_,
    new_n23256_, new_n23257_, new_n23258_, new_n23259_, new_n23260_,
    new_n23261_, new_n23262_, new_n23263_, new_n23264_, new_n23265_,
    new_n23266_, new_n23267_, new_n23268_, new_n23269_, new_n23270_,
    new_n23271_, new_n23272_, new_n23273_, new_n23274_, new_n23275_,
    new_n23276_, new_n23277_, new_n23278_, new_n23279_, new_n23280_,
    new_n23281_, new_n23282_, new_n23283_, new_n23284_, new_n23285_,
    new_n23286_, new_n23287_, new_n23288_, new_n23289_, new_n23290_,
    new_n23291_, new_n23292_, new_n23293_, new_n23294_, new_n23295_,
    new_n23296_, new_n23297_, new_n23298_, new_n23299_, new_n23300_,
    new_n23301_, new_n23302_, new_n23303_, new_n23304_, new_n23305_,
    new_n23306_, new_n23307_, new_n23308_, new_n23309_, new_n23310_,
    new_n23311_, new_n23312_, new_n23313_, new_n23314_, new_n23315_,
    new_n23316_, new_n23317_, new_n23318_, new_n23319_, new_n23320_,
    new_n23321_, new_n23322_, new_n23323_, new_n23324_, new_n23325_,
    new_n23326_, new_n23327_, new_n23328_, new_n23329_, new_n23330_,
    new_n23331_, new_n23332_, new_n23333_, new_n23334_, new_n23335_,
    new_n23336_, new_n23337_, new_n23338_, new_n23339_, new_n23340_,
    new_n23341_, new_n23342_, new_n23343_, new_n23344_, new_n23345_,
    new_n23346_, new_n23347_, new_n23348_, new_n23349_, new_n23350_,
    new_n23351_, new_n23352_, new_n23353_, new_n23354_, new_n23355_,
    new_n23356_, new_n23357_, new_n23358_, new_n23359_, new_n23360_,
    new_n23361_, new_n23362_, new_n23363_, new_n23364_, new_n23365_,
    new_n23366_, new_n23367_, new_n23368_, new_n23369_, new_n23370_,
    new_n23371_, new_n23372_, new_n23373_, new_n23374_, new_n23375_,
    new_n23376_, new_n23377_, new_n23378_, new_n23379_, new_n23380_,
    new_n23381_, new_n23382_, new_n23383_, new_n23384_, new_n23385_,
    new_n23386_, new_n23387_, new_n23388_, new_n23389_, new_n23390_,
    new_n23391_, new_n23392_, new_n23393_, new_n23394_, new_n23395_,
    new_n23396_, new_n23397_, new_n23398_, new_n23399_, new_n23400_,
    new_n23401_, new_n23402_, new_n23403_, new_n23404_, new_n23405_,
    new_n23406_, new_n23407_, new_n23408_, new_n23409_, new_n23410_,
    new_n23411_, new_n23412_, new_n23413_, new_n23414_, new_n23415_,
    new_n23416_, new_n23417_, new_n23418_, new_n23419_, new_n23420_,
    new_n23421_, new_n23422_, new_n23423_, new_n23424_, new_n23425_,
    new_n23426_, new_n23427_, new_n23428_, new_n23429_, new_n23430_,
    new_n23431_, new_n23432_, new_n23433_, new_n23434_, new_n23435_,
    new_n23436_, new_n23437_, new_n23438_, new_n23439_, new_n23440_,
    new_n23441_, new_n23442_, new_n23443_, new_n23444_, new_n23445_,
    new_n23446_, new_n23447_, new_n23448_, new_n23449_, new_n23450_,
    new_n23451_, new_n23452_, new_n23453_, new_n23454_, new_n23455_,
    new_n23456_, new_n23457_, new_n23458_, new_n23459_, new_n23460_,
    new_n23461_, new_n23462_, new_n23463_, new_n23464_, new_n23465_,
    new_n23466_, new_n23467_, new_n23468_, new_n23469_, new_n23470_,
    new_n23471_, new_n23472_, new_n23473_, new_n23474_, new_n23475_,
    new_n23476_, new_n23477_, new_n23478_, new_n23479_, new_n23480_,
    new_n23481_, new_n23482_, new_n23483_, new_n23484_, new_n23485_,
    new_n23486_, new_n23487_, new_n23488_, new_n23489_, new_n23490_,
    new_n23491_, new_n23492_, new_n23493_, new_n23494_, new_n23495_,
    new_n23496_, new_n23497_, new_n23498_, new_n23499_, new_n23500_,
    new_n23501_, new_n23502_, new_n23503_, new_n23504_, new_n23505_,
    new_n23506_, new_n23507_, new_n23508_, new_n23509_, new_n23510_,
    new_n23511_, new_n23512_, new_n23513_, new_n23514_, new_n23515_,
    new_n23516_, new_n23517_, new_n23518_, new_n23519_, new_n23520_,
    new_n23521_, new_n23522_, new_n23523_, new_n23524_, new_n23525_,
    new_n23526_, new_n23527_, new_n23528_, new_n23529_, new_n23530_,
    new_n23531_, new_n23532_, new_n23533_, new_n23534_, new_n23535_,
    new_n23536_, new_n23537_, new_n23538_, new_n23539_, new_n23540_,
    new_n23541_, new_n23542_, new_n23543_, new_n23544_, new_n23545_,
    new_n23546_, new_n23547_, new_n23548_, new_n23549_, new_n23550_,
    new_n23551_, new_n23552_, new_n23553_, new_n23554_, new_n23555_,
    new_n23556_, new_n23557_, new_n23558_, new_n23559_, new_n23560_,
    new_n23561_, new_n23562_, new_n23563_, new_n23564_, new_n23565_,
    new_n23566_, new_n23567_, new_n23568_, new_n23569_, new_n23570_,
    new_n23571_, new_n23572_, new_n23573_, new_n23574_, new_n23575_,
    new_n23576_, new_n23577_, new_n23578_, new_n23579_, new_n23580_,
    new_n23581_, new_n23582_, new_n23583_, new_n23584_, new_n23585_,
    new_n23586_, new_n23587_, new_n23588_, new_n23589_, new_n23590_,
    new_n23591_, new_n23592_, new_n23593_, new_n23594_, new_n23595_,
    new_n23596_, new_n23597_, new_n23598_, new_n23599_, new_n23600_,
    new_n23601_, new_n23602_, new_n23603_, new_n23604_, new_n23605_,
    new_n23606_, new_n23607_, new_n23608_, new_n23609_, new_n23610_,
    new_n23611_, new_n23612_, new_n23613_, new_n23614_, new_n23615_,
    new_n23616_, new_n23617_, new_n23618_, new_n23619_, new_n23620_,
    new_n23621_, new_n23622_, new_n23624_, new_n23625_, new_n23626_,
    new_n23627_, new_n23628_, new_n23629_, new_n23630_, new_n23631_,
    new_n23632_, new_n23633_, new_n23634_, new_n23635_, new_n23636_,
    new_n23637_, new_n23638_, new_n23639_, new_n23640_, new_n23641_,
    new_n23642_, new_n23643_, new_n23644_, new_n23645_, new_n23646_,
    new_n23647_, new_n23648_, new_n23649_, new_n23650_, new_n23651_,
    new_n23652_, new_n23653_, new_n23654_, new_n23655_, new_n23656_,
    new_n23657_, new_n23658_, new_n23659_, new_n23660_, new_n23661_,
    new_n23662_, new_n23663_, new_n23664_, new_n23665_, new_n23666_,
    new_n23667_, new_n23668_, new_n23669_, new_n23670_, new_n23671_,
    new_n23672_, new_n23673_, new_n23674_, new_n23675_, new_n23676_,
    new_n23677_, new_n23678_, new_n23679_, new_n23680_, new_n23681_,
    new_n23682_, new_n23683_, new_n23684_, new_n23685_, new_n23686_,
    new_n23687_, new_n23688_, new_n23689_, new_n23690_, new_n23691_,
    new_n23692_, new_n23693_, new_n23694_, new_n23695_, new_n23696_,
    new_n23697_, new_n23698_, new_n23699_, new_n23700_, new_n23701_,
    new_n23702_, new_n23703_, new_n23704_, new_n23705_, new_n23706_,
    new_n23707_, new_n23708_, new_n23709_, new_n23710_, new_n23711_,
    new_n23712_, new_n23713_, new_n23714_, new_n23715_, new_n23716_,
    new_n23717_, new_n23718_, new_n23719_, new_n23720_, new_n23721_,
    new_n23722_, new_n23723_, new_n23724_, new_n23725_, new_n23726_,
    new_n23727_, new_n23728_, new_n23729_, new_n23730_, new_n23731_,
    new_n23732_, new_n23733_, new_n23734_, new_n23735_, new_n23736_,
    new_n23737_, new_n23738_, new_n23739_, new_n23740_, new_n23741_,
    new_n23742_, new_n23743_, new_n23744_, new_n23745_, new_n23746_,
    new_n23747_, new_n23748_, new_n23749_, new_n23750_, new_n23751_,
    new_n23752_, new_n23753_, new_n23754_, new_n23755_, new_n23756_,
    new_n23757_, new_n23758_, new_n23759_, new_n23760_, new_n23761_,
    new_n23762_, new_n23763_, new_n23764_, new_n23765_, new_n23766_,
    new_n23767_, new_n23768_, new_n23769_, new_n23770_, new_n23771_,
    new_n23772_, new_n23773_, new_n23774_, new_n23775_, new_n23776_,
    new_n23777_, new_n23778_, new_n23779_, new_n23780_, new_n23781_,
    new_n23782_, new_n23783_, new_n23784_, new_n23785_, new_n23786_,
    new_n23787_, new_n23788_, new_n23789_, new_n23790_, new_n23791_,
    new_n23792_, new_n23793_, new_n23794_, new_n23795_, new_n23796_,
    new_n23797_, new_n23798_, new_n23799_, new_n23800_, new_n23801_,
    new_n23802_, new_n23803_, new_n23804_, new_n23805_, new_n23806_,
    new_n23807_, new_n23808_, new_n23809_, new_n23810_, new_n23811_,
    new_n23812_, new_n23813_, new_n23814_, new_n23815_, new_n23816_,
    new_n23817_, new_n23818_, new_n23819_, new_n23820_, new_n23821_,
    new_n23822_, new_n23823_, new_n23824_, new_n23825_, new_n23826_,
    new_n23827_, new_n23828_, new_n23829_, new_n23830_, new_n23831_,
    new_n23832_, new_n23833_, new_n23834_, new_n23835_, new_n23836_,
    new_n23837_, new_n23838_, new_n23839_, new_n23840_, new_n23841_,
    new_n23842_, new_n23843_, new_n23844_, new_n23845_, new_n23846_,
    new_n23847_, new_n23848_, new_n23849_, new_n23850_, new_n23851_,
    new_n23852_, new_n23853_, new_n23854_, new_n23855_, new_n23856_,
    new_n23857_, new_n23858_, new_n23859_, new_n23860_, new_n23861_,
    new_n23862_, new_n23863_, new_n23864_, new_n23865_, new_n23866_,
    new_n23867_, new_n23868_, new_n23869_, new_n23870_, new_n23871_,
    new_n23872_, new_n23873_, new_n23874_, new_n23875_, new_n23876_,
    new_n23877_, new_n23878_, new_n23879_, new_n23880_, new_n23881_,
    new_n23882_, new_n23883_, new_n23884_, new_n23885_, new_n23886_,
    new_n23887_, new_n23888_, new_n23889_, new_n23890_, new_n23891_,
    new_n23892_, new_n23893_, new_n23894_, new_n23895_, new_n23896_,
    new_n23897_, new_n23898_, new_n23899_, new_n23900_, new_n23901_,
    new_n23902_, new_n23903_, new_n23904_, new_n23905_, new_n23906_,
    new_n23907_, new_n23908_, new_n23909_, new_n23910_, new_n23911_,
    new_n23912_, new_n23913_, new_n23914_, new_n23915_, new_n23916_,
    new_n23917_, new_n23918_, new_n23919_, new_n23920_, new_n23921_,
    new_n23922_, new_n23923_, new_n23924_, new_n23925_, new_n23926_,
    new_n23927_, new_n23928_, new_n23929_, new_n23930_, new_n23931_,
    new_n23932_, new_n23933_, new_n23934_, new_n23935_, new_n23936_,
    new_n23937_, new_n23938_, new_n23939_, new_n23940_, new_n23941_,
    new_n23942_, new_n23943_, new_n23944_, new_n23945_, new_n23946_,
    new_n23947_, new_n23948_, new_n23949_, new_n23950_, new_n23951_,
    new_n23952_, new_n23953_, new_n23954_, new_n23955_, new_n23956_,
    new_n23957_, new_n23958_, new_n23959_, new_n23960_, new_n23961_,
    new_n23962_, new_n23963_, new_n23964_, new_n23965_, new_n23966_,
    new_n23967_, new_n23968_, new_n23969_, new_n23970_, new_n23971_,
    new_n23972_, new_n23973_, new_n23974_, new_n23975_, new_n23976_,
    new_n23977_, new_n23978_, new_n23979_, new_n23980_, new_n23981_,
    new_n23982_, new_n23983_, new_n23984_, new_n23985_, new_n23986_,
    new_n23987_, new_n23988_, new_n23989_, new_n23990_, new_n23991_,
    new_n23992_, new_n23993_, new_n23994_, new_n23995_, new_n23996_,
    new_n23997_, new_n23998_, new_n23999_, new_n24000_, new_n24001_,
    new_n24002_, new_n24003_, new_n24004_, new_n24005_, new_n24006_,
    new_n24007_, new_n24008_, new_n24009_, new_n24010_, new_n24011_,
    new_n24012_, new_n24013_, new_n24014_, new_n24015_, new_n24016_,
    new_n24017_, new_n24018_, new_n24019_, new_n24020_, new_n24021_,
    new_n24022_, new_n24023_, new_n24024_, new_n24025_, new_n24026_,
    new_n24027_, new_n24028_, new_n24029_, new_n24030_, new_n24031_,
    new_n24032_, new_n24033_, new_n24034_, new_n24035_, new_n24036_,
    new_n24037_, new_n24038_, new_n24039_, new_n24040_, new_n24041_,
    new_n24042_, new_n24043_, new_n24044_, new_n24045_, new_n24046_,
    new_n24047_, new_n24048_, new_n24049_, new_n24050_, new_n24051_,
    new_n24052_, new_n24053_, new_n24054_, new_n24055_, new_n24056_,
    new_n24057_, new_n24058_, new_n24059_, new_n24060_, new_n24061_,
    new_n24062_, new_n24063_, new_n24064_, new_n24065_, new_n24066_,
    new_n24067_, new_n24068_, new_n24069_, new_n24070_, new_n24071_,
    new_n24072_, new_n24073_, new_n24074_, new_n24075_, new_n24076_,
    new_n24077_, new_n24078_, new_n24079_, new_n24080_, new_n24081_,
    new_n24082_, new_n24083_, new_n24084_, new_n24085_, new_n24086_,
    new_n24087_, new_n24088_, new_n24089_, new_n24090_, new_n24091_,
    new_n24092_, new_n24093_, new_n24094_, new_n24095_, new_n24096_,
    new_n24097_, new_n24098_, new_n24099_, new_n24100_, new_n24101_,
    new_n24102_, new_n24103_, new_n24104_, new_n24105_, new_n24106_,
    new_n24107_, new_n24108_, new_n24109_, new_n24110_, new_n24111_,
    new_n24112_, new_n24113_, new_n24114_, new_n24115_, new_n24116_,
    new_n24117_, new_n24118_, new_n24119_, new_n24120_, new_n24121_,
    new_n24122_, new_n24123_, new_n24124_, new_n24125_, new_n24126_,
    new_n24127_, new_n24128_, new_n24129_, new_n24130_, new_n24131_,
    new_n24132_, new_n24133_, new_n24134_, new_n24135_, new_n24136_,
    new_n24137_, new_n24138_, new_n24139_, new_n24140_, new_n24141_,
    new_n24142_, new_n24143_, new_n24144_, new_n24145_, new_n24146_,
    new_n24147_, new_n24148_, new_n24149_, new_n24150_, new_n24151_,
    new_n24152_, new_n24153_, new_n24154_, new_n24155_, new_n24156_,
    new_n24157_, new_n24158_, new_n24159_, new_n24160_, new_n24161_,
    new_n24162_, new_n24163_, new_n24164_, new_n24165_, new_n24166_,
    new_n24167_, new_n24168_, new_n24169_, new_n24170_, new_n24171_,
    new_n24172_, new_n24173_, new_n24174_, new_n24175_, new_n24176_,
    new_n24177_, new_n24178_, new_n24179_, new_n24180_, new_n24181_,
    new_n24182_, new_n24183_, new_n24184_, new_n24185_, new_n24186_,
    new_n24187_, new_n24188_, new_n24189_, new_n24190_, new_n24191_,
    new_n24192_, new_n24193_, new_n24194_, new_n24195_, new_n24196_,
    new_n24197_, new_n24198_, new_n24199_, new_n24200_, new_n24201_,
    new_n24202_, new_n24203_, new_n24204_, new_n24205_, new_n24206_,
    new_n24207_, new_n24208_, new_n24209_, new_n24210_, new_n24211_,
    new_n24212_, new_n24213_, new_n24214_, new_n24215_, new_n24216_,
    new_n24217_, new_n24218_, new_n24219_, new_n24220_, new_n24221_,
    new_n24222_, new_n24223_, new_n24224_, new_n24225_, new_n24226_,
    new_n24227_, new_n24228_, new_n24229_, new_n24230_, new_n24231_,
    new_n24232_, new_n24233_, new_n24234_, new_n24235_, new_n24236_,
    new_n24237_, new_n24238_, new_n24239_, new_n24240_, new_n24241_,
    new_n24242_, new_n24243_, new_n24244_, new_n24245_, new_n24246_,
    new_n24247_, new_n24248_, new_n24249_, new_n24250_, new_n24251_,
    new_n24252_, new_n24253_, new_n24254_, new_n24255_, new_n24256_,
    new_n24257_, new_n24258_, new_n24259_, new_n24260_, new_n24261_,
    new_n24262_, new_n24263_, new_n24264_, new_n24265_, new_n24266_,
    new_n24267_, new_n24268_, new_n24269_, new_n24270_, new_n24271_,
    new_n24272_, new_n24273_, new_n24274_, new_n24275_, new_n24276_,
    new_n24277_, new_n24278_, new_n24279_, new_n24280_, new_n24281_,
    new_n24282_, new_n24283_, new_n24284_, new_n24285_, new_n24286_,
    new_n24287_, new_n24288_, new_n24289_, new_n24290_, new_n24291_,
    new_n24292_, new_n24293_, new_n24294_, new_n24295_, new_n24296_,
    new_n24297_, new_n24298_, new_n24299_, new_n24300_, new_n24301_,
    new_n24302_, new_n24303_, new_n24304_, new_n24305_, new_n24306_,
    new_n24307_, new_n24308_, new_n24309_, new_n24310_, new_n24311_,
    new_n24312_, new_n24313_, new_n24314_, new_n24315_, new_n24316_,
    new_n24317_, new_n24318_, new_n24319_, new_n24320_, new_n24321_,
    new_n24322_, new_n24323_, new_n24324_, new_n24325_, new_n24326_,
    new_n24327_, new_n24328_, new_n24329_, new_n24330_, new_n24331_,
    new_n24332_, new_n24333_, new_n24334_, new_n24335_, new_n24336_,
    new_n24337_, new_n24338_, new_n24339_, new_n24340_, new_n24341_,
    new_n24342_, new_n24343_, new_n24344_, new_n24345_, new_n24346_,
    new_n24347_, new_n24348_, new_n24349_, new_n24350_, new_n24351_,
    new_n24352_, new_n24353_, new_n24354_, new_n24355_, new_n24356_,
    new_n24357_, new_n24358_, new_n24359_, new_n24360_, new_n24361_,
    new_n24362_, new_n24363_, new_n24364_, new_n24365_, new_n24366_,
    new_n24367_, new_n24368_, new_n24369_, new_n24370_, new_n24371_,
    new_n24372_, new_n24373_, new_n24374_, new_n24375_, new_n24376_,
    new_n24377_, new_n24378_, new_n24379_, new_n24380_, new_n24381_,
    new_n24383_, new_n24384_, new_n24385_, new_n24386_, new_n24387_,
    new_n24388_, new_n24389_, new_n24390_, new_n24391_, new_n24392_,
    new_n24393_, new_n24394_, new_n24395_, new_n24396_, new_n24397_,
    new_n24398_, new_n24399_, new_n24400_, new_n24401_, new_n24402_,
    new_n24403_, new_n24404_, new_n24405_, new_n24406_, new_n24407_,
    new_n24408_, new_n24409_, new_n24410_, new_n24411_, new_n24412_,
    new_n24413_, new_n24414_, new_n24415_, new_n24416_, new_n24417_,
    new_n24418_, new_n24419_, new_n24420_, new_n24421_, new_n24422_,
    new_n24423_, new_n24424_, new_n24425_, new_n24426_, new_n24427_,
    new_n24428_, new_n24429_, new_n24430_, new_n24431_, new_n24432_,
    new_n24433_, new_n24434_, new_n24435_, new_n24436_, new_n24437_,
    new_n24438_, new_n24439_, new_n24440_, new_n24441_, new_n24442_,
    new_n24443_, new_n24444_, new_n24445_, new_n24446_, new_n24447_,
    new_n24448_, new_n24449_, new_n24450_, new_n24451_, new_n24452_,
    new_n24453_, new_n24454_, new_n24455_, new_n24456_, new_n24457_,
    new_n24458_, new_n24459_, new_n24460_, new_n24461_, new_n24462_,
    new_n24463_, new_n24464_, new_n24465_, new_n24466_, new_n24467_,
    new_n24468_, new_n24469_, new_n24470_, new_n24471_, new_n24472_,
    new_n24473_, new_n24474_, new_n24475_, new_n24476_, new_n24477_,
    new_n24478_, new_n24479_, new_n24480_, new_n24481_, new_n24482_,
    new_n24483_, new_n24484_, new_n24485_, new_n24486_, new_n24487_,
    new_n24488_, new_n24489_, new_n24490_, new_n24491_, new_n24492_,
    new_n24493_, new_n24494_, new_n24495_, new_n24496_, new_n24497_,
    new_n24498_, new_n24499_, new_n24500_, new_n24501_, new_n24502_,
    new_n24503_, new_n24504_, new_n24505_, new_n24506_, new_n24507_,
    new_n24508_, new_n24509_, new_n24510_, new_n24511_, new_n24512_,
    new_n24513_, new_n24514_, new_n24515_, new_n24516_, new_n24517_,
    new_n24518_, new_n24519_, new_n24520_, new_n24521_, new_n24522_,
    new_n24523_, new_n24524_, new_n24525_, new_n24526_, new_n24527_,
    new_n24528_, new_n24529_, new_n24530_, new_n24531_, new_n24532_,
    new_n24533_, new_n24534_, new_n24535_, new_n24536_, new_n24537_,
    new_n24538_, new_n24539_, new_n24540_, new_n24541_, new_n24542_,
    new_n24543_, new_n24544_, new_n24545_, new_n24546_, new_n24547_,
    new_n24548_, new_n24549_, new_n24550_, new_n24551_, new_n24552_,
    new_n24553_, new_n24554_, new_n24555_, new_n24556_, new_n24557_,
    new_n24558_, new_n24559_, new_n24560_, new_n24561_, new_n24562_,
    new_n24563_, new_n24564_, new_n24565_, new_n24566_, new_n24567_,
    new_n24568_, new_n24569_, new_n24570_, new_n24571_, new_n24572_,
    new_n24573_, new_n24574_, new_n24575_, new_n24576_, new_n24577_,
    new_n24578_, new_n24579_, new_n24580_, new_n24581_, new_n24582_,
    new_n24583_, new_n24584_, new_n24585_, new_n24586_, new_n24587_,
    new_n24588_, new_n24589_, new_n24590_, new_n24591_, new_n24592_,
    new_n24593_, new_n24594_, new_n24595_, new_n24596_, new_n24597_,
    new_n24598_, new_n24599_, new_n24600_, new_n24601_, new_n24602_,
    new_n24603_, new_n24604_, new_n24605_, new_n24606_, new_n24607_,
    new_n24608_, new_n24609_, new_n24610_, new_n24611_, new_n24612_,
    new_n24613_, new_n24614_, new_n24615_, new_n24616_, new_n24617_,
    new_n24618_, new_n24619_, new_n24620_, new_n24621_, new_n24622_,
    new_n24623_, new_n24624_, new_n24625_, new_n24626_, new_n24627_,
    new_n24628_, new_n24629_, new_n24630_, new_n24631_, new_n24632_,
    new_n24633_, new_n24634_, new_n24635_, new_n24636_, new_n24637_,
    new_n24638_, new_n24639_, new_n24640_, new_n24641_, new_n24642_,
    new_n24643_, new_n24644_, new_n24645_, new_n24646_, new_n24647_,
    new_n24648_, new_n24649_, new_n24650_, new_n24651_, new_n24652_,
    new_n24653_, new_n24654_, new_n24655_, new_n24656_, new_n24657_,
    new_n24658_, new_n24659_, new_n24660_, new_n24661_, new_n24662_,
    new_n24663_, new_n24664_, new_n24665_, new_n24666_, new_n24667_,
    new_n24668_, new_n24669_, new_n24670_, new_n24671_, new_n24672_,
    new_n24673_, new_n24674_, new_n24675_, new_n24676_, new_n24677_,
    new_n24678_, new_n24679_, new_n24680_, new_n24681_, new_n24682_,
    new_n24683_, new_n24684_, new_n24685_, new_n24686_, new_n24687_,
    new_n24688_, new_n24689_, new_n24690_, new_n24691_, new_n24692_,
    new_n24693_, new_n24694_, new_n24695_, new_n24696_, new_n24697_,
    new_n24698_, new_n24699_, new_n24700_, new_n24701_, new_n24702_,
    new_n24703_, new_n24704_, new_n24705_, new_n24706_, new_n24707_,
    new_n24708_, new_n24709_, new_n24710_, new_n24711_, new_n24712_,
    new_n24713_, new_n24714_, new_n24715_, new_n24716_, new_n24717_,
    new_n24718_, new_n24719_, new_n24720_, new_n24721_, new_n24722_,
    new_n24723_, new_n24724_, new_n24725_, new_n24726_, new_n24727_,
    new_n24728_, new_n24729_, new_n24730_, new_n24731_, new_n24732_,
    new_n24733_, new_n24734_, new_n24735_, new_n24736_, new_n24737_,
    new_n24738_, new_n24739_, new_n24740_, new_n24741_, new_n24742_,
    new_n24743_, new_n24744_, new_n24745_, new_n24746_, new_n24747_,
    new_n24748_, new_n24749_, new_n24750_, new_n24751_, new_n24752_,
    new_n24753_, new_n24754_, new_n24755_, new_n24756_, new_n24757_,
    new_n24758_, new_n24759_, new_n24760_, new_n24761_, new_n24762_,
    new_n24763_, new_n24764_, new_n24765_, new_n24766_, new_n24767_,
    new_n24768_, new_n24769_, new_n24770_, new_n24771_, new_n24772_,
    new_n24773_, new_n24774_, new_n24775_, new_n24776_, new_n24777_,
    new_n24778_, new_n24779_, new_n24780_, new_n24781_, new_n24782_,
    new_n24783_, new_n24784_, new_n24785_, new_n24786_, new_n24787_,
    new_n24788_, new_n24789_, new_n24790_, new_n24791_, new_n24792_,
    new_n24793_, new_n24794_, new_n24795_, new_n24796_, new_n24797_,
    new_n24798_, new_n24799_, new_n24800_, new_n24801_, new_n24802_,
    new_n24803_, new_n24804_, new_n24805_, new_n24806_, new_n24807_,
    new_n24808_, new_n24809_, new_n24810_, new_n24811_, new_n24812_,
    new_n24813_, new_n24814_, new_n24815_, new_n24816_, new_n24817_,
    new_n24818_, new_n24819_, new_n24820_, new_n24821_, new_n24822_,
    new_n24823_, new_n24824_, new_n24825_, new_n24826_, new_n24827_,
    new_n24828_, new_n24829_, new_n24830_, new_n24831_, new_n24832_,
    new_n24833_, new_n24834_, new_n24835_, new_n24836_, new_n24837_,
    new_n24838_, new_n24839_, new_n24840_, new_n24841_, new_n24842_,
    new_n24843_, new_n24844_, new_n24845_, new_n24846_, new_n24847_,
    new_n24848_, new_n24849_, new_n24850_, new_n24851_, new_n24852_,
    new_n24853_, new_n24854_, new_n24855_, new_n24856_, new_n24857_,
    new_n24858_, new_n24859_, new_n24860_, new_n24861_, new_n24862_,
    new_n24863_, new_n24864_, new_n24865_, new_n24866_, new_n24867_,
    new_n24868_, new_n24869_, new_n24870_, new_n24871_, new_n24872_,
    new_n24873_, new_n24874_, new_n24875_, new_n24876_, new_n24877_,
    new_n24878_, new_n24879_, new_n24880_, new_n24881_, new_n24882_,
    new_n24883_, new_n24884_, new_n24885_, new_n24886_, new_n24887_,
    new_n24888_, new_n24889_, new_n24890_, new_n24891_, new_n24892_,
    new_n24893_, new_n24894_, new_n24895_, new_n24896_, new_n24897_,
    new_n24898_, new_n24899_, new_n24900_, new_n24901_, new_n24902_,
    new_n24903_, new_n24904_, new_n24905_, new_n24906_, new_n24907_,
    new_n24908_, new_n24909_, new_n24910_, new_n24911_, new_n24912_,
    new_n24913_, new_n24914_, new_n24915_, new_n24916_, new_n24917_,
    new_n24918_, new_n24919_, new_n24920_, new_n24921_, new_n24922_,
    new_n24923_, new_n24924_, new_n24925_, new_n24926_, new_n24927_,
    new_n24928_, new_n24929_, new_n24930_, new_n24931_, new_n24932_,
    new_n24933_, new_n24934_, new_n24935_, new_n24936_, new_n24937_,
    new_n24938_, new_n24939_, new_n24940_, new_n24941_, new_n24942_,
    new_n24943_, new_n24944_, new_n24945_, new_n24946_, new_n24947_,
    new_n24948_, new_n24949_, new_n24950_, new_n24951_, new_n24952_,
    new_n24953_, new_n24954_, new_n24955_, new_n24956_, new_n24957_,
    new_n24958_, new_n24959_, new_n24960_, new_n24961_, new_n24962_,
    new_n24963_, new_n24964_, new_n24965_, new_n24966_, new_n24967_,
    new_n24968_, new_n24969_, new_n24970_, new_n24971_, new_n24972_,
    new_n24973_, new_n24974_, new_n24975_, new_n24976_, new_n24977_,
    new_n24978_, new_n24979_, new_n24980_, new_n24981_, new_n24982_,
    new_n24983_, new_n24984_, new_n24985_, new_n24986_, new_n24987_,
    new_n24988_, new_n24989_, new_n24990_, new_n24991_, new_n24992_,
    new_n24993_, new_n24994_, new_n24995_, new_n24996_, new_n24997_,
    new_n24998_, new_n24999_, new_n25000_, new_n25001_, new_n25002_,
    new_n25003_, new_n25004_, new_n25005_, new_n25006_, new_n25007_,
    new_n25008_, new_n25009_, new_n25010_, new_n25011_, new_n25012_,
    new_n25013_, new_n25014_, new_n25015_, new_n25016_, new_n25017_,
    new_n25018_, new_n25019_, new_n25020_, new_n25021_, new_n25022_,
    new_n25023_, new_n25024_, new_n25025_, new_n25026_, new_n25027_,
    new_n25028_, new_n25029_, new_n25030_, new_n25031_, new_n25032_,
    new_n25033_, new_n25034_, new_n25035_, new_n25036_, new_n25037_,
    new_n25038_, new_n25039_, new_n25040_, new_n25041_, new_n25042_,
    new_n25043_, new_n25044_, new_n25045_, new_n25046_, new_n25047_,
    new_n25048_, new_n25049_, new_n25050_, new_n25051_, new_n25052_,
    new_n25053_, new_n25054_, new_n25055_, new_n25056_, new_n25057_,
    new_n25058_, new_n25059_, new_n25060_, new_n25061_, new_n25062_,
    new_n25063_, new_n25064_, new_n25065_, new_n25066_, new_n25067_,
    new_n25068_, new_n25069_, new_n25070_, new_n25071_, new_n25072_,
    new_n25073_, new_n25074_, new_n25075_, new_n25076_, new_n25077_,
    new_n25078_, new_n25079_, new_n25080_, new_n25081_, new_n25082_,
    new_n25083_, new_n25084_, new_n25085_, new_n25086_, new_n25087_,
    new_n25088_, new_n25089_, new_n25090_, new_n25091_, new_n25092_,
    new_n25093_, new_n25094_, new_n25095_, new_n25096_, new_n25097_,
    new_n25098_, new_n25099_, new_n25100_, new_n25101_, new_n25102_,
    new_n25103_, new_n25104_, new_n25105_, new_n25106_, new_n25107_,
    new_n25108_, new_n25109_, new_n25110_, new_n25111_, new_n25112_,
    new_n25113_, new_n25114_, new_n25115_, new_n25116_, new_n25117_,
    new_n25118_, new_n25119_, new_n25120_, new_n25121_, new_n25122_,
    new_n25123_, new_n25124_, new_n25125_, new_n25126_, new_n25127_,
    new_n25128_, new_n25129_, new_n25130_, new_n25131_, new_n25132_,
    new_n25133_, new_n25134_, new_n25135_, new_n25136_, new_n25137_,
    new_n25138_, new_n25139_, new_n25140_, new_n25141_, new_n25142_,
    new_n25143_, new_n25144_, new_n25145_, new_n25146_, new_n25147_,
    new_n25148_, new_n25149_, new_n25150_, new_n25151_, new_n25152_,
    new_n25153_, new_n25154_, new_n25155_, new_n25156_, new_n25157_,
    new_n25158_, new_n25159_, new_n25160_, new_n25161_, new_n25162_,
    new_n25163_, new_n25164_, new_n25165_, new_n25166_, new_n25167_,
    new_n25168_, new_n25169_, new_n25170_, new_n25171_, new_n25172_,
    new_n25173_, new_n25174_, new_n25175_, new_n25176_, new_n25177_,
    new_n25178_, new_n25179_, new_n25180_, new_n25181_, new_n25182_,
    new_n25183_, new_n25184_, new_n25185_, new_n25186_, new_n25187_,
    new_n25188_, new_n25189_, new_n25190_, new_n25191_, new_n25192_,
    new_n25193_, new_n25194_, new_n25195_, new_n25196_, new_n25197_,
    new_n25198_, new_n25199_, new_n25200_, new_n25201_, new_n25202_,
    new_n25203_, new_n25204_, new_n25205_, new_n25206_, new_n25207_,
    new_n25208_, new_n25209_, new_n25211_, new_n25212_, new_n25213_,
    new_n25214_, new_n25215_, new_n25216_, new_n25217_, new_n25218_,
    new_n25219_, new_n25220_, new_n25221_, new_n25222_, new_n25223_,
    new_n25224_, new_n25225_, new_n25226_, new_n25227_, new_n25228_,
    new_n25229_, new_n25230_, new_n25231_, new_n25232_, new_n25233_,
    new_n25234_, new_n25235_, new_n25236_, new_n25237_, new_n25238_,
    new_n25239_, new_n25240_, new_n25241_, new_n25242_, new_n25243_,
    new_n25244_, new_n25245_, new_n25246_, new_n25247_, new_n25248_,
    new_n25249_, new_n25250_, new_n25251_, new_n25252_, new_n25253_,
    new_n25254_, new_n25255_, new_n25256_, new_n25257_, new_n25258_,
    new_n25259_, new_n25260_, new_n25261_, new_n25262_, new_n25263_,
    new_n25264_, new_n25265_, new_n25266_, new_n25267_, new_n25268_,
    new_n25269_, new_n25270_, new_n25271_, new_n25272_, new_n25273_,
    new_n25274_, new_n25275_, new_n25276_, new_n25277_, new_n25278_,
    new_n25279_, new_n25280_, new_n25281_, new_n25282_, new_n25283_,
    new_n25284_, new_n25285_, new_n25286_, new_n25287_, new_n25288_,
    new_n25289_, new_n25290_, new_n25291_, new_n25292_, new_n25293_,
    new_n25294_, new_n25295_, new_n25296_, new_n25297_, new_n25298_,
    new_n25299_, new_n25300_, new_n25301_, new_n25302_, new_n25303_,
    new_n25304_, new_n25305_, new_n25306_, new_n25307_, new_n25308_,
    new_n25309_, new_n25310_, new_n25311_, new_n25312_, new_n25313_,
    new_n25314_, new_n25315_, new_n25316_, new_n25317_, new_n25318_,
    new_n25319_, new_n25320_, new_n25321_, new_n25322_, new_n25323_,
    new_n25324_, new_n25325_, new_n25326_, new_n25327_, new_n25328_,
    new_n25329_, new_n25330_, new_n25331_, new_n25332_, new_n25333_,
    new_n25334_, new_n25335_, new_n25336_, new_n25337_, new_n25338_,
    new_n25339_, new_n25340_, new_n25341_, new_n25342_, new_n25343_,
    new_n25344_, new_n25345_, new_n25346_, new_n25347_, new_n25348_,
    new_n25349_, new_n25350_, new_n25351_, new_n25352_, new_n25353_,
    new_n25354_, new_n25355_, new_n25356_, new_n25357_, new_n25358_,
    new_n25359_, new_n25360_, new_n25361_, new_n25362_, new_n25363_,
    new_n25364_, new_n25365_, new_n25366_, new_n25367_, new_n25368_,
    new_n25369_, new_n25370_, new_n25371_, new_n25372_, new_n25373_,
    new_n25374_, new_n25375_, new_n25376_, new_n25377_, new_n25378_,
    new_n25379_, new_n25380_, new_n25381_, new_n25382_, new_n25383_,
    new_n25384_, new_n25385_, new_n25386_, new_n25387_, new_n25388_,
    new_n25389_, new_n25390_, new_n25391_, new_n25392_, new_n25393_,
    new_n25394_, new_n25395_, new_n25396_, new_n25397_, new_n25398_,
    new_n25399_, new_n25400_, new_n25401_, new_n25402_, new_n25403_,
    new_n25404_, new_n25405_, new_n25406_, new_n25407_, new_n25408_,
    new_n25409_, new_n25410_, new_n25411_, new_n25412_, new_n25413_,
    new_n25414_, new_n25415_, new_n25416_, new_n25417_, new_n25418_,
    new_n25419_, new_n25420_, new_n25421_, new_n25422_, new_n25423_,
    new_n25424_, new_n25425_, new_n25426_, new_n25427_, new_n25428_,
    new_n25429_, new_n25430_, new_n25431_, new_n25432_, new_n25433_,
    new_n25434_, new_n25435_, new_n25436_, new_n25437_, new_n25438_,
    new_n25439_, new_n25440_, new_n25441_, new_n25442_, new_n25443_,
    new_n25444_, new_n25445_, new_n25446_, new_n25447_, new_n25448_,
    new_n25449_, new_n25450_, new_n25451_, new_n25452_, new_n25453_,
    new_n25454_, new_n25455_, new_n25456_, new_n25457_, new_n25458_,
    new_n25459_, new_n25460_, new_n25461_, new_n25462_, new_n25463_,
    new_n25464_, new_n25465_, new_n25466_, new_n25467_, new_n25468_,
    new_n25469_, new_n25470_, new_n25471_, new_n25472_, new_n25473_,
    new_n25474_, new_n25475_, new_n25476_, new_n25477_, new_n25478_,
    new_n25479_, new_n25480_, new_n25481_, new_n25482_, new_n25483_,
    new_n25484_, new_n25485_, new_n25486_, new_n25487_, new_n25488_,
    new_n25489_, new_n25490_, new_n25491_, new_n25492_, new_n25493_,
    new_n25494_, new_n25495_, new_n25496_, new_n25497_, new_n25498_,
    new_n25499_, new_n25500_, new_n25501_, new_n25502_, new_n25503_,
    new_n25504_, new_n25505_, new_n25506_, new_n25507_, new_n25508_,
    new_n25509_, new_n25510_, new_n25511_, new_n25512_, new_n25513_,
    new_n25514_, new_n25515_, new_n25516_, new_n25517_, new_n25518_,
    new_n25519_, new_n25520_, new_n25521_, new_n25522_, new_n25523_,
    new_n25524_, new_n25525_, new_n25526_, new_n25527_, new_n25528_,
    new_n25529_, new_n25530_, new_n25531_, new_n25532_, new_n25533_,
    new_n25534_, new_n25535_, new_n25536_, new_n25537_, new_n25538_,
    new_n25539_, new_n25540_, new_n25541_, new_n25542_, new_n25543_,
    new_n25544_, new_n25545_, new_n25546_, new_n25547_, new_n25548_,
    new_n25549_, new_n25550_, new_n25551_, new_n25552_, new_n25553_,
    new_n25554_, new_n25555_, new_n25556_, new_n25557_, new_n25558_,
    new_n25559_, new_n25560_, new_n25561_, new_n25562_, new_n25563_,
    new_n25564_, new_n25565_, new_n25566_, new_n25567_, new_n25568_,
    new_n25569_, new_n25570_, new_n25571_, new_n25572_, new_n25573_,
    new_n25574_, new_n25575_, new_n25576_, new_n25577_, new_n25578_,
    new_n25579_, new_n25580_, new_n25581_, new_n25582_, new_n25583_,
    new_n25584_, new_n25585_, new_n25586_, new_n25587_, new_n25588_,
    new_n25589_, new_n25590_, new_n25591_, new_n25592_, new_n25593_,
    new_n25594_, new_n25595_, new_n25596_, new_n25597_, new_n25598_,
    new_n25599_, new_n25600_, new_n25601_, new_n25602_, new_n25603_,
    new_n25604_, new_n25605_, new_n25606_, new_n25607_, new_n25608_,
    new_n25609_, new_n25610_, new_n25611_, new_n25612_, new_n25613_,
    new_n25614_, new_n25615_, new_n25616_, new_n25617_, new_n25618_,
    new_n25619_, new_n25620_, new_n25621_, new_n25622_, new_n25623_,
    new_n25624_, new_n25625_, new_n25626_, new_n25627_, new_n25628_,
    new_n25629_, new_n25630_, new_n25631_, new_n25632_, new_n25633_,
    new_n25634_, new_n25635_, new_n25636_, new_n25637_, new_n25638_,
    new_n25639_, new_n25640_, new_n25641_, new_n25642_, new_n25643_,
    new_n25644_, new_n25645_, new_n25646_, new_n25647_, new_n25648_,
    new_n25649_, new_n25650_, new_n25651_, new_n25652_, new_n25653_,
    new_n25654_, new_n25655_, new_n25656_, new_n25657_, new_n25658_,
    new_n25659_, new_n25660_, new_n25661_, new_n25662_, new_n25663_,
    new_n25664_, new_n25665_, new_n25666_, new_n25667_, new_n25668_,
    new_n25669_, new_n25670_, new_n25671_, new_n25672_, new_n25673_,
    new_n25674_, new_n25675_, new_n25676_, new_n25677_, new_n25678_,
    new_n25679_, new_n25680_, new_n25681_, new_n25682_, new_n25683_,
    new_n25684_, new_n25685_, new_n25686_, new_n25687_, new_n25688_,
    new_n25689_, new_n25690_, new_n25691_, new_n25692_, new_n25693_,
    new_n25694_, new_n25695_, new_n25696_, new_n25697_, new_n25698_,
    new_n25699_, new_n25700_, new_n25701_, new_n25702_, new_n25703_,
    new_n25704_, new_n25705_, new_n25706_, new_n25707_, new_n25708_,
    new_n25709_, new_n25710_, new_n25711_, new_n25712_, new_n25713_,
    new_n25714_, new_n25715_, new_n25716_, new_n25717_, new_n25718_,
    new_n25719_, new_n25720_, new_n25721_, new_n25722_, new_n25723_,
    new_n25724_, new_n25725_, new_n25726_, new_n25727_, new_n25728_,
    new_n25729_, new_n25730_, new_n25731_, new_n25732_, new_n25733_,
    new_n25734_, new_n25735_, new_n25736_, new_n25737_, new_n25738_,
    new_n25739_, new_n25740_, new_n25741_, new_n25742_, new_n25743_,
    new_n25744_, new_n25745_, new_n25746_, new_n25747_, new_n25748_,
    new_n25749_, new_n25750_, new_n25751_, new_n25752_, new_n25753_,
    new_n25754_, new_n25755_, new_n25756_, new_n25757_, new_n25758_,
    new_n25759_, new_n25760_, new_n25761_, new_n25762_, new_n25763_,
    new_n25764_, new_n25765_, new_n25766_, new_n25767_, new_n25768_,
    new_n25769_, new_n25770_, new_n25771_, new_n25772_, new_n25773_,
    new_n25774_, new_n25775_, new_n25776_, new_n25777_, new_n25778_,
    new_n25779_, new_n25780_, new_n25781_, new_n25782_, new_n25783_,
    new_n25784_, new_n25785_, new_n25786_, new_n25787_, new_n25788_,
    new_n25789_, new_n25790_, new_n25791_, new_n25792_, new_n25793_,
    new_n25794_, new_n25795_, new_n25796_, new_n25797_, new_n25798_,
    new_n25799_, new_n25800_, new_n25801_, new_n25802_, new_n25803_,
    new_n25804_, new_n25805_, new_n25806_, new_n25807_, new_n25808_,
    new_n25809_, new_n25810_, new_n25811_, new_n25812_, new_n25813_,
    new_n25814_, new_n25815_, new_n25816_, new_n25817_, new_n25818_,
    new_n25819_, new_n25820_, new_n25821_, new_n25822_, new_n25823_,
    new_n25824_, new_n25825_, new_n25826_, new_n25827_, new_n25828_,
    new_n25829_, new_n25830_, new_n25831_, new_n25832_, new_n25833_,
    new_n25834_, new_n25835_, new_n25836_, new_n25837_, new_n25838_,
    new_n25839_, new_n25840_, new_n25841_, new_n25842_, new_n25843_,
    new_n25844_, new_n25845_, new_n25846_, new_n25847_, new_n25848_,
    new_n25849_, new_n25850_, new_n25851_, new_n25852_, new_n25853_,
    new_n25854_, new_n25855_, new_n25856_, new_n25857_, new_n25858_,
    new_n25859_, new_n25860_, new_n25861_, new_n25862_, new_n25863_,
    new_n25864_, new_n25865_, new_n25866_, new_n25867_, new_n25868_,
    new_n25869_, new_n25870_, new_n25871_, new_n25872_, new_n25873_,
    new_n25874_, new_n25875_, new_n25876_, new_n25877_, new_n25878_,
    new_n25879_, new_n25880_, new_n25881_, new_n25882_, new_n25883_,
    new_n25884_, new_n25885_, new_n25886_, new_n25887_, new_n25888_,
    new_n25889_, new_n25890_, new_n25891_, new_n25892_, new_n25893_,
    new_n25894_, new_n25895_, new_n25896_, new_n25897_, new_n25898_,
    new_n25899_, new_n25900_, new_n25901_, new_n25902_, new_n25903_,
    new_n25904_, new_n25905_, new_n25906_, new_n25907_, new_n25908_,
    new_n25909_, new_n25910_, new_n25911_, new_n25912_, new_n25913_,
    new_n25914_, new_n25915_, new_n25916_, new_n25917_, new_n25918_;
  NOR2X1   g00000(.A(\a[127] ), .B(\a[126] ), .Y(new_n193_));
  OR2X1    g00001(.A(\a[125] ), .B(\a[124] ), .Y(new_n194_));
  MX2X1    g00002(.A(new_n194_), .B(\a[127] ), .S0(\a[126] ), .Y(\asqrt[62] ));
  INVX1    g00003(.A(new_n193_), .Y(\asqrt[63] ));
  INVX1    g00004(.A(\a[127] ), .Y(new_n197_));
  NOR2X1   g00005(.A(\a[125] ), .B(\a[124] ), .Y(new_n198_));
  MX2X1    g00006(.A(new_n198_), .B(new_n197_), .S0(\a[126] ), .Y(new_n199_));
  OR2X1    g00007(.A(\a[123] ), .B(\a[122] ), .Y(new_n200_));
  MX2X1    g00008(.A(new_n200_), .B(new_n199_), .S0(\a[124] ), .Y(new_n201_));
  INVX1    g00009(.A(\a[124] ), .Y(new_n202_));
  INVX1    g00010(.A(\a[125] ), .Y(new_n203_));
  AOI21X1  g00011(.A0(\asqrt[62] ), .A1(new_n202_), .B0(new_n203_), .Y(new_n204_));
  INVX1    g00012(.A(\a[126] ), .Y(new_n205_));
  NOR3X1   g00013(.A(new_n194_), .B(new_n197_), .C(new_n205_), .Y(new_n206_));
  NOR3X1   g00014(.A(new_n206_), .B(new_n204_), .C(new_n201_), .Y(new_n207_));
  OR2X1    g00015(.A(new_n207_), .B(\asqrt[63] ), .Y(new_n208_));
  NOR2X1   g00016(.A(\a[123] ), .B(\a[122] ), .Y(new_n209_));
  MX2X1    g00017(.A(new_n209_), .B(\asqrt[62] ), .S0(\a[124] ), .Y(new_n210_));
  OAI21X1  g00018(.A0(new_n199_), .A1(\a[124] ), .B0(\a[125] ), .Y(new_n211_));
  NAND3X1  g00019(.A(new_n198_), .B(\a[127] ), .C(\a[126] ), .Y(new_n212_));
  AOI21X1  g00020(.A0(new_n212_), .A1(new_n211_), .B0(new_n210_), .Y(new_n213_));
  OAI21X1  g00021(.A0(new_n194_), .A1(new_n205_), .B0(\a[127] ), .Y(new_n214_));
  AOI21X1  g00022(.A0(new_n194_), .A1(new_n205_), .B0(new_n214_), .Y(new_n215_));
  NOR2X1   g00023(.A(new_n215_), .B(new_n213_), .Y(new_n216_));
  AND2X1   g00024(.A(new_n216_), .B(new_n208_), .Y(new_n217_));
  INVX1    g00025(.A(\a[122] ), .Y(new_n218_));
  AOI21X1  g00026(.A0(new_n216_), .A1(new_n208_), .B0(new_n218_), .Y(new_n219_));
  NOR3X1   g00027(.A(\a[122] ), .B(\a[121] ), .C(\a[120] ), .Y(new_n220_));
  OAI21X1  g00028(.A0(new_n220_), .A1(new_n219_), .B0(\asqrt[62] ), .Y(new_n221_));
  OAI21X1  g00029(.A0(\a[125] ), .A1(\a[124] ), .B0(new_n205_), .Y(new_n222_));
  AOI21X1  g00030(.A0(\a[127] ), .A1(\a[126] ), .B0(new_n220_), .Y(new_n223_));
  NAND2X1  g00031(.A(new_n223_), .B(new_n222_), .Y(new_n224_));
  NOR2X1   g00032(.A(new_n224_), .B(new_n219_), .Y(new_n225_));
  INVX1    g00033(.A(\a[123] ), .Y(new_n226_));
  NAND3X1  g00034(.A(new_n212_), .B(new_n211_), .C(new_n210_), .Y(new_n227_));
  AND2X1   g00035(.A(new_n227_), .B(new_n193_), .Y(new_n228_));
  OR2X1    g00036(.A(new_n215_), .B(new_n213_), .Y(new_n229_));
  OAI21X1  g00037(.A0(new_n229_), .A1(new_n228_), .B0(new_n209_), .Y(new_n230_));
  AOI21X1  g00038(.A0(new_n216_), .A1(new_n208_), .B0(\a[122] ), .Y(new_n231_));
  OAI21X1  g00039(.A0(new_n231_), .A1(new_n226_), .B0(new_n230_), .Y(new_n232_));
  OAI21X1  g00040(.A0(new_n232_), .A1(new_n225_), .B0(new_n221_), .Y(new_n233_));
  AOI21X1  g00041(.A0(new_n216_), .A1(new_n208_), .B0(new_n200_), .Y(new_n234_));
  NOR4X1   g00042(.A(new_n215_), .B(new_n213_), .C(new_n228_), .D(new_n199_), .Y(new_n235_));
  OAI21X1  g00043(.A0(new_n235_), .A1(new_n234_), .B0(\a[124] ), .Y(new_n236_));
  OR4X1    g00044(.A(new_n215_), .B(new_n213_), .C(new_n228_), .D(new_n199_), .Y(new_n237_));
  NAND3X1  g00045(.A(new_n237_), .B(new_n230_), .C(new_n202_), .Y(new_n238_));
  AOI21X1  g00046(.A0(new_n216_), .A1(new_n208_), .B0(new_n227_), .Y(new_n239_));
  OR2X1    g00047(.A(new_n239_), .B(new_n213_), .Y(new_n240_));
  AOI21X1  g00048(.A0(new_n238_), .A1(new_n236_), .B0(new_n240_), .Y(new_n241_));
  AOI21X1  g00049(.A0(new_n241_), .A1(new_n233_), .B0(\asqrt[63] ), .Y(new_n242_));
  AOI21X1  g00050(.A0(new_n237_), .A1(new_n230_), .B0(new_n202_), .Y(new_n243_));
  NOR3X1   g00051(.A(new_n235_), .B(new_n234_), .C(\a[124] ), .Y(new_n244_));
  OR2X1    g00052(.A(new_n244_), .B(new_n243_), .Y(new_n245_));
  AND2X1   g00053(.A(new_n212_), .B(new_n211_), .Y(new_n246_));
  OAI21X1  g00054(.A0(new_n229_), .A1(new_n228_), .B0(new_n246_), .Y(new_n247_));
  OR2X1    g00055(.A(new_n207_), .B(new_n193_), .Y(new_n248_));
  AOI21X1  g00056(.A0(new_n247_), .A1(new_n201_), .B0(new_n248_), .Y(new_n249_));
  NOR4X1   g00057(.A(new_n215_), .B(new_n246_), .C(new_n201_), .D(new_n193_), .Y(new_n250_));
  NOR2X1   g00058(.A(new_n250_), .B(new_n249_), .Y(new_n251_));
  OAI21X1  g00059(.A0(new_n245_), .A1(new_n233_), .B0(new_n251_), .Y(new_n252_));
  OR2X1    g00060(.A(new_n252_), .B(new_n242_), .Y(\asqrt[60] ));
  INVX1    g00061(.A(new_n217_), .Y(\asqrt[61] ));
  INVX1    g00062(.A(\a[120] ), .Y(new_n255_));
  OAI21X1  g00063(.A0(new_n229_), .A1(new_n228_), .B0(\a[122] ), .Y(new_n256_));
  INVX1    g00064(.A(new_n220_), .Y(new_n257_));
  AOI21X1  g00065(.A0(new_n257_), .A1(new_n256_), .B0(new_n199_), .Y(new_n258_));
  OR2X1    g00066(.A(new_n224_), .B(new_n219_), .Y(new_n259_));
  OAI21X1  g00067(.A0(new_n229_), .A1(new_n228_), .B0(new_n218_), .Y(new_n260_));
  AOI21X1  g00068(.A0(new_n260_), .A1(\a[123] ), .B0(new_n234_), .Y(new_n261_));
  AOI21X1  g00069(.A0(new_n261_), .A1(new_n259_), .B0(new_n258_), .Y(new_n262_));
  NOR2X1   g00070(.A(new_n239_), .B(new_n213_), .Y(new_n263_));
  OAI21X1  g00071(.A0(new_n244_), .A1(new_n243_), .B0(new_n263_), .Y(new_n264_));
  OAI21X1  g00072(.A0(new_n264_), .A1(new_n262_), .B0(new_n193_), .Y(new_n265_));
  NOR2X1   g00073(.A(new_n244_), .B(new_n243_), .Y(new_n266_));
  OR2X1    g00074(.A(new_n250_), .B(new_n249_), .Y(new_n267_));
  AOI21X1  g00075(.A0(new_n266_), .A1(new_n262_), .B0(new_n267_), .Y(new_n268_));
  AOI21X1  g00076(.A0(new_n268_), .A1(new_n265_), .B0(new_n255_), .Y(new_n269_));
  NOR3X1   g00077(.A(\a[120] ), .B(\a[119] ), .C(\a[118] ), .Y(new_n270_));
  OR2X1    g00078(.A(new_n270_), .B(new_n269_), .Y(new_n271_));
  OAI21X1  g00079(.A0(new_n252_), .A1(new_n242_), .B0(new_n255_), .Y(new_n272_));
  NOR2X1   g00080(.A(\a[121] ), .B(\a[120] ), .Y(new_n273_));
  INVX1    g00081(.A(new_n273_), .Y(new_n274_));
  AOI21X1  g00082(.A0(new_n268_), .A1(new_n265_), .B0(new_n274_), .Y(new_n275_));
  AOI21X1  g00083(.A0(new_n272_), .A1(\a[121] ), .B0(new_n275_), .Y(new_n276_));
  OR4X1    g00084(.A(new_n270_), .B(new_n215_), .C(new_n213_), .D(new_n228_), .Y(new_n277_));
  OR2X1    g00085(.A(new_n277_), .B(new_n269_), .Y(new_n278_));
  AOI22X1  g00086(.A0(new_n278_), .A1(new_n276_), .B0(new_n271_), .B1(\asqrt[61] ), .Y(new_n279_));
  OR2X1    g00087(.A(new_n279_), .B(new_n199_), .Y(new_n280_));
  AND2X1   g00088(.A(new_n278_), .B(new_n276_), .Y(new_n281_));
  NOR2X1   g00089(.A(new_n270_), .B(new_n269_), .Y(new_n282_));
  OAI21X1  g00090(.A0(new_n282_), .A1(new_n217_), .B0(new_n199_), .Y(new_n283_));
  OAI21X1  g00091(.A0(new_n252_), .A1(new_n242_), .B0(new_n273_), .Y(new_n284_));
  AND2X1   g00092(.A(new_n266_), .B(new_n262_), .Y(new_n285_));
  OR2X1    g00093(.A(new_n250_), .B(new_n217_), .Y(new_n286_));
  OR4X1    g00094(.A(new_n286_), .B(new_n249_), .C(new_n285_), .D(new_n242_), .Y(new_n287_));
  AOI21X1  g00095(.A0(new_n287_), .A1(new_n284_), .B0(new_n218_), .Y(new_n288_));
  NOR4X1   g00096(.A(new_n286_), .B(new_n249_), .C(new_n285_), .D(new_n242_), .Y(new_n289_));
  NOR3X1   g00097(.A(new_n289_), .B(new_n275_), .C(\a[122] ), .Y(new_n290_));
  OAI22X1  g00098(.A0(new_n290_), .A1(new_n288_), .B0(new_n283_), .B1(new_n281_), .Y(new_n291_));
  AND2X1   g00099(.A(new_n268_), .B(new_n265_), .Y(new_n292_));
  NOR4X1   g00100(.A(new_n292_), .B(new_n261_), .C(new_n225_), .D(new_n258_), .Y(new_n293_));
  AND2X1   g00101(.A(new_n259_), .B(new_n221_), .Y(new_n294_));
  AOI21X1  g00102(.A0(new_n294_), .A1(\asqrt[60] ), .B0(new_n232_), .Y(new_n295_));
  NOR2X1   g00103(.A(new_n266_), .B(new_n262_), .Y(new_n296_));
  AOI21X1  g00104(.A0(new_n296_), .A1(\asqrt[60] ), .B0(new_n285_), .Y(new_n297_));
  OAI21X1  g00105(.A0(new_n295_), .A1(new_n293_), .B0(new_n297_), .Y(new_n298_));
  AOI21X1  g00106(.A0(new_n291_), .A1(new_n280_), .B0(new_n298_), .Y(new_n299_));
  INVX1    g00107(.A(\a[121] ), .Y(new_n300_));
  AOI21X1  g00108(.A0(new_n268_), .A1(new_n265_), .B0(\a[120] ), .Y(new_n301_));
  OAI21X1  g00109(.A0(new_n301_), .A1(new_n300_), .B0(new_n284_), .Y(new_n302_));
  NOR2X1   g00110(.A(new_n277_), .B(new_n269_), .Y(new_n303_));
  OAI22X1  g00111(.A0(new_n303_), .A1(new_n302_), .B0(new_n282_), .B1(new_n217_), .Y(new_n304_));
  OR2X1    g00112(.A(new_n295_), .B(new_n293_), .Y(new_n305_));
  AOI21X1  g00113(.A0(new_n304_), .A1(\asqrt[62] ), .B0(new_n305_), .Y(new_n306_));
  AOI21X1  g00114(.A0(new_n268_), .A1(new_n265_), .B0(new_n233_), .Y(new_n307_));
  AOI21X1  g00115(.A0(new_n266_), .A1(new_n262_), .B0(new_n193_), .Y(new_n308_));
  OAI21X1  g00116(.A0(new_n307_), .A1(new_n266_), .B0(new_n308_), .Y(new_n309_));
  OR4X1    g00117(.A(new_n250_), .B(new_n249_), .C(new_n244_), .D(new_n243_), .Y(new_n310_));
  AOI21X1  g00118(.A0(new_n266_), .A1(new_n262_), .B0(new_n310_), .Y(new_n311_));
  AND2X1   g00119(.A(new_n311_), .B(new_n265_), .Y(new_n312_));
  INVX1    g00120(.A(new_n312_), .Y(new_n313_));
  NAND2X1  g00121(.A(new_n313_), .B(new_n309_), .Y(new_n314_));
  AOI21X1  g00122(.A0(new_n306_), .A1(new_n291_), .B0(new_n314_), .Y(new_n315_));
  OAI21X1  g00123(.A0(new_n299_), .A1(\asqrt[63] ), .B0(new_n315_), .Y(\asqrt[59] ));
  AND2X1   g00124(.A(new_n304_), .B(\asqrt[62] ), .Y(new_n317_));
  NAND2X1  g00125(.A(new_n278_), .B(new_n276_), .Y(new_n318_));
  AOI21X1  g00126(.A0(new_n271_), .A1(\asqrt[61] ), .B0(\asqrt[62] ), .Y(new_n319_));
  NOR2X1   g00127(.A(new_n290_), .B(new_n288_), .Y(new_n320_));
  AOI21X1  g00128(.A0(new_n319_), .A1(new_n318_), .B0(new_n320_), .Y(new_n321_));
  AND2X1   g00129(.A(new_n297_), .B(new_n305_), .Y(new_n322_));
  OAI21X1  g00130(.A0(new_n321_), .A1(new_n317_), .B0(new_n322_), .Y(new_n323_));
  NOR2X1   g00131(.A(new_n295_), .B(new_n293_), .Y(new_n324_));
  OAI21X1  g00132(.A0(new_n279_), .A1(new_n199_), .B0(new_n324_), .Y(new_n325_));
  AND2X1   g00133(.A(new_n313_), .B(new_n309_), .Y(new_n326_));
  OAI21X1  g00134(.A0(new_n325_), .A1(new_n321_), .B0(new_n326_), .Y(new_n327_));
  AOI21X1  g00135(.A0(new_n323_), .A1(new_n193_), .B0(new_n327_), .Y(new_n328_));
  NOR2X1   g00136(.A(\a[117] ), .B(\a[116] ), .Y(new_n329_));
  INVX1    g00137(.A(new_n329_), .Y(new_n330_));
  MX2X1    g00138(.A(new_n330_), .B(new_n328_), .S0(\a[118] ), .Y(new_n331_));
  OR2X1    g00139(.A(new_n331_), .B(new_n292_), .Y(new_n332_));
  INVX1    g00140(.A(\a[118] ), .Y(new_n333_));
  NOR3X1   g00141(.A(\a[118] ), .B(\a[117] ), .C(\a[116] ), .Y(new_n334_));
  OR2X1    g00142(.A(new_n334_), .B(new_n250_), .Y(new_n335_));
  NOR4X1   g00143(.A(new_n335_), .B(new_n249_), .C(new_n285_), .D(new_n242_), .Y(new_n336_));
  OAI21X1  g00144(.A0(new_n328_), .A1(new_n333_), .B0(new_n336_), .Y(new_n337_));
  OAI21X1  g00145(.A0(new_n328_), .A1(\a[118] ), .B0(\a[119] ), .Y(new_n338_));
  NOR2X1   g00146(.A(\a[119] ), .B(\a[118] ), .Y(new_n339_));
  INVX1    g00147(.A(new_n339_), .Y(new_n340_));
  OR2X1    g00148(.A(new_n328_), .B(new_n340_), .Y(new_n341_));
  NAND3X1  g00149(.A(new_n341_), .B(new_n338_), .C(new_n337_), .Y(new_n342_));
  AOI21X1  g00150(.A0(new_n342_), .A1(new_n332_), .B0(new_n217_), .Y(new_n343_));
  MX2X1    g00151(.A(new_n329_), .B(\asqrt[59] ), .S0(\a[118] ), .Y(new_n344_));
  AOI21X1  g00152(.A0(new_n344_), .A1(\asqrt[60] ), .B0(\asqrt[61] ), .Y(new_n345_));
  OR2X1    g00153(.A(new_n307_), .B(new_n266_), .Y(new_n346_));
  AND2X1   g00154(.A(new_n308_), .B(new_n346_), .Y(new_n347_));
  NOR3X1   g00155(.A(new_n312_), .B(new_n347_), .C(new_n292_), .Y(new_n348_));
  OAI21X1  g00156(.A0(new_n325_), .A1(new_n321_), .B0(new_n348_), .Y(new_n349_));
  AOI21X1  g00157(.A0(new_n323_), .A1(new_n193_), .B0(new_n349_), .Y(new_n350_));
  AOI21X1  g00158(.A0(\asqrt[59] ), .A1(new_n339_), .B0(new_n350_), .Y(new_n351_));
  OR2X1    g00159(.A(new_n351_), .B(new_n255_), .Y(new_n352_));
  AND2X1   g00160(.A(\asqrt[59] ), .B(new_n339_), .Y(new_n353_));
  OR2X1    g00161(.A(new_n350_), .B(\a[120] ), .Y(new_n354_));
  OR2X1    g00162(.A(new_n354_), .B(new_n353_), .Y(new_n355_));
  AOI22X1  g00163(.A0(new_n355_), .A1(new_n352_), .B0(new_n345_), .B1(new_n342_), .Y(new_n356_));
  OAI21X1  g00164(.A0(new_n356_), .A1(new_n343_), .B0(\asqrt[62] ), .Y(new_n357_));
  NOR3X1   g00165(.A(new_n356_), .B(new_n343_), .C(\asqrt[62] ), .Y(new_n358_));
  AOI21X1  g00166(.A0(new_n271_), .A1(\asqrt[61] ), .B0(new_n303_), .Y(new_n359_));
  NAND3X1  g00167(.A(new_n359_), .B(\asqrt[59] ), .C(new_n302_), .Y(new_n360_));
  INVX1    g00168(.A(new_n359_), .Y(new_n361_));
  OAI21X1  g00169(.A0(new_n361_), .A1(new_n328_), .B0(new_n276_), .Y(new_n362_));
  AND2X1   g00170(.A(new_n362_), .B(new_n360_), .Y(new_n363_));
  OAI21X1  g00171(.A0(new_n363_), .A1(new_n358_), .B0(new_n357_), .Y(new_n364_));
  OAI21X1  g00172(.A0(new_n283_), .A1(new_n281_), .B0(new_n320_), .Y(new_n365_));
  NOR3X1   g00173(.A(new_n365_), .B(new_n328_), .C(new_n317_), .Y(new_n366_));
  AOI22X1  g00174(.A0(new_n319_), .A1(new_n318_), .B0(new_n304_), .B1(\asqrt[62] ), .Y(new_n367_));
  AOI21X1  g00175(.A0(new_n367_), .A1(\asqrt[59] ), .B0(new_n320_), .Y(new_n368_));
  OR2X1    g00176(.A(new_n368_), .B(new_n366_), .Y(new_n369_));
  AND2X1   g00177(.A(new_n306_), .B(new_n291_), .Y(new_n370_));
  AOI21X1  g00178(.A0(new_n291_), .A1(new_n280_), .B0(new_n324_), .Y(new_n371_));
  AOI21X1  g00179(.A0(new_n371_), .A1(\asqrt[59] ), .B0(new_n370_), .Y(new_n372_));
  AND2X1   g00180(.A(new_n372_), .B(new_n369_), .Y(new_n373_));
  AOI21X1  g00181(.A0(new_n373_), .A1(new_n364_), .B0(\asqrt[63] ), .Y(new_n374_));
  AND2X1   g00182(.A(new_n344_), .B(\asqrt[60] ), .Y(new_n375_));
  INVX1    g00183(.A(new_n336_), .Y(new_n376_));
  AOI21X1  g00184(.A0(\asqrt[59] ), .A1(\a[118] ), .B0(new_n376_), .Y(new_n377_));
  INVX1    g00185(.A(\a[119] ), .Y(new_n378_));
  AOI21X1  g00186(.A0(\asqrt[59] ), .A1(new_n333_), .B0(new_n378_), .Y(new_n379_));
  NOR3X1   g00187(.A(new_n353_), .B(new_n379_), .C(new_n377_), .Y(new_n380_));
  OAI21X1  g00188(.A0(new_n380_), .A1(new_n375_), .B0(\asqrt[61] ), .Y(new_n381_));
  OAI21X1  g00189(.A0(new_n331_), .A1(new_n292_), .B0(new_n217_), .Y(new_n382_));
  OAI22X1  g00190(.A0(new_n354_), .A1(new_n353_), .B0(new_n351_), .B1(new_n255_), .Y(new_n383_));
  OAI21X1  g00191(.A0(new_n382_), .A1(new_n380_), .B0(new_n383_), .Y(new_n384_));
  NAND3X1  g00192(.A(new_n384_), .B(new_n381_), .C(new_n199_), .Y(new_n385_));
  INVX1    g00193(.A(new_n363_), .Y(new_n386_));
  AND2X1   g00194(.A(new_n386_), .B(new_n385_), .Y(new_n387_));
  AOI21X1  g00195(.A0(new_n384_), .A1(new_n381_), .B0(new_n199_), .Y(new_n388_));
  OR2X1    g00196(.A(new_n369_), .B(new_n388_), .Y(new_n389_));
  AND2X1   g00197(.A(new_n291_), .B(new_n280_), .Y(new_n390_));
  AOI21X1  g00198(.A0(\asqrt[59] ), .A1(new_n390_), .B0(new_n324_), .Y(new_n391_));
  NOR3X1   g00199(.A(new_n391_), .B(new_n370_), .C(new_n193_), .Y(new_n392_));
  AND2X1   g00200(.A(new_n323_), .B(new_n193_), .Y(new_n393_));
  OR4X1    g00201(.A(new_n312_), .B(new_n347_), .C(new_n295_), .D(new_n293_), .Y(new_n394_));
  NOR3X1   g00202(.A(new_n394_), .B(new_n370_), .C(new_n393_), .Y(new_n395_));
  NOR2X1   g00203(.A(new_n395_), .B(new_n392_), .Y(new_n396_));
  OAI21X1  g00204(.A0(new_n389_), .A1(new_n387_), .B0(new_n396_), .Y(new_n397_));
  OR2X1    g00205(.A(new_n397_), .B(new_n374_), .Y(\asqrt[58] ));
  INVX1    g00206(.A(\asqrt[58] ), .Y(new_n399_));
  INVX1    g00207(.A(\a[116] ), .Y(new_n400_));
  AOI21X1  g00208(.A0(new_n386_), .A1(new_n385_), .B0(new_n388_), .Y(new_n401_));
  INVX1    g00209(.A(new_n373_), .Y(new_n402_));
  OAI21X1  g00210(.A0(new_n402_), .A1(new_n401_), .B0(new_n193_), .Y(new_n403_));
  NAND2X1  g00211(.A(new_n386_), .B(new_n385_), .Y(new_n404_));
  NOR2X1   g00212(.A(new_n369_), .B(new_n388_), .Y(new_n405_));
  INVX1    g00213(.A(new_n396_), .Y(new_n406_));
  AOI21X1  g00214(.A0(new_n405_), .A1(new_n404_), .B0(new_n406_), .Y(new_n407_));
  AOI21X1  g00215(.A0(new_n407_), .A1(new_n403_), .B0(new_n400_), .Y(new_n408_));
  NOR3X1   g00216(.A(\a[116] ), .B(\a[115] ), .C(\a[114] ), .Y(new_n409_));
  OR2X1    g00217(.A(new_n409_), .B(new_n408_), .Y(new_n410_));
  NOR4X1   g00218(.A(new_n409_), .B(new_n312_), .C(new_n347_), .D(new_n370_), .Y(new_n411_));
  OAI21X1  g00219(.A0(new_n299_), .A1(\asqrt[63] ), .B0(new_n411_), .Y(new_n412_));
  OR2X1    g00220(.A(new_n412_), .B(new_n408_), .Y(new_n413_));
  OAI21X1  g00221(.A0(new_n397_), .A1(new_n374_), .B0(new_n400_), .Y(new_n414_));
  AOI21X1  g00222(.A0(new_n407_), .A1(new_n403_), .B0(new_n330_), .Y(new_n415_));
  AOI21X1  g00223(.A0(new_n414_), .A1(\a[117] ), .B0(new_n415_), .Y(new_n416_));
  AOI22X1  g00224(.A0(new_n416_), .A1(new_n413_), .B0(new_n410_), .B1(\asqrt[59] ), .Y(new_n417_));
  OR2X1    g00225(.A(new_n417_), .B(new_n292_), .Y(new_n418_));
  AND2X1   g00226(.A(new_n416_), .B(new_n413_), .Y(new_n419_));
  NOR2X1   g00227(.A(new_n409_), .B(new_n408_), .Y(new_n420_));
  OAI21X1  g00228(.A0(new_n420_), .A1(new_n328_), .B0(new_n292_), .Y(new_n421_));
  OAI21X1  g00229(.A0(new_n397_), .A1(new_n374_), .B0(new_n329_), .Y(new_n422_));
  AND2X1   g00230(.A(new_n405_), .B(new_n404_), .Y(new_n423_));
  OR2X1    g00231(.A(new_n395_), .B(new_n328_), .Y(new_n424_));
  OR4X1    g00232(.A(new_n424_), .B(new_n392_), .C(new_n423_), .D(new_n374_), .Y(new_n425_));
  AOI21X1  g00233(.A0(new_n425_), .A1(new_n422_), .B0(new_n333_), .Y(new_n426_));
  NOR4X1   g00234(.A(new_n424_), .B(new_n392_), .C(new_n423_), .D(new_n374_), .Y(new_n427_));
  NOR3X1   g00235(.A(new_n427_), .B(new_n415_), .C(\a[118] ), .Y(new_n428_));
  OR2X1    g00236(.A(new_n428_), .B(new_n426_), .Y(new_n429_));
  OAI21X1  g00237(.A0(new_n421_), .A1(new_n419_), .B0(new_n429_), .Y(new_n430_));
  AOI21X1  g00238(.A0(new_n430_), .A1(new_n418_), .B0(new_n217_), .Y(new_n431_));
  AND2X1   g00239(.A(new_n341_), .B(new_n338_), .Y(new_n432_));
  NOR3X1   g00240(.A(new_n432_), .B(new_n377_), .C(new_n375_), .Y(new_n433_));
  OAI21X1  g00241(.A0(new_n397_), .A1(new_n374_), .B0(new_n433_), .Y(new_n434_));
  NAND3X1  g00242(.A(\asqrt[58] ), .B(new_n337_), .C(new_n332_), .Y(new_n435_));
  NAND2X1  g00243(.A(new_n435_), .B(new_n432_), .Y(new_n436_));
  NOR2X1   g00244(.A(new_n412_), .B(new_n408_), .Y(new_n437_));
  INVX1    g00245(.A(\a[117] ), .Y(new_n438_));
  AOI21X1  g00246(.A0(new_n407_), .A1(new_n403_), .B0(\a[116] ), .Y(new_n439_));
  OAI21X1  g00247(.A0(new_n439_), .A1(new_n438_), .B0(new_n422_), .Y(new_n440_));
  OAI22X1  g00248(.A0(new_n440_), .A1(new_n437_), .B0(new_n420_), .B1(new_n328_), .Y(new_n441_));
  AOI21X1  g00249(.A0(new_n441_), .A1(\asqrt[60] ), .B0(\asqrt[61] ), .Y(new_n442_));
  AOI22X1  g00250(.A0(new_n442_), .A1(new_n430_), .B0(new_n436_), .B1(new_n434_), .Y(new_n443_));
  OAI21X1  g00251(.A0(new_n443_), .A1(new_n431_), .B0(\asqrt[62] ), .Y(new_n444_));
  AND2X1   g00252(.A(new_n345_), .B(new_n342_), .Y(new_n445_));
  NOR3X1   g00253(.A(new_n383_), .B(new_n445_), .C(new_n343_), .Y(new_n446_));
  NOR2X1   g00254(.A(new_n445_), .B(new_n343_), .Y(new_n447_));
  OAI21X1  g00255(.A0(new_n397_), .A1(new_n374_), .B0(new_n447_), .Y(new_n448_));
  AOI22X1  g00256(.A0(new_n448_), .A1(new_n383_), .B0(new_n446_), .B1(\asqrt[58] ), .Y(new_n449_));
  NOR3X1   g00257(.A(new_n443_), .B(new_n431_), .C(\asqrt[62] ), .Y(new_n450_));
  OAI21X1  g00258(.A0(new_n450_), .A1(new_n449_), .B0(new_n444_), .Y(new_n451_));
  NOR4X1   g00259(.A(new_n399_), .B(new_n386_), .C(new_n358_), .D(new_n388_), .Y(new_n452_));
  AND2X1   g00260(.A(new_n385_), .B(new_n357_), .Y(new_n453_));
  AOI21X1  g00261(.A0(new_n453_), .A1(\asqrt[58] ), .B0(new_n363_), .Y(new_n454_));
  OR2X1    g00262(.A(new_n454_), .B(new_n452_), .Y(new_n455_));
  INVX1    g00263(.A(new_n369_), .Y(new_n456_));
  NOR2X1   g00264(.A(new_n456_), .B(new_n401_), .Y(new_n457_));
  AOI21X1  g00265(.A0(new_n457_), .A1(\asqrt[58] ), .B0(new_n423_), .Y(new_n458_));
  AND2X1   g00266(.A(new_n458_), .B(new_n455_), .Y(new_n459_));
  AOI21X1  g00267(.A0(new_n459_), .A1(new_n451_), .B0(\asqrt[63] ), .Y(new_n460_));
  NOR2X1   g00268(.A(new_n450_), .B(new_n449_), .Y(new_n461_));
  AND2X1   g00269(.A(new_n441_), .B(\asqrt[60] ), .Y(new_n462_));
  NAND2X1  g00270(.A(new_n416_), .B(new_n413_), .Y(new_n463_));
  AOI21X1  g00271(.A0(new_n410_), .A1(\asqrt[59] ), .B0(\asqrt[60] ), .Y(new_n464_));
  NOR2X1   g00272(.A(new_n428_), .B(new_n426_), .Y(new_n465_));
  AOI21X1  g00273(.A0(new_n464_), .A1(new_n463_), .B0(new_n465_), .Y(new_n466_));
  OAI21X1  g00274(.A0(new_n466_), .A1(new_n462_), .B0(\asqrt[61] ), .Y(new_n467_));
  NAND2X1  g00275(.A(new_n436_), .B(new_n434_), .Y(new_n468_));
  OAI21X1  g00276(.A0(new_n417_), .A1(new_n292_), .B0(new_n217_), .Y(new_n469_));
  OAI21X1  g00277(.A0(new_n469_), .A1(new_n466_), .B0(new_n468_), .Y(new_n470_));
  AOI21X1  g00278(.A0(new_n470_), .A1(new_n467_), .B0(new_n199_), .Y(new_n471_));
  OR2X1    g00279(.A(new_n455_), .B(new_n471_), .Y(new_n472_));
  AOI21X1  g00280(.A0(\asqrt[58] ), .A1(new_n369_), .B0(new_n364_), .Y(new_n473_));
  OAI21X1  g00281(.A0(new_n456_), .A1(new_n401_), .B0(\asqrt[63] ), .Y(new_n474_));
  NOR2X1   g00282(.A(new_n474_), .B(new_n473_), .Y(new_n475_));
  NOR4X1   g00283(.A(new_n395_), .B(new_n392_), .C(new_n368_), .D(new_n366_), .Y(new_n476_));
  OAI21X1  g00284(.A0(new_n389_), .A1(new_n387_), .B0(new_n476_), .Y(new_n477_));
  NOR2X1   g00285(.A(new_n477_), .B(new_n374_), .Y(new_n478_));
  NOR2X1   g00286(.A(new_n478_), .B(new_n475_), .Y(new_n479_));
  OAI21X1  g00287(.A0(new_n472_), .A1(new_n461_), .B0(new_n479_), .Y(new_n480_));
  NOR2X1   g00288(.A(new_n480_), .B(new_n460_), .Y(new_n481_));
  OR2X1    g00289(.A(new_n480_), .B(new_n460_), .Y(\asqrt[57] ));
  NOR2X1   g00290(.A(\a[113] ), .B(\a[112] ), .Y(new_n483_));
  MX2X1    g00291(.A(new_n483_), .B(\asqrt[57] ), .S0(\a[114] ), .Y(new_n484_));
  OAI21X1  g00292(.A0(new_n480_), .A1(new_n460_), .B0(\a[114] ), .Y(new_n485_));
  NOR3X1   g00293(.A(\a[114] ), .B(\a[113] ), .C(\a[112] ), .Y(new_n486_));
  OR2X1    g00294(.A(new_n486_), .B(new_n395_), .Y(new_n487_));
  NOR4X1   g00295(.A(new_n487_), .B(new_n392_), .C(new_n423_), .D(new_n374_), .Y(new_n488_));
  NAND2X1  g00296(.A(new_n488_), .B(new_n485_), .Y(new_n489_));
  INVX1    g00297(.A(\a[114] ), .Y(new_n490_));
  OAI21X1  g00298(.A0(new_n480_), .A1(new_n460_), .B0(new_n490_), .Y(new_n491_));
  NOR2X1   g00299(.A(\a[115] ), .B(\a[114] ), .Y(new_n492_));
  INVX1    g00300(.A(new_n492_), .Y(new_n493_));
  INVX1    g00301(.A(new_n449_), .Y(new_n494_));
  NAND3X1  g00302(.A(new_n470_), .B(new_n467_), .C(new_n199_), .Y(new_n495_));
  AOI21X1  g00303(.A0(new_n495_), .A1(new_n494_), .B0(new_n471_), .Y(new_n496_));
  INVX1    g00304(.A(new_n459_), .Y(new_n497_));
  OAI21X1  g00305(.A0(new_n497_), .A1(new_n496_), .B0(new_n193_), .Y(new_n498_));
  OR2X1    g00306(.A(new_n450_), .B(new_n449_), .Y(new_n499_));
  NOR2X1   g00307(.A(new_n455_), .B(new_n471_), .Y(new_n500_));
  INVX1    g00308(.A(new_n479_), .Y(new_n501_));
  AOI21X1  g00309(.A0(new_n500_), .A1(new_n499_), .B0(new_n501_), .Y(new_n502_));
  AOI21X1  g00310(.A0(new_n502_), .A1(new_n498_), .B0(new_n493_), .Y(new_n503_));
  AOI21X1  g00311(.A0(new_n491_), .A1(\a[115] ), .B0(new_n503_), .Y(new_n504_));
  AOI22X1  g00312(.A0(new_n504_), .A1(new_n489_), .B0(new_n484_), .B1(\asqrt[58] ), .Y(new_n505_));
  OR2X1    g00313(.A(new_n505_), .B(new_n328_), .Y(new_n506_));
  AND2X1   g00314(.A(new_n504_), .B(new_n489_), .Y(new_n507_));
  AOI21X1  g00315(.A0(\asqrt[57] ), .A1(\a[114] ), .B0(new_n486_), .Y(new_n508_));
  OAI21X1  g00316(.A0(new_n508_), .A1(new_n399_), .B0(new_n328_), .Y(new_n509_));
  OAI21X1  g00317(.A0(new_n480_), .A1(new_n460_), .B0(new_n492_), .Y(new_n510_));
  AOI21X1  g00318(.A0(new_n407_), .A1(new_n403_), .B0(new_n478_), .Y(new_n511_));
  OAI21X1  g00319(.A0(new_n474_), .A1(new_n473_), .B0(new_n511_), .Y(new_n512_));
  AOI21X1  g00320(.A0(new_n500_), .A1(new_n499_), .B0(new_n512_), .Y(new_n513_));
  NAND2X1  g00321(.A(new_n513_), .B(new_n498_), .Y(new_n514_));
  AOI21X1  g00322(.A0(new_n514_), .A1(new_n510_), .B0(new_n400_), .Y(new_n515_));
  AOI21X1  g00323(.A0(new_n513_), .A1(new_n498_), .B0(\a[116] ), .Y(new_n516_));
  AND2X1   g00324(.A(new_n516_), .B(new_n510_), .Y(new_n517_));
  OR2X1    g00325(.A(new_n517_), .B(new_n515_), .Y(new_n518_));
  OAI21X1  g00326(.A0(new_n509_), .A1(new_n507_), .B0(new_n518_), .Y(new_n519_));
  AOI21X1  g00327(.A0(new_n519_), .A1(new_n506_), .B0(new_n292_), .Y(new_n520_));
  AOI21X1  g00328(.A0(new_n410_), .A1(\asqrt[59] ), .B0(new_n437_), .Y(new_n521_));
  AND2X1   g00329(.A(new_n521_), .B(new_n440_), .Y(new_n522_));
  OAI21X1  g00330(.A0(new_n480_), .A1(new_n460_), .B0(new_n521_), .Y(new_n523_));
  AOI22X1  g00331(.A0(new_n523_), .A1(new_n416_), .B0(new_n522_), .B1(\asqrt[57] ), .Y(new_n524_));
  AND2X1   g00332(.A(new_n488_), .B(new_n485_), .Y(new_n525_));
  INVX1    g00333(.A(\a[115] ), .Y(new_n526_));
  AOI21X1  g00334(.A0(new_n502_), .A1(new_n498_), .B0(\a[114] ), .Y(new_n527_));
  OAI21X1  g00335(.A0(new_n527_), .A1(new_n526_), .B0(new_n510_), .Y(new_n528_));
  OAI22X1  g00336(.A0(new_n528_), .A1(new_n525_), .B0(new_n508_), .B1(new_n399_), .Y(new_n529_));
  AOI21X1  g00337(.A0(new_n529_), .A1(\asqrt[59] ), .B0(\asqrt[60] ), .Y(new_n530_));
  AOI21X1  g00338(.A0(new_n530_), .A1(new_n519_), .B0(new_n524_), .Y(new_n531_));
  OAI21X1  g00339(.A0(new_n531_), .A1(new_n520_), .B0(\asqrt[61] ), .Y(new_n532_));
  AOI21X1  g00340(.A0(new_n464_), .A1(new_n463_), .B0(new_n429_), .Y(new_n533_));
  AND2X1   g00341(.A(new_n533_), .B(new_n418_), .Y(new_n534_));
  AOI22X1  g00342(.A0(new_n464_), .A1(new_n463_), .B0(new_n441_), .B1(\asqrt[60] ), .Y(new_n535_));
  OAI21X1  g00343(.A0(new_n480_), .A1(new_n460_), .B0(new_n535_), .Y(new_n536_));
  AOI22X1  g00344(.A0(new_n536_), .A1(new_n429_), .B0(new_n534_), .B1(\asqrt[57] ), .Y(new_n537_));
  NOR3X1   g00345(.A(new_n531_), .B(new_n520_), .C(\asqrt[61] ), .Y(new_n538_));
  OAI21X1  g00346(.A0(new_n538_), .A1(new_n537_), .B0(new_n532_), .Y(new_n539_));
  AND2X1   g00347(.A(new_n539_), .B(\asqrt[62] ), .Y(new_n540_));
  INVX1    g00348(.A(new_n537_), .Y(new_n541_));
  AND2X1   g00349(.A(new_n529_), .B(\asqrt[59] ), .Y(new_n542_));
  OR2X1    g00350(.A(new_n528_), .B(new_n525_), .Y(new_n543_));
  AOI21X1  g00351(.A0(new_n484_), .A1(\asqrt[58] ), .B0(\asqrt[59] ), .Y(new_n544_));
  NOR2X1   g00352(.A(new_n517_), .B(new_n515_), .Y(new_n545_));
  AOI21X1  g00353(.A0(new_n544_), .A1(new_n543_), .B0(new_n545_), .Y(new_n546_));
  OAI21X1  g00354(.A0(new_n546_), .A1(new_n542_), .B0(\asqrt[60] ), .Y(new_n547_));
  INVX1    g00355(.A(new_n524_), .Y(new_n548_));
  OAI21X1  g00356(.A0(new_n505_), .A1(new_n328_), .B0(new_n292_), .Y(new_n549_));
  OAI21X1  g00357(.A0(new_n549_), .A1(new_n546_), .B0(new_n548_), .Y(new_n550_));
  NAND3X1  g00358(.A(new_n550_), .B(new_n547_), .C(new_n217_), .Y(new_n551_));
  NAND2X1  g00359(.A(new_n551_), .B(new_n541_), .Y(new_n552_));
  AND2X1   g00360(.A(new_n442_), .B(new_n430_), .Y(new_n553_));
  NOR3X1   g00361(.A(new_n553_), .B(new_n468_), .C(new_n431_), .Y(new_n554_));
  NOR2X1   g00362(.A(new_n553_), .B(new_n431_), .Y(new_n555_));
  OAI21X1  g00363(.A0(new_n480_), .A1(new_n460_), .B0(new_n555_), .Y(new_n556_));
  AOI22X1  g00364(.A0(new_n556_), .A1(new_n468_), .B0(new_n554_), .B1(\asqrt[57] ), .Y(new_n557_));
  AOI21X1  g00365(.A0(new_n550_), .A1(new_n547_), .B0(new_n217_), .Y(new_n558_));
  NOR2X1   g00366(.A(new_n558_), .B(\asqrt[62] ), .Y(new_n559_));
  AOI21X1  g00367(.A0(new_n559_), .A1(new_n552_), .B0(new_n557_), .Y(new_n560_));
  NOR4X1   g00368(.A(new_n481_), .B(new_n450_), .C(new_n494_), .D(new_n471_), .Y(new_n561_));
  NAND3X1  g00369(.A(\asqrt[57] ), .B(new_n495_), .C(new_n444_), .Y(new_n562_));
  AND2X1   g00370(.A(new_n562_), .B(new_n494_), .Y(new_n563_));
  AND2X1   g00371(.A(new_n500_), .B(new_n499_), .Y(new_n564_));
  AND2X1   g00372(.A(new_n455_), .B(new_n451_), .Y(new_n565_));
  AOI21X1  g00373(.A0(new_n565_), .A1(\asqrt[57] ), .B0(new_n564_), .Y(new_n566_));
  OAI21X1  g00374(.A0(new_n563_), .A1(new_n561_), .B0(new_n566_), .Y(new_n567_));
  INVX1    g00375(.A(new_n567_), .Y(new_n568_));
  OAI21X1  g00376(.A0(new_n560_), .A1(new_n540_), .B0(new_n568_), .Y(new_n569_));
  AOI21X1  g00377(.A0(new_n551_), .A1(new_n541_), .B0(new_n558_), .Y(new_n570_));
  AOI21X1  g00378(.A0(new_n562_), .A1(new_n494_), .B0(new_n561_), .Y(new_n571_));
  OAI21X1  g00379(.A0(new_n570_), .A1(new_n199_), .B0(new_n571_), .Y(new_n572_));
  OAI21X1  g00380(.A0(new_n480_), .A1(new_n460_), .B0(new_n455_), .Y(new_n573_));
  AND2X1   g00381(.A(new_n573_), .B(new_n496_), .Y(new_n574_));
  NOR3X1   g00382(.A(new_n574_), .B(new_n565_), .C(new_n193_), .Y(new_n575_));
  INVX1    g00383(.A(new_n564_), .Y(new_n576_));
  NOR4X1   g00384(.A(new_n478_), .B(new_n475_), .C(new_n454_), .D(new_n452_), .Y(new_n577_));
  NAND3X1  g00385(.A(new_n577_), .B(new_n576_), .C(new_n498_), .Y(new_n578_));
  INVX1    g00386(.A(new_n578_), .Y(new_n579_));
  NOR2X1   g00387(.A(new_n579_), .B(new_n575_), .Y(new_n580_));
  OAI21X1  g00388(.A0(new_n572_), .A1(new_n560_), .B0(new_n580_), .Y(new_n581_));
  AOI21X1  g00389(.A0(new_n569_), .A1(new_n193_), .B0(new_n581_), .Y(new_n582_));
  OR2X1    g00390(.A(new_n570_), .B(new_n199_), .Y(new_n583_));
  AND2X1   g00391(.A(new_n551_), .B(new_n541_), .Y(new_n584_));
  INVX1    g00392(.A(new_n557_), .Y(new_n585_));
  OR2X1    g00393(.A(new_n558_), .B(\asqrt[62] ), .Y(new_n586_));
  OAI21X1  g00394(.A0(new_n586_), .A1(new_n584_), .B0(new_n585_), .Y(new_n587_));
  AOI21X1  g00395(.A0(new_n587_), .A1(new_n583_), .B0(new_n567_), .Y(new_n588_));
  INVX1    g00396(.A(new_n571_), .Y(new_n589_));
  AOI21X1  g00397(.A0(new_n539_), .A1(\asqrt[62] ), .B0(new_n589_), .Y(new_n590_));
  INVX1    g00398(.A(new_n580_), .Y(new_n591_));
  AOI21X1  g00399(.A0(new_n590_), .A1(new_n587_), .B0(new_n591_), .Y(new_n592_));
  OAI21X1  g00400(.A0(new_n588_), .A1(\asqrt[63] ), .B0(new_n592_), .Y(\asqrt[56] ));
  NOR2X1   g00401(.A(\a[111] ), .B(\a[110] ), .Y(new_n594_));
  MX2X1    g00402(.A(new_n594_), .B(\asqrt[56] ), .S0(\a[112] ), .Y(new_n595_));
  AND2X1   g00403(.A(new_n595_), .B(\asqrt[57] ), .Y(new_n596_));
  INVX1    g00404(.A(\a[112] ), .Y(new_n597_));
  INVX1    g00405(.A(\a[113] ), .Y(new_n598_));
  AOI21X1  g00406(.A0(\asqrt[56] ), .A1(new_n597_), .B0(new_n598_), .Y(new_n599_));
  AND2X1   g00407(.A(\asqrt[56] ), .B(new_n483_), .Y(new_n600_));
  NOR3X1   g00408(.A(\a[112] ), .B(\a[111] ), .C(\a[110] ), .Y(new_n601_));
  NOR3X1   g00409(.A(new_n601_), .B(new_n478_), .C(new_n475_), .Y(new_n602_));
  NAND3X1  g00410(.A(new_n602_), .B(new_n576_), .C(new_n498_), .Y(new_n603_));
  AOI21X1  g00411(.A0(\asqrt[56] ), .A1(\a[112] ), .B0(new_n603_), .Y(new_n604_));
  NOR3X1   g00412(.A(new_n604_), .B(new_n600_), .C(new_n599_), .Y(new_n605_));
  OAI21X1  g00413(.A0(new_n605_), .A1(new_n596_), .B0(\asqrt[58] ), .Y(new_n606_));
  INVX1    g00414(.A(new_n594_), .Y(new_n607_));
  MX2X1    g00415(.A(new_n607_), .B(new_n582_), .S0(\a[112] ), .Y(new_n608_));
  OAI21X1  g00416(.A0(new_n608_), .A1(new_n481_), .B0(new_n399_), .Y(new_n609_));
  NOR3X1   g00417(.A(new_n579_), .B(new_n575_), .C(new_n481_), .Y(new_n610_));
  OAI21X1  g00418(.A0(new_n572_), .A1(new_n560_), .B0(new_n610_), .Y(new_n611_));
  AOI21X1  g00419(.A0(new_n569_), .A1(new_n193_), .B0(new_n611_), .Y(new_n612_));
  AOI21X1  g00420(.A0(\asqrt[56] ), .A1(new_n483_), .B0(new_n612_), .Y(new_n613_));
  OR2X1    g00421(.A(new_n612_), .B(\a[114] ), .Y(new_n614_));
  OAI22X1  g00422(.A0(new_n614_), .A1(new_n600_), .B0(new_n613_), .B1(new_n490_), .Y(new_n615_));
  OAI21X1  g00423(.A0(new_n609_), .A1(new_n605_), .B0(new_n615_), .Y(new_n616_));
  AOI21X1  g00424(.A0(new_n616_), .A1(new_n606_), .B0(new_n328_), .Y(new_n617_));
  AOI21X1  g00425(.A0(new_n484_), .A1(\asqrt[58] ), .B0(new_n525_), .Y(new_n618_));
  NAND3X1  g00426(.A(new_n618_), .B(\asqrt[56] ), .C(new_n528_), .Y(new_n619_));
  INVX1    g00427(.A(new_n618_), .Y(new_n620_));
  OAI21X1  g00428(.A0(new_n620_), .A1(new_n582_), .B0(new_n504_), .Y(new_n621_));
  AND2X1   g00429(.A(new_n621_), .B(new_n619_), .Y(new_n622_));
  INVX1    g00430(.A(new_n622_), .Y(new_n623_));
  NAND3X1  g00431(.A(new_n616_), .B(new_n606_), .C(new_n328_), .Y(new_n624_));
  AOI21X1  g00432(.A0(new_n624_), .A1(new_n623_), .B0(new_n617_), .Y(new_n625_));
  OR2X1    g00433(.A(new_n625_), .B(new_n292_), .Y(new_n626_));
  AND2X1   g00434(.A(new_n624_), .B(new_n623_), .Y(new_n627_));
  OAI21X1  g00435(.A0(new_n509_), .A1(new_n507_), .B0(new_n545_), .Y(new_n628_));
  NOR3X1   g00436(.A(new_n628_), .B(new_n582_), .C(new_n542_), .Y(new_n629_));
  OAI22X1  g00437(.A0(new_n509_), .A1(new_n507_), .B0(new_n505_), .B1(new_n328_), .Y(new_n630_));
  OR2X1    g00438(.A(new_n630_), .B(new_n582_), .Y(new_n631_));
  AOI21X1  g00439(.A0(new_n631_), .A1(new_n518_), .B0(new_n629_), .Y(new_n632_));
  INVX1    g00440(.A(new_n632_), .Y(new_n633_));
  OR2X1    g00441(.A(new_n617_), .B(\asqrt[60] ), .Y(new_n634_));
  OAI21X1  g00442(.A0(new_n634_), .A1(new_n627_), .B0(new_n633_), .Y(new_n635_));
  AOI21X1  g00443(.A0(new_n635_), .A1(new_n626_), .B0(new_n217_), .Y(new_n636_));
  AND2X1   g00444(.A(new_n530_), .B(new_n519_), .Y(new_n637_));
  OR4X1    g00445(.A(new_n582_), .B(new_n637_), .C(new_n548_), .D(new_n520_), .Y(new_n638_));
  OR2X1    g00446(.A(new_n637_), .B(new_n520_), .Y(new_n639_));
  OAI21X1  g00447(.A0(new_n639_), .A1(new_n582_), .B0(new_n548_), .Y(new_n640_));
  AND2X1   g00448(.A(new_n640_), .B(new_n638_), .Y(new_n641_));
  OR2X1    g00449(.A(new_n608_), .B(new_n481_), .Y(new_n642_));
  OAI21X1  g00450(.A0(new_n582_), .A1(\a[112] ), .B0(\a[113] ), .Y(new_n643_));
  INVX1    g00451(.A(new_n483_), .Y(new_n644_));
  OR2X1    g00452(.A(new_n582_), .B(new_n644_), .Y(new_n645_));
  INVX1    g00453(.A(new_n603_), .Y(new_n646_));
  OAI21X1  g00454(.A0(new_n582_), .A1(new_n597_), .B0(new_n646_), .Y(new_n647_));
  NAND3X1  g00455(.A(new_n647_), .B(new_n645_), .C(new_n643_), .Y(new_n648_));
  AOI21X1  g00456(.A0(new_n648_), .A1(new_n642_), .B0(new_n399_), .Y(new_n649_));
  AOI21X1  g00457(.A0(new_n595_), .A1(\asqrt[57] ), .B0(\asqrt[58] ), .Y(new_n650_));
  OR2X1    g00458(.A(new_n613_), .B(new_n490_), .Y(new_n651_));
  OR2X1    g00459(.A(new_n614_), .B(new_n600_), .Y(new_n652_));
  AOI22X1  g00460(.A0(new_n652_), .A1(new_n651_), .B0(new_n650_), .B1(new_n648_), .Y(new_n653_));
  OAI21X1  g00461(.A0(new_n653_), .A1(new_n649_), .B0(\asqrt[59] ), .Y(new_n654_));
  NOR3X1   g00462(.A(new_n653_), .B(new_n649_), .C(\asqrt[59] ), .Y(new_n655_));
  OAI21X1  g00463(.A0(new_n655_), .A1(new_n622_), .B0(new_n654_), .Y(new_n656_));
  AOI21X1  g00464(.A0(new_n656_), .A1(\asqrt[60] ), .B0(\asqrt[61] ), .Y(new_n657_));
  AOI21X1  g00465(.A0(new_n657_), .A1(new_n635_), .B0(new_n641_), .Y(new_n658_));
  OAI21X1  g00466(.A0(new_n658_), .A1(new_n636_), .B0(\asqrt[62] ), .Y(new_n659_));
  NAND3X1  g00467(.A(new_n551_), .B(new_n537_), .C(new_n532_), .Y(new_n660_));
  NOR3X1   g00468(.A(new_n582_), .B(new_n538_), .C(new_n558_), .Y(new_n661_));
  OAI22X1  g00469(.A0(new_n661_), .A1(new_n537_), .B0(new_n660_), .B1(new_n582_), .Y(new_n662_));
  INVX1    g00470(.A(new_n662_), .Y(new_n663_));
  NOR3X1   g00471(.A(new_n658_), .B(new_n636_), .C(\asqrt[62] ), .Y(new_n664_));
  OAI21X1  g00472(.A0(new_n664_), .A1(new_n663_), .B0(new_n659_), .Y(new_n665_));
  AND2X1   g00473(.A(new_n559_), .B(new_n552_), .Y(new_n666_));
  NOR4X1   g00474(.A(new_n582_), .B(new_n666_), .C(new_n585_), .D(new_n540_), .Y(new_n667_));
  AOI22X1  g00475(.A0(new_n559_), .A1(new_n552_), .B0(new_n539_), .B1(\asqrt[62] ), .Y(new_n668_));
  AOI21X1  g00476(.A0(new_n668_), .A1(\asqrt[56] ), .B0(new_n557_), .Y(new_n669_));
  NOR2X1   g00477(.A(new_n669_), .B(new_n667_), .Y(new_n670_));
  INVX1    g00478(.A(new_n670_), .Y(new_n671_));
  AND2X1   g00479(.A(new_n590_), .B(new_n587_), .Y(new_n672_));
  AOI21X1  g00480(.A0(new_n587_), .A1(new_n583_), .B0(new_n571_), .Y(new_n673_));
  AOI21X1  g00481(.A0(new_n673_), .A1(\asqrt[56] ), .B0(new_n672_), .Y(new_n674_));
  AND2X1   g00482(.A(new_n674_), .B(new_n671_), .Y(new_n675_));
  AOI21X1  g00483(.A0(new_n675_), .A1(new_n665_), .B0(\asqrt[63] ), .Y(new_n676_));
  AND2X1   g00484(.A(new_n656_), .B(\asqrt[60] ), .Y(new_n677_));
  NAND2X1  g00485(.A(new_n624_), .B(new_n623_), .Y(new_n678_));
  NOR2X1   g00486(.A(new_n617_), .B(\asqrt[60] ), .Y(new_n679_));
  AOI21X1  g00487(.A0(new_n679_), .A1(new_n678_), .B0(new_n632_), .Y(new_n680_));
  OAI21X1  g00488(.A0(new_n680_), .A1(new_n677_), .B0(\asqrt[61] ), .Y(new_n681_));
  INVX1    g00489(.A(new_n641_), .Y(new_n682_));
  OAI21X1  g00490(.A0(new_n625_), .A1(new_n292_), .B0(new_n217_), .Y(new_n683_));
  OAI21X1  g00491(.A0(new_n683_), .A1(new_n680_), .B0(new_n682_), .Y(new_n684_));
  NAND3X1  g00492(.A(new_n684_), .B(new_n681_), .C(new_n199_), .Y(new_n685_));
  AND2X1   g00493(.A(new_n685_), .B(new_n662_), .Y(new_n686_));
  AOI21X1  g00494(.A0(new_n684_), .A1(new_n681_), .B0(new_n199_), .Y(new_n687_));
  OR2X1    g00495(.A(new_n671_), .B(new_n687_), .Y(new_n688_));
  NAND2X1  g00496(.A(new_n587_), .B(new_n583_), .Y(new_n689_));
  AOI21X1  g00497(.A0(\asqrt[56] ), .A1(new_n589_), .B0(new_n689_), .Y(new_n690_));
  NOR3X1   g00498(.A(new_n690_), .B(new_n673_), .C(new_n193_), .Y(new_n691_));
  AND2X1   g00499(.A(new_n569_), .B(new_n193_), .Y(new_n692_));
  OR4X1    g00500(.A(new_n579_), .B(new_n575_), .C(new_n563_), .D(new_n561_), .Y(new_n693_));
  NOR3X1   g00501(.A(new_n693_), .B(new_n672_), .C(new_n692_), .Y(new_n694_));
  NOR2X1   g00502(.A(new_n694_), .B(new_n691_), .Y(new_n695_));
  OAI21X1  g00503(.A0(new_n688_), .A1(new_n686_), .B0(new_n695_), .Y(new_n696_));
  NOR2X1   g00504(.A(new_n696_), .B(new_n676_), .Y(new_n697_));
  INVX1    g00505(.A(new_n697_), .Y(\asqrt[55] ));
  NOR2X1   g00506(.A(\a[109] ), .B(\a[108] ), .Y(new_n699_));
  INVX1    g00507(.A(new_n699_), .Y(new_n700_));
  MX2X1    g00508(.A(new_n700_), .B(new_n697_), .S0(\a[110] ), .Y(new_n701_));
  INVX1    g00509(.A(\a[110] ), .Y(new_n702_));
  AOI21X1  g00510(.A0(new_n685_), .A1(new_n662_), .B0(new_n687_), .Y(new_n703_));
  INVX1    g00511(.A(new_n675_), .Y(new_n704_));
  OAI21X1  g00512(.A0(new_n704_), .A1(new_n703_), .B0(new_n193_), .Y(new_n705_));
  NAND2X1  g00513(.A(new_n685_), .B(new_n662_), .Y(new_n706_));
  NOR2X1   g00514(.A(new_n671_), .B(new_n687_), .Y(new_n707_));
  INVX1    g00515(.A(new_n695_), .Y(new_n708_));
  AOI21X1  g00516(.A0(new_n707_), .A1(new_n706_), .B0(new_n708_), .Y(new_n709_));
  AOI21X1  g00517(.A0(new_n709_), .A1(new_n705_), .B0(new_n702_), .Y(new_n710_));
  NAND2X1  g00518(.A(new_n699_), .B(new_n702_), .Y(new_n711_));
  NAND2X1  g00519(.A(new_n711_), .B(new_n578_), .Y(new_n712_));
  OR2X1    g00520(.A(new_n712_), .B(new_n575_), .Y(new_n713_));
  NOR4X1   g00521(.A(new_n713_), .B(new_n710_), .C(new_n672_), .D(new_n692_), .Y(new_n714_));
  INVX1    g00522(.A(\a[111] ), .Y(new_n715_));
  AOI21X1  g00523(.A0(new_n709_), .A1(new_n705_), .B0(\a[110] ), .Y(new_n716_));
  OAI21X1  g00524(.A0(new_n696_), .A1(new_n676_), .B0(new_n594_), .Y(new_n717_));
  OAI21X1  g00525(.A0(new_n716_), .A1(new_n715_), .B0(new_n717_), .Y(new_n718_));
  OAI22X1  g00526(.A0(new_n718_), .A1(new_n714_), .B0(new_n701_), .B1(new_n582_), .Y(new_n719_));
  AND2X1   g00527(.A(new_n719_), .B(\asqrt[57] ), .Y(new_n720_));
  OR4X1    g00528(.A(new_n713_), .B(new_n710_), .C(new_n672_), .D(new_n692_), .Y(new_n721_));
  OAI21X1  g00529(.A0(new_n696_), .A1(new_n676_), .B0(new_n702_), .Y(new_n722_));
  AOI21X1  g00530(.A0(new_n709_), .A1(new_n705_), .B0(new_n607_), .Y(new_n723_));
  AOI21X1  g00531(.A0(new_n722_), .A1(\a[111] ), .B0(new_n723_), .Y(new_n724_));
  NAND2X1  g00532(.A(new_n724_), .B(new_n721_), .Y(new_n725_));
  OAI21X1  g00533(.A0(new_n697_), .A1(new_n702_), .B0(new_n711_), .Y(new_n726_));
  AOI21X1  g00534(.A0(new_n726_), .A1(\asqrt[56] ), .B0(\asqrt[57] ), .Y(new_n727_));
  AND2X1   g00535(.A(new_n707_), .B(new_n706_), .Y(new_n728_));
  OR2X1    g00536(.A(new_n694_), .B(new_n582_), .Y(new_n729_));
  OR4X1    g00537(.A(new_n729_), .B(new_n691_), .C(new_n728_), .D(new_n676_), .Y(new_n730_));
  AOI21X1  g00538(.A0(new_n730_), .A1(new_n717_), .B0(new_n597_), .Y(new_n731_));
  NOR4X1   g00539(.A(new_n729_), .B(new_n691_), .C(new_n728_), .D(new_n676_), .Y(new_n732_));
  NOR3X1   g00540(.A(new_n732_), .B(new_n723_), .C(\a[112] ), .Y(new_n733_));
  NOR2X1   g00541(.A(new_n733_), .B(new_n731_), .Y(new_n734_));
  AOI21X1  g00542(.A0(new_n727_), .A1(new_n725_), .B0(new_n734_), .Y(new_n735_));
  OAI21X1  g00543(.A0(new_n735_), .A1(new_n720_), .B0(\asqrt[58] ), .Y(new_n736_));
  AOI22X1  g00544(.A0(new_n724_), .A1(new_n721_), .B0(new_n726_), .B1(\asqrt[56] ), .Y(new_n737_));
  OAI21X1  g00545(.A0(new_n737_), .A1(new_n481_), .B0(new_n399_), .Y(new_n738_));
  AND2X1   g00546(.A(new_n645_), .B(new_n643_), .Y(new_n739_));
  NOR3X1   g00547(.A(new_n604_), .B(new_n739_), .C(new_n596_), .Y(new_n740_));
  OAI21X1  g00548(.A0(new_n696_), .A1(new_n676_), .B0(new_n740_), .Y(new_n741_));
  AOI21X1  g00549(.A0(new_n595_), .A1(\asqrt[57] ), .B0(new_n604_), .Y(new_n742_));
  OAI21X1  g00550(.A0(new_n696_), .A1(new_n676_), .B0(new_n742_), .Y(new_n743_));
  NAND2X1  g00551(.A(new_n743_), .B(new_n739_), .Y(new_n744_));
  NAND2X1  g00552(.A(new_n744_), .B(new_n741_), .Y(new_n745_));
  OAI21X1  g00553(.A0(new_n738_), .A1(new_n735_), .B0(new_n745_), .Y(new_n746_));
  AOI21X1  g00554(.A0(new_n746_), .A1(new_n736_), .B0(new_n328_), .Y(new_n747_));
  AND2X1   g00555(.A(new_n650_), .B(new_n648_), .Y(new_n748_));
  NOR3X1   g00556(.A(new_n615_), .B(new_n748_), .C(new_n649_), .Y(new_n749_));
  OAI21X1  g00557(.A0(new_n696_), .A1(new_n676_), .B0(new_n749_), .Y(new_n750_));
  NOR2X1   g00558(.A(new_n748_), .B(new_n649_), .Y(new_n751_));
  OAI21X1  g00559(.A0(new_n696_), .A1(new_n676_), .B0(new_n751_), .Y(new_n752_));
  NAND2X1  g00560(.A(new_n752_), .B(new_n615_), .Y(new_n753_));
  AND2X1   g00561(.A(new_n753_), .B(new_n750_), .Y(new_n754_));
  INVX1    g00562(.A(new_n754_), .Y(new_n755_));
  NAND3X1  g00563(.A(new_n746_), .B(new_n736_), .C(new_n328_), .Y(new_n756_));
  AOI21X1  g00564(.A0(new_n756_), .A1(new_n755_), .B0(new_n747_), .Y(new_n757_));
  OR2X1    g00565(.A(new_n757_), .B(new_n292_), .Y(new_n758_));
  OR2X1    g00566(.A(new_n737_), .B(new_n481_), .Y(new_n759_));
  AND2X1   g00567(.A(new_n724_), .B(new_n721_), .Y(new_n760_));
  OAI21X1  g00568(.A0(new_n701_), .A1(new_n582_), .B0(new_n481_), .Y(new_n761_));
  OR2X1    g00569(.A(new_n733_), .B(new_n731_), .Y(new_n762_));
  OAI21X1  g00570(.A0(new_n761_), .A1(new_n760_), .B0(new_n762_), .Y(new_n763_));
  AOI21X1  g00571(.A0(new_n763_), .A1(new_n759_), .B0(new_n399_), .Y(new_n764_));
  AOI21X1  g00572(.A0(new_n719_), .A1(\asqrt[57] ), .B0(\asqrt[58] ), .Y(new_n765_));
  AOI22X1  g00573(.A0(new_n744_), .A1(new_n741_), .B0(new_n765_), .B1(new_n763_), .Y(new_n766_));
  NOR3X1   g00574(.A(new_n766_), .B(new_n764_), .C(\asqrt[59] ), .Y(new_n767_));
  NOR2X1   g00575(.A(new_n767_), .B(new_n754_), .Y(new_n768_));
  NOR3X1   g00576(.A(new_n655_), .B(new_n623_), .C(new_n617_), .Y(new_n769_));
  OAI21X1  g00577(.A0(new_n696_), .A1(new_n676_), .B0(new_n769_), .Y(new_n770_));
  NOR3X1   g00578(.A(new_n697_), .B(new_n655_), .C(new_n617_), .Y(new_n771_));
  OR2X1    g00579(.A(new_n771_), .B(new_n622_), .Y(new_n772_));
  AND2X1   g00580(.A(new_n772_), .B(new_n770_), .Y(new_n773_));
  INVX1    g00581(.A(new_n773_), .Y(new_n774_));
  OR2X1    g00582(.A(new_n747_), .B(\asqrt[60] ), .Y(new_n775_));
  OAI21X1  g00583(.A0(new_n775_), .A1(new_n768_), .B0(new_n774_), .Y(new_n776_));
  AOI21X1  g00584(.A0(new_n776_), .A1(new_n758_), .B0(new_n217_), .Y(new_n777_));
  AOI21X1  g00585(.A0(new_n679_), .A1(new_n678_), .B0(new_n633_), .Y(new_n778_));
  AND2X1   g00586(.A(new_n778_), .B(new_n626_), .Y(new_n779_));
  AOI22X1  g00587(.A0(new_n679_), .A1(new_n678_), .B0(new_n656_), .B1(\asqrt[60] ), .Y(new_n780_));
  AOI21X1  g00588(.A0(new_n780_), .A1(\asqrt[55] ), .B0(new_n632_), .Y(new_n781_));
  AOI21X1  g00589(.A0(new_n779_), .A1(\asqrt[55] ), .B0(new_n781_), .Y(new_n782_));
  OAI21X1  g00590(.A0(new_n766_), .A1(new_n764_), .B0(\asqrt[59] ), .Y(new_n783_));
  OAI21X1  g00591(.A0(new_n767_), .A1(new_n754_), .B0(new_n783_), .Y(new_n784_));
  AOI21X1  g00592(.A0(new_n784_), .A1(\asqrt[60] ), .B0(\asqrt[61] ), .Y(new_n785_));
  AOI21X1  g00593(.A0(new_n785_), .A1(new_n776_), .B0(new_n782_), .Y(new_n786_));
  OAI21X1  g00594(.A0(new_n786_), .A1(new_n777_), .B0(\asqrt[62] ), .Y(new_n787_));
  AND2X1   g00595(.A(new_n657_), .B(new_n635_), .Y(new_n788_));
  NOR3X1   g00596(.A(new_n788_), .B(new_n682_), .C(new_n636_), .Y(new_n789_));
  NOR3X1   g00597(.A(new_n697_), .B(new_n788_), .C(new_n636_), .Y(new_n790_));
  NOR2X1   g00598(.A(new_n790_), .B(new_n641_), .Y(new_n791_));
  AOI21X1  g00599(.A0(new_n789_), .A1(\asqrt[55] ), .B0(new_n791_), .Y(new_n792_));
  NOR3X1   g00600(.A(new_n786_), .B(new_n777_), .C(\asqrt[62] ), .Y(new_n793_));
  OAI21X1  g00601(.A0(new_n793_), .A1(new_n792_), .B0(new_n787_), .Y(new_n794_));
  NOR4X1   g00602(.A(new_n697_), .B(new_n664_), .C(new_n662_), .D(new_n687_), .Y(new_n795_));
  NAND3X1  g00603(.A(\asqrt[55] ), .B(new_n685_), .C(new_n659_), .Y(new_n796_));
  AOI21X1  g00604(.A0(new_n796_), .A1(new_n662_), .B0(new_n795_), .Y(new_n797_));
  INVX1    g00605(.A(new_n797_), .Y(new_n798_));
  NOR2X1   g00606(.A(new_n670_), .B(new_n703_), .Y(new_n799_));
  AOI21X1  g00607(.A0(new_n799_), .A1(\asqrt[55] ), .B0(new_n728_), .Y(new_n800_));
  AND2X1   g00608(.A(new_n800_), .B(new_n798_), .Y(new_n801_));
  AOI21X1  g00609(.A0(new_n801_), .A1(new_n794_), .B0(\asqrt[63] ), .Y(new_n802_));
  NOR2X1   g00610(.A(new_n793_), .B(new_n792_), .Y(new_n803_));
  NAND2X1  g00611(.A(new_n797_), .B(new_n787_), .Y(new_n804_));
  AOI21X1  g00612(.A0(new_n709_), .A1(new_n705_), .B0(new_n670_), .Y(new_n805_));
  AOI21X1  g00613(.A0(new_n671_), .A1(new_n665_), .B0(new_n193_), .Y(new_n806_));
  OAI21X1  g00614(.A0(new_n805_), .A1(new_n665_), .B0(new_n806_), .Y(new_n807_));
  NOR4X1   g00615(.A(new_n694_), .B(new_n691_), .C(new_n669_), .D(new_n667_), .Y(new_n808_));
  OAI21X1  g00616(.A0(new_n688_), .A1(new_n686_), .B0(new_n808_), .Y(new_n809_));
  NOR2X1   g00617(.A(new_n809_), .B(new_n676_), .Y(new_n810_));
  INVX1    g00618(.A(new_n810_), .Y(new_n811_));
  AND2X1   g00619(.A(new_n811_), .B(new_n807_), .Y(new_n812_));
  OAI21X1  g00620(.A0(new_n804_), .A1(new_n803_), .B0(new_n812_), .Y(new_n813_));
  OR2X1    g00621(.A(new_n813_), .B(new_n802_), .Y(\asqrt[54] ));
  NOR2X1   g00622(.A(\a[107] ), .B(\a[106] ), .Y(new_n815_));
  MX2X1    g00623(.A(new_n815_), .B(\asqrt[54] ), .S0(\a[108] ), .Y(new_n816_));
  OAI21X1  g00624(.A0(new_n813_), .A1(new_n802_), .B0(\a[108] ), .Y(new_n817_));
  NOR3X1   g00625(.A(\a[108] ), .B(\a[107] ), .C(\a[106] ), .Y(new_n818_));
  OR2X1    g00626(.A(new_n818_), .B(new_n694_), .Y(new_n819_));
  NOR4X1   g00627(.A(new_n819_), .B(new_n691_), .C(new_n728_), .D(new_n676_), .Y(new_n820_));
  NAND2X1  g00628(.A(new_n820_), .B(new_n817_), .Y(new_n821_));
  INVX1    g00629(.A(\a[108] ), .Y(new_n822_));
  OAI21X1  g00630(.A0(new_n813_), .A1(new_n802_), .B0(new_n822_), .Y(new_n823_));
  AND2X1   g00631(.A(new_n784_), .B(\asqrt[60] ), .Y(new_n824_));
  OR2X1    g00632(.A(new_n767_), .B(new_n754_), .Y(new_n825_));
  NOR2X1   g00633(.A(new_n747_), .B(\asqrt[60] ), .Y(new_n826_));
  AOI21X1  g00634(.A0(new_n826_), .A1(new_n825_), .B0(new_n773_), .Y(new_n827_));
  OAI21X1  g00635(.A0(new_n827_), .A1(new_n824_), .B0(\asqrt[61] ), .Y(new_n828_));
  INVX1    g00636(.A(new_n782_), .Y(new_n829_));
  OAI21X1  g00637(.A0(new_n757_), .A1(new_n292_), .B0(new_n217_), .Y(new_n830_));
  OAI21X1  g00638(.A0(new_n830_), .A1(new_n827_), .B0(new_n829_), .Y(new_n831_));
  AOI21X1  g00639(.A0(new_n831_), .A1(new_n828_), .B0(new_n199_), .Y(new_n832_));
  INVX1    g00640(.A(new_n792_), .Y(new_n833_));
  NAND3X1  g00641(.A(new_n831_), .B(new_n828_), .C(new_n199_), .Y(new_n834_));
  AOI21X1  g00642(.A0(new_n834_), .A1(new_n833_), .B0(new_n832_), .Y(new_n835_));
  INVX1    g00643(.A(new_n801_), .Y(new_n836_));
  OAI21X1  g00644(.A0(new_n836_), .A1(new_n835_), .B0(new_n193_), .Y(new_n837_));
  OR2X1    g00645(.A(new_n793_), .B(new_n792_), .Y(new_n838_));
  AND2X1   g00646(.A(new_n797_), .B(new_n787_), .Y(new_n839_));
  INVX1    g00647(.A(new_n812_), .Y(new_n840_));
  AOI21X1  g00648(.A0(new_n839_), .A1(new_n838_), .B0(new_n840_), .Y(new_n841_));
  AOI21X1  g00649(.A0(new_n841_), .A1(new_n837_), .B0(new_n700_), .Y(new_n842_));
  AOI21X1  g00650(.A0(new_n823_), .A1(\a[109] ), .B0(new_n842_), .Y(new_n843_));
  AOI22X1  g00651(.A0(new_n843_), .A1(new_n821_), .B0(new_n816_), .B1(\asqrt[55] ), .Y(new_n844_));
  OR2X1    g00652(.A(new_n844_), .B(new_n582_), .Y(new_n845_));
  AND2X1   g00653(.A(new_n843_), .B(new_n821_), .Y(new_n846_));
  AOI21X1  g00654(.A0(\asqrt[54] ), .A1(\a[108] ), .B0(new_n818_), .Y(new_n847_));
  OAI21X1  g00655(.A0(new_n847_), .A1(new_n697_), .B0(new_n582_), .Y(new_n848_));
  OAI21X1  g00656(.A0(new_n813_), .A1(new_n802_), .B0(new_n699_), .Y(new_n849_));
  INVX1    g00657(.A(new_n807_), .Y(new_n850_));
  NOR3X1   g00658(.A(new_n810_), .B(new_n850_), .C(new_n697_), .Y(new_n851_));
  OAI21X1  g00659(.A0(new_n804_), .A1(new_n803_), .B0(new_n851_), .Y(new_n852_));
  OR2X1    g00660(.A(new_n852_), .B(new_n802_), .Y(new_n853_));
  AOI21X1  g00661(.A0(new_n853_), .A1(new_n849_), .B0(new_n702_), .Y(new_n854_));
  OAI21X1  g00662(.A0(new_n852_), .A1(new_n802_), .B0(new_n702_), .Y(new_n855_));
  NOR2X1   g00663(.A(new_n855_), .B(new_n842_), .Y(new_n856_));
  OR2X1    g00664(.A(new_n856_), .B(new_n854_), .Y(new_n857_));
  OAI21X1  g00665(.A0(new_n848_), .A1(new_n846_), .B0(new_n857_), .Y(new_n858_));
  AOI21X1  g00666(.A0(new_n858_), .A1(new_n845_), .B0(new_n481_), .Y(new_n859_));
  AOI21X1  g00667(.A0(new_n726_), .A1(\asqrt[56] ), .B0(new_n714_), .Y(new_n860_));
  AND2X1   g00668(.A(new_n860_), .B(new_n718_), .Y(new_n861_));
  OAI21X1  g00669(.A0(new_n813_), .A1(new_n802_), .B0(new_n860_), .Y(new_n862_));
  AOI22X1  g00670(.A0(new_n862_), .A1(new_n724_), .B0(new_n861_), .B1(\asqrt[54] ), .Y(new_n863_));
  AND2X1   g00671(.A(new_n820_), .B(new_n817_), .Y(new_n864_));
  INVX1    g00672(.A(\a[109] ), .Y(new_n865_));
  AOI21X1  g00673(.A0(new_n841_), .A1(new_n837_), .B0(\a[108] ), .Y(new_n866_));
  OAI21X1  g00674(.A0(new_n866_), .A1(new_n865_), .B0(new_n849_), .Y(new_n867_));
  OAI22X1  g00675(.A0(new_n867_), .A1(new_n864_), .B0(new_n847_), .B1(new_n697_), .Y(new_n868_));
  AOI21X1  g00676(.A0(new_n868_), .A1(\asqrt[56] ), .B0(\asqrt[57] ), .Y(new_n869_));
  AOI21X1  g00677(.A0(new_n869_), .A1(new_n858_), .B0(new_n863_), .Y(new_n870_));
  OAI21X1  g00678(.A0(new_n870_), .A1(new_n859_), .B0(\asqrt[58] ), .Y(new_n871_));
  AOI21X1  g00679(.A0(new_n727_), .A1(new_n725_), .B0(new_n762_), .Y(new_n872_));
  AND2X1   g00680(.A(new_n872_), .B(new_n759_), .Y(new_n873_));
  AOI22X1  g00681(.A0(new_n727_), .A1(new_n725_), .B0(new_n719_), .B1(\asqrt[57] ), .Y(new_n874_));
  OAI21X1  g00682(.A0(new_n813_), .A1(new_n802_), .B0(new_n874_), .Y(new_n875_));
  AOI22X1  g00683(.A0(new_n875_), .A1(new_n762_), .B0(new_n873_), .B1(\asqrt[54] ), .Y(new_n876_));
  NOR3X1   g00684(.A(new_n870_), .B(new_n859_), .C(\asqrt[58] ), .Y(new_n877_));
  OAI21X1  g00685(.A0(new_n877_), .A1(new_n876_), .B0(new_n871_), .Y(new_n878_));
  AND2X1   g00686(.A(new_n878_), .B(\asqrt[59] ), .Y(new_n879_));
  INVX1    g00687(.A(new_n876_), .Y(new_n880_));
  AND2X1   g00688(.A(new_n868_), .B(\asqrt[56] ), .Y(new_n881_));
  NAND2X1  g00689(.A(new_n843_), .B(new_n821_), .Y(new_n882_));
  AOI21X1  g00690(.A0(new_n816_), .A1(\asqrt[55] ), .B0(\asqrt[56] ), .Y(new_n883_));
  NOR2X1   g00691(.A(new_n856_), .B(new_n854_), .Y(new_n884_));
  AOI21X1  g00692(.A0(new_n883_), .A1(new_n882_), .B0(new_n884_), .Y(new_n885_));
  OAI21X1  g00693(.A0(new_n885_), .A1(new_n881_), .B0(\asqrt[57] ), .Y(new_n886_));
  INVX1    g00694(.A(new_n863_), .Y(new_n887_));
  OAI21X1  g00695(.A0(new_n844_), .A1(new_n582_), .B0(new_n481_), .Y(new_n888_));
  OAI21X1  g00696(.A0(new_n888_), .A1(new_n885_), .B0(new_n887_), .Y(new_n889_));
  NAND3X1  g00697(.A(new_n889_), .B(new_n886_), .C(new_n399_), .Y(new_n890_));
  NAND2X1  g00698(.A(new_n890_), .B(new_n880_), .Y(new_n891_));
  AOI21X1  g00699(.A0(new_n889_), .A1(new_n886_), .B0(new_n399_), .Y(new_n892_));
  NOR2X1   g00700(.A(new_n892_), .B(\asqrt[59] ), .Y(new_n893_));
  AND2X1   g00701(.A(new_n765_), .B(new_n763_), .Y(new_n894_));
  NOR3X1   g00702(.A(new_n745_), .B(new_n894_), .C(new_n764_), .Y(new_n895_));
  NOR2X1   g00703(.A(new_n894_), .B(new_n764_), .Y(new_n896_));
  OAI21X1  g00704(.A0(new_n813_), .A1(new_n802_), .B0(new_n896_), .Y(new_n897_));
  AOI22X1  g00705(.A0(new_n897_), .A1(new_n745_), .B0(new_n895_), .B1(\asqrt[54] ), .Y(new_n898_));
  AOI21X1  g00706(.A0(new_n893_), .A1(new_n891_), .B0(new_n898_), .Y(new_n899_));
  OAI21X1  g00707(.A0(new_n899_), .A1(new_n879_), .B0(\asqrt[60] ), .Y(new_n900_));
  NAND4X1  g00708(.A(\asqrt[54] ), .B(new_n756_), .C(new_n754_), .D(new_n783_), .Y(new_n901_));
  NOR2X1   g00709(.A(new_n813_), .B(new_n802_), .Y(new_n902_));
  NOR3X1   g00710(.A(new_n902_), .B(new_n767_), .C(new_n747_), .Y(new_n903_));
  OAI21X1  g00711(.A0(new_n903_), .A1(new_n754_), .B0(new_n901_), .Y(new_n904_));
  AOI21X1  g00712(.A0(new_n890_), .A1(new_n880_), .B0(new_n892_), .Y(new_n905_));
  OAI21X1  g00713(.A0(new_n905_), .A1(new_n328_), .B0(new_n292_), .Y(new_n906_));
  OAI21X1  g00714(.A0(new_n906_), .A1(new_n899_), .B0(new_n904_), .Y(new_n907_));
  AOI21X1  g00715(.A0(new_n907_), .A1(new_n900_), .B0(new_n217_), .Y(new_n908_));
  AND2X1   g00716(.A(new_n826_), .B(new_n825_), .Y(new_n909_));
  NOR3X1   g00717(.A(new_n909_), .B(new_n774_), .C(new_n824_), .Y(new_n910_));
  AOI22X1  g00718(.A0(new_n826_), .A1(new_n825_), .B0(new_n784_), .B1(\asqrt[60] ), .Y(new_n911_));
  AOI21X1  g00719(.A0(new_n911_), .A1(\asqrt[54] ), .B0(new_n773_), .Y(new_n912_));
  AOI21X1  g00720(.A0(new_n910_), .A1(\asqrt[54] ), .B0(new_n912_), .Y(new_n913_));
  INVX1    g00721(.A(new_n913_), .Y(new_n914_));
  NAND3X1  g00722(.A(new_n907_), .B(new_n900_), .C(new_n217_), .Y(new_n915_));
  AOI21X1  g00723(.A0(new_n915_), .A1(new_n914_), .B0(new_n908_), .Y(new_n916_));
  OR2X1    g00724(.A(new_n916_), .B(new_n199_), .Y(new_n917_));
  AND2X1   g00725(.A(new_n915_), .B(new_n914_), .Y(new_n918_));
  AND2X1   g00726(.A(new_n785_), .B(new_n776_), .Y(new_n919_));
  NOR3X1   g00727(.A(new_n919_), .B(new_n829_), .C(new_n777_), .Y(new_n920_));
  NOR2X1   g00728(.A(new_n919_), .B(new_n777_), .Y(new_n921_));
  AOI21X1  g00729(.A0(new_n921_), .A1(\asqrt[54] ), .B0(new_n782_), .Y(new_n922_));
  AOI21X1  g00730(.A0(new_n920_), .A1(\asqrt[54] ), .B0(new_n922_), .Y(new_n923_));
  INVX1    g00731(.A(new_n923_), .Y(new_n924_));
  OR2X1    g00732(.A(new_n908_), .B(\asqrt[62] ), .Y(new_n925_));
  OAI21X1  g00733(.A0(new_n925_), .A1(new_n918_), .B0(new_n924_), .Y(new_n926_));
  NAND3X1  g00734(.A(new_n834_), .B(new_n792_), .C(new_n787_), .Y(new_n927_));
  AOI21X1  g00735(.A0(new_n841_), .A1(new_n837_), .B0(new_n927_), .Y(new_n928_));
  NAND3X1  g00736(.A(\asqrt[54] ), .B(new_n834_), .C(new_n787_), .Y(new_n929_));
  AOI21X1  g00737(.A0(new_n929_), .A1(new_n833_), .B0(new_n928_), .Y(new_n930_));
  INVX1    g00738(.A(new_n930_), .Y(new_n931_));
  AND2X1   g00739(.A(new_n798_), .B(new_n794_), .Y(new_n932_));
  AOI22X1  g00740(.A0(new_n932_), .A1(\asqrt[54] ), .B0(new_n839_), .B1(new_n838_), .Y(new_n933_));
  AND2X1   g00741(.A(new_n933_), .B(new_n931_), .Y(new_n934_));
  INVX1    g00742(.A(new_n934_), .Y(new_n935_));
  AOI21X1  g00743(.A0(new_n926_), .A1(new_n917_), .B0(new_n935_), .Y(new_n936_));
  OR2X1    g00744(.A(new_n905_), .B(new_n328_), .Y(new_n937_));
  AND2X1   g00745(.A(new_n890_), .B(new_n880_), .Y(new_n938_));
  OR2X1    g00746(.A(new_n892_), .B(\asqrt[59] ), .Y(new_n939_));
  INVX1    g00747(.A(new_n898_), .Y(new_n940_));
  OAI21X1  g00748(.A0(new_n939_), .A1(new_n938_), .B0(new_n940_), .Y(new_n941_));
  AOI21X1  g00749(.A0(new_n941_), .A1(new_n937_), .B0(new_n292_), .Y(new_n942_));
  INVX1    g00750(.A(new_n904_), .Y(new_n943_));
  AOI21X1  g00751(.A0(new_n878_), .A1(\asqrt[59] ), .B0(\asqrt[60] ), .Y(new_n944_));
  AOI21X1  g00752(.A0(new_n944_), .A1(new_n941_), .B0(new_n943_), .Y(new_n945_));
  OAI21X1  g00753(.A0(new_n945_), .A1(new_n942_), .B0(\asqrt[61] ), .Y(new_n946_));
  NOR3X1   g00754(.A(new_n945_), .B(new_n942_), .C(\asqrt[61] ), .Y(new_n947_));
  OAI21X1  g00755(.A0(new_n947_), .A1(new_n913_), .B0(new_n946_), .Y(new_n948_));
  AOI21X1  g00756(.A0(new_n948_), .A1(\asqrt[62] ), .B0(new_n931_), .Y(new_n949_));
  AOI21X1  g00757(.A0(new_n841_), .A1(new_n837_), .B0(new_n797_), .Y(new_n950_));
  AOI21X1  g00758(.A0(new_n798_), .A1(new_n794_), .B0(new_n193_), .Y(new_n951_));
  OAI21X1  g00759(.A0(new_n950_), .A1(new_n794_), .B0(new_n951_), .Y(new_n952_));
  OR2X1    g00760(.A(new_n804_), .B(new_n803_), .Y(new_n953_));
  AND2X1   g00761(.A(new_n796_), .B(new_n662_), .Y(new_n954_));
  NOR4X1   g00762(.A(new_n810_), .B(new_n850_), .C(new_n954_), .D(new_n795_), .Y(new_n955_));
  NAND3X1  g00763(.A(new_n955_), .B(new_n953_), .C(new_n837_), .Y(new_n956_));
  AND2X1   g00764(.A(new_n956_), .B(new_n952_), .Y(new_n957_));
  INVX1    g00765(.A(new_n957_), .Y(new_n958_));
  AOI21X1  g00766(.A0(new_n949_), .A1(new_n926_), .B0(new_n958_), .Y(new_n959_));
  OAI21X1  g00767(.A0(new_n936_), .A1(\asqrt[63] ), .B0(new_n959_), .Y(\asqrt[53] ));
  AND2X1   g00768(.A(new_n948_), .B(\asqrt[62] ), .Y(new_n961_));
  NAND2X1  g00769(.A(new_n915_), .B(new_n914_), .Y(new_n962_));
  NOR2X1   g00770(.A(new_n908_), .B(\asqrt[62] ), .Y(new_n963_));
  AOI21X1  g00771(.A0(new_n963_), .A1(new_n962_), .B0(new_n923_), .Y(new_n964_));
  OAI21X1  g00772(.A0(new_n964_), .A1(new_n961_), .B0(new_n934_), .Y(new_n965_));
  OAI21X1  g00773(.A0(new_n916_), .A1(new_n199_), .B0(new_n930_), .Y(new_n966_));
  OAI21X1  g00774(.A0(new_n966_), .A1(new_n964_), .B0(new_n957_), .Y(new_n967_));
  AOI21X1  g00775(.A0(new_n965_), .A1(new_n193_), .B0(new_n967_), .Y(new_n968_));
  NOR2X1   g00776(.A(\a[105] ), .B(\a[104] ), .Y(new_n969_));
  INVX1    g00777(.A(new_n969_), .Y(new_n970_));
  MX2X1    g00778(.A(new_n970_), .B(new_n968_), .S0(\a[106] ), .Y(new_n971_));
  OR2X1    g00779(.A(new_n971_), .B(new_n902_), .Y(new_n972_));
  INVX1    g00780(.A(\a[106] ), .Y(new_n973_));
  NOR3X1   g00781(.A(\a[106] ), .B(\a[105] ), .C(\a[104] ), .Y(new_n974_));
  NOR3X1   g00782(.A(new_n974_), .B(new_n810_), .C(new_n850_), .Y(new_n975_));
  NAND3X1  g00783(.A(new_n975_), .B(new_n953_), .C(new_n837_), .Y(new_n976_));
  INVX1    g00784(.A(new_n976_), .Y(new_n977_));
  OAI21X1  g00785(.A0(new_n968_), .A1(new_n973_), .B0(new_n977_), .Y(new_n978_));
  OAI21X1  g00786(.A0(new_n968_), .A1(\a[106] ), .B0(\a[107] ), .Y(new_n979_));
  INVX1    g00787(.A(new_n815_), .Y(new_n980_));
  OR2X1    g00788(.A(new_n968_), .B(new_n980_), .Y(new_n981_));
  NAND3X1  g00789(.A(new_n981_), .B(new_n979_), .C(new_n978_), .Y(new_n982_));
  AOI21X1  g00790(.A0(new_n982_), .A1(new_n972_), .B0(new_n697_), .Y(new_n983_));
  MX2X1    g00791(.A(new_n969_), .B(\asqrt[53] ), .S0(\a[106] ), .Y(new_n984_));
  AOI21X1  g00792(.A0(new_n984_), .A1(\asqrt[54] ), .B0(\asqrt[55] ), .Y(new_n985_));
  NAND3X1  g00793(.A(new_n956_), .B(new_n952_), .C(\asqrt[54] ), .Y(new_n986_));
  INVX1    g00794(.A(new_n986_), .Y(new_n987_));
  OAI21X1  g00795(.A0(new_n966_), .A1(new_n964_), .B0(new_n987_), .Y(new_n988_));
  AOI21X1  g00796(.A0(new_n965_), .A1(new_n193_), .B0(new_n988_), .Y(new_n989_));
  AOI21X1  g00797(.A0(\asqrt[53] ), .A1(new_n815_), .B0(new_n989_), .Y(new_n990_));
  OR2X1    g00798(.A(new_n990_), .B(new_n822_), .Y(new_n991_));
  AND2X1   g00799(.A(\asqrt[53] ), .B(new_n815_), .Y(new_n992_));
  OR2X1    g00800(.A(new_n989_), .B(\a[108] ), .Y(new_n993_));
  OR2X1    g00801(.A(new_n993_), .B(new_n992_), .Y(new_n994_));
  AOI22X1  g00802(.A0(new_n994_), .A1(new_n991_), .B0(new_n985_), .B1(new_n982_), .Y(new_n995_));
  OAI21X1  g00803(.A0(new_n995_), .A1(new_n983_), .B0(\asqrt[56] ), .Y(new_n996_));
  AOI21X1  g00804(.A0(new_n816_), .A1(\asqrt[55] ), .B0(new_n864_), .Y(new_n997_));
  NAND3X1  g00805(.A(new_n997_), .B(\asqrt[53] ), .C(new_n867_), .Y(new_n998_));
  INVX1    g00806(.A(new_n997_), .Y(new_n999_));
  OAI21X1  g00807(.A0(new_n999_), .A1(new_n968_), .B0(new_n843_), .Y(new_n1000_));
  AND2X1   g00808(.A(new_n1000_), .B(new_n998_), .Y(new_n1001_));
  NOR3X1   g00809(.A(new_n995_), .B(new_n983_), .C(\asqrt[56] ), .Y(new_n1002_));
  OAI21X1  g00810(.A0(new_n1002_), .A1(new_n1001_), .B0(new_n996_), .Y(new_n1003_));
  AND2X1   g00811(.A(new_n1003_), .B(\asqrt[57] ), .Y(new_n1004_));
  INVX1    g00812(.A(new_n1001_), .Y(new_n1005_));
  AND2X1   g00813(.A(new_n984_), .B(\asqrt[54] ), .Y(new_n1006_));
  AOI21X1  g00814(.A0(\asqrt[53] ), .A1(\a[106] ), .B0(new_n976_), .Y(new_n1007_));
  INVX1    g00815(.A(\a[107] ), .Y(new_n1008_));
  AOI21X1  g00816(.A0(\asqrt[53] ), .A1(new_n973_), .B0(new_n1008_), .Y(new_n1009_));
  NOR3X1   g00817(.A(new_n992_), .B(new_n1009_), .C(new_n1007_), .Y(new_n1010_));
  OAI21X1  g00818(.A0(new_n1010_), .A1(new_n1006_), .B0(\asqrt[55] ), .Y(new_n1011_));
  OAI21X1  g00819(.A0(new_n971_), .A1(new_n902_), .B0(new_n697_), .Y(new_n1012_));
  OAI22X1  g00820(.A0(new_n993_), .A1(new_n992_), .B0(new_n990_), .B1(new_n822_), .Y(new_n1013_));
  OAI21X1  g00821(.A0(new_n1012_), .A1(new_n1010_), .B0(new_n1013_), .Y(new_n1014_));
  NAND3X1  g00822(.A(new_n1014_), .B(new_n1011_), .C(new_n582_), .Y(new_n1015_));
  NAND2X1  g00823(.A(new_n1015_), .B(new_n1005_), .Y(new_n1016_));
  OAI21X1  g00824(.A0(new_n848_), .A1(new_n846_), .B0(new_n884_), .Y(new_n1017_));
  NOR3X1   g00825(.A(new_n1017_), .B(new_n968_), .C(new_n881_), .Y(new_n1018_));
  OAI22X1  g00826(.A0(new_n848_), .A1(new_n846_), .B0(new_n844_), .B1(new_n582_), .Y(new_n1019_));
  OR2X1    g00827(.A(new_n1019_), .B(new_n968_), .Y(new_n1020_));
  AOI21X1  g00828(.A0(new_n1020_), .A1(new_n857_), .B0(new_n1018_), .Y(new_n1021_));
  AOI21X1  g00829(.A0(new_n1014_), .A1(new_n1011_), .B0(new_n582_), .Y(new_n1022_));
  NOR2X1   g00830(.A(new_n1022_), .B(\asqrt[57] ), .Y(new_n1023_));
  AOI21X1  g00831(.A0(new_n1023_), .A1(new_n1016_), .B0(new_n1021_), .Y(new_n1024_));
  OAI21X1  g00832(.A0(new_n1024_), .A1(new_n1004_), .B0(\asqrt[58] ), .Y(new_n1025_));
  AND2X1   g00833(.A(new_n869_), .B(new_n858_), .Y(new_n1026_));
  NOR4X1   g00834(.A(new_n968_), .B(new_n1026_), .C(new_n887_), .D(new_n859_), .Y(new_n1027_));
  OR2X1    g00835(.A(new_n1026_), .B(new_n859_), .Y(new_n1028_));
  OR2X1    g00836(.A(new_n1028_), .B(new_n968_), .Y(new_n1029_));
  AOI21X1  g00837(.A0(new_n1029_), .A1(new_n887_), .B0(new_n1027_), .Y(new_n1030_));
  INVX1    g00838(.A(new_n1030_), .Y(new_n1031_));
  AOI21X1  g00839(.A0(new_n1015_), .A1(new_n1005_), .B0(new_n1022_), .Y(new_n1032_));
  OAI21X1  g00840(.A0(new_n1032_), .A1(new_n481_), .B0(new_n399_), .Y(new_n1033_));
  OAI21X1  g00841(.A0(new_n1033_), .A1(new_n1024_), .B0(new_n1031_), .Y(new_n1034_));
  AOI21X1  g00842(.A0(new_n1034_), .A1(new_n1025_), .B0(new_n328_), .Y(new_n1035_));
  NAND3X1  g00843(.A(new_n890_), .B(new_n876_), .C(new_n871_), .Y(new_n1036_));
  NOR3X1   g00844(.A(new_n968_), .B(new_n877_), .C(new_n892_), .Y(new_n1037_));
  OAI22X1  g00845(.A0(new_n1037_), .A1(new_n876_), .B0(new_n1036_), .B1(new_n968_), .Y(new_n1038_));
  NAND3X1  g00846(.A(new_n1034_), .B(new_n1025_), .C(new_n328_), .Y(new_n1039_));
  AOI21X1  g00847(.A0(new_n1039_), .A1(new_n1038_), .B0(new_n1035_), .Y(new_n1040_));
  OR2X1    g00848(.A(new_n1040_), .B(new_n292_), .Y(new_n1041_));
  AND2X1   g00849(.A(new_n1039_), .B(new_n1038_), .Y(new_n1042_));
  OR2X1    g00850(.A(new_n1035_), .B(\asqrt[60] ), .Y(new_n1043_));
  AND2X1   g00851(.A(new_n893_), .B(new_n891_), .Y(new_n1044_));
  NOR4X1   g00852(.A(new_n968_), .B(new_n940_), .C(new_n1044_), .D(new_n879_), .Y(new_n1045_));
  AOI22X1  g00853(.A0(new_n893_), .A1(new_n891_), .B0(new_n878_), .B1(\asqrt[59] ), .Y(new_n1046_));
  AOI21X1  g00854(.A0(new_n1046_), .A1(\asqrt[53] ), .B0(new_n898_), .Y(new_n1047_));
  NOR2X1   g00855(.A(new_n1047_), .B(new_n1045_), .Y(new_n1048_));
  INVX1    g00856(.A(new_n1048_), .Y(new_n1049_));
  OAI21X1  g00857(.A0(new_n1043_), .A1(new_n1042_), .B0(new_n1049_), .Y(new_n1050_));
  AOI21X1  g00858(.A0(new_n1050_), .A1(new_n1041_), .B0(new_n217_), .Y(new_n1051_));
  AND2X1   g00859(.A(new_n944_), .B(new_n941_), .Y(new_n1052_));
  NOR4X1   g00860(.A(new_n968_), .B(new_n1052_), .C(new_n904_), .D(new_n942_), .Y(new_n1053_));
  NOR2X1   g00861(.A(new_n1052_), .B(new_n942_), .Y(new_n1054_));
  AOI21X1  g00862(.A0(new_n1054_), .A1(\asqrt[53] ), .B0(new_n943_), .Y(new_n1055_));
  NOR2X1   g00863(.A(new_n1055_), .B(new_n1053_), .Y(new_n1056_));
  OR2X1    g00864(.A(new_n1032_), .B(new_n481_), .Y(new_n1057_));
  AND2X1   g00865(.A(new_n1015_), .B(new_n1005_), .Y(new_n1058_));
  INVX1    g00866(.A(new_n1021_), .Y(new_n1059_));
  OR2X1    g00867(.A(new_n1022_), .B(\asqrt[57] ), .Y(new_n1060_));
  OAI21X1  g00868(.A0(new_n1060_), .A1(new_n1058_), .B0(new_n1059_), .Y(new_n1061_));
  AOI21X1  g00869(.A0(new_n1061_), .A1(new_n1057_), .B0(new_n399_), .Y(new_n1062_));
  AOI21X1  g00870(.A0(new_n1003_), .A1(\asqrt[57] ), .B0(\asqrt[58] ), .Y(new_n1063_));
  AOI21X1  g00871(.A0(new_n1063_), .A1(new_n1061_), .B0(new_n1030_), .Y(new_n1064_));
  OAI21X1  g00872(.A0(new_n1064_), .A1(new_n1062_), .B0(\asqrt[59] ), .Y(new_n1065_));
  INVX1    g00873(.A(new_n1038_), .Y(new_n1066_));
  NOR3X1   g00874(.A(new_n1064_), .B(new_n1062_), .C(\asqrt[59] ), .Y(new_n1067_));
  OAI21X1  g00875(.A0(new_n1067_), .A1(new_n1066_), .B0(new_n1065_), .Y(new_n1068_));
  AOI21X1  g00876(.A0(new_n1068_), .A1(\asqrt[60] ), .B0(\asqrt[61] ), .Y(new_n1069_));
  AOI21X1  g00877(.A0(new_n1069_), .A1(new_n1050_), .B0(new_n1056_), .Y(new_n1070_));
  OAI21X1  g00878(.A0(new_n1070_), .A1(new_n1051_), .B0(\asqrt[62] ), .Y(new_n1071_));
  NAND3X1  g00879(.A(new_n915_), .B(new_n913_), .C(new_n946_), .Y(new_n1072_));
  NOR3X1   g00880(.A(new_n968_), .B(new_n947_), .C(new_n908_), .Y(new_n1073_));
  OAI22X1  g00881(.A0(new_n1073_), .A1(new_n913_), .B0(new_n1072_), .B1(new_n968_), .Y(new_n1074_));
  INVX1    g00882(.A(new_n1074_), .Y(new_n1075_));
  NOR3X1   g00883(.A(new_n1070_), .B(new_n1051_), .C(\asqrt[62] ), .Y(new_n1076_));
  OAI21X1  g00884(.A0(new_n1076_), .A1(new_n1075_), .B0(new_n1071_), .Y(new_n1077_));
  OAI21X1  g00885(.A0(new_n925_), .A1(new_n918_), .B0(new_n923_), .Y(new_n1078_));
  NOR3X1   g00886(.A(new_n1078_), .B(new_n968_), .C(new_n961_), .Y(new_n1079_));
  AOI22X1  g00887(.A0(new_n963_), .A1(new_n962_), .B0(new_n948_), .B1(\asqrt[62] ), .Y(new_n1080_));
  AOI21X1  g00888(.A0(new_n1080_), .A1(\asqrt[53] ), .B0(new_n923_), .Y(new_n1081_));
  NOR2X1   g00889(.A(new_n1081_), .B(new_n1079_), .Y(new_n1082_));
  INVX1    g00890(.A(new_n1082_), .Y(new_n1083_));
  AND2X1   g00891(.A(new_n949_), .B(new_n926_), .Y(new_n1084_));
  AOI21X1  g00892(.A0(new_n926_), .A1(new_n917_), .B0(new_n930_), .Y(new_n1085_));
  AOI21X1  g00893(.A0(new_n1085_), .A1(\asqrt[53] ), .B0(new_n1084_), .Y(new_n1086_));
  AND2X1   g00894(.A(new_n1086_), .B(new_n1083_), .Y(new_n1087_));
  AOI21X1  g00895(.A0(new_n1087_), .A1(new_n1077_), .B0(\asqrt[63] ), .Y(new_n1088_));
  AND2X1   g00896(.A(new_n1068_), .B(\asqrt[60] ), .Y(new_n1089_));
  NAND2X1  g00897(.A(new_n1039_), .B(new_n1038_), .Y(new_n1090_));
  NOR2X1   g00898(.A(new_n1035_), .B(\asqrt[60] ), .Y(new_n1091_));
  AOI21X1  g00899(.A0(new_n1091_), .A1(new_n1090_), .B0(new_n1048_), .Y(new_n1092_));
  OAI21X1  g00900(.A0(new_n1092_), .A1(new_n1089_), .B0(\asqrt[61] ), .Y(new_n1093_));
  INVX1    g00901(.A(new_n1056_), .Y(new_n1094_));
  OAI21X1  g00902(.A0(new_n1040_), .A1(new_n292_), .B0(new_n217_), .Y(new_n1095_));
  OAI21X1  g00903(.A0(new_n1095_), .A1(new_n1092_), .B0(new_n1094_), .Y(new_n1096_));
  NAND3X1  g00904(.A(new_n1096_), .B(new_n1093_), .C(new_n199_), .Y(new_n1097_));
  AND2X1   g00905(.A(new_n1097_), .B(new_n1074_), .Y(new_n1098_));
  NAND2X1  g00906(.A(new_n1082_), .B(new_n1071_), .Y(new_n1099_));
  NAND2X1  g00907(.A(new_n926_), .B(new_n917_), .Y(new_n1100_));
  AOI21X1  g00908(.A0(\asqrt[53] ), .A1(new_n931_), .B0(new_n1100_), .Y(new_n1101_));
  NOR3X1   g00909(.A(new_n1101_), .B(new_n1085_), .C(new_n193_), .Y(new_n1102_));
  AND2X1   g00910(.A(new_n965_), .B(new_n193_), .Y(new_n1103_));
  OAI21X1  g00911(.A0(new_n927_), .A1(new_n902_), .B0(new_n956_), .Y(new_n1104_));
  AOI21X1  g00912(.A0(new_n929_), .A1(new_n833_), .B0(new_n1104_), .Y(new_n1105_));
  NAND2X1  g00913(.A(new_n1105_), .B(new_n952_), .Y(new_n1106_));
  OR2X1    g00914(.A(new_n1106_), .B(new_n1084_), .Y(new_n1107_));
  NOR2X1   g00915(.A(new_n1107_), .B(new_n1103_), .Y(new_n1108_));
  NOR2X1   g00916(.A(new_n1108_), .B(new_n1102_), .Y(new_n1109_));
  OAI21X1  g00917(.A0(new_n1099_), .A1(new_n1098_), .B0(new_n1109_), .Y(new_n1110_));
  NOR2X1   g00918(.A(new_n1110_), .B(new_n1088_), .Y(new_n1111_));
  INVX1    g00919(.A(\a[104] ), .Y(new_n1112_));
  NOR2X1   g00920(.A(\a[103] ), .B(\a[102] ), .Y(new_n1113_));
  NAND2X1  g00921(.A(new_n1113_), .B(new_n1112_), .Y(new_n1114_));
  OAI21X1  g00922(.A0(new_n1111_), .A1(new_n1112_), .B0(new_n1114_), .Y(new_n1115_));
  AOI21X1  g00923(.A0(new_n1096_), .A1(new_n1093_), .B0(new_n199_), .Y(new_n1116_));
  AOI21X1  g00924(.A0(new_n1097_), .A1(new_n1074_), .B0(new_n1116_), .Y(new_n1117_));
  INVX1    g00925(.A(new_n1087_), .Y(new_n1118_));
  OAI21X1  g00926(.A0(new_n1118_), .A1(new_n1117_), .B0(new_n193_), .Y(new_n1119_));
  NAND2X1  g00927(.A(new_n1097_), .B(new_n1074_), .Y(new_n1120_));
  AND2X1   g00928(.A(new_n1082_), .B(new_n1071_), .Y(new_n1121_));
  INVX1    g00929(.A(new_n1109_), .Y(new_n1122_));
  AOI21X1  g00930(.A0(new_n1121_), .A1(new_n1120_), .B0(new_n1122_), .Y(new_n1123_));
  AOI21X1  g00931(.A0(new_n1123_), .A1(new_n1119_), .B0(new_n1112_), .Y(new_n1124_));
  NAND3X1  g00932(.A(new_n1114_), .B(new_n956_), .C(new_n952_), .Y(new_n1125_));
  OR4X1    g00933(.A(new_n1125_), .B(new_n1124_), .C(new_n1084_), .D(new_n1103_), .Y(new_n1126_));
  OAI21X1  g00934(.A0(new_n1110_), .A1(new_n1088_), .B0(new_n1112_), .Y(new_n1127_));
  AOI21X1  g00935(.A0(new_n1123_), .A1(new_n1119_), .B0(new_n970_), .Y(new_n1128_));
  AOI21X1  g00936(.A0(new_n1127_), .A1(\a[105] ), .B0(new_n1128_), .Y(new_n1129_));
  AOI22X1  g00937(.A0(new_n1129_), .A1(new_n1126_), .B0(new_n1115_), .B1(\asqrt[53] ), .Y(new_n1130_));
  OR2X1    g00938(.A(new_n1130_), .B(new_n902_), .Y(new_n1131_));
  AND2X1   g00939(.A(new_n1129_), .B(new_n1126_), .Y(new_n1132_));
  INVX1    g00940(.A(new_n1113_), .Y(new_n1133_));
  MX2X1    g00941(.A(new_n1133_), .B(new_n1111_), .S0(\a[104] ), .Y(new_n1134_));
  OAI21X1  g00942(.A0(new_n1134_), .A1(new_n968_), .B0(new_n902_), .Y(new_n1135_));
  OAI21X1  g00943(.A0(new_n1110_), .A1(new_n1088_), .B0(new_n969_), .Y(new_n1136_));
  AND2X1   g00944(.A(new_n1121_), .B(new_n1120_), .Y(new_n1137_));
  OAI21X1  g00945(.A0(new_n1107_), .A1(new_n1103_), .B0(\asqrt[53] ), .Y(new_n1138_));
  OR4X1    g00946(.A(new_n1138_), .B(new_n1102_), .C(new_n1137_), .D(new_n1088_), .Y(new_n1139_));
  AOI21X1  g00947(.A0(new_n1139_), .A1(new_n1136_), .B0(new_n973_), .Y(new_n1140_));
  NOR4X1   g00948(.A(new_n1138_), .B(new_n1102_), .C(new_n1137_), .D(new_n1088_), .Y(new_n1141_));
  NOR3X1   g00949(.A(new_n1141_), .B(new_n1128_), .C(\a[106] ), .Y(new_n1142_));
  OR2X1    g00950(.A(new_n1142_), .B(new_n1140_), .Y(new_n1143_));
  OAI21X1  g00951(.A0(new_n1135_), .A1(new_n1132_), .B0(new_n1143_), .Y(new_n1144_));
  AOI21X1  g00952(.A0(new_n1144_), .A1(new_n1131_), .B0(new_n697_), .Y(new_n1145_));
  AND2X1   g00953(.A(new_n981_), .B(new_n979_), .Y(new_n1146_));
  NOR3X1   g00954(.A(new_n1146_), .B(new_n1007_), .C(new_n1006_), .Y(new_n1147_));
  OAI21X1  g00955(.A0(new_n1110_), .A1(new_n1088_), .B0(new_n1147_), .Y(new_n1148_));
  AOI21X1  g00956(.A0(new_n984_), .A1(\asqrt[54] ), .B0(new_n1007_), .Y(new_n1149_));
  OAI21X1  g00957(.A0(new_n1110_), .A1(new_n1088_), .B0(new_n1149_), .Y(new_n1150_));
  NAND2X1  g00958(.A(new_n1150_), .B(new_n1146_), .Y(new_n1151_));
  NOR4X1   g00959(.A(new_n1125_), .B(new_n1124_), .C(new_n1084_), .D(new_n1103_), .Y(new_n1152_));
  INVX1    g00960(.A(\a[105] ), .Y(new_n1153_));
  AOI21X1  g00961(.A0(new_n1123_), .A1(new_n1119_), .B0(\a[104] ), .Y(new_n1154_));
  OAI21X1  g00962(.A0(new_n1154_), .A1(new_n1153_), .B0(new_n1136_), .Y(new_n1155_));
  OAI22X1  g00963(.A0(new_n1155_), .A1(new_n1152_), .B0(new_n1134_), .B1(new_n968_), .Y(new_n1156_));
  AOI21X1  g00964(.A0(new_n1156_), .A1(\asqrt[54] ), .B0(\asqrt[55] ), .Y(new_n1157_));
  AOI22X1  g00965(.A0(new_n1157_), .A1(new_n1144_), .B0(new_n1151_), .B1(new_n1148_), .Y(new_n1158_));
  OAI21X1  g00966(.A0(new_n1158_), .A1(new_n1145_), .B0(\asqrt[56] ), .Y(new_n1159_));
  AND2X1   g00967(.A(new_n985_), .B(new_n982_), .Y(new_n1160_));
  NOR3X1   g00968(.A(new_n1013_), .B(new_n1160_), .C(new_n983_), .Y(new_n1161_));
  OAI21X1  g00969(.A0(new_n1110_), .A1(new_n1088_), .B0(new_n1161_), .Y(new_n1162_));
  NOR2X1   g00970(.A(new_n1160_), .B(new_n983_), .Y(new_n1163_));
  OAI21X1  g00971(.A0(new_n1110_), .A1(new_n1088_), .B0(new_n1163_), .Y(new_n1164_));
  NAND2X1  g00972(.A(new_n1164_), .B(new_n1013_), .Y(new_n1165_));
  AND2X1   g00973(.A(new_n1165_), .B(new_n1162_), .Y(new_n1166_));
  NOR3X1   g00974(.A(new_n1158_), .B(new_n1145_), .C(\asqrt[56] ), .Y(new_n1167_));
  OAI21X1  g00975(.A0(new_n1167_), .A1(new_n1166_), .B0(new_n1159_), .Y(new_n1168_));
  AND2X1   g00976(.A(new_n1168_), .B(\asqrt[57] ), .Y(new_n1169_));
  OR2X1    g00977(.A(new_n1167_), .B(new_n1166_), .Y(new_n1170_));
  NOR3X1   g00978(.A(new_n1002_), .B(new_n1005_), .C(new_n1022_), .Y(new_n1171_));
  OAI21X1  g00979(.A0(new_n1110_), .A1(new_n1088_), .B0(new_n1171_), .Y(new_n1172_));
  NOR3X1   g00980(.A(new_n1111_), .B(new_n1002_), .C(new_n1022_), .Y(new_n1173_));
  OR2X1    g00981(.A(new_n1173_), .B(new_n1001_), .Y(new_n1174_));
  AND2X1   g00982(.A(new_n1174_), .B(new_n1172_), .Y(new_n1175_));
  AND2X1   g00983(.A(new_n1156_), .B(\asqrt[54] ), .Y(new_n1176_));
  NAND2X1  g00984(.A(new_n1129_), .B(new_n1126_), .Y(new_n1177_));
  AOI21X1  g00985(.A0(new_n1115_), .A1(\asqrt[53] ), .B0(\asqrt[54] ), .Y(new_n1178_));
  NOR2X1   g00986(.A(new_n1142_), .B(new_n1140_), .Y(new_n1179_));
  AOI21X1  g00987(.A0(new_n1178_), .A1(new_n1177_), .B0(new_n1179_), .Y(new_n1180_));
  OAI21X1  g00988(.A0(new_n1180_), .A1(new_n1176_), .B0(\asqrt[55] ), .Y(new_n1181_));
  NAND2X1  g00989(.A(new_n1151_), .B(new_n1148_), .Y(new_n1182_));
  OAI21X1  g00990(.A0(new_n1130_), .A1(new_n902_), .B0(new_n697_), .Y(new_n1183_));
  OAI21X1  g00991(.A0(new_n1183_), .A1(new_n1180_), .B0(new_n1182_), .Y(new_n1184_));
  AOI21X1  g00992(.A0(new_n1184_), .A1(new_n1181_), .B0(new_n582_), .Y(new_n1185_));
  NOR2X1   g00993(.A(new_n1185_), .B(\asqrt[57] ), .Y(new_n1186_));
  AOI21X1  g00994(.A0(new_n1186_), .A1(new_n1170_), .B0(new_n1175_), .Y(new_n1187_));
  OAI21X1  g00995(.A0(new_n1187_), .A1(new_n1169_), .B0(\asqrt[58] ), .Y(new_n1188_));
  INVX1    g00996(.A(new_n1111_), .Y(\asqrt[52] ));
  AOI21X1  g00997(.A0(new_n1023_), .A1(new_n1016_), .B0(new_n1059_), .Y(new_n1190_));
  AND2X1   g00998(.A(new_n1190_), .B(new_n1057_), .Y(new_n1191_));
  AOI22X1  g00999(.A0(new_n1023_), .A1(new_n1016_), .B0(new_n1003_), .B1(\asqrt[57] ), .Y(new_n1192_));
  AOI21X1  g01000(.A0(new_n1192_), .A1(\asqrt[52] ), .B0(new_n1021_), .Y(new_n1193_));
  AOI21X1  g01001(.A0(new_n1191_), .A1(\asqrt[52] ), .B0(new_n1193_), .Y(new_n1194_));
  INVX1    g01002(.A(new_n1194_), .Y(new_n1195_));
  INVX1    g01003(.A(new_n1166_), .Y(new_n1196_));
  NAND3X1  g01004(.A(new_n1184_), .B(new_n1181_), .C(new_n582_), .Y(new_n1197_));
  AOI21X1  g01005(.A0(new_n1197_), .A1(new_n1196_), .B0(new_n1185_), .Y(new_n1198_));
  OAI21X1  g01006(.A0(new_n1198_), .A1(new_n481_), .B0(new_n399_), .Y(new_n1199_));
  OAI21X1  g01007(.A0(new_n1199_), .A1(new_n1187_), .B0(new_n1195_), .Y(new_n1200_));
  AOI21X1  g01008(.A0(new_n1200_), .A1(new_n1188_), .B0(new_n328_), .Y(new_n1201_));
  AND2X1   g01009(.A(new_n1063_), .B(new_n1061_), .Y(new_n1202_));
  NOR3X1   g01010(.A(new_n1202_), .B(new_n1031_), .C(new_n1062_), .Y(new_n1203_));
  NOR3X1   g01011(.A(new_n1111_), .B(new_n1202_), .C(new_n1062_), .Y(new_n1204_));
  NOR2X1   g01012(.A(new_n1204_), .B(new_n1030_), .Y(new_n1205_));
  AOI21X1  g01013(.A0(new_n1203_), .A1(\asqrt[52] ), .B0(new_n1205_), .Y(new_n1206_));
  INVX1    g01014(.A(new_n1206_), .Y(new_n1207_));
  NAND3X1  g01015(.A(new_n1200_), .B(new_n1188_), .C(new_n328_), .Y(new_n1208_));
  AOI21X1  g01016(.A0(new_n1208_), .A1(new_n1207_), .B0(new_n1201_), .Y(new_n1209_));
  OR2X1    g01017(.A(new_n1209_), .B(new_n292_), .Y(new_n1210_));
  OR2X1    g01018(.A(new_n1198_), .B(new_n481_), .Y(new_n1211_));
  NOR2X1   g01019(.A(new_n1167_), .B(new_n1166_), .Y(new_n1212_));
  INVX1    g01020(.A(new_n1175_), .Y(new_n1213_));
  OR2X1    g01021(.A(new_n1185_), .B(\asqrt[57] ), .Y(new_n1214_));
  OAI21X1  g01022(.A0(new_n1214_), .A1(new_n1212_), .B0(new_n1213_), .Y(new_n1215_));
  AOI21X1  g01023(.A0(new_n1215_), .A1(new_n1211_), .B0(new_n399_), .Y(new_n1216_));
  AOI21X1  g01024(.A0(new_n1168_), .A1(\asqrt[57] ), .B0(\asqrt[58] ), .Y(new_n1217_));
  AOI21X1  g01025(.A0(new_n1217_), .A1(new_n1215_), .B0(new_n1194_), .Y(new_n1218_));
  NOR3X1   g01026(.A(new_n1218_), .B(new_n1216_), .C(\asqrt[59] ), .Y(new_n1219_));
  NOR2X1   g01027(.A(new_n1219_), .B(new_n1206_), .Y(new_n1220_));
  OR4X1    g01028(.A(new_n1111_), .B(new_n1067_), .C(new_n1038_), .D(new_n1035_), .Y(new_n1221_));
  NAND2X1  g01029(.A(new_n1039_), .B(new_n1065_), .Y(new_n1222_));
  OAI21X1  g01030(.A0(new_n1222_), .A1(new_n1111_), .B0(new_n1038_), .Y(new_n1223_));
  AND2X1   g01031(.A(new_n1223_), .B(new_n1221_), .Y(new_n1224_));
  INVX1    g01032(.A(new_n1224_), .Y(new_n1225_));
  OAI21X1  g01033(.A0(new_n1218_), .A1(new_n1216_), .B0(\asqrt[59] ), .Y(new_n1226_));
  NAND2X1  g01034(.A(new_n1226_), .B(new_n292_), .Y(new_n1227_));
  OAI21X1  g01035(.A0(new_n1227_), .A1(new_n1220_), .B0(new_n1225_), .Y(new_n1228_));
  AOI21X1  g01036(.A0(new_n1228_), .A1(new_n1210_), .B0(new_n217_), .Y(new_n1229_));
  OAI21X1  g01037(.A0(new_n1219_), .A1(new_n1206_), .B0(new_n1226_), .Y(new_n1230_));
  AOI21X1  g01038(.A0(new_n1230_), .A1(\asqrt[60] ), .B0(\asqrt[61] ), .Y(new_n1231_));
  AND2X1   g01039(.A(new_n1091_), .B(new_n1090_), .Y(new_n1232_));
  NOR3X1   g01040(.A(new_n1049_), .B(new_n1232_), .C(new_n1089_), .Y(new_n1233_));
  NOR3X1   g01041(.A(new_n1111_), .B(new_n1232_), .C(new_n1089_), .Y(new_n1234_));
  NOR2X1   g01042(.A(new_n1234_), .B(new_n1048_), .Y(new_n1235_));
  AOI21X1  g01043(.A0(new_n1233_), .A1(\asqrt[52] ), .B0(new_n1235_), .Y(new_n1236_));
  AOI21X1  g01044(.A0(new_n1231_), .A1(new_n1228_), .B0(new_n1236_), .Y(new_n1237_));
  OAI21X1  g01045(.A0(new_n1237_), .A1(new_n1229_), .B0(\asqrt[62] ), .Y(new_n1238_));
  AND2X1   g01046(.A(new_n1069_), .B(new_n1050_), .Y(new_n1239_));
  NOR3X1   g01047(.A(new_n1239_), .B(new_n1094_), .C(new_n1051_), .Y(new_n1240_));
  NOR3X1   g01048(.A(new_n1111_), .B(new_n1239_), .C(new_n1051_), .Y(new_n1241_));
  NOR2X1   g01049(.A(new_n1241_), .B(new_n1056_), .Y(new_n1242_));
  AOI21X1  g01050(.A0(new_n1240_), .A1(\asqrt[52] ), .B0(new_n1242_), .Y(new_n1243_));
  NOR3X1   g01051(.A(new_n1237_), .B(new_n1229_), .C(\asqrt[62] ), .Y(new_n1244_));
  OAI21X1  g01052(.A0(new_n1244_), .A1(new_n1243_), .B0(new_n1238_), .Y(new_n1245_));
  NOR4X1   g01053(.A(new_n1111_), .B(new_n1076_), .C(new_n1074_), .D(new_n1116_), .Y(new_n1246_));
  NAND3X1  g01054(.A(\asqrt[52] ), .B(new_n1097_), .C(new_n1071_), .Y(new_n1247_));
  AOI21X1  g01055(.A0(new_n1247_), .A1(new_n1074_), .B0(new_n1246_), .Y(new_n1248_));
  INVX1    g01056(.A(new_n1248_), .Y(new_n1249_));
  AND2X1   g01057(.A(new_n1083_), .B(new_n1077_), .Y(new_n1250_));
  AOI21X1  g01058(.A0(new_n1250_), .A1(\asqrt[52] ), .B0(new_n1137_), .Y(new_n1251_));
  AND2X1   g01059(.A(new_n1251_), .B(new_n1249_), .Y(new_n1252_));
  AOI21X1  g01060(.A0(new_n1252_), .A1(new_n1245_), .B0(\asqrt[63] ), .Y(new_n1253_));
  INVX1    g01061(.A(new_n1243_), .Y(new_n1254_));
  AND2X1   g01062(.A(new_n1230_), .B(\asqrt[60] ), .Y(new_n1255_));
  OR2X1    g01063(.A(new_n1219_), .B(new_n1206_), .Y(new_n1256_));
  AND2X1   g01064(.A(new_n1226_), .B(new_n292_), .Y(new_n1257_));
  AOI21X1  g01065(.A0(new_n1257_), .A1(new_n1256_), .B0(new_n1224_), .Y(new_n1258_));
  OAI21X1  g01066(.A0(new_n1258_), .A1(new_n1255_), .B0(\asqrt[61] ), .Y(new_n1259_));
  OAI21X1  g01067(.A0(new_n1209_), .A1(new_n292_), .B0(new_n217_), .Y(new_n1260_));
  INVX1    g01068(.A(new_n1236_), .Y(new_n1261_));
  OAI21X1  g01069(.A0(new_n1260_), .A1(new_n1258_), .B0(new_n1261_), .Y(new_n1262_));
  NAND3X1  g01070(.A(new_n1262_), .B(new_n1259_), .C(new_n199_), .Y(new_n1263_));
  AND2X1   g01071(.A(new_n1263_), .B(new_n1254_), .Y(new_n1264_));
  AOI21X1  g01072(.A0(new_n1262_), .A1(new_n1259_), .B0(new_n199_), .Y(new_n1265_));
  OR2X1    g01073(.A(new_n1249_), .B(new_n1265_), .Y(new_n1266_));
  AOI21X1  g01074(.A0(new_n1123_), .A1(new_n1119_), .B0(new_n1082_), .Y(new_n1267_));
  AOI21X1  g01075(.A0(new_n1083_), .A1(new_n1077_), .B0(new_n193_), .Y(new_n1268_));
  OAI21X1  g01076(.A0(new_n1267_), .A1(new_n1077_), .B0(new_n1268_), .Y(new_n1269_));
  NOR4X1   g01077(.A(new_n1108_), .B(new_n1102_), .C(new_n1081_), .D(new_n1079_), .Y(new_n1270_));
  OAI21X1  g01078(.A0(new_n1099_), .A1(new_n1098_), .B0(new_n1270_), .Y(new_n1271_));
  NOR2X1   g01079(.A(new_n1271_), .B(new_n1088_), .Y(new_n1272_));
  INVX1    g01080(.A(new_n1272_), .Y(new_n1273_));
  AND2X1   g01081(.A(new_n1273_), .B(new_n1269_), .Y(new_n1274_));
  OAI21X1  g01082(.A0(new_n1266_), .A1(new_n1264_), .B0(new_n1274_), .Y(new_n1275_));
  OR2X1    g01083(.A(new_n1275_), .B(new_n1253_), .Y(\asqrt[51] ));
  NOR2X1   g01084(.A(new_n1275_), .B(new_n1253_), .Y(new_n1277_));
  NOR2X1   g01085(.A(\a[101] ), .B(\a[100] ), .Y(new_n1278_));
  INVX1    g01086(.A(new_n1278_), .Y(new_n1279_));
  MX2X1    g01087(.A(new_n1279_), .B(new_n1277_), .S0(\a[102] ), .Y(new_n1280_));
  OAI21X1  g01088(.A0(new_n1275_), .A1(new_n1253_), .B0(\a[102] ), .Y(new_n1281_));
  OAI22X1  g01089(.A0(new_n1279_), .A1(\a[102] ), .B0(new_n1107_), .B1(new_n1103_), .Y(new_n1282_));
  NOR4X1   g01090(.A(new_n1282_), .B(new_n1102_), .C(new_n1137_), .D(new_n1088_), .Y(new_n1283_));
  AND2X1   g01091(.A(new_n1283_), .B(new_n1281_), .Y(new_n1284_));
  INVX1    g01092(.A(\a[103] ), .Y(new_n1285_));
  AOI21X1  g01093(.A0(new_n1263_), .A1(new_n1254_), .B0(new_n1265_), .Y(new_n1286_));
  INVX1    g01094(.A(new_n1252_), .Y(new_n1287_));
  OAI21X1  g01095(.A0(new_n1287_), .A1(new_n1286_), .B0(new_n193_), .Y(new_n1288_));
  NAND2X1  g01096(.A(new_n1263_), .B(new_n1254_), .Y(new_n1289_));
  NOR2X1   g01097(.A(new_n1249_), .B(new_n1265_), .Y(new_n1290_));
  INVX1    g01098(.A(new_n1274_), .Y(new_n1291_));
  AOI21X1  g01099(.A0(new_n1290_), .A1(new_n1289_), .B0(new_n1291_), .Y(new_n1292_));
  AOI21X1  g01100(.A0(new_n1292_), .A1(new_n1288_), .B0(\a[102] ), .Y(new_n1293_));
  OAI21X1  g01101(.A0(new_n1275_), .A1(new_n1253_), .B0(new_n1113_), .Y(new_n1294_));
  OAI21X1  g01102(.A0(new_n1293_), .A1(new_n1285_), .B0(new_n1294_), .Y(new_n1295_));
  OAI22X1  g01103(.A0(new_n1295_), .A1(new_n1284_), .B0(new_n1280_), .B1(new_n1111_), .Y(new_n1296_));
  AND2X1   g01104(.A(new_n1296_), .B(\asqrt[53] ), .Y(new_n1297_));
  NAND2X1  g01105(.A(new_n1283_), .B(new_n1281_), .Y(new_n1298_));
  INVX1    g01106(.A(\a[102] ), .Y(new_n1299_));
  OAI21X1  g01107(.A0(new_n1275_), .A1(new_n1253_), .B0(new_n1299_), .Y(new_n1300_));
  AOI21X1  g01108(.A0(new_n1292_), .A1(new_n1288_), .B0(new_n1133_), .Y(new_n1301_));
  AOI21X1  g01109(.A0(new_n1300_), .A1(\a[103] ), .B0(new_n1301_), .Y(new_n1302_));
  NAND2X1  g01110(.A(new_n1302_), .B(new_n1298_), .Y(new_n1303_));
  MX2X1    g01111(.A(new_n1278_), .B(\asqrt[51] ), .S0(\a[102] ), .Y(new_n1304_));
  AOI21X1  g01112(.A0(new_n1304_), .A1(\asqrt[52] ), .B0(\asqrt[53] ), .Y(new_n1305_));
  INVX1    g01113(.A(new_n1269_), .Y(new_n1306_));
  NOR3X1   g01114(.A(new_n1272_), .B(new_n1306_), .C(new_n1111_), .Y(new_n1307_));
  OAI21X1  g01115(.A0(new_n1266_), .A1(new_n1264_), .B0(new_n1307_), .Y(new_n1308_));
  OR2X1    g01116(.A(new_n1308_), .B(new_n1253_), .Y(new_n1309_));
  AOI21X1  g01117(.A0(new_n1309_), .A1(new_n1294_), .B0(new_n1112_), .Y(new_n1310_));
  OAI21X1  g01118(.A0(new_n1308_), .A1(new_n1253_), .B0(new_n1112_), .Y(new_n1311_));
  NOR2X1   g01119(.A(new_n1311_), .B(new_n1301_), .Y(new_n1312_));
  NOR2X1   g01120(.A(new_n1312_), .B(new_n1310_), .Y(new_n1313_));
  AOI21X1  g01121(.A0(new_n1305_), .A1(new_n1303_), .B0(new_n1313_), .Y(new_n1314_));
  OAI21X1  g01122(.A0(new_n1314_), .A1(new_n1297_), .B0(\asqrt[54] ), .Y(new_n1315_));
  AOI21X1  g01123(.A0(new_n1115_), .A1(\asqrt[53] ), .B0(new_n1152_), .Y(new_n1316_));
  AND2X1   g01124(.A(new_n1316_), .B(new_n1155_), .Y(new_n1317_));
  OAI21X1  g01125(.A0(new_n1275_), .A1(new_n1253_), .B0(new_n1316_), .Y(new_n1318_));
  AOI22X1  g01126(.A0(new_n1318_), .A1(new_n1129_), .B0(new_n1317_), .B1(\asqrt[51] ), .Y(new_n1319_));
  INVX1    g01127(.A(new_n1319_), .Y(new_n1320_));
  AOI22X1  g01128(.A0(new_n1302_), .A1(new_n1298_), .B0(new_n1304_), .B1(\asqrt[52] ), .Y(new_n1321_));
  OAI21X1  g01129(.A0(new_n1321_), .A1(new_n968_), .B0(new_n902_), .Y(new_n1322_));
  OAI21X1  g01130(.A0(new_n1322_), .A1(new_n1314_), .B0(new_n1320_), .Y(new_n1323_));
  AOI21X1  g01131(.A0(new_n1323_), .A1(new_n1315_), .B0(new_n697_), .Y(new_n1324_));
  AOI21X1  g01132(.A0(new_n1178_), .A1(new_n1177_), .B0(new_n1143_), .Y(new_n1325_));
  AND2X1   g01133(.A(new_n1325_), .B(new_n1131_), .Y(new_n1326_));
  AOI22X1  g01134(.A0(new_n1178_), .A1(new_n1177_), .B0(new_n1156_), .B1(\asqrt[54] ), .Y(new_n1327_));
  OAI21X1  g01135(.A0(new_n1275_), .A1(new_n1253_), .B0(new_n1327_), .Y(new_n1328_));
  AOI22X1  g01136(.A0(new_n1328_), .A1(new_n1143_), .B0(new_n1326_), .B1(\asqrt[51] ), .Y(new_n1329_));
  INVX1    g01137(.A(new_n1329_), .Y(new_n1330_));
  NAND3X1  g01138(.A(new_n1323_), .B(new_n1315_), .C(new_n697_), .Y(new_n1331_));
  AOI21X1  g01139(.A0(new_n1331_), .A1(new_n1330_), .B0(new_n1324_), .Y(new_n1332_));
  OR2X1    g01140(.A(new_n1332_), .B(new_n582_), .Y(new_n1333_));
  OR2X1    g01141(.A(new_n1321_), .B(new_n968_), .Y(new_n1334_));
  AND2X1   g01142(.A(new_n1302_), .B(new_n1298_), .Y(new_n1335_));
  OAI21X1  g01143(.A0(new_n1280_), .A1(new_n1111_), .B0(new_n968_), .Y(new_n1336_));
  OR2X1    g01144(.A(new_n1312_), .B(new_n1310_), .Y(new_n1337_));
  OAI21X1  g01145(.A0(new_n1336_), .A1(new_n1335_), .B0(new_n1337_), .Y(new_n1338_));
  AOI21X1  g01146(.A0(new_n1338_), .A1(new_n1334_), .B0(new_n902_), .Y(new_n1339_));
  AOI21X1  g01147(.A0(new_n1296_), .A1(\asqrt[53] ), .B0(\asqrt[54] ), .Y(new_n1340_));
  AOI21X1  g01148(.A0(new_n1340_), .A1(new_n1338_), .B0(new_n1319_), .Y(new_n1341_));
  NOR3X1   g01149(.A(new_n1341_), .B(new_n1339_), .C(\asqrt[55] ), .Y(new_n1342_));
  NOR2X1   g01150(.A(new_n1342_), .B(new_n1329_), .Y(new_n1343_));
  AND2X1   g01151(.A(new_n1157_), .B(new_n1144_), .Y(new_n1344_));
  NOR3X1   g01152(.A(new_n1344_), .B(new_n1182_), .C(new_n1145_), .Y(new_n1345_));
  NOR2X1   g01153(.A(new_n1344_), .B(new_n1145_), .Y(new_n1346_));
  OAI21X1  g01154(.A0(new_n1275_), .A1(new_n1253_), .B0(new_n1346_), .Y(new_n1347_));
  AOI22X1  g01155(.A0(new_n1347_), .A1(new_n1182_), .B0(new_n1345_), .B1(\asqrt[51] ), .Y(new_n1348_));
  INVX1    g01156(.A(new_n1348_), .Y(new_n1349_));
  OAI21X1  g01157(.A0(new_n1341_), .A1(new_n1339_), .B0(\asqrt[55] ), .Y(new_n1350_));
  NAND2X1  g01158(.A(new_n1350_), .B(new_n582_), .Y(new_n1351_));
  OAI21X1  g01159(.A0(new_n1351_), .A1(new_n1343_), .B0(new_n1349_), .Y(new_n1352_));
  AOI21X1  g01160(.A0(new_n1352_), .A1(new_n1333_), .B0(new_n481_), .Y(new_n1353_));
  NAND4X1  g01161(.A(\asqrt[51] ), .B(new_n1197_), .C(new_n1166_), .D(new_n1159_), .Y(new_n1354_));
  NOR3X1   g01162(.A(new_n1277_), .B(new_n1167_), .C(new_n1185_), .Y(new_n1355_));
  OAI21X1  g01163(.A0(new_n1355_), .A1(new_n1166_), .B0(new_n1354_), .Y(new_n1356_));
  INVX1    g01164(.A(new_n1356_), .Y(new_n1357_));
  OAI21X1  g01165(.A0(new_n1342_), .A1(new_n1329_), .B0(new_n1350_), .Y(new_n1358_));
  AOI21X1  g01166(.A0(new_n1358_), .A1(\asqrt[56] ), .B0(\asqrt[57] ), .Y(new_n1359_));
  AOI21X1  g01167(.A0(new_n1359_), .A1(new_n1352_), .B0(new_n1357_), .Y(new_n1360_));
  OAI21X1  g01168(.A0(new_n1360_), .A1(new_n1353_), .B0(\asqrt[58] ), .Y(new_n1361_));
  AND2X1   g01169(.A(new_n1186_), .B(new_n1170_), .Y(new_n1362_));
  NOR3X1   g01170(.A(new_n1362_), .B(new_n1213_), .C(new_n1169_), .Y(new_n1363_));
  AOI22X1  g01171(.A0(new_n1186_), .A1(new_n1170_), .B0(new_n1168_), .B1(\asqrt[57] ), .Y(new_n1364_));
  AOI21X1  g01172(.A0(new_n1364_), .A1(\asqrt[51] ), .B0(new_n1175_), .Y(new_n1365_));
  AOI21X1  g01173(.A0(new_n1363_), .A1(\asqrt[51] ), .B0(new_n1365_), .Y(new_n1366_));
  NOR3X1   g01174(.A(new_n1360_), .B(new_n1353_), .C(\asqrt[58] ), .Y(new_n1367_));
  OAI21X1  g01175(.A0(new_n1367_), .A1(new_n1366_), .B0(new_n1361_), .Y(new_n1368_));
  AND2X1   g01176(.A(new_n1368_), .B(\asqrt[59] ), .Y(new_n1369_));
  INVX1    g01177(.A(new_n1366_), .Y(new_n1370_));
  AND2X1   g01178(.A(new_n1358_), .B(\asqrt[56] ), .Y(new_n1371_));
  OR2X1    g01179(.A(new_n1342_), .B(new_n1329_), .Y(new_n1372_));
  AND2X1   g01180(.A(new_n1350_), .B(new_n582_), .Y(new_n1373_));
  AOI21X1  g01181(.A0(new_n1373_), .A1(new_n1372_), .B0(new_n1348_), .Y(new_n1374_));
  OAI21X1  g01182(.A0(new_n1374_), .A1(new_n1371_), .B0(\asqrt[57] ), .Y(new_n1375_));
  OAI21X1  g01183(.A0(new_n1332_), .A1(new_n582_), .B0(new_n481_), .Y(new_n1376_));
  OAI21X1  g01184(.A0(new_n1376_), .A1(new_n1374_), .B0(new_n1356_), .Y(new_n1377_));
  NAND3X1  g01185(.A(new_n1377_), .B(new_n1375_), .C(new_n399_), .Y(new_n1378_));
  NAND2X1  g01186(.A(new_n1378_), .B(new_n1370_), .Y(new_n1379_));
  AND2X1   g01187(.A(new_n1217_), .B(new_n1215_), .Y(new_n1380_));
  NOR3X1   g01188(.A(new_n1380_), .B(new_n1195_), .C(new_n1216_), .Y(new_n1381_));
  NOR2X1   g01189(.A(new_n1380_), .B(new_n1216_), .Y(new_n1382_));
  AOI21X1  g01190(.A0(new_n1382_), .A1(\asqrt[51] ), .B0(new_n1194_), .Y(new_n1383_));
  AOI21X1  g01191(.A0(new_n1381_), .A1(\asqrt[51] ), .B0(new_n1383_), .Y(new_n1384_));
  AOI21X1  g01192(.A0(new_n1377_), .A1(new_n1375_), .B0(new_n399_), .Y(new_n1385_));
  NOR2X1   g01193(.A(new_n1385_), .B(\asqrt[59] ), .Y(new_n1386_));
  AOI21X1  g01194(.A0(new_n1386_), .A1(new_n1379_), .B0(new_n1384_), .Y(new_n1387_));
  OAI21X1  g01195(.A0(new_n1387_), .A1(new_n1369_), .B0(\asqrt[60] ), .Y(new_n1388_));
  OR4X1    g01196(.A(new_n1277_), .B(new_n1219_), .C(new_n1207_), .D(new_n1201_), .Y(new_n1389_));
  OR2X1    g01197(.A(new_n1219_), .B(new_n1201_), .Y(new_n1390_));
  OAI21X1  g01198(.A0(new_n1390_), .A1(new_n1277_), .B0(new_n1207_), .Y(new_n1391_));
  AND2X1   g01199(.A(new_n1391_), .B(new_n1389_), .Y(new_n1392_));
  INVX1    g01200(.A(new_n1392_), .Y(new_n1393_));
  AOI21X1  g01201(.A0(new_n1378_), .A1(new_n1370_), .B0(new_n1385_), .Y(new_n1394_));
  OAI21X1  g01202(.A0(new_n1394_), .A1(new_n328_), .B0(new_n292_), .Y(new_n1395_));
  OAI21X1  g01203(.A0(new_n1395_), .A1(new_n1387_), .B0(new_n1393_), .Y(new_n1396_));
  AOI21X1  g01204(.A0(new_n1396_), .A1(new_n1388_), .B0(new_n217_), .Y(new_n1397_));
  AOI21X1  g01205(.A0(new_n1257_), .A1(new_n1256_), .B0(new_n1225_), .Y(new_n1398_));
  AND2X1   g01206(.A(new_n1398_), .B(new_n1210_), .Y(new_n1399_));
  AOI22X1  g01207(.A0(new_n1257_), .A1(new_n1256_), .B0(new_n1230_), .B1(\asqrt[60] ), .Y(new_n1400_));
  AOI21X1  g01208(.A0(new_n1400_), .A1(\asqrt[51] ), .B0(new_n1224_), .Y(new_n1401_));
  AOI21X1  g01209(.A0(new_n1399_), .A1(\asqrt[51] ), .B0(new_n1401_), .Y(new_n1402_));
  INVX1    g01210(.A(new_n1402_), .Y(new_n1403_));
  NAND3X1  g01211(.A(new_n1396_), .B(new_n1388_), .C(new_n217_), .Y(new_n1404_));
  AOI21X1  g01212(.A0(new_n1404_), .A1(new_n1403_), .B0(new_n1397_), .Y(new_n1405_));
  OR2X1    g01213(.A(new_n1405_), .B(new_n199_), .Y(new_n1406_));
  AND2X1   g01214(.A(new_n1404_), .B(new_n1403_), .Y(new_n1407_));
  OR2X1    g01215(.A(new_n1397_), .B(\asqrt[62] ), .Y(new_n1408_));
  AND2X1   g01216(.A(new_n1231_), .B(new_n1228_), .Y(new_n1409_));
  NOR3X1   g01217(.A(new_n1261_), .B(new_n1409_), .C(new_n1229_), .Y(new_n1410_));
  NOR2X1   g01218(.A(new_n1409_), .B(new_n1229_), .Y(new_n1411_));
  AOI21X1  g01219(.A0(new_n1411_), .A1(\asqrt[51] ), .B0(new_n1236_), .Y(new_n1412_));
  AOI21X1  g01220(.A0(new_n1410_), .A1(\asqrt[51] ), .B0(new_n1412_), .Y(new_n1413_));
  INVX1    g01221(.A(new_n1413_), .Y(new_n1414_));
  OAI21X1  g01222(.A0(new_n1408_), .A1(new_n1407_), .B0(new_n1414_), .Y(new_n1415_));
  OR4X1    g01223(.A(new_n1277_), .B(new_n1244_), .C(new_n1254_), .D(new_n1265_), .Y(new_n1416_));
  OR2X1    g01224(.A(new_n1244_), .B(new_n1265_), .Y(new_n1417_));
  OAI21X1  g01225(.A0(new_n1417_), .A1(new_n1277_), .B0(new_n1254_), .Y(new_n1418_));
  AND2X1   g01226(.A(new_n1418_), .B(new_n1416_), .Y(new_n1419_));
  INVX1    g01227(.A(new_n1419_), .Y(new_n1420_));
  NOR2X1   g01228(.A(new_n1248_), .B(new_n1286_), .Y(new_n1421_));
  AOI22X1  g01229(.A0(new_n1421_), .A1(\asqrt[51] ), .B0(new_n1290_), .B1(new_n1289_), .Y(new_n1422_));
  AND2X1   g01230(.A(new_n1422_), .B(new_n1420_), .Y(new_n1423_));
  INVX1    g01231(.A(new_n1423_), .Y(new_n1424_));
  AOI21X1  g01232(.A0(new_n1415_), .A1(new_n1406_), .B0(new_n1424_), .Y(new_n1425_));
  OR2X1    g01233(.A(new_n1394_), .B(new_n328_), .Y(new_n1426_));
  AND2X1   g01234(.A(new_n1378_), .B(new_n1370_), .Y(new_n1427_));
  INVX1    g01235(.A(new_n1384_), .Y(new_n1428_));
  OR2X1    g01236(.A(new_n1385_), .B(\asqrt[59] ), .Y(new_n1429_));
  OAI21X1  g01237(.A0(new_n1429_), .A1(new_n1427_), .B0(new_n1428_), .Y(new_n1430_));
  AOI21X1  g01238(.A0(new_n1430_), .A1(new_n1426_), .B0(new_n292_), .Y(new_n1431_));
  AOI21X1  g01239(.A0(new_n1368_), .A1(\asqrt[59] ), .B0(\asqrt[60] ), .Y(new_n1432_));
  AOI21X1  g01240(.A0(new_n1432_), .A1(new_n1430_), .B0(new_n1392_), .Y(new_n1433_));
  OAI21X1  g01241(.A0(new_n1433_), .A1(new_n1431_), .B0(\asqrt[61] ), .Y(new_n1434_));
  NOR3X1   g01242(.A(new_n1433_), .B(new_n1431_), .C(\asqrt[61] ), .Y(new_n1435_));
  OAI21X1  g01243(.A0(new_n1435_), .A1(new_n1402_), .B0(new_n1434_), .Y(new_n1436_));
  AOI21X1  g01244(.A0(new_n1436_), .A1(\asqrt[62] ), .B0(new_n1420_), .Y(new_n1437_));
  AOI21X1  g01245(.A0(new_n1292_), .A1(new_n1288_), .B0(new_n1248_), .Y(new_n1438_));
  AOI21X1  g01246(.A0(new_n1249_), .A1(new_n1245_), .B0(new_n193_), .Y(new_n1439_));
  OAI21X1  g01247(.A0(new_n1438_), .A1(new_n1245_), .B0(new_n1439_), .Y(new_n1440_));
  OR2X1    g01248(.A(new_n1266_), .B(new_n1264_), .Y(new_n1441_));
  AND2X1   g01249(.A(new_n1247_), .B(new_n1074_), .Y(new_n1442_));
  NOR4X1   g01250(.A(new_n1272_), .B(new_n1306_), .C(new_n1442_), .D(new_n1246_), .Y(new_n1443_));
  NAND3X1  g01251(.A(new_n1443_), .B(new_n1441_), .C(new_n1288_), .Y(new_n1444_));
  AND2X1   g01252(.A(new_n1444_), .B(new_n1440_), .Y(new_n1445_));
  INVX1    g01253(.A(new_n1445_), .Y(new_n1446_));
  AOI21X1  g01254(.A0(new_n1437_), .A1(new_n1415_), .B0(new_n1446_), .Y(new_n1447_));
  OAI21X1  g01255(.A0(new_n1425_), .A1(\asqrt[63] ), .B0(new_n1447_), .Y(\asqrt[50] ));
  NOR2X1   g01256(.A(\a[99] ), .B(\a[98] ), .Y(new_n1449_));
  MX2X1    g01257(.A(new_n1449_), .B(\asqrt[50] ), .S0(\a[100] ), .Y(new_n1450_));
  AND2X1   g01258(.A(new_n1450_), .B(\asqrt[51] ), .Y(new_n1451_));
  NOR3X1   g01259(.A(\a[100] ), .B(\a[99] ), .C(\a[98] ), .Y(new_n1452_));
  NOR3X1   g01260(.A(new_n1452_), .B(new_n1272_), .C(new_n1306_), .Y(new_n1453_));
  NAND3X1  g01261(.A(new_n1453_), .B(new_n1441_), .C(new_n1288_), .Y(new_n1454_));
  AOI21X1  g01262(.A0(\asqrt[50] ), .A1(\a[100] ), .B0(new_n1454_), .Y(new_n1455_));
  INVX1    g01263(.A(\a[100] ), .Y(new_n1456_));
  INVX1    g01264(.A(\a[101] ), .Y(new_n1457_));
  AOI21X1  g01265(.A0(\asqrt[50] ), .A1(new_n1456_), .B0(new_n1457_), .Y(new_n1458_));
  AND2X1   g01266(.A(\asqrt[50] ), .B(new_n1278_), .Y(new_n1459_));
  NOR3X1   g01267(.A(new_n1459_), .B(new_n1458_), .C(new_n1455_), .Y(new_n1460_));
  OAI21X1  g01268(.A0(new_n1460_), .A1(new_n1451_), .B0(\asqrt[52] ), .Y(new_n1461_));
  AND2X1   g01269(.A(new_n1436_), .B(\asqrt[62] ), .Y(new_n1462_));
  NAND2X1  g01270(.A(new_n1404_), .B(new_n1403_), .Y(new_n1463_));
  NOR2X1   g01271(.A(new_n1397_), .B(\asqrt[62] ), .Y(new_n1464_));
  AOI21X1  g01272(.A0(new_n1464_), .A1(new_n1463_), .B0(new_n1413_), .Y(new_n1465_));
  OAI21X1  g01273(.A0(new_n1465_), .A1(new_n1462_), .B0(new_n1423_), .Y(new_n1466_));
  OAI21X1  g01274(.A0(new_n1405_), .A1(new_n199_), .B0(new_n1419_), .Y(new_n1467_));
  OAI21X1  g01275(.A0(new_n1467_), .A1(new_n1465_), .B0(new_n1445_), .Y(new_n1468_));
  AOI21X1  g01276(.A0(new_n1466_), .A1(new_n193_), .B0(new_n1468_), .Y(new_n1469_));
  INVX1    g01277(.A(new_n1449_), .Y(new_n1470_));
  MX2X1    g01278(.A(new_n1470_), .B(new_n1469_), .S0(\a[100] ), .Y(new_n1471_));
  OAI21X1  g01279(.A0(new_n1471_), .A1(new_n1277_), .B0(new_n1111_), .Y(new_n1472_));
  NAND3X1  g01280(.A(new_n1444_), .B(new_n1440_), .C(\asqrt[51] ), .Y(new_n1473_));
  INVX1    g01281(.A(new_n1473_), .Y(new_n1474_));
  OAI21X1  g01282(.A0(new_n1467_), .A1(new_n1465_), .B0(new_n1474_), .Y(new_n1475_));
  AOI21X1  g01283(.A0(new_n1466_), .A1(new_n193_), .B0(new_n1475_), .Y(new_n1476_));
  AOI21X1  g01284(.A0(\asqrt[50] ), .A1(new_n1278_), .B0(new_n1476_), .Y(new_n1477_));
  OR2X1    g01285(.A(new_n1476_), .B(\a[102] ), .Y(new_n1478_));
  OAI22X1  g01286(.A0(new_n1478_), .A1(new_n1459_), .B0(new_n1477_), .B1(new_n1299_), .Y(new_n1479_));
  OAI21X1  g01287(.A0(new_n1472_), .A1(new_n1460_), .B0(new_n1479_), .Y(new_n1480_));
  AOI21X1  g01288(.A0(new_n1480_), .A1(new_n1461_), .B0(new_n968_), .Y(new_n1481_));
  AOI21X1  g01289(.A0(new_n1304_), .A1(\asqrt[52] ), .B0(new_n1284_), .Y(new_n1482_));
  NAND3X1  g01290(.A(new_n1482_), .B(\asqrt[50] ), .C(new_n1295_), .Y(new_n1483_));
  INVX1    g01291(.A(new_n1482_), .Y(new_n1484_));
  OAI21X1  g01292(.A0(new_n1484_), .A1(new_n1469_), .B0(new_n1302_), .Y(new_n1485_));
  AND2X1   g01293(.A(new_n1485_), .B(new_n1483_), .Y(new_n1486_));
  INVX1    g01294(.A(new_n1486_), .Y(new_n1487_));
  NAND3X1  g01295(.A(new_n1480_), .B(new_n1461_), .C(new_n968_), .Y(new_n1488_));
  AOI21X1  g01296(.A0(new_n1488_), .A1(new_n1487_), .B0(new_n1481_), .Y(new_n1489_));
  OR2X1    g01297(.A(new_n1489_), .B(new_n902_), .Y(new_n1490_));
  AND2X1   g01298(.A(new_n1488_), .B(new_n1487_), .Y(new_n1491_));
  OAI21X1  g01299(.A0(new_n1336_), .A1(new_n1335_), .B0(new_n1313_), .Y(new_n1492_));
  NOR3X1   g01300(.A(new_n1492_), .B(new_n1469_), .C(new_n1297_), .Y(new_n1493_));
  OAI22X1  g01301(.A0(new_n1336_), .A1(new_n1335_), .B0(new_n1321_), .B1(new_n968_), .Y(new_n1494_));
  OR2X1    g01302(.A(new_n1494_), .B(new_n1469_), .Y(new_n1495_));
  AOI21X1  g01303(.A0(new_n1495_), .A1(new_n1337_), .B0(new_n1493_), .Y(new_n1496_));
  INVX1    g01304(.A(new_n1496_), .Y(new_n1497_));
  OR2X1    g01305(.A(new_n1481_), .B(\asqrt[54] ), .Y(new_n1498_));
  OAI21X1  g01306(.A0(new_n1498_), .A1(new_n1491_), .B0(new_n1497_), .Y(new_n1499_));
  AOI21X1  g01307(.A0(new_n1499_), .A1(new_n1490_), .B0(new_n697_), .Y(new_n1500_));
  AND2X1   g01308(.A(new_n1340_), .B(new_n1338_), .Y(new_n1501_));
  NOR4X1   g01309(.A(new_n1469_), .B(new_n1501_), .C(new_n1320_), .D(new_n1339_), .Y(new_n1502_));
  OR2X1    g01310(.A(new_n1501_), .B(new_n1339_), .Y(new_n1503_));
  OR2X1    g01311(.A(new_n1503_), .B(new_n1469_), .Y(new_n1504_));
  AOI21X1  g01312(.A0(new_n1504_), .A1(new_n1320_), .B0(new_n1502_), .Y(new_n1505_));
  OR2X1    g01313(.A(new_n1471_), .B(new_n1277_), .Y(new_n1506_));
  INVX1    g01314(.A(new_n1454_), .Y(new_n1507_));
  OAI21X1  g01315(.A0(new_n1469_), .A1(new_n1456_), .B0(new_n1507_), .Y(new_n1508_));
  OAI21X1  g01316(.A0(new_n1469_), .A1(\a[100] ), .B0(\a[101] ), .Y(new_n1509_));
  OR2X1    g01317(.A(new_n1469_), .B(new_n1279_), .Y(new_n1510_));
  NAND3X1  g01318(.A(new_n1510_), .B(new_n1509_), .C(new_n1508_), .Y(new_n1511_));
  AOI21X1  g01319(.A0(new_n1511_), .A1(new_n1506_), .B0(new_n1111_), .Y(new_n1512_));
  AOI21X1  g01320(.A0(new_n1450_), .A1(\asqrt[51] ), .B0(\asqrt[52] ), .Y(new_n1513_));
  OR2X1    g01321(.A(new_n1477_), .B(new_n1299_), .Y(new_n1514_));
  OR2X1    g01322(.A(new_n1478_), .B(new_n1459_), .Y(new_n1515_));
  AOI22X1  g01323(.A0(new_n1515_), .A1(new_n1514_), .B0(new_n1513_), .B1(new_n1511_), .Y(new_n1516_));
  OAI21X1  g01324(.A0(new_n1516_), .A1(new_n1512_), .B0(\asqrt[53] ), .Y(new_n1517_));
  NOR3X1   g01325(.A(new_n1516_), .B(new_n1512_), .C(\asqrt[53] ), .Y(new_n1518_));
  OAI21X1  g01326(.A0(new_n1518_), .A1(new_n1486_), .B0(new_n1517_), .Y(new_n1519_));
  AOI21X1  g01327(.A0(new_n1519_), .A1(\asqrt[54] ), .B0(\asqrt[55] ), .Y(new_n1520_));
  AOI21X1  g01328(.A0(new_n1520_), .A1(new_n1499_), .B0(new_n1505_), .Y(new_n1521_));
  OAI21X1  g01329(.A0(new_n1521_), .A1(new_n1500_), .B0(\asqrt[56] ), .Y(new_n1522_));
  NOR3X1   g01330(.A(new_n1342_), .B(new_n1330_), .C(new_n1324_), .Y(new_n1523_));
  NOR2X1   g01331(.A(new_n1342_), .B(new_n1324_), .Y(new_n1524_));
  AOI21X1  g01332(.A0(new_n1524_), .A1(\asqrt[50] ), .B0(new_n1329_), .Y(new_n1525_));
  AOI21X1  g01333(.A0(new_n1523_), .A1(\asqrt[50] ), .B0(new_n1525_), .Y(new_n1526_));
  NOR3X1   g01334(.A(new_n1521_), .B(new_n1500_), .C(\asqrt[56] ), .Y(new_n1527_));
  OAI21X1  g01335(.A0(new_n1527_), .A1(new_n1526_), .B0(new_n1522_), .Y(new_n1528_));
  AND2X1   g01336(.A(new_n1528_), .B(\asqrt[57] ), .Y(new_n1529_));
  INVX1    g01337(.A(new_n1526_), .Y(new_n1530_));
  AND2X1   g01338(.A(new_n1519_), .B(\asqrt[54] ), .Y(new_n1531_));
  NAND2X1  g01339(.A(new_n1488_), .B(new_n1487_), .Y(new_n1532_));
  NOR2X1   g01340(.A(new_n1481_), .B(\asqrt[54] ), .Y(new_n1533_));
  AOI21X1  g01341(.A0(new_n1533_), .A1(new_n1532_), .B0(new_n1496_), .Y(new_n1534_));
  OAI21X1  g01342(.A0(new_n1534_), .A1(new_n1531_), .B0(\asqrt[55] ), .Y(new_n1535_));
  INVX1    g01343(.A(new_n1505_), .Y(new_n1536_));
  OAI21X1  g01344(.A0(new_n1489_), .A1(new_n902_), .B0(new_n697_), .Y(new_n1537_));
  OAI21X1  g01345(.A0(new_n1537_), .A1(new_n1534_), .B0(new_n1536_), .Y(new_n1538_));
  NAND3X1  g01346(.A(new_n1538_), .B(new_n1535_), .C(new_n582_), .Y(new_n1539_));
  NAND2X1  g01347(.A(new_n1539_), .B(new_n1530_), .Y(new_n1540_));
  AND2X1   g01348(.A(new_n1373_), .B(new_n1372_), .Y(new_n1541_));
  NOR4X1   g01349(.A(new_n1469_), .B(new_n1541_), .C(new_n1349_), .D(new_n1371_), .Y(new_n1542_));
  AOI22X1  g01350(.A0(new_n1373_), .A1(new_n1372_), .B0(new_n1358_), .B1(\asqrt[56] ), .Y(new_n1543_));
  AOI21X1  g01351(.A0(new_n1543_), .A1(\asqrt[50] ), .B0(new_n1348_), .Y(new_n1544_));
  NOR2X1   g01352(.A(new_n1544_), .B(new_n1542_), .Y(new_n1545_));
  AOI21X1  g01353(.A0(new_n1538_), .A1(new_n1535_), .B0(new_n582_), .Y(new_n1546_));
  NOR2X1   g01354(.A(new_n1546_), .B(\asqrt[57] ), .Y(new_n1547_));
  AOI21X1  g01355(.A0(new_n1547_), .A1(new_n1540_), .B0(new_n1545_), .Y(new_n1548_));
  OAI21X1  g01356(.A0(new_n1548_), .A1(new_n1529_), .B0(\asqrt[58] ), .Y(new_n1549_));
  AND2X1   g01357(.A(new_n1359_), .B(new_n1352_), .Y(new_n1550_));
  NOR4X1   g01358(.A(new_n1469_), .B(new_n1550_), .C(new_n1356_), .D(new_n1353_), .Y(new_n1551_));
  NOR2X1   g01359(.A(new_n1550_), .B(new_n1353_), .Y(new_n1552_));
  AOI21X1  g01360(.A0(new_n1552_), .A1(\asqrt[50] ), .B0(new_n1357_), .Y(new_n1553_));
  NOR2X1   g01361(.A(new_n1553_), .B(new_n1551_), .Y(new_n1554_));
  INVX1    g01362(.A(new_n1554_), .Y(new_n1555_));
  AOI21X1  g01363(.A0(new_n1539_), .A1(new_n1530_), .B0(new_n1546_), .Y(new_n1556_));
  OAI21X1  g01364(.A0(new_n1556_), .A1(new_n481_), .B0(new_n399_), .Y(new_n1557_));
  OAI21X1  g01365(.A0(new_n1557_), .A1(new_n1548_), .B0(new_n1555_), .Y(new_n1558_));
  AOI21X1  g01366(.A0(new_n1558_), .A1(new_n1549_), .B0(new_n328_), .Y(new_n1559_));
  NAND3X1  g01367(.A(new_n1378_), .B(new_n1366_), .C(new_n1361_), .Y(new_n1560_));
  NOR3X1   g01368(.A(new_n1469_), .B(new_n1367_), .C(new_n1385_), .Y(new_n1561_));
  OAI22X1  g01369(.A0(new_n1561_), .A1(new_n1366_), .B0(new_n1560_), .B1(new_n1469_), .Y(new_n1562_));
  NAND3X1  g01370(.A(new_n1558_), .B(new_n1549_), .C(new_n328_), .Y(new_n1563_));
  AOI21X1  g01371(.A0(new_n1563_), .A1(new_n1562_), .B0(new_n1559_), .Y(new_n1564_));
  OR2X1    g01372(.A(new_n1564_), .B(new_n292_), .Y(new_n1565_));
  AND2X1   g01373(.A(new_n1563_), .B(new_n1562_), .Y(new_n1566_));
  OAI21X1  g01374(.A0(new_n1429_), .A1(new_n1427_), .B0(new_n1384_), .Y(new_n1567_));
  NOR3X1   g01375(.A(new_n1567_), .B(new_n1469_), .C(new_n1369_), .Y(new_n1568_));
  AOI22X1  g01376(.A0(new_n1386_), .A1(new_n1379_), .B0(new_n1368_), .B1(\asqrt[59] ), .Y(new_n1569_));
  AOI21X1  g01377(.A0(new_n1569_), .A1(\asqrt[50] ), .B0(new_n1384_), .Y(new_n1570_));
  NOR2X1   g01378(.A(new_n1570_), .B(new_n1568_), .Y(new_n1571_));
  INVX1    g01379(.A(new_n1571_), .Y(new_n1572_));
  OR2X1    g01380(.A(new_n1556_), .B(new_n481_), .Y(new_n1573_));
  AND2X1   g01381(.A(new_n1539_), .B(new_n1530_), .Y(new_n1574_));
  INVX1    g01382(.A(new_n1545_), .Y(new_n1575_));
  OR2X1    g01383(.A(new_n1546_), .B(\asqrt[57] ), .Y(new_n1576_));
  OAI21X1  g01384(.A0(new_n1576_), .A1(new_n1574_), .B0(new_n1575_), .Y(new_n1577_));
  AOI21X1  g01385(.A0(new_n1577_), .A1(new_n1573_), .B0(new_n399_), .Y(new_n1578_));
  AOI21X1  g01386(.A0(new_n1528_), .A1(\asqrt[57] ), .B0(\asqrt[58] ), .Y(new_n1579_));
  AOI21X1  g01387(.A0(new_n1579_), .A1(new_n1577_), .B0(new_n1554_), .Y(new_n1580_));
  OAI21X1  g01388(.A0(new_n1580_), .A1(new_n1578_), .B0(\asqrt[59] ), .Y(new_n1581_));
  NAND2X1  g01389(.A(new_n1581_), .B(new_n292_), .Y(new_n1582_));
  OAI21X1  g01390(.A0(new_n1582_), .A1(new_n1566_), .B0(new_n1572_), .Y(new_n1583_));
  AOI21X1  g01391(.A0(new_n1583_), .A1(new_n1565_), .B0(new_n217_), .Y(new_n1584_));
  AND2X1   g01392(.A(new_n1432_), .B(new_n1430_), .Y(new_n1585_));
  NOR4X1   g01393(.A(new_n1469_), .B(new_n1585_), .C(new_n1393_), .D(new_n1431_), .Y(new_n1586_));
  NOR2X1   g01394(.A(new_n1585_), .B(new_n1431_), .Y(new_n1587_));
  AOI21X1  g01395(.A0(new_n1587_), .A1(\asqrt[50] ), .B0(new_n1392_), .Y(new_n1588_));
  NOR2X1   g01396(.A(new_n1588_), .B(new_n1586_), .Y(new_n1589_));
  INVX1    g01397(.A(new_n1562_), .Y(new_n1590_));
  NOR3X1   g01398(.A(new_n1580_), .B(new_n1578_), .C(\asqrt[59] ), .Y(new_n1591_));
  OAI21X1  g01399(.A0(new_n1591_), .A1(new_n1590_), .B0(new_n1581_), .Y(new_n1592_));
  AOI21X1  g01400(.A0(new_n1592_), .A1(\asqrt[60] ), .B0(\asqrt[61] ), .Y(new_n1593_));
  AOI21X1  g01401(.A0(new_n1593_), .A1(new_n1583_), .B0(new_n1589_), .Y(new_n1594_));
  OAI21X1  g01402(.A0(new_n1594_), .A1(new_n1584_), .B0(\asqrt[62] ), .Y(new_n1595_));
  NAND3X1  g01403(.A(new_n1404_), .B(new_n1402_), .C(new_n1434_), .Y(new_n1596_));
  NOR3X1   g01404(.A(new_n1469_), .B(new_n1435_), .C(new_n1397_), .Y(new_n1597_));
  OAI22X1  g01405(.A0(new_n1597_), .A1(new_n1402_), .B0(new_n1596_), .B1(new_n1469_), .Y(new_n1598_));
  INVX1    g01406(.A(new_n1598_), .Y(new_n1599_));
  NOR3X1   g01407(.A(new_n1594_), .B(new_n1584_), .C(\asqrt[62] ), .Y(new_n1600_));
  OAI21X1  g01408(.A0(new_n1600_), .A1(new_n1599_), .B0(new_n1595_), .Y(new_n1601_));
  AND2X1   g01409(.A(new_n1464_), .B(new_n1463_), .Y(new_n1602_));
  NOR4X1   g01410(.A(new_n1469_), .B(new_n1414_), .C(new_n1602_), .D(new_n1462_), .Y(new_n1603_));
  AOI22X1  g01411(.A0(new_n1464_), .A1(new_n1463_), .B0(new_n1436_), .B1(\asqrt[62] ), .Y(new_n1604_));
  AOI21X1  g01412(.A0(new_n1604_), .A1(\asqrt[50] ), .B0(new_n1413_), .Y(new_n1605_));
  NOR2X1   g01413(.A(new_n1605_), .B(new_n1603_), .Y(new_n1606_));
  INVX1    g01414(.A(new_n1606_), .Y(new_n1607_));
  AND2X1   g01415(.A(new_n1437_), .B(new_n1415_), .Y(new_n1608_));
  AOI21X1  g01416(.A0(new_n1415_), .A1(new_n1406_), .B0(new_n1419_), .Y(new_n1609_));
  AOI21X1  g01417(.A0(new_n1609_), .A1(\asqrt[50] ), .B0(new_n1608_), .Y(new_n1610_));
  AND2X1   g01418(.A(new_n1610_), .B(new_n1607_), .Y(new_n1611_));
  AOI21X1  g01419(.A0(new_n1611_), .A1(new_n1601_), .B0(\asqrt[63] ), .Y(new_n1612_));
  AND2X1   g01420(.A(new_n1592_), .B(\asqrt[60] ), .Y(new_n1613_));
  NAND2X1  g01421(.A(new_n1563_), .B(new_n1562_), .Y(new_n1614_));
  AND2X1   g01422(.A(new_n1581_), .B(new_n292_), .Y(new_n1615_));
  AOI21X1  g01423(.A0(new_n1615_), .A1(new_n1614_), .B0(new_n1571_), .Y(new_n1616_));
  OAI21X1  g01424(.A0(new_n1616_), .A1(new_n1613_), .B0(\asqrt[61] ), .Y(new_n1617_));
  INVX1    g01425(.A(new_n1589_), .Y(new_n1618_));
  OAI21X1  g01426(.A0(new_n1564_), .A1(new_n292_), .B0(new_n217_), .Y(new_n1619_));
  OAI21X1  g01427(.A0(new_n1619_), .A1(new_n1616_), .B0(new_n1618_), .Y(new_n1620_));
  NAND3X1  g01428(.A(new_n1620_), .B(new_n1617_), .C(new_n199_), .Y(new_n1621_));
  AND2X1   g01429(.A(new_n1621_), .B(new_n1598_), .Y(new_n1622_));
  NAND2X1  g01430(.A(new_n1606_), .B(new_n1595_), .Y(new_n1623_));
  NAND2X1  g01431(.A(new_n1415_), .B(new_n1406_), .Y(new_n1624_));
  AOI21X1  g01432(.A0(\asqrt[50] ), .A1(new_n1420_), .B0(new_n1624_), .Y(new_n1625_));
  NOR3X1   g01433(.A(new_n1625_), .B(new_n1609_), .C(new_n193_), .Y(new_n1626_));
  AND2X1   g01434(.A(new_n1466_), .B(new_n193_), .Y(new_n1627_));
  NAND4X1  g01435(.A(new_n1444_), .B(new_n1440_), .C(new_n1418_), .D(new_n1416_), .Y(new_n1628_));
  NOR3X1   g01436(.A(new_n1628_), .B(new_n1608_), .C(new_n1627_), .Y(new_n1629_));
  NOR2X1   g01437(.A(new_n1629_), .B(new_n1626_), .Y(new_n1630_));
  OAI21X1  g01438(.A0(new_n1623_), .A1(new_n1622_), .B0(new_n1630_), .Y(new_n1631_));
  NOR2X1   g01439(.A(new_n1631_), .B(new_n1612_), .Y(new_n1632_));
  NOR2X1   g01440(.A(\a[97] ), .B(\a[96] ), .Y(new_n1633_));
  INVX1    g01441(.A(new_n1633_), .Y(new_n1634_));
  MX2X1    g01442(.A(new_n1634_), .B(new_n1632_), .S0(\a[98] ), .Y(new_n1635_));
  INVX1    g01443(.A(\a[98] ), .Y(new_n1636_));
  AOI21X1  g01444(.A0(new_n1620_), .A1(new_n1617_), .B0(new_n199_), .Y(new_n1637_));
  AOI21X1  g01445(.A0(new_n1621_), .A1(new_n1598_), .B0(new_n1637_), .Y(new_n1638_));
  INVX1    g01446(.A(new_n1611_), .Y(new_n1639_));
  OAI21X1  g01447(.A0(new_n1639_), .A1(new_n1638_), .B0(new_n193_), .Y(new_n1640_));
  NAND2X1  g01448(.A(new_n1621_), .B(new_n1598_), .Y(new_n1641_));
  AND2X1   g01449(.A(new_n1606_), .B(new_n1595_), .Y(new_n1642_));
  INVX1    g01450(.A(new_n1630_), .Y(new_n1643_));
  AOI21X1  g01451(.A0(new_n1642_), .A1(new_n1641_), .B0(new_n1643_), .Y(new_n1644_));
  AOI21X1  g01452(.A0(new_n1644_), .A1(new_n1640_), .B0(new_n1636_), .Y(new_n1645_));
  NAND2X1  g01453(.A(new_n1633_), .B(new_n1636_), .Y(new_n1646_));
  NAND3X1  g01454(.A(new_n1646_), .B(new_n1444_), .C(new_n1440_), .Y(new_n1647_));
  NOR4X1   g01455(.A(new_n1647_), .B(new_n1645_), .C(new_n1608_), .D(new_n1627_), .Y(new_n1648_));
  INVX1    g01456(.A(\a[99] ), .Y(new_n1649_));
  AOI21X1  g01457(.A0(new_n1644_), .A1(new_n1640_), .B0(\a[98] ), .Y(new_n1650_));
  OAI21X1  g01458(.A0(new_n1631_), .A1(new_n1612_), .B0(new_n1449_), .Y(new_n1651_));
  OAI21X1  g01459(.A0(new_n1650_), .A1(new_n1649_), .B0(new_n1651_), .Y(new_n1652_));
  OAI22X1  g01460(.A0(new_n1652_), .A1(new_n1648_), .B0(new_n1635_), .B1(new_n1469_), .Y(new_n1653_));
  AND2X1   g01461(.A(new_n1653_), .B(\asqrt[51] ), .Y(new_n1654_));
  OR4X1    g01462(.A(new_n1647_), .B(new_n1645_), .C(new_n1608_), .D(new_n1627_), .Y(new_n1655_));
  OAI21X1  g01463(.A0(new_n1631_), .A1(new_n1612_), .B0(new_n1636_), .Y(new_n1656_));
  AOI21X1  g01464(.A0(new_n1644_), .A1(new_n1640_), .B0(new_n1470_), .Y(new_n1657_));
  AOI21X1  g01465(.A0(new_n1656_), .A1(\a[99] ), .B0(new_n1657_), .Y(new_n1658_));
  NAND2X1  g01466(.A(new_n1658_), .B(new_n1655_), .Y(new_n1659_));
  OAI21X1  g01467(.A0(new_n1632_), .A1(new_n1636_), .B0(new_n1646_), .Y(new_n1660_));
  AOI21X1  g01468(.A0(new_n1660_), .A1(\asqrt[50] ), .B0(\asqrt[51] ), .Y(new_n1661_));
  AND2X1   g01469(.A(new_n1642_), .B(new_n1641_), .Y(new_n1662_));
  OR2X1    g01470(.A(new_n1629_), .B(new_n1469_), .Y(new_n1663_));
  OR4X1    g01471(.A(new_n1663_), .B(new_n1626_), .C(new_n1662_), .D(new_n1612_), .Y(new_n1664_));
  AOI21X1  g01472(.A0(new_n1664_), .A1(new_n1651_), .B0(new_n1456_), .Y(new_n1665_));
  NOR4X1   g01473(.A(new_n1663_), .B(new_n1626_), .C(new_n1662_), .D(new_n1612_), .Y(new_n1666_));
  NOR3X1   g01474(.A(new_n1666_), .B(new_n1657_), .C(\a[100] ), .Y(new_n1667_));
  NOR2X1   g01475(.A(new_n1667_), .B(new_n1665_), .Y(new_n1668_));
  AOI21X1  g01476(.A0(new_n1661_), .A1(new_n1659_), .B0(new_n1668_), .Y(new_n1669_));
  OAI21X1  g01477(.A0(new_n1669_), .A1(new_n1654_), .B0(\asqrt[52] ), .Y(new_n1670_));
  AND2X1   g01478(.A(new_n1510_), .B(new_n1509_), .Y(new_n1671_));
  NOR3X1   g01479(.A(new_n1671_), .B(new_n1455_), .C(new_n1451_), .Y(new_n1672_));
  OAI21X1  g01480(.A0(new_n1631_), .A1(new_n1612_), .B0(new_n1672_), .Y(new_n1673_));
  AOI21X1  g01481(.A0(new_n1450_), .A1(\asqrt[51] ), .B0(new_n1455_), .Y(new_n1674_));
  OAI21X1  g01482(.A0(new_n1631_), .A1(new_n1612_), .B0(new_n1674_), .Y(new_n1675_));
  NAND2X1  g01483(.A(new_n1675_), .B(new_n1671_), .Y(new_n1676_));
  NAND2X1  g01484(.A(new_n1676_), .B(new_n1673_), .Y(new_n1677_));
  AOI22X1  g01485(.A0(new_n1658_), .A1(new_n1655_), .B0(new_n1660_), .B1(\asqrt[50] ), .Y(new_n1678_));
  OAI21X1  g01486(.A0(new_n1678_), .A1(new_n1277_), .B0(new_n1111_), .Y(new_n1679_));
  OAI21X1  g01487(.A0(new_n1679_), .A1(new_n1669_), .B0(new_n1677_), .Y(new_n1680_));
  AOI21X1  g01488(.A0(new_n1680_), .A1(new_n1670_), .B0(new_n968_), .Y(new_n1681_));
  AND2X1   g01489(.A(new_n1513_), .B(new_n1511_), .Y(new_n1682_));
  NOR3X1   g01490(.A(new_n1479_), .B(new_n1682_), .C(new_n1512_), .Y(new_n1683_));
  OAI21X1  g01491(.A0(new_n1631_), .A1(new_n1612_), .B0(new_n1683_), .Y(new_n1684_));
  NOR2X1   g01492(.A(new_n1682_), .B(new_n1512_), .Y(new_n1685_));
  OAI21X1  g01493(.A0(new_n1631_), .A1(new_n1612_), .B0(new_n1685_), .Y(new_n1686_));
  NAND2X1  g01494(.A(new_n1686_), .B(new_n1479_), .Y(new_n1687_));
  AND2X1   g01495(.A(new_n1687_), .B(new_n1684_), .Y(new_n1688_));
  INVX1    g01496(.A(new_n1688_), .Y(new_n1689_));
  NAND3X1  g01497(.A(new_n1680_), .B(new_n1670_), .C(new_n968_), .Y(new_n1690_));
  AOI21X1  g01498(.A0(new_n1690_), .A1(new_n1689_), .B0(new_n1681_), .Y(new_n1691_));
  OR2X1    g01499(.A(new_n1691_), .B(new_n902_), .Y(new_n1692_));
  OR2X1    g01500(.A(new_n1678_), .B(new_n1277_), .Y(new_n1693_));
  AND2X1   g01501(.A(new_n1658_), .B(new_n1655_), .Y(new_n1694_));
  OAI21X1  g01502(.A0(new_n1635_), .A1(new_n1469_), .B0(new_n1277_), .Y(new_n1695_));
  OR2X1    g01503(.A(new_n1667_), .B(new_n1665_), .Y(new_n1696_));
  OAI21X1  g01504(.A0(new_n1695_), .A1(new_n1694_), .B0(new_n1696_), .Y(new_n1697_));
  AOI21X1  g01505(.A0(new_n1697_), .A1(new_n1693_), .B0(new_n1111_), .Y(new_n1698_));
  AOI21X1  g01506(.A0(new_n1653_), .A1(\asqrt[51] ), .B0(\asqrt[52] ), .Y(new_n1699_));
  AOI22X1  g01507(.A0(new_n1699_), .A1(new_n1697_), .B0(new_n1676_), .B1(new_n1673_), .Y(new_n1700_));
  NOR3X1   g01508(.A(new_n1700_), .B(new_n1698_), .C(\asqrt[53] ), .Y(new_n1701_));
  NOR2X1   g01509(.A(new_n1701_), .B(new_n1688_), .Y(new_n1702_));
  NOR3X1   g01510(.A(new_n1518_), .B(new_n1487_), .C(new_n1481_), .Y(new_n1703_));
  OAI21X1  g01511(.A0(new_n1631_), .A1(new_n1612_), .B0(new_n1703_), .Y(new_n1704_));
  NOR3X1   g01512(.A(new_n1632_), .B(new_n1518_), .C(new_n1481_), .Y(new_n1705_));
  OR2X1    g01513(.A(new_n1705_), .B(new_n1486_), .Y(new_n1706_));
  AND2X1   g01514(.A(new_n1706_), .B(new_n1704_), .Y(new_n1707_));
  INVX1    g01515(.A(new_n1707_), .Y(new_n1708_));
  OR2X1    g01516(.A(new_n1681_), .B(\asqrt[54] ), .Y(new_n1709_));
  OAI21X1  g01517(.A0(new_n1709_), .A1(new_n1702_), .B0(new_n1708_), .Y(new_n1710_));
  AOI21X1  g01518(.A0(new_n1710_), .A1(new_n1692_), .B0(new_n697_), .Y(new_n1711_));
  INVX1    g01519(.A(new_n1632_), .Y(\asqrt[49] ));
  AOI21X1  g01520(.A0(new_n1533_), .A1(new_n1532_), .B0(new_n1497_), .Y(new_n1713_));
  AND2X1   g01521(.A(new_n1713_), .B(new_n1490_), .Y(new_n1714_));
  AOI22X1  g01522(.A0(new_n1533_), .A1(new_n1532_), .B0(new_n1519_), .B1(\asqrt[54] ), .Y(new_n1715_));
  AOI21X1  g01523(.A0(new_n1715_), .A1(\asqrt[49] ), .B0(new_n1496_), .Y(new_n1716_));
  AOI21X1  g01524(.A0(new_n1714_), .A1(\asqrt[49] ), .B0(new_n1716_), .Y(new_n1717_));
  OAI21X1  g01525(.A0(new_n1700_), .A1(new_n1698_), .B0(\asqrt[53] ), .Y(new_n1718_));
  OAI21X1  g01526(.A0(new_n1701_), .A1(new_n1688_), .B0(new_n1718_), .Y(new_n1719_));
  AOI21X1  g01527(.A0(new_n1719_), .A1(\asqrt[54] ), .B0(\asqrt[55] ), .Y(new_n1720_));
  AOI21X1  g01528(.A0(new_n1720_), .A1(new_n1710_), .B0(new_n1717_), .Y(new_n1721_));
  OAI21X1  g01529(.A0(new_n1721_), .A1(new_n1711_), .B0(\asqrt[56] ), .Y(new_n1722_));
  AND2X1   g01530(.A(new_n1520_), .B(new_n1499_), .Y(new_n1723_));
  NOR3X1   g01531(.A(new_n1723_), .B(new_n1536_), .C(new_n1500_), .Y(new_n1724_));
  NOR3X1   g01532(.A(new_n1632_), .B(new_n1723_), .C(new_n1500_), .Y(new_n1725_));
  NOR2X1   g01533(.A(new_n1725_), .B(new_n1505_), .Y(new_n1726_));
  AOI21X1  g01534(.A0(new_n1724_), .A1(\asqrt[49] ), .B0(new_n1726_), .Y(new_n1727_));
  NOR3X1   g01535(.A(new_n1721_), .B(new_n1711_), .C(\asqrt[56] ), .Y(new_n1728_));
  OAI21X1  g01536(.A0(new_n1728_), .A1(new_n1727_), .B0(new_n1722_), .Y(new_n1729_));
  AND2X1   g01537(.A(new_n1729_), .B(\asqrt[57] ), .Y(new_n1730_));
  INVX1    g01538(.A(new_n1727_), .Y(new_n1731_));
  AND2X1   g01539(.A(new_n1719_), .B(\asqrt[54] ), .Y(new_n1732_));
  OR2X1    g01540(.A(new_n1701_), .B(new_n1688_), .Y(new_n1733_));
  NOR2X1   g01541(.A(new_n1681_), .B(\asqrt[54] ), .Y(new_n1734_));
  AOI21X1  g01542(.A0(new_n1734_), .A1(new_n1733_), .B0(new_n1707_), .Y(new_n1735_));
  OAI21X1  g01543(.A0(new_n1735_), .A1(new_n1732_), .B0(\asqrt[55] ), .Y(new_n1736_));
  INVX1    g01544(.A(new_n1717_), .Y(new_n1737_));
  OAI21X1  g01545(.A0(new_n1691_), .A1(new_n902_), .B0(new_n697_), .Y(new_n1738_));
  OAI21X1  g01546(.A0(new_n1738_), .A1(new_n1735_), .B0(new_n1737_), .Y(new_n1739_));
  NAND3X1  g01547(.A(new_n1739_), .B(new_n1736_), .C(new_n582_), .Y(new_n1740_));
  NAND2X1  g01548(.A(new_n1740_), .B(new_n1731_), .Y(new_n1741_));
  OR4X1    g01549(.A(new_n1632_), .B(new_n1527_), .C(new_n1530_), .D(new_n1546_), .Y(new_n1742_));
  NAND2X1  g01550(.A(new_n1539_), .B(new_n1522_), .Y(new_n1743_));
  OAI21X1  g01551(.A0(new_n1743_), .A1(new_n1632_), .B0(new_n1530_), .Y(new_n1744_));
  AND2X1   g01552(.A(new_n1744_), .B(new_n1742_), .Y(new_n1745_));
  AND2X1   g01553(.A(new_n1722_), .B(new_n481_), .Y(new_n1746_));
  AOI21X1  g01554(.A0(new_n1746_), .A1(new_n1741_), .B0(new_n1745_), .Y(new_n1747_));
  OAI21X1  g01555(.A0(new_n1747_), .A1(new_n1730_), .B0(\asqrt[58] ), .Y(new_n1748_));
  AND2X1   g01556(.A(new_n1547_), .B(new_n1540_), .Y(new_n1749_));
  NOR3X1   g01557(.A(new_n1749_), .B(new_n1575_), .C(new_n1529_), .Y(new_n1750_));
  NOR3X1   g01558(.A(new_n1632_), .B(new_n1749_), .C(new_n1529_), .Y(new_n1751_));
  NOR2X1   g01559(.A(new_n1751_), .B(new_n1545_), .Y(new_n1752_));
  AOI21X1  g01560(.A0(new_n1750_), .A1(\asqrt[49] ), .B0(new_n1752_), .Y(new_n1753_));
  INVX1    g01561(.A(new_n1753_), .Y(new_n1754_));
  AOI21X1  g01562(.A0(new_n1739_), .A1(new_n1736_), .B0(new_n582_), .Y(new_n1755_));
  AOI21X1  g01563(.A0(new_n1740_), .A1(new_n1731_), .B0(new_n1755_), .Y(new_n1756_));
  OAI21X1  g01564(.A0(new_n1756_), .A1(new_n481_), .B0(new_n399_), .Y(new_n1757_));
  OAI21X1  g01565(.A0(new_n1757_), .A1(new_n1747_), .B0(new_n1754_), .Y(new_n1758_));
  AOI21X1  g01566(.A0(new_n1758_), .A1(new_n1748_), .B0(new_n328_), .Y(new_n1759_));
  AND2X1   g01567(.A(new_n1579_), .B(new_n1577_), .Y(new_n1760_));
  NOR3X1   g01568(.A(new_n1760_), .B(new_n1555_), .C(new_n1578_), .Y(new_n1761_));
  NOR3X1   g01569(.A(new_n1632_), .B(new_n1760_), .C(new_n1578_), .Y(new_n1762_));
  NOR2X1   g01570(.A(new_n1762_), .B(new_n1554_), .Y(new_n1763_));
  AOI21X1  g01571(.A0(new_n1761_), .A1(\asqrt[49] ), .B0(new_n1763_), .Y(new_n1764_));
  INVX1    g01572(.A(new_n1764_), .Y(new_n1765_));
  NAND3X1  g01573(.A(new_n1758_), .B(new_n1748_), .C(new_n328_), .Y(new_n1766_));
  AOI21X1  g01574(.A0(new_n1766_), .A1(new_n1765_), .B0(new_n1759_), .Y(new_n1767_));
  OR2X1    g01575(.A(new_n1767_), .B(new_n292_), .Y(new_n1768_));
  AND2X1   g01576(.A(new_n1766_), .B(new_n1765_), .Y(new_n1769_));
  OR4X1    g01577(.A(new_n1632_), .B(new_n1591_), .C(new_n1562_), .D(new_n1559_), .Y(new_n1770_));
  OR2X1    g01578(.A(new_n1591_), .B(new_n1559_), .Y(new_n1771_));
  OAI21X1  g01579(.A0(new_n1771_), .A1(new_n1632_), .B0(new_n1562_), .Y(new_n1772_));
  AND2X1   g01580(.A(new_n1772_), .B(new_n1770_), .Y(new_n1773_));
  INVX1    g01581(.A(new_n1773_), .Y(new_n1774_));
  OR2X1    g01582(.A(new_n1759_), .B(\asqrt[60] ), .Y(new_n1775_));
  OAI21X1  g01583(.A0(new_n1775_), .A1(new_n1769_), .B0(new_n1774_), .Y(new_n1776_));
  AOI21X1  g01584(.A0(new_n1776_), .A1(new_n1768_), .B0(new_n217_), .Y(new_n1777_));
  AOI21X1  g01585(.A0(new_n1615_), .A1(new_n1614_), .B0(new_n1572_), .Y(new_n1778_));
  AND2X1   g01586(.A(new_n1778_), .B(new_n1565_), .Y(new_n1779_));
  AOI22X1  g01587(.A0(new_n1615_), .A1(new_n1614_), .B0(new_n1592_), .B1(\asqrt[60] ), .Y(new_n1780_));
  AOI21X1  g01588(.A0(new_n1780_), .A1(\asqrt[49] ), .B0(new_n1571_), .Y(new_n1781_));
  AOI21X1  g01589(.A0(new_n1779_), .A1(\asqrt[49] ), .B0(new_n1781_), .Y(new_n1782_));
  OR2X1    g01590(.A(new_n1756_), .B(new_n481_), .Y(new_n1783_));
  AND2X1   g01591(.A(new_n1740_), .B(new_n1731_), .Y(new_n1784_));
  INVX1    g01592(.A(new_n1745_), .Y(new_n1785_));
  NAND2X1  g01593(.A(new_n1722_), .B(new_n481_), .Y(new_n1786_));
  OAI21X1  g01594(.A0(new_n1786_), .A1(new_n1784_), .B0(new_n1785_), .Y(new_n1787_));
  AOI21X1  g01595(.A0(new_n1787_), .A1(new_n1783_), .B0(new_n399_), .Y(new_n1788_));
  AOI21X1  g01596(.A0(new_n1729_), .A1(\asqrt[57] ), .B0(\asqrt[58] ), .Y(new_n1789_));
  AOI21X1  g01597(.A0(new_n1789_), .A1(new_n1787_), .B0(new_n1753_), .Y(new_n1790_));
  OAI21X1  g01598(.A0(new_n1790_), .A1(new_n1788_), .B0(\asqrt[59] ), .Y(new_n1791_));
  NOR3X1   g01599(.A(new_n1790_), .B(new_n1788_), .C(\asqrt[59] ), .Y(new_n1792_));
  OAI21X1  g01600(.A0(new_n1792_), .A1(new_n1764_), .B0(new_n1791_), .Y(new_n1793_));
  AOI21X1  g01601(.A0(new_n1793_), .A1(\asqrt[60] ), .B0(\asqrt[61] ), .Y(new_n1794_));
  AOI21X1  g01602(.A0(new_n1794_), .A1(new_n1776_), .B0(new_n1782_), .Y(new_n1795_));
  OAI21X1  g01603(.A0(new_n1795_), .A1(new_n1777_), .B0(\asqrt[62] ), .Y(new_n1796_));
  AND2X1   g01604(.A(new_n1593_), .B(new_n1583_), .Y(new_n1797_));
  NOR3X1   g01605(.A(new_n1797_), .B(new_n1618_), .C(new_n1584_), .Y(new_n1798_));
  NOR3X1   g01606(.A(new_n1632_), .B(new_n1797_), .C(new_n1584_), .Y(new_n1799_));
  NOR2X1   g01607(.A(new_n1799_), .B(new_n1589_), .Y(new_n1800_));
  AOI21X1  g01608(.A0(new_n1798_), .A1(\asqrt[49] ), .B0(new_n1800_), .Y(new_n1801_));
  NOR3X1   g01609(.A(new_n1795_), .B(new_n1777_), .C(\asqrt[62] ), .Y(new_n1802_));
  OAI21X1  g01610(.A0(new_n1802_), .A1(new_n1801_), .B0(new_n1796_), .Y(new_n1803_));
  NOR4X1   g01611(.A(new_n1632_), .B(new_n1600_), .C(new_n1598_), .D(new_n1637_), .Y(new_n1804_));
  NAND3X1  g01612(.A(\asqrt[49] ), .B(new_n1621_), .C(new_n1595_), .Y(new_n1805_));
  AOI21X1  g01613(.A0(new_n1805_), .A1(new_n1598_), .B0(new_n1804_), .Y(new_n1806_));
  INVX1    g01614(.A(new_n1806_), .Y(new_n1807_));
  NOR2X1   g01615(.A(new_n1606_), .B(new_n1638_), .Y(new_n1808_));
  AOI21X1  g01616(.A0(new_n1808_), .A1(\asqrt[49] ), .B0(new_n1662_), .Y(new_n1809_));
  AND2X1   g01617(.A(new_n1809_), .B(new_n1807_), .Y(new_n1810_));
  AOI21X1  g01618(.A0(new_n1810_), .A1(new_n1803_), .B0(\asqrt[63] ), .Y(new_n1811_));
  INVX1    g01619(.A(new_n1801_), .Y(new_n1812_));
  AND2X1   g01620(.A(new_n1793_), .B(\asqrt[60] ), .Y(new_n1813_));
  NAND2X1  g01621(.A(new_n1766_), .B(new_n1765_), .Y(new_n1814_));
  NOR2X1   g01622(.A(new_n1759_), .B(\asqrt[60] ), .Y(new_n1815_));
  AOI21X1  g01623(.A0(new_n1815_), .A1(new_n1814_), .B0(new_n1773_), .Y(new_n1816_));
  OAI21X1  g01624(.A0(new_n1816_), .A1(new_n1813_), .B0(\asqrt[61] ), .Y(new_n1817_));
  INVX1    g01625(.A(new_n1782_), .Y(new_n1818_));
  OAI21X1  g01626(.A0(new_n1767_), .A1(new_n292_), .B0(new_n217_), .Y(new_n1819_));
  OAI21X1  g01627(.A0(new_n1819_), .A1(new_n1816_), .B0(new_n1818_), .Y(new_n1820_));
  NAND3X1  g01628(.A(new_n1820_), .B(new_n1817_), .C(new_n199_), .Y(new_n1821_));
  AND2X1   g01629(.A(new_n1821_), .B(new_n1812_), .Y(new_n1822_));
  AOI21X1  g01630(.A0(new_n1820_), .A1(new_n1817_), .B0(new_n199_), .Y(new_n1823_));
  OR2X1    g01631(.A(new_n1807_), .B(new_n1823_), .Y(new_n1824_));
  AOI21X1  g01632(.A0(new_n1644_), .A1(new_n1640_), .B0(new_n1606_), .Y(new_n1825_));
  AOI21X1  g01633(.A0(new_n1607_), .A1(new_n1601_), .B0(new_n193_), .Y(new_n1826_));
  OAI21X1  g01634(.A0(new_n1825_), .A1(new_n1601_), .B0(new_n1826_), .Y(new_n1827_));
  NOR4X1   g01635(.A(new_n1629_), .B(new_n1626_), .C(new_n1605_), .D(new_n1603_), .Y(new_n1828_));
  OAI21X1  g01636(.A0(new_n1623_), .A1(new_n1622_), .B0(new_n1828_), .Y(new_n1829_));
  NOR2X1   g01637(.A(new_n1829_), .B(new_n1612_), .Y(new_n1830_));
  INVX1    g01638(.A(new_n1830_), .Y(new_n1831_));
  AND2X1   g01639(.A(new_n1831_), .B(new_n1827_), .Y(new_n1832_));
  OAI21X1  g01640(.A0(new_n1824_), .A1(new_n1822_), .B0(new_n1832_), .Y(new_n1833_));
  NOR2X1   g01641(.A(new_n1833_), .B(new_n1811_), .Y(new_n1834_));
  OR2X1    g01642(.A(new_n1833_), .B(new_n1811_), .Y(\asqrt[48] ));
  NOR3X1   g01643(.A(\a[96] ), .B(\a[95] ), .C(\a[94] ), .Y(new_n1836_));
  AOI21X1  g01644(.A0(\asqrt[48] ), .A1(\a[96] ), .B0(new_n1836_), .Y(new_n1837_));
  INVX1    g01645(.A(\a[97] ), .Y(new_n1838_));
  AOI21X1  g01646(.A0(new_n1821_), .A1(new_n1812_), .B0(new_n1823_), .Y(new_n1839_));
  INVX1    g01647(.A(new_n1810_), .Y(new_n1840_));
  OAI21X1  g01648(.A0(new_n1840_), .A1(new_n1839_), .B0(new_n193_), .Y(new_n1841_));
  NAND2X1  g01649(.A(new_n1821_), .B(new_n1812_), .Y(new_n1842_));
  NOR2X1   g01650(.A(new_n1807_), .B(new_n1823_), .Y(new_n1843_));
  INVX1    g01651(.A(new_n1832_), .Y(new_n1844_));
  AOI21X1  g01652(.A0(new_n1843_), .A1(new_n1842_), .B0(new_n1844_), .Y(new_n1845_));
  AOI21X1  g01653(.A0(new_n1845_), .A1(new_n1841_), .B0(\a[96] ), .Y(new_n1846_));
  OAI21X1  g01654(.A0(new_n1833_), .A1(new_n1811_), .B0(new_n1633_), .Y(new_n1847_));
  OAI21X1  g01655(.A0(new_n1846_), .A1(new_n1838_), .B0(new_n1847_), .Y(new_n1848_));
  OAI21X1  g01656(.A0(new_n1833_), .A1(new_n1811_), .B0(\a[96] ), .Y(new_n1849_));
  OR2X1    g01657(.A(new_n1836_), .B(new_n1629_), .Y(new_n1850_));
  NOR4X1   g01658(.A(new_n1850_), .B(new_n1626_), .C(new_n1662_), .D(new_n1612_), .Y(new_n1851_));
  AND2X1   g01659(.A(new_n1851_), .B(new_n1849_), .Y(new_n1852_));
  OAI22X1  g01660(.A0(new_n1852_), .A1(new_n1848_), .B0(new_n1837_), .B1(new_n1632_), .Y(new_n1853_));
  AND2X1   g01661(.A(new_n1853_), .B(\asqrt[50] ), .Y(new_n1854_));
  INVX1    g01662(.A(\a[96] ), .Y(new_n1855_));
  OAI21X1  g01663(.A0(new_n1833_), .A1(new_n1811_), .B0(new_n1855_), .Y(new_n1856_));
  AOI21X1  g01664(.A0(new_n1845_), .A1(new_n1841_), .B0(new_n1634_), .Y(new_n1857_));
  AOI21X1  g01665(.A0(new_n1856_), .A1(\a[97] ), .B0(new_n1857_), .Y(new_n1858_));
  NAND2X1  g01666(.A(new_n1851_), .B(new_n1849_), .Y(new_n1859_));
  NAND2X1  g01667(.A(new_n1859_), .B(new_n1858_), .Y(new_n1860_));
  NOR2X1   g01668(.A(\a[95] ), .B(\a[94] ), .Y(new_n1861_));
  MX2X1    g01669(.A(new_n1861_), .B(\asqrt[48] ), .S0(\a[96] ), .Y(new_n1862_));
  AOI21X1  g01670(.A0(new_n1862_), .A1(\asqrt[49] ), .B0(\asqrt[50] ), .Y(new_n1863_));
  INVX1    g01671(.A(new_n1827_), .Y(new_n1864_));
  NOR3X1   g01672(.A(new_n1830_), .B(new_n1864_), .C(new_n1632_), .Y(new_n1865_));
  OAI21X1  g01673(.A0(new_n1824_), .A1(new_n1822_), .B0(new_n1865_), .Y(new_n1866_));
  OR2X1    g01674(.A(new_n1866_), .B(new_n1811_), .Y(new_n1867_));
  AOI21X1  g01675(.A0(new_n1867_), .A1(new_n1847_), .B0(new_n1636_), .Y(new_n1868_));
  OAI21X1  g01676(.A0(new_n1866_), .A1(new_n1811_), .B0(new_n1636_), .Y(new_n1869_));
  NOR2X1   g01677(.A(new_n1869_), .B(new_n1857_), .Y(new_n1870_));
  NOR2X1   g01678(.A(new_n1870_), .B(new_n1868_), .Y(new_n1871_));
  AOI21X1  g01679(.A0(new_n1863_), .A1(new_n1860_), .B0(new_n1871_), .Y(new_n1872_));
  OAI21X1  g01680(.A0(new_n1872_), .A1(new_n1854_), .B0(\asqrt[51] ), .Y(new_n1873_));
  AOI21X1  g01681(.A0(new_n1660_), .A1(\asqrt[50] ), .B0(new_n1648_), .Y(new_n1874_));
  AND2X1   g01682(.A(new_n1874_), .B(new_n1652_), .Y(new_n1875_));
  OAI21X1  g01683(.A0(new_n1833_), .A1(new_n1811_), .B0(new_n1874_), .Y(new_n1876_));
  AOI22X1  g01684(.A0(new_n1876_), .A1(new_n1658_), .B0(new_n1875_), .B1(\asqrt[48] ), .Y(new_n1877_));
  INVX1    g01685(.A(new_n1877_), .Y(new_n1878_));
  AOI22X1  g01686(.A0(new_n1859_), .A1(new_n1858_), .B0(new_n1862_), .B1(\asqrt[49] ), .Y(new_n1879_));
  OAI21X1  g01687(.A0(new_n1879_), .A1(new_n1469_), .B0(new_n1277_), .Y(new_n1880_));
  OAI21X1  g01688(.A0(new_n1880_), .A1(new_n1872_), .B0(new_n1878_), .Y(new_n1881_));
  AOI21X1  g01689(.A0(new_n1881_), .A1(new_n1873_), .B0(new_n1111_), .Y(new_n1882_));
  AOI21X1  g01690(.A0(new_n1661_), .A1(new_n1659_), .B0(new_n1696_), .Y(new_n1883_));
  AND2X1   g01691(.A(new_n1883_), .B(new_n1693_), .Y(new_n1884_));
  AOI22X1  g01692(.A0(new_n1661_), .A1(new_n1659_), .B0(new_n1653_), .B1(\asqrt[51] ), .Y(new_n1885_));
  OAI21X1  g01693(.A0(new_n1833_), .A1(new_n1811_), .B0(new_n1885_), .Y(new_n1886_));
  AOI22X1  g01694(.A0(new_n1886_), .A1(new_n1696_), .B0(new_n1884_), .B1(\asqrt[48] ), .Y(new_n1887_));
  INVX1    g01695(.A(new_n1887_), .Y(new_n1888_));
  NAND3X1  g01696(.A(new_n1881_), .B(new_n1873_), .C(new_n1111_), .Y(new_n1889_));
  AOI21X1  g01697(.A0(new_n1889_), .A1(new_n1888_), .B0(new_n1882_), .Y(new_n1890_));
  OR2X1    g01698(.A(new_n1890_), .B(new_n968_), .Y(new_n1891_));
  AND2X1   g01699(.A(new_n1889_), .B(new_n1888_), .Y(new_n1892_));
  AND2X1   g01700(.A(new_n1699_), .B(new_n1697_), .Y(new_n1893_));
  NOR3X1   g01701(.A(new_n1893_), .B(new_n1677_), .C(new_n1698_), .Y(new_n1894_));
  NOR2X1   g01702(.A(new_n1893_), .B(new_n1698_), .Y(new_n1895_));
  OAI21X1  g01703(.A0(new_n1833_), .A1(new_n1811_), .B0(new_n1895_), .Y(new_n1896_));
  AOI22X1  g01704(.A0(new_n1896_), .A1(new_n1677_), .B0(new_n1894_), .B1(\asqrt[48] ), .Y(new_n1897_));
  INVX1    g01705(.A(new_n1897_), .Y(new_n1898_));
  OR2X1    g01706(.A(new_n1882_), .B(\asqrt[53] ), .Y(new_n1899_));
  OAI21X1  g01707(.A0(new_n1899_), .A1(new_n1892_), .B0(new_n1898_), .Y(new_n1900_));
  AOI21X1  g01708(.A0(new_n1900_), .A1(new_n1891_), .B0(new_n902_), .Y(new_n1901_));
  NAND4X1  g01709(.A(\asqrt[48] ), .B(new_n1690_), .C(new_n1688_), .D(new_n1718_), .Y(new_n1902_));
  NOR3X1   g01710(.A(new_n1834_), .B(new_n1701_), .C(new_n1681_), .Y(new_n1903_));
  OAI21X1  g01711(.A0(new_n1903_), .A1(new_n1688_), .B0(new_n1902_), .Y(new_n1904_));
  INVX1    g01712(.A(new_n1904_), .Y(new_n1905_));
  OR2X1    g01713(.A(new_n1879_), .B(new_n1469_), .Y(new_n1906_));
  AND2X1   g01714(.A(new_n1859_), .B(new_n1858_), .Y(new_n1907_));
  OAI21X1  g01715(.A0(new_n1837_), .A1(new_n1632_), .B0(new_n1469_), .Y(new_n1908_));
  OR2X1    g01716(.A(new_n1870_), .B(new_n1868_), .Y(new_n1909_));
  OAI21X1  g01717(.A0(new_n1908_), .A1(new_n1907_), .B0(new_n1909_), .Y(new_n1910_));
  AOI21X1  g01718(.A0(new_n1910_), .A1(new_n1906_), .B0(new_n1277_), .Y(new_n1911_));
  AOI21X1  g01719(.A0(new_n1853_), .A1(\asqrt[50] ), .B0(\asqrt[51] ), .Y(new_n1912_));
  AOI21X1  g01720(.A0(new_n1912_), .A1(new_n1910_), .B0(new_n1877_), .Y(new_n1913_));
  OAI21X1  g01721(.A0(new_n1913_), .A1(new_n1911_), .B0(\asqrt[52] ), .Y(new_n1914_));
  NOR3X1   g01722(.A(new_n1913_), .B(new_n1911_), .C(\asqrt[52] ), .Y(new_n1915_));
  OAI21X1  g01723(.A0(new_n1915_), .A1(new_n1887_), .B0(new_n1914_), .Y(new_n1916_));
  AOI21X1  g01724(.A0(new_n1916_), .A1(\asqrt[53] ), .B0(\asqrt[54] ), .Y(new_n1917_));
  AOI21X1  g01725(.A0(new_n1917_), .A1(new_n1900_), .B0(new_n1905_), .Y(new_n1918_));
  OAI21X1  g01726(.A0(new_n1918_), .A1(new_n1901_), .B0(\asqrt[55] ), .Y(new_n1919_));
  AND2X1   g01727(.A(new_n1734_), .B(new_n1733_), .Y(new_n1920_));
  NOR3X1   g01728(.A(new_n1920_), .B(new_n1708_), .C(new_n1732_), .Y(new_n1921_));
  AOI22X1  g01729(.A0(new_n1734_), .A1(new_n1733_), .B0(new_n1719_), .B1(\asqrt[54] ), .Y(new_n1922_));
  AOI21X1  g01730(.A0(new_n1922_), .A1(\asqrt[48] ), .B0(new_n1707_), .Y(new_n1923_));
  AOI21X1  g01731(.A0(new_n1921_), .A1(\asqrt[48] ), .B0(new_n1923_), .Y(new_n1924_));
  NOR3X1   g01732(.A(new_n1918_), .B(new_n1901_), .C(\asqrt[55] ), .Y(new_n1925_));
  OAI21X1  g01733(.A0(new_n1925_), .A1(new_n1924_), .B0(new_n1919_), .Y(new_n1926_));
  AND2X1   g01734(.A(new_n1926_), .B(\asqrt[56] ), .Y(new_n1927_));
  INVX1    g01735(.A(new_n1924_), .Y(new_n1928_));
  AND2X1   g01736(.A(new_n1916_), .B(\asqrt[53] ), .Y(new_n1929_));
  NAND2X1  g01737(.A(new_n1889_), .B(new_n1888_), .Y(new_n1930_));
  NOR2X1   g01738(.A(new_n1882_), .B(\asqrt[53] ), .Y(new_n1931_));
  AOI21X1  g01739(.A0(new_n1931_), .A1(new_n1930_), .B0(new_n1897_), .Y(new_n1932_));
  OAI21X1  g01740(.A0(new_n1932_), .A1(new_n1929_), .B0(\asqrt[54] ), .Y(new_n1933_));
  OAI21X1  g01741(.A0(new_n1890_), .A1(new_n968_), .B0(new_n902_), .Y(new_n1934_));
  OAI21X1  g01742(.A0(new_n1934_), .A1(new_n1932_), .B0(new_n1904_), .Y(new_n1935_));
  NAND3X1  g01743(.A(new_n1935_), .B(new_n1933_), .C(new_n697_), .Y(new_n1936_));
  NAND2X1  g01744(.A(new_n1936_), .B(new_n1928_), .Y(new_n1937_));
  AND2X1   g01745(.A(new_n1720_), .B(new_n1710_), .Y(new_n1938_));
  NOR3X1   g01746(.A(new_n1938_), .B(new_n1737_), .C(new_n1711_), .Y(new_n1939_));
  NOR2X1   g01747(.A(new_n1938_), .B(new_n1711_), .Y(new_n1940_));
  AOI21X1  g01748(.A0(new_n1940_), .A1(\asqrt[48] ), .B0(new_n1717_), .Y(new_n1941_));
  AOI21X1  g01749(.A0(new_n1939_), .A1(\asqrt[48] ), .B0(new_n1941_), .Y(new_n1942_));
  AOI21X1  g01750(.A0(new_n1935_), .A1(new_n1933_), .B0(new_n697_), .Y(new_n1943_));
  NOR2X1   g01751(.A(new_n1943_), .B(\asqrt[56] ), .Y(new_n1944_));
  AOI21X1  g01752(.A0(new_n1944_), .A1(new_n1937_), .B0(new_n1942_), .Y(new_n1945_));
  OAI21X1  g01753(.A0(new_n1945_), .A1(new_n1927_), .B0(\asqrt[57] ), .Y(new_n1946_));
  OR4X1    g01754(.A(new_n1834_), .B(new_n1728_), .C(new_n1731_), .D(new_n1755_), .Y(new_n1947_));
  OR2X1    g01755(.A(new_n1728_), .B(new_n1755_), .Y(new_n1948_));
  OAI21X1  g01756(.A0(new_n1948_), .A1(new_n1834_), .B0(new_n1731_), .Y(new_n1949_));
  AND2X1   g01757(.A(new_n1949_), .B(new_n1947_), .Y(new_n1950_));
  INVX1    g01758(.A(new_n1950_), .Y(new_n1951_));
  AOI21X1  g01759(.A0(new_n1936_), .A1(new_n1928_), .B0(new_n1943_), .Y(new_n1952_));
  OAI21X1  g01760(.A0(new_n1952_), .A1(new_n582_), .B0(new_n481_), .Y(new_n1953_));
  OAI21X1  g01761(.A0(new_n1953_), .A1(new_n1945_), .B0(new_n1951_), .Y(new_n1954_));
  AOI21X1  g01762(.A0(new_n1954_), .A1(new_n1946_), .B0(new_n399_), .Y(new_n1955_));
  AOI21X1  g01763(.A0(new_n1746_), .A1(new_n1741_), .B0(new_n1785_), .Y(new_n1956_));
  AND2X1   g01764(.A(new_n1956_), .B(new_n1783_), .Y(new_n1957_));
  AOI22X1  g01765(.A0(new_n1746_), .A1(new_n1741_), .B0(new_n1729_), .B1(\asqrt[57] ), .Y(new_n1958_));
  AOI21X1  g01766(.A0(new_n1958_), .A1(\asqrt[48] ), .B0(new_n1745_), .Y(new_n1959_));
  AOI21X1  g01767(.A0(new_n1957_), .A1(\asqrt[48] ), .B0(new_n1959_), .Y(new_n1960_));
  INVX1    g01768(.A(new_n1960_), .Y(new_n1961_));
  NAND3X1  g01769(.A(new_n1954_), .B(new_n1946_), .C(new_n399_), .Y(new_n1962_));
  AOI21X1  g01770(.A0(new_n1962_), .A1(new_n1961_), .B0(new_n1955_), .Y(new_n1963_));
  OR2X1    g01771(.A(new_n1963_), .B(new_n328_), .Y(new_n1964_));
  AND2X1   g01772(.A(new_n1962_), .B(new_n1961_), .Y(new_n1965_));
  AND2X1   g01773(.A(new_n1789_), .B(new_n1787_), .Y(new_n1966_));
  NOR3X1   g01774(.A(new_n1966_), .B(new_n1754_), .C(new_n1788_), .Y(new_n1967_));
  NOR2X1   g01775(.A(new_n1966_), .B(new_n1788_), .Y(new_n1968_));
  AOI21X1  g01776(.A0(new_n1968_), .A1(\asqrt[48] ), .B0(new_n1753_), .Y(new_n1969_));
  AOI21X1  g01777(.A0(new_n1967_), .A1(\asqrt[48] ), .B0(new_n1969_), .Y(new_n1970_));
  INVX1    g01778(.A(new_n1970_), .Y(new_n1971_));
  OR2X1    g01779(.A(new_n1955_), .B(\asqrt[59] ), .Y(new_n1972_));
  OAI21X1  g01780(.A0(new_n1972_), .A1(new_n1965_), .B0(new_n1971_), .Y(new_n1973_));
  AOI21X1  g01781(.A0(new_n1973_), .A1(new_n1964_), .B0(new_n292_), .Y(new_n1974_));
  OR4X1    g01782(.A(new_n1834_), .B(new_n1792_), .C(new_n1765_), .D(new_n1759_), .Y(new_n1975_));
  NAND2X1  g01783(.A(new_n1766_), .B(new_n1791_), .Y(new_n1976_));
  OAI21X1  g01784(.A0(new_n1976_), .A1(new_n1834_), .B0(new_n1765_), .Y(new_n1977_));
  AND2X1   g01785(.A(new_n1977_), .B(new_n1975_), .Y(new_n1978_));
  OR2X1    g01786(.A(new_n1952_), .B(new_n582_), .Y(new_n1979_));
  AND2X1   g01787(.A(new_n1936_), .B(new_n1928_), .Y(new_n1980_));
  INVX1    g01788(.A(new_n1942_), .Y(new_n1981_));
  OR2X1    g01789(.A(new_n1943_), .B(\asqrt[56] ), .Y(new_n1982_));
  OAI21X1  g01790(.A0(new_n1982_), .A1(new_n1980_), .B0(new_n1981_), .Y(new_n1983_));
  AOI21X1  g01791(.A0(new_n1983_), .A1(new_n1979_), .B0(new_n481_), .Y(new_n1984_));
  AOI21X1  g01792(.A0(new_n1926_), .A1(\asqrt[56] ), .B0(\asqrt[57] ), .Y(new_n1985_));
  AOI21X1  g01793(.A0(new_n1985_), .A1(new_n1983_), .B0(new_n1950_), .Y(new_n1986_));
  OAI21X1  g01794(.A0(new_n1986_), .A1(new_n1984_), .B0(\asqrt[58] ), .Y(new_n1987_));
  NOR3X1   g01795(.A(new_n1986_), .B(new_n1984_), .C(\asqrt[58] ), .Y(new_n1988_));
  OAI21X1  g01796(.A0(new_n1988_), .A1(new_n1960_), .B0(new_n1987_), .Y(new_n1989_));
  AOI21X1  g01797(.A0(new_n1989_), .A1(\asqrt[59] ), .B0(\asqrt[60] ), .Y(new_n1990_));
  AOI21X1  g01798(.A0(new_n1990_), .A1(new_n1973_), .B0(new_n1978_), .Y(new_n1991_));
  OAI21X1  g01799(.A0(new_n1991_), .A1(new_n1974_), .B0(\asqrt[61] ), .Y(new_n1992_));
  AND2X1   g01800(.A(new_n1815_), .B(new_n1814_), .Y(new_n1993_));
  NOR3X1   g01801(.A(new_n1993_), .B(new_n1774_), .C(new_n1813_), .Y(new_n1994_));
  AOI22X1  g01802(.A0(new_n1815_), .A1(new_n1814_), .B0(new_n1793_), .B1(\asqrt[60] ), .Y(new_n1995_));
  AOI21X1  g01803(.A0(new_n1995_), .A1(\asqrt[48] ), .B0(new_n1773_), .Y(new_n1996_));
  AOI21X1  g01804(.A0(new_n1994_), .A1(\asqrt[48] ), .B0(new_n1996_), .Y(new_n1997_));
  NOR3X1   g01805(.A(new_n1991_), .B(new_n1974_), .C(\asqrt[61] ), .Y(new_n1998_));
  OAI21X1  g01806(.A0(new_n1998_), .A1(new_n1997_), .B0(new_n1992_), .Y(new_n1999_));
  AND2X1   g01807(.A(new_n1999_), .B(\asqrt[62] ), .Y(new_n2000_));
  INVX1    g01808(.A(new_n1997_), .Y(new_n2001_));
  AND2X1   g01809(.A(new_n1989_), .B(\asqrt[59] ), .Y(new_n2002_));
  NAND2X1  g01810(.A(new_n1962_), .B(new_n1961_), .Y(new_n2003_));
  NOR2X1   g01811(.A(new_n1955_), .B(\asqrt[59] ), .Y(new_n2004_));
  AOI21X1  g01812(.A0(new_n2004_), .A1(new_n2003_), .B0(new_n1970_), .Y(new_n2005_));
  OAI21X1  g01813(.A0(new_n2005_), .A1(new_n2002_), .B0(\asqrt[60] ), .Y(new_n2006_));
  INVX1    g01814(.A(new_n1978_), .Y(new_n2007_));
  OAI21X1  g01815(.A0(new_n1963_), .A1(new_n328_), .B0(new_n292_), .Y(new_n2008_));
  OAI21X1  g01816(.A0(new_n2008_), .A1(new_n2005_), .B0(new_n2007_), .Y(new_n2009_));
  NAND3X1  g01817(.A(new_n2009_), .B(new_n2006_), .C(new_n217_), .Y(new_n2010_));
  NAND2X1  g01818(.A(new_n2010_), .B(new_n2001_), .Y(new_n2011_));
  AND2X1   g01819(.A(new_n1794_), .B(new_n1776_), .Y(new_n2012_));
  NOR3X1   g01820(.A(new_n2012_), .B(new_n1818_), .C(new_n1777_), .Y(new_n2013_));
  NOR2X1   g01821(.A(new_n2012_), .B(new_n1777_), .Y(new_n2014_));
  AOI21X1  g01822(.A0(new_n2014_), .A1(\asqrt[48] ), .B0(new_n1782_), .Y(new_n2015_));
  AOI21X1  g01823(.A0(new_n2013_), .A1(\asqrt[48] ), .B0(new_n2015_), .Y(new_n2016_));
  AOI21X1  g01824(.A0(new_n2009_), .A1(new_n2006_), .B0(new_n217_), .Y(new_n2017_));
  NOR2X1   g01825(.A(new_n2017_), .B(\asqrt[62] ), .Y(new_n2018_));
  AOI21X1  g01826(.A0(new_n2018_), .A1(new_n2011_), .B0(new_n2016_), .Y(new_n2019_));
  OR4X1    g01827(.A(new_n1834_), .B(new_n1802_), .C(new_n1812_), .D(new_n1823_), .Y(new_n2020_));
  NAND2X1  g01828(.A(new_n1821_), .B(new_n1796_), .Y(new_n2021_));
  OAI21X1  g01829(.A0(new_n2021_), .A1(new_n1834_), .B0(new_n1812_), .Y(new_n2022_));
  AND2X1   g01830(.A(new_n2022_), .B(new_n2020_), .Y(new_n2023_));
  INVX1    g01831(.A(new_n2023_), .Y(new_n2024_));
  NOR2X1   g01832(.A(new_n1806_), .B(new_n1839_), .Y(new_n2025_));
  AOI22X1  g01833(.A0(new_n2025_), .A1(\asqrt[48] ), .B0(new_n1843_), .B1(new_n1842_), .Y(new_n2026_));
  AND2X1   g01834(.A(new_n2026_), .B(new_n2024_), .Y(new_n2027_));
  OAI21X1  g01835(.A0(new_n2019_), .A1(new_n2000_), .B0(new_n2027_), .Y(new_n2028_));
  AOI21X1  g01836(.A0(new_n2010_), .A1(new_n2001_), .B0(new_n2017_), .Y(new_n2029_));
  OAI21X1  g01837(.A0(new_n2029_), .A1(new_n199_), .B0(new_n2023_), .Y(new_n2030_));
  AOI21X1  g01838(.A0(new_n1845_), .A1(new_n1841_), .B0(new_n1806_), .Y(new_n2031_));
  AOI21X1  g01839(.A0(new_n1807_), .A1(new_n1803_), .B0(new_n193_), .Y(new_n2032_));
  OAI21X1  g01840(.A0(new_n2031_), .A1(new_n1803_), .B0(new_n2032_), .Y(new_n2033_));
  OR2X1    g01841(.A(new_n1824_), .B(new_n1822_), .Y(new_n2034_));
  AND2X1   g01842(.A(new_n1805_), .B(new_n1598_), .Y(new_n2035_));
  NOR4X1   g01843(.A(new_n1830_), .B(new_n1864_), .C(new_n2035_), .D(new_n1804_), .Y(new_n2036_));
  NAND3X1  g01844(.A(new_n2036_), .B(new_n2034_), .C(new_n1841_), .Y(new_n2037_));
  AND2X1   g01845(.A(new_n2037_), .B(new_n2033_), .Y(new_n2038_));
  OAI21X1  g01846(.A0(new_n2030_), .A1(new_n2019_), .B0(new_n2038_), .Y(new_n2039_));
  AOI21X1  g01847(.A0(new_n2028_), .A1(new_n193_), .B0(new_n2039_), .Y(new_n2040_));
  NOR2X1   g01848(.A(\a[93] ), .B(\a[92] ), .Y(new_n2041_));
  INVX1    g01849(.A(new_n2041_), .Y(new_n2042_));
  MX2X1    g01850(.A(new_n2042_), .B(new_n2040_), .S0(\a[94] ), .Y(new_n2043_));
  OR2X1    g01851(.A(new_n2043_), .B(new_n1834_), .Y(new_n2044_));
  INVX1    g01852(.A(\a[94] ), .Y(new_n2045_));
  NOR3X1   g01853(.A(\a[94] ), .B(\a[93] ), .C(\a[92] ), .Y(new_n2046_));
  NOR3X1   g01854(.A(new_n2046_), .B(new_n1830_), .C(new_n1864_), .Y(new_n2047_));
  NAND3X1  g01855(.A(new_n2047_), .B(new_n2034_), .C(new_n1841_), .Y(new_n2048_));
  INVX1    g01856(.A(new_n2048_), .Y(new_n2049_));
  OAI21X1  g01857(.A0(new_n2040_), .A1(new_n2045_), .B0(new_n2049_), .Y(new_n2050_));
  OAI21X1  g01858(.A0(new_n2040_), .A1(\a[94] ), .B0(\a[95] ), .Y(new_n2051_));
  INVX1    g01859(.A(new_n1861_), .Y(new_n2052_));
  OR2X1    g01860(.A(new_n2040_), .B(new_n2052_), .Y(new_n2053_));
  NAND3X1  g01861(.A(new_n2053_), .B(new_n2051_), .C(new_n2050_), .Y(new_n2054_));
  AOI21X1  g01862(.A0(new_n2054_), .A1(new_n2044_), .B0(new_n1632_), .Y(new_n2055_));
  OR2X1    g01863(.A(new_n2029_), .B(new_n199_), .Y(new_n2056_));
  AND2X1   g01864(.A(new_n2010_), .B(new_n2001_), .Y(new_n2057_));
  INVX1    g01865(.A(new_n2016_), .Y(new_n2058_));
  OR2X1    g01866(.A(new_n2017_), .B(\asqrt[62] ), .Y(new_n2059_));
  OAI21X1  g01867(.A0(new_n2059_), .A1(new_n2057_), .B0(new_n2058_), .Y(new_n2060_));
  INVX1    g01868(.A(new_n2027_), .Y(new_n2061_));
  AOI21X1  g01869(.A0(new_n2060_), .A1(new_n2056_), .B0(new_n2061_), .Y(new_n2062_));
  AOI21X1  g01870(.A0(new_n1999_), .A1(\asqrt[62] ), .B0(new_n2024_), .Y(new_n2063_));
  INVX1    g01871(.A(new_n2038_), .Y(new_n2064_));
  AOI21X1  g01872(.A0(new_n2063_), .A1(new_n2060_), .B0(new_n2064_), .Y(new_n2065_));
  OAI21X1  g01873(.A0(new_n2062_), .A1(\asqrt[63] ), .B0(new_n2065_), .Y(\asqrt[47] ));
  MX2X1    g01874(.A(new_n2041_), .B(\asqrt[47] ), .S0(\a[94] ), .Y(new_n2067_));
  AOI21X1  g01875(.A0(new_n2067_), .A1(\asqrt[48] ), .B0(\asqrt[49] ), .Y(new_n2068_));
  NAND3X1  g01876(.A(new_n2037_), .B(new_n2033_), .C(\asqrt[48] ), .Y(new_n2069_));
  INVX1    g01877(.A(new_n2069_), .Y(new_n2070_));
  OAI21X1  g01878(.A0(new_n2030_), .A1(new_n2019_), .B0(new_n2070_), .Y(new_n2071_));
  AOI21X1  g01879(.A0(new_n2028_), .A1(new_n193_), .B0(new_n2071_), .Y(new_n2072_));
  AOI21X1  g01880(.A0(\asqrt[47] ), .A1(new_n1861_), .B0(new_n2072_), .Y(new_n2073_));
  OR2X1    g01881(.A(new_n2073_), .B(new_n1855_), .Y(new_n2074_));
  AND2X1   g01882(.A(\asqrt[47] ), .B(new_n1861_), .Y(new_n2075_));
  OR2X1    g01883(.A(new_n2072_), .B(\a[96] ), .Y(new_n2076_));
  OR2X1    g01884(.A(new_n2076_), .B(new_n2075_), .Y(new_n2077_));
  AOI22X1  g01885(.A0(new_n2077_), .A1(new_n2074_), .B0(new_n2068_), .B1(new_n2054_), .Y(new_n2078_));
  OAI21X1  g01886(.A0(new_n2078_), .A1(new_n2055_), .B0(\asqrt[50] ), .Y(new_n2079_));
  NOR3X1   g01887(.A(new_n2078_), .B(new_n2055_), .C(\asqrt[50] ), .Y(new_n2080_));
  AOI21X1  g01888(.A0(new_n1862_), .A1(\asqrt[49] ), .B0(new_n1852_), .Y(new_n2081_));
  NAND3X1  g01889(.A(new_n2081_), .B(\asqrt[47] ), .C(new_n1848_), .Y(new_n2082_));
  INVX1    g01890(.A(new_n2081_), .Y(new_n2083_));
  OAI21X1  g01891(.A0(new_n2083_), .A1(new_n2040_), .B0(new_n1858_), .Y(new_n2084_));
  AND2X1   g01892(.A(new_n2084_), .B(new_n2082_), .Y(new_n2085_));
  OAI21X1  g01893(.A0(new_n2085_), .A1(new_n2080_), .B0(new_n2079_), .Y(new_n2086_));
  AND2X1   g01894(.A(new_n2086_), .B(\asqrt[51] ), .Y(new_n2087_));
  AND2X1   g01895(.A(new_n2067_), .B(\asqrt[48] ), .Y(new_n2088_));
  AOI21X1  g01896(.A0(\asqrt[47] ), .A1(\a[94] ), .B0(new_n2048_), .Y(new_n2089_));
  INVX1    g01897(.A(\a[95] ), .Y(new_n2090_));
  AOI21X1  g01898(.A0(\asqrt[47] ), .A1(new_n2045_), .B0(new_n2090_), .Y(new_n2091_));
  NOR3X1   g01899(.A(new_n2075_), .B(new_n2091_), .C(new_n2089_), .Y(new_n2092_));
  OAI21X1  g01900(.A0(new_n2092_), .A1(new_n2088_), .B0(\asqrt[49] ), .Y(new_n2093_));
  OAI21X1  g01901(.A0(new_n2043_), .A1(new_n1834_), .B0(new_n1632_), .Y(new_n2094_));
  OAI22X1  g01902(.A0(new_n2076_), .A1(new_n2075_), .B0(new_n2073_), .B1(new_n1855_), .Y(new_n2095_));
  OAI21X1  g01903(.A0(new_n2094_), .A1(new_n2092_), .B0(new_n2095_), .Y(new_n2096_));
  NAND3X1  g01904(.A(new_n2096_), .B(new_n2093_), .C(new_n1469_), .Y(new_n2097_));
  INVX1    g01905(.A(new_n2085_), .Y(new_n2098_));
  NAND2X1  g01906(.A(new_n2098_), .B(new_n2097_), .Y(new_n2099_));
  OAI21X1  g01907(.A0(new_n1908_), .A1(new_n1907_), .B0(new_n1871_), .Y(new_n2100_));
  NOR3X1   g01908(.A(new_n2100_), .B(new_n2040_), .C(new_n1854_), .Y(new_n2101_));
  OAI22X1  g01909(.A0(new_n1908_), .A1(new_n1907_), .B0(new_n1879_), .B1(new_n1469_), .Y(new_n2102_));
  OR2X1    g01910(.A(new_n2102_), .B(new_n2040_), .Y(new_n2103_));
  AOI21X1  g01911(.A0(new_n2103_), .A1(new_n1909_), .B0(new_n2101_), .Y(new_n2104_));
  AOI21X1  g01912(.A0(new_n2096_), .A1(new_n2093_), .B0(new_n1469_), .Y(new_n2105_));
  NOR2X1   g01913(.A(new_n2105_), .B(\asqrt[51] ), .Y(new_n2106_));
  AOI21X1  g01914(.A0(new_n2106_), .A1(new_n2099_), .B0(new_n2104_), .Y(new_n2107_));
  OAI21X1  g01915(.A0(new_n2107_), .A1(new_n2087_), .B0(\asqrt[52] ), .Y(new_n2108_));
  AND2X1   g01916(.A(new_n1912_), .B(new_n1910_), .Y(new_n2109_));
  NOR4X1   g01917(.A(new_n2040_), .B(new_n2109_), .C(new_n1878_), .D(new_n1911_), .Y(new_n2110_));
  OR2X1    g01918(.A(new_n2109_), .B(new_n1911_), .Y(new_n2111_));
  OR2X1    g01919(.A(new_n2111_), .B(new_n2040_), .Y(new_n2112_));
  AOI21X1  g01920(.A0(new_n2112_), .A1(new_n1878_), .B0(new_n2110_), .Y(new_n2113_));
  INVX1    g01921(.A(new_n2113_), .Y(new_n2114_));
  AOI21X1  g01922(.A0(new_n2098_), .A1(new_n2097_), .B0(new_n2105_), .Y(new_n2115_));
  OAI21X1  g01923(.A0(new_n2115_), .A1(new_n1277_), .B0(new_n1111_), .Y(new_n2116_));
  OAI21X1  g01924(.A0(new_n2116_), .A1(new_n2107_), .B0(new_n2114_), .Y(new_n2117_));
  AOI21X1  g01925(.A0(new_n2117_), .A1(new_n2108_), .B0(new_n968_), .Y(new_n2118_));
  NAND3X1  g01926(.A(new_n1889_), .B(new_n1887_), .C(new_n1914_), .Y(new_n2119_));
  NOR3X1   g01927(.A(new_n2040_), .B(new_n1915_), .C(new_n1882_), .Y(new_n2120_));
  OAI22X1  g01928(.A0(new_n2120_), .A1(new_n1887_), .B0(new_n2119_), .B1(new_n2040_), .Y(new_n2121_));
  NAND3X1  g01929(.A(new_n2117_), .B(new_n2108_), .C(new_n968_), .Y(new_n2122_));
  AOI21X1  g01930(.A0(new_n2122_), .A1(new_n2121_), .B0(new_n2118_), .Y(new_n2123_));
  OR2X1    g01931(.A(new_n2123_), .B(new_n902_), .Y(new_n2124_));
  AND2X1   g01932(.A(new_n2122_), .B(new_n2121_), .Y(new_n2125_));
  AND2X1   g01933(.A(new_n1931_), .B(new_n1930_), .Y(new_n2126_));
  NOR4X1   g01934(.A(new_n2040_), .B(new_n2126_), .C(new_n1898_), .D(new_n1929_), .Y(new_n2127_));
  AOI22X1  g01935(.A0(new_n1931_), .A1(new_n1930_), .B0(new_n1916_), .B1(\asqrt[53] ), .Y(new_n2128_));
  AOI21X1  g01936(.A0(new_n2128_), .A1(\asqrt[47] ), .B0(new_n1897_), .Y(new_n2129_));
  NOR2X1   g01937(.A(new_n2129_), .B(new_n2127_), .Y(new_n2130_));
  INVX1    g01938(.A(new_n2130_), .Y(new_n2131_));
  OR2X1    g01939(.A(new_n2118_), .B(\asqrt[54] ), .Y(new_n2132_));
  OAI21X1  g01940(.A0(new_n2132_), .A1(new_n2125_), .B0(new_n2131_), .Y(new_n2133_));
  AOI21X1  g01941(.A0(new_n2133_), .A1(new_n2124_), .B0(new_n697_), .Y(new_n2134_));
  AND2X1   g01942(.A(new_n1917_), .B(new_n1900_), .Y(new_n2135_));
  NOR4X1   g01943(.A(new_n2040_), .B(new_n2135_), .C(new_n1904_), .D(new_n1901_), .Y(new_n2136_));
  NOR2X1   g01944(.A(new_n2135_), .B(new_n1901_), .Y(new_n2137_));
  AOI21X1  g01945(.A0(new_n2137_), .A1(\asqrt[47] ), .B0(new_n1905_), .Y(new_n2138_));
  NOR2X1   g01946(.A(new_n2138_), .B(new_n2136_), .Y(new_n2139_));
  OR2X1    g01947(.A(new_n2115_), .B(new_n1277_), .Y(new_n2140_));
  AND2X1   g01948(.A(new_n2098_), .B(new_n2097_), .Y(new_n2141_));
  INVX1    g01949(.A(new_n2104_), .Y(new_n2142_));
  OR2X1    g01950(.A(new_n2105_), .B(\asqrt[51] ), .Y(new_n2143_));
  OAI21X1  g01951(.A0(new_n2143_), .A1(new_n2141_), .B0(new_n2142_), .Y(new_n2144_));
  AOI21X1  g01952(.A0(new_n2144_), .A1(new_n2140_), .B0(new_n1111_), .Y(new_n2145_));
  AOI21X1  g01953(.A0(new_n2086_), .A1(\asqrt[51] ), .B0(\asqrt[52] ), .Y(new_n2146_));
  AOI21X1  g01954(.A0(new_n2146_), .A1(new_n2144_), .B0(new_n2113_), .Y(new_n2147_));
  OAI21X1  g01955(.A0(new_n2147_), .A1(new_n2145_), .B0(\asqrt[53] ), .Y(new_n2148_));
  INVX1    g01956(.A(new_n2121_), .Y(new_n2149_));
  NOR3X1   g01957(.A(new_n2147_), .B(new_n2145_), .C(\asqrt[53] ), .Y(new_n2150_));
  OAI21X1  g01958(.A0(new_n2150_), .A1(new_n2149_), .B0(new_n2148_), .Y(new_n2151_));
  AOI21X1  g01959(.A0(new_n2151_), .A1(\asqrt[54] ), .B0(\asqrt[55] ), .Y(new_n2152_));
  AOI21X1  g01960(.A0(new_n2152_), .A1(new_n2133_), .B0(new_n2139_), .Y(new_n2153_));
  OAI21X1  g01961(.A0(new_n2153_), .A1(new_n2134_), .B0(\asqrt[56] ), .Y(new_n2154_));
  NAND3X1  g01962(.A(new_n1936_), .B(new_n1924_), .C(new_n1919_), .Y(new_n2155_));
  NOR3X1   g01963(.A(new_n2040_), .B(new_n1925_), .C(new_n1943_), .Y(new_n2156_));
  OAI22X1  g01964(.A0(new_n2156_), .A1(new_n1924_), .B0(new_n2155_), .B1(new_n2040_), .Y(new_n2157_));
  INVX1    g01965(.A(new_n2157_), .Y(new_n2158_));
  NOR3X1   g01966(.A(new_n2153_), .B(new_n2134_), .C(\asqrt[56] ), .Y(new_n2159_));
  OAI21X1  g01967(.A0(new_n2159_), .A1(new_n2158_), .B0(new_n2154_), .Y(new_n2160_));
  AND2X1   g01968(.A(new_n2160_), .B(\asqrt[57] ), .Y(new_n2161_));
  AND2X1   g01969(.A(new_n2151_), .B(\asqrt[54] ), .Y(new_n2162_));
  NAND2X1  g01970(.A(new_n2122_), .B(new_n2121_), .Y(new_n2163_));
  NOR2X1   g01971(.A(new_n2118_), .B(\asqrt[54] ), .Y(new_n2164_));
  AOI21X1  g01972(.A0(new_n2164_), .A1(new_n2163_), .B0(new_n2130_), .Y(new_n2165_));
  OAI21X1  g01973(.A0(new_n2165_), .A1(new_n2162_), .B0(\asqrt[55] ), .Y(new_n2166_));
  INVX1    g01974(.A(new_n2139_), .Y(new_n2167_));
  OAI21X1  g01975(.A0(new_n2123_), .A1(new_n902_), .B0(new_n697_), .Y(new_n2168_));
  OAI21X1  g01976(.A0(new_n2168_), .A1(new_n2165_), .B0(new_n2167_), .Y(new_n2169_));
  NAND3X1  g01977(.A(new_n2169_), .B(new_n2166_), .C(new_n582_), .Y(new_n2170_));
  NAND2X1  g01978(.A(new_n2170_), .B(new_n2157_), .Y(new_n2171_));
  OAI21X1  g01979(.A0(new_n1982_), .A1(new_n1980_), .B0(new_n1942_), .Y(new_n2172_));
  NOR3X1   g01980(.A(new_n2172_), .B(new_n2040_), .C(new_n1927_), .Y(new_n2173_));
  AOI22X1  g01981(.A0(new_n1944_), .A1(new_n1937_), .B0(new_n1926_), .B1(\asqrt[56] ), .Y(new_n2174_));
  AOI21X1  g01982(.A0(new_n2174_), .A1(\asqrt[47] ), .B0(new_n1942_), .Y(new_n2175_));
  NOR2X1   g01983(.A(new_n2175_), .B(new_n2173_), .Y(new_n2176_));
  AND2X1   g01984(.A(new_n2154_), .B(new_n481_), .Y(new_n2177_));
  AOI21X1  g01985(.A0(new_n2177_), .A1(new_n2171_), .B0(new_n2176_), .Y(new_n2178_));
  OAI21X1  g01986(.A0(new_n2178_), .A1(new_n2161_), .B0(\asqrt[58] ), .Y(new_n2179_));
  AND2X1   g01987(.A(new_n1985_), .B(new_n1983_), .Y(new_n2180_));
  NOR4X1   g01988(.A(new_n2040_), .B(new_n2180_), .C(new_n1951_), .D(new_n1984_), .Y(new_n2181_));
  NOR2X1   g01989(.A(new_n2180_), .B(new_n1984_), .Y(new_n2182_));
  AOI21X1  g01990(.A0(new_n2182_), .A1(\asqrt[47] ), .B0(new_n1950_), .Y(new_n2183_));
  NOR2X1   g01991(.A(new_n2183_), .B(new_n2181_), .Y(new_n2184_));
  INVX1    g01992(.A(new_n2184_), .Y(new_n2185_));
  AOI21X1  g01993(.A0(new_n2169_), .A1(new_n2166_), .B0(new_n582_), .Y(new_n2186_));
  AOI21X1  g01994(.A0(new_n2170_), .A1(new_n2157_), .B0(new_n2186_), .Y(new_n2187_));
  OAI21X1  g01995(.A0(new_n2187_), .A1(new_n481_), .B0(new_n399_), .Y(new_n2188_));
  OAI21X1  g01996(.A0(new_n2188_), .A1(new_n2178_), .B0(new_n2185_), .Y(new_n2189_));
  AOI21X1  g01997(.A0(new_n2189_), .A1(new_n2179_), .B0(new_n328_), .Y(new_n2190_));
  NAND3X1  g01998(.A(new_n1962_), .B(new_n1960_), .C(new_n1987_), .Y(new_n2191_));
  NOR3X1   g01999(.A(new_n2040_), .B(new_n1988_), .C(new_n1955_), .Y(new_n2192_));
  OAI22X1  g02000(.A0(new_n2192_), .A1(new_n1960_), .B0(new_n2191_), .B1(new_n2040_), .Y(new_n2193_));
  NAND3X1  g02001(.A(new_n2189_), .B(new_n2179_), .C(new_n328_), .Y(new_n2194_));
  AOI21X1  g02002(.A0(new_n2194_), .A1(new_n2193_), .B0(new_n2190_), .Y(new_n2195_));
  OR2X1    g02003(.A(new_n2195_), .B(new_n292_), .Y(new_n2196_));
  AND2X1   g02004(.A(new_n2194_), .B(new_n2193_), .Y(new_n2197_));
  AND2X1   g02005(.A(new_n2004_), .B(new_n2003_), .Y(new_n2198_));
  NOR4X1   g02006(.A(new_n2040_), .B(new_n2198_), .C(new_n1971_), .D(new_n2002_), .Y(new_n2199_));
  AOI22X1  g02007(.A0(new_n2004_), .A1(new_n2003_), .B0(new_n1989_), .B1(\asqrt[59] ), .Y(new_n2200_));
  AOI21X1  g02008(.A0(new_n2200_), .A1(\asqrt[47] ), .B0(new_n1970_), .Y(new_n2201_));
  NOR2X1   g02009(.A(new_n2201_), .B(new_n2199_), .Y(new_n2202_));
  INVX1    g02010(.A(new_n2202_), .Y(new_n2203_));
  OR2X1    g02011(.A(new_n2187_), .B(new_n481_), .Y(new_n2204_));
  AND2X1   g02012(.A(new_n2170_), .B(new_n2157_), .Y(new_n2205_));
  INVX1    g02013(.A(new_n2176_), .Y(new_n2206_));
  NAND2X1  g02014(.A(new_n2154_), .B(new_n481_), .Y(new_n2207_));
  OAI21X1  g02015(.A0(new_n2207_), .A1(new_n2205_), .B0(new_n2206_), .Y(new_n2208_));
  AOI21X1  g02016(.A0(new_n2208_), .A1(new_n2204_), .B0(new_n399_), .Y(new_n2209_));
  AOI21X1  g02017(.A0(new_n2160_), .A1(\asqrt[57] ), .B0(\asqrt[58] ), .Y(new_n2210_));
  AOI21X1  g02018(.A0(new_n2210_), .A1(new_n2208_), .B0(new_n2184_), .Y(new_n2211_));
  OAI21X1  g02019(.A0(new_n2211_), .A1(new_n2209_), .B0(\asqrt[59] ), .Y(new_n2212_));
  NAND2X1  g02020(.A(new_n2212_), .B(new_n292_), .Y(new_n2213_));
  OAI21X1  g02021(.A0(new_n2213_), .A1(new_n2197_), .B0(new_n2203_), .Y(new_n2214_));
  AOI21X1  g02022(.A0(new_n2214_), .A1(new_n2196_), .B0(new_n217_), .Y(new_n2215_));
  AND2X1   g02023(.A(new_n1990_), .B(new_n1973_), .Y(new_n2216_));
  NOR4X1   g02024(.A(new_n2040_), .B(new_n2216_), .C(new_n2007_), .D(new_n1974_), .Y(new_n2217_));
  NOR2X1   g02025(.A(new_n2216_), .B(new_n1974_), .Y(new_n2218_));
  AOI21X1  g02026(.A0(new_n2218_), .A1(\asqrt[47] ), .B0(new_n1978_), .Y(new_n2219_));
  NOR2X1   g02027(.A(new_n2219_), .B(new_n2217_), .Y(new_n2220_));
  INVX1    g02028(.A(new_n2193_), .Y(new_n2221_));
  NOR3X1   g02029(.A(new_n2211_), .B(new_n2209_), .C(\asqrt[59] ), .Y(new_n2222_));
  OAI21X1  g02030(.A0(new_n2222_), .A1(new_n2221_), .B0(new_n2212_), .Y(new_n2223_));
  AOI21X1  g02031(.A0(new_n2223_), .A1(\asqrt[60] ), .B0(\asqrt[61] ), .Y(new_n2224_));
  AOI21X1  g02032(.A0(new_n2224_), .A1(new_n2214_), .B0(new_n2220_), .Y(new_n2225_));
  OAI21X1  g02033(.A0(new_n2225_), .A1(new_n2215_), .B0(\asqrt[62] ), .Y(new_n2226_));
  NAND3X1  g02034(.A(new_n2010_), .B(new_n1997_), .C(new_n1992_), .Y(new_n2227_));
  NOR3X1   g02035(.A(new_n2040_), .B(new_n1998_), .C(new_n2017_), .Y(new_n2228_));
  OAI22X1  g02036(.A0(new_n2228_), .A1(new_n1997_), .B0(new_n2227_), .B1(new_n2040_), .Y(new_n2229_));
  INVX1    g02037(.A(new_n2229_), .Y(new_n2230_));
  NOR3X1   g02038(.A(new_n2225_), .B(new_n2215_), .C(\asqrt[62] ), .Y(new_n2231_));
  OAI21X1  g02039(.A0(new_n2231_), .A1(new_n2230_), .B0(new_n2226_), .Y(new_n2232_));
  OAI21X1  g02040(.A0(new_n2059_), .A1(new_n2057_), .B0(new_n2016_), .Y(new_n2233_));
  NOR3X1   g02041(.A(new_n2233_), .B(new_n2040_), .C(new_n2000_), .Y(new_n2234_));
  AOI22X1  g02042(.A0(new_n2018_), .A1(new_n2011_), .B0(new_n1999_), .B1(\asqrt[62] ), .Y(new_n2235_));
  AOI21X1  g02043(.A0(new_n2235_), .A1(\asqrt[47] ), .B0(new_n2016_), .Y(new_n2236_));
  NOR2X1   g02044(.A(new_n2236_), .B(new_n2234_), .Y(new_n2237_));
  INVX1    g02045(.A(new_n2237_), .Y(new_n2238_));
  AND2X1   g02046(.A(new_n2063_), .B(new_n2060_), .Y(new_n2239_));
  AOI21X1  g02047(.A0(new_n2060_), .A1(new_n2056_), .B0(new_n2023_), .Y(new_n2240_));
  AOI21X1  g02048(.A0(new_n2240_), .A1(\asqrt[47] ), .B0(new_n2239_), .Y(new_n2241_));
  AND2X1   g02049(.A(new_n2241_), .B(new_n2238_), .Y(new_n2242_));
  AOI21X1  g02050(.A0(new_n2242_), .A1(new_n2232_), .B0(\asqrt[63] ), .Y(new_n2243_));
  AND2X1   g02051(.A(new_n2223_), .B(\asqrt[60] ), .Y(new_n2244_));
  NAND2X1  g02052(.A(new_n2194_), .B(new_n2193_), .Y(new_n2245_));
  AND2X1   g02053(.A(new_n2212_), .B(new_n292_), .Y(new_n2246_));
  AOI21X1  g02054(.A0(new_n2246_), .A1(new_n2245_), .B0(new_n2202_), .Y(new_n2247_));
  OAI21X1  g02055(.A0(new_n2247_), .A1(new_n2244_), .B0(\asqrt[61] ), .Y(new_n2248_));
  INVX1    g02056(.A(new_n2220_), .Y(new_n2249_));
  OAI21X1  g02057(.A0(new_n2195_), .A1(new_n292_), .B0(new_n217_), .Y(new_n2250_));
  OAI21X1  g02058(.A0(new_n2250_), .A1(new_n2247_), .B0(new_n2249_), .Y(new_n2251_));
  NAND3X1  g02059(.A(new_n2251_), .B(new_n2248_), .C(new_n199_), .Y(new_n2252_));
  AND2X1   g02060(.A(new_n2252_), .B(new_n2229_), .Y(new_n2253_));
  NAND2X1  g02061(.A(new_n2237_), .B(new_n2226_), .Y(new_n2254_));
  NAND2X1  g02062(.A(new_n2060_), .B(new_n2056_), .Y(new_n2255_));
  AOI21X1  g02063(.A0(\asqrt[47] ), .A1(new_n2024_), .B0(new_n2255_), .Y(new_n2256_));
  NOR3X1   g02064(.A(new_n2256_), .B(new_n2240_), .C(new_n193_), .Y(new_n2257_));
  AND2X1   g02065(.A(new_n2028_), .B(new_n193_), .Y(new_n2258_));
  NAND4X1  g02066(.A(new_n2037_), .B(new_n2033_), .C(new_n2022_), .D(new_n2020_), .Y(new_n2259_));
  NOR3X1   g02067(.A(new_n2259_), .B(new_n2239_), .C(new_n2258_), .Y(new_n2260_));
  NOR2X1   g02068(.A(new_n2260_), .B(new_n2257_), .Y(new_n2261_));
  OAI21X1  g02069(.A0(new_n2254_), .A1(new_n2253_), .B0(new_n2261_), .Y(new_n2262_));
  NOR2X1   g02070(.A(new_n2262_), .B(new_n2243_), .Y(new_n2263_));
  INVX1    g02071(.A(new_n2263_), .Y(\asqrt[46] ));
  INVX1    g02072(.A(\a[92] ), .Y(new_n2265_));
  NOR2X1   g02073(.A(\a[91] ), .B(\a[90] ), .Y(new_n2266_));
  NAND2X1  g02074(.A(new_n2266_), .B(new_n2265_), .Y(new_n2267_));
  OAI21X1  g02075(.A0(new_n2263_), .A1(new_n2265_), .B0(new_n2267_), .Y(new_n2268_));
  AOI21X1  g02076(.A0(new_n2251_), .A1(new_n2248_), .B0(new_n199_), .Y(new_n2269_));
  AOI21X1  g02077(.A0(new_n2252_), .A1(new_n2229_), .B0(new_n2269_), .Y(new_n2270_));
  INVX1    g02078(.A(new_n2242_), .Y(new_n2271_));
  OAI21X1  g02079(.A0(new_n2271_), .A1(new_n2270_), .B0(new_n193_), .Y(new_n2272_));
  NAND2X1  g02080(.A(new_n2252_), .B(new_n2229_), .Y(new_n2273_));
  AND2X1   g02081(.A(new_n2237_), .B(new_n2226_), .Y(new_n2274_));
  INVX1    g02082(.A(new_n2261_), .Y(new_n2275_));
  AOI21X1  g02083(.A0(new_n2274_), .A1(new_n2273_), .B0(new_n2275_), .Y(new_n2276_));
  AOI21X1  g02084(.A0(new_n2276_), .A1(new_n2272_), .B0(new_n2265_), .Y(new_n2277_));
  NAND3X1  g02085(.A(new_n2267_), .B(new_n2037_), .C(new_n2033_), .Y(new_n2278_));
  OR4X1    g02086(.A(new_n2278_), .B(new_n2277_), .C(new_n2239_), .D(new_n2258_), .Y(new_n2279_));
  OAI21X1  g02087(.A0(new_n2262_), .A1(new_n2243_), .B0(new_n2265_), .Y(new_n2280_));
  AOI21X1  g02088(.A0(new_n2276_), .A1(new_n2272_), .B0(new_n2042_), .Y(new_n2281_));
  AOI21X1  g02089(.A0(new_n2280_), .A1(\a[93] ), .B0(new_n2281_), .Y(new_n2282_));
  AOI22X1  g02090(.A0(new_n2282_), .A1(new_n2279_), .B0(new_n2268_), .B1(\asqrt[47] ), .Y(new_n2283_));
  OR2X1    g02091(.A(new_n2283_), .B(new_n1834_), .Y(new_n2284_));
  AND2X1   g02092(.A(new_n2282_), .B(new_n2279_), .Y(new_n2285_));
  INVX1    g02093(.A(new_n2266_), .Y(new_n2286_));
  MX2X1    g02094(.A(new_n2286_), .B(new_n2263_), .S0(\a[92] ), .Y(new_n2287_));
  OAI21X1  g02095(.A0(new_n2287_), .A1(new_n2040_), .B0(new_n1834_), .Y(new_n2288_));
  OAI21X1  g02096(.A0(new_n2262_), .A1(new_n2243_), .B0(new_n2041_), .Y(new_n2289_));
  AND2X1   g02097(.A(new_n2274_), .B(new_n2273_), .Y(new_n2290_));
  OR2X1    g02098(.A(new_n2260_), .B(new_n2040_), .Y(new_n2291_));
  OR4X1    g02099(.A(new_n2291_), .B(new_n2257_), .C(new_n2290_), .D(new_n2243_), .Y(new_n2292_));
  AOI21X1  g02100(.A0(new_n2292_), .A1(new_n2289_), .B0(new_n2045_), .Y(new_n2293_));
  NOR4X1   g02101(.A(new_n2291_), .B(new_n2257_), .C(new_n2290_), .D(new_n2243_), .Y(new_n2294_));
  NOR3X1   g02102(.A(new_n2294_), .B(new_n2281_), .C(\a[94] ), .Y(new_n2295_));
  OR2X1    g02103(.A(new_n2295_), .B(new_n2293_), .Y(new_n2296_));
  OAI21X1  g02104(.A0(new_n2288_), .A1(new_n2285_), .B0(new_n2296_), .Y(new_n2297_));
  AOI21X1  g02105(.A0(new_n2297_), .A1(new_n2284_), .B0(new_n1632_), .Y(new_n2298_));
  AND2X1   g02106(.A(new_n2053_), .B(new_n2051_), .Y(new_n2299_));
  NOR3X1   g02107(.A(new_n2299_), .B(new_n2089_), .C(new_n2088_), .Y(new_n2300_));
  OAI21X1  g02108(.A0(new_n2262_), .A1(new_n2243_), .B0(new_n2300_), .Y(new_n2301_));
  AOI21X1  g02109(.A0(new_n2067_), .A1(\asqrt[48] ), .B0(new_n2089_), .Y(new_n2302_));
  OAI21X1  g02110(.A0(new_n2262_), .A1(new_n2243_), .B0(new_n2302_), .Y(new_n2303_));
  NAND2X1  g02111(.A(new_n2303_), .B(new_n2299_), .Y(new_n2304_));
  NOR4X1   g02112(.A(new_n2278_), .B(new_n2277_), .C(new_n2239_), .D(new_n2258_), .Y(new_n2305_));
  INVX1    g02113(.A(\a[93] ), .Y(new_n2306_));
  AOI21X1  g02114(.A0(new_n2276_), .A1(new_n2272_), .B0(\a[92] ), .Y(new_n2307_));
  OAI21X1  g02115(.A0(new_n2307_), .A1(new_n2306_), .B0(new_n2289_), .Y(new_n2308_));
  OAI22X1  g02116(.A0(new_n2308_), .A1(new_n2305_), .B0(new_n2287_), .B1(new_n2040_), .Y(new_n2309_));
  AOI21X1  g02117(.A0(new_n2309_), .A1(\asqrt[48] ), .B0(\asqrt[49] ), .Y(new_n2310_));
  AOI22X1  g02118(.A0(new_n2310_), .A1(new_n2297_), .B0(new_n2304_), .B1(new_n2301_), .Y(new_n2311_));
  OAI21X1  g02119(.A0(new_n2311_), .A1(new_n2298_), .B0(\asqrt[50] ), .Y(new_n2312_));
  AND2X1   g02120(.A(new_n2068_), .B(new_n2054_), .Y(new_n2313_));
  NOR3X1   g02121(.A(new_n2095_), .B(new_n2313_), .C(new_n2055_), .Y(new_n2314_));
  OAI21X1  g02122(.A0(new_n2262_), .A1(new_n2243_), .B0(new_n2314_), .Y(new_n2315_));
  NOR2X1   g02123(.A(new_n2313_), .B(new_n2055_), .Y(new_n2316_));
  OAI21X1  g02124(.A0(new_n2262_), .A1(new_n2243_), .B0(new_n2316_), .Y(new_n2317_));
  NAND2X1  g02125(.A(new_n2317_), .B(new_n2095_), .Y(new_n2318_));
  AND2X1   g02126(.A(new_n2318_), .B(new_n2315_), .Y(new_n2319_));
  NOR3X1   g02127(.A(new_n2311_), .B(new_n2298_), .C(\asqrt[50] ), .Y(new_n2320_));
  OAI21X1  g02128(.A0(new_n2320_), .A1(new_n2319_), .B0(new_n2312_), .Y(new_n2321_));
  AND2X1   g02129(.A(new_n2321_), .B(\asqrt[51] ), .Y(new_n2322_));
  OR2X1    g02130(.A(new_n2320_), .B(new_n2319_), .Y(new_n2323_));
  AND2X1   g02131(.A(new_n2309_), .B(\asqrt[48] ), .Y(new_n2324_));
  NAND2X1  g02132(.A(new_n2282_), .B(new_n2279_), .Y(new_n2325_));
  AOI21X1  g02133(.A0(new_n2268_), .A1(\asqrt[47] ), .B0(\asqrt[48] ), .Y(new_n2326_));
  NOR2X1   g02134(.A(new_n2295_), .B(new_n2293_), .Y(new_n2327_));
  AOI21X1  g02135(.A0(new_n2326_), .A1(new_n2325_), .B0(new_n2327_), .Y(new_n2328_));
  OAI21X1  g02136(.A0(new_n2328_), .A1(new_n2324_), .B0(\asqrt[49] ), .Y(new_n2329_));
  NAND2X1  g02137(.A(new_n2304_), .B(new_n2301_), .Y(new_n2330_));
  OAI21X1  g02138(.A0(new_n2283_), .A1(new_n1834_), .B0(new_n1632_), .Y(new_n2331_));
  OAI21X1  g02139(.A0(new_n2331_), .A1(new_n2328_), .B0(new_n2330_), .Y(new_n2332_));
  AOI21X1  g02140(.A0(new_n2332_), .A1(new_n2329_), .B0(new_n1469_), .Y(new_n2333_));
  NOR2X1   g02141(.A(new_n2333_), .B(\asqrt[51] ), .Y(new_n2334_));
  NOR3X1   g02142(.A(new_n2098_), .B(new_n2080_), .C(new_n2105_), .Y(new_n2335_));
  OAI21X1  g02143(.A0(new_n2262_), .A1(new_n2243_), .B0(new_n2335_), .Y(new_n2336_));
  NOR3X1   g02144(.A(new_n2263_), .B(new_n2080_), .C(new_n2105_), .Y(new_n2337_));
  OR2X1    g02145(.A(new_n2337_), .B(new_n2085_), .Y(new_n2338_));
  AND2X1   g02146(.A(new_n2338_), .B(new_n2336_), .Y(new_n2339_));
  AOI21X1  g02147(.A0(new_n2334_), .A1(new_n2323_), .B0(new_n2339_), .Y(new_n2340_));
  OAI21X1  g02148(.A0(new_n2340_), .A1(new_n2322_), .B0(\asqrt[52] ), .Y(new_n2341_));
  AOI21X1  g02149(.A0(new_n2106_), .A1(new_n2099_), .B0(new_n2142_), .Y(new_n2342_));
  AND2X1   g02150(.A(new_n2342_), .B(new_n2140_), .Y(new_n2343_));
  AOI22X1  g02151(.A0(new_n2106_), .A1(new_n2099_), .B0(new_n2086_), .B1(\asqrt[51] ), .Y(new_n2344_));
  AOI21X1  g02152(.A0(new_n2344_), .A1(\asqrt[46] ), .B0(new_n2104_), .Y(new_n2345_));
  AOI21X1  g02153(.A0(new_n2343_), .A1(\asqrt[46] ), .B0(new_n2345_), .Y(new_n2346_));
  INVX1    g02154(.A(new_n2346_), .Y(new_n2347_));
  INVX1    g02155(.A(new_n2319_), .Y(new_n2348_));
  NAND3X1  g02156(.A(new_n2332_), .B(new_n2329_), .C(new_n1469_), .Y(new_n2349_));
  AOI21X1  g02157(.A0(new_n2349_), .A1(new_n2348_), .B0(new_n2333_), .Y(new_n2350_));
  OAI21X1  g02158(.A0(new_n2350_), .A1(new_n1277_), .B0(new_n1111_), .Y(new_n2351_));
  OAI21X1  g02159(.A0(new_n2351_), .A1(new_n2340_), .B0(new_n2347_), .Y(new_n2352_));
  AOI21X1  g02160(.A0(new_n2352_), .A1(new_n2341_), .B0(new_n968_), .Y(new_n2353_));
  AND2X1   g02161(.A(new_n2146_), .B(new_n2144_), .Y(new_n2354_));
  NOR3X1   g02162(.A(new_n2354_), .B(new_n2114_), .C(new_n2145_), .Y(new_n2355_));
  NOR3X1   g02163(.A(new_n2263_), .B(new_n2354_), .C(new_n2145_), .Y(new_n2356_));
  NOR2X1   g02164(.A(new_n2356_), .B(new_n2113_), .Y(new_n2357_));
  AOI21X1  g02165(.A0(new_n2355_), .A1(\asqrt[46] ), .B0(new_n2357_), .Y(new_n2358_));
  INVX1    g02166(.A(new_n2358_), .Y(new_n2359_));
  NAND3X1  g02167(.A(new_n2352_), .B(new_n2341_), .C(new_n968_), .Y(new_n2360_));
  AOI21X1  g02168(.A0(new_n2360_), .A1(new_n2359_), .B0(new_n2353_), .Y(new_n2361_));
  OR2X1    g02169(.A(new_n2361_), .B(new_n902_), .Y(new_n2362_));
  AND2X1   g02170(.A(new_n2360_), .B(new_n2359_), .Y(new_n2363_));
  OR4X1    g02171(.A(new_n2263_), .B(new_n2150_), .C(new_n2121_), .D(new_n2118_), .Y(new_n2364_));
  NAND2X1  g02172(.A(new_n2122_), .B(new_n2148_), .Y(new_n2365_));
  OAI21X1  g02173(.A0(new_n2365_), .A1(new_n2263_), .B0(new_n2121_), .Y(new_n2366_));
  AND2X1   g02174(.A(new_n2366_), .B(new_n2364_), .Y(new_n2367_));
  INVX1    g02175(.A(new_n2367_), .Y(new_n2368_));
  OR2X1    g02176(.A(new_n2350_), .B(new_n1277_), .Y(new_n2369_));
  NOR2X1   g02177(.A(new_n2320_), .B(new_n2319_), .Y(new_n2370_));
  OR2X1    g02178(.A(new_n2333_), .B(\asqrt[51] ), .Y(new_n2371_));
  INVX1    g02179(.A(new_n2339_), .Y(new_n2372_));
  OAI21X1  g02180(.A0(new_n2371_), .A1(new_n2370_), .B0(new_n2372_), .Y(new_n2373_));
  AOI21X1  g02181(.A0(new_n2373_), .A1(new_n2369_), .B0(new_n1111_), .Y(new_n2374_));
  AOI21X1  g02182(.A0(new_n2321_), .A1(\asqrt[51] ), .B0(\asqrt[52] ), .Y(new_n2375_));
  AOI21X1  g02183(.A0(new_n2375_), .A1(new_n2373_), .B0(new_n2346_), .Y(new_n2376_));
  OAI21X1  g02184(.A0(new_n2376_), .A1(new_n2374_), .B0(\asqrt[53] ), .Y(new_n2377_));
  NAND2X1  g02185(.A(new_n2377_), .B(new_n902_), .Y(new_n2378_));
  OAI21X1  g02186(.A0(new_n2378_), .A1(new_n2363_), .B0(new_n2368_), .Y(new_n2379_));
  AOI21X1  g02187(.A0(new_n2379_), .A1(new_n2362_), .B0(new_n697_), .Y(new_n2380_));
  AND2X1   g02188(.A(new_n2164_), .B(new_n2163_), .Y(new_n2381_));
  NOR3X1   g02189(.A(new_n2381_), .B(new_n2131_), .C(new_n2162_), .Y(new_n2382_));
  NOR3X1   g02190(.A(new_n2263_), .B(new_n2381_), .C(new_n2162_), .Y(new_n2383_));
  NOR2X1   g02191(.A(new_n2383_), .B(new_n2130_), .Y(new_n2384_));
  AOI21X1  g02192(.A0(new_n2382_), .A1(\asqrt[46] ), .B0(new_n2384_), .Y(new_n2385_));
  NOR3X1   g02193(.A(new_n2376_), .B(new_n2374_), .C(\asqrt[53] ), .Y(new_n2386_));
  OAI21X1  g02194(.A0(new_n2386_), .A1(new_n2358_), .B0(new_n2377_), .Y(new_n2387_));
  AOI21X1  g02195(.A0(new_n2387_), .A1(\asqrt[54] ), .B0(\asqrt[55] ), .Y(new_n2388_));
  AOI21X1  g02196(.A0(new_n2388_), .A1(new_n2379_), .B0(new_n2385_), .Y(new_n2389_));
  OAI21X1  g02197(.A0(new_n2389_), .A1(new_n2380_), .B0(\asqrt[56] ), .Y(new_n2390_));
  AND2X1   g02198(.A(new_n2152_), .B(new_n2133_), .Y(new_n2391_));
  NOR3X1   g02199(.A(new_n2391_), .B(new_n2167_), .C(new_n2134_), .Y(new_n2392_));
  NOR3X1   g02200(.A(new_n2263_), .B(new_n2391_), .C(new_n2134_), .Y(new_n2393_));
  NOR2X1   g02201(.A(new_n2393_), .B(new_n2139_), .Y(new_n2394_));
  AOI21X1  g02202(.A0(new_n2392_), .A1(\asqrt[46] ), .B0(new_n2394_), .Y(new_n2395_));
  NOR3X1   g02203(.A(new_n2389_), .B(new_n2380_), .C(\asqrt[56] ), .Y(new_n2396_));
  OAI21X1  g02204(.A0(new_n2396_), .A1(new_n2395_), .B0(new_n2390_), .Y(new_n2397_));
  AND2X1   g02205(.A(new_n2397_), .B(\asqrt[57] ), .Y(new_n2398_));
  INVX1    g02206(.A(new_n2395_), .Y(new_n2399_));
  AND2X1   g02207(.A(new_n2387_), .B(\asqrt[54] ), .Y(new_n2400_));
  OR2X1    g02208(.A(new_n2386_), .B(new_n2358_), .Y(new_n2401_));
  AND2X1   g02209(.A(new_n2377_), .B(new_n902_), .Y(new_n2402_));
  AOI21X1  g02210(.A0(new_n2402_), .A1(new_n2401_), .B0(new_n2367_), .Y(new_n2403_));
  OAI21X1  g02211(.A0(new_n2403_), .A1(new_n2400_), .B0(\asqrt[55] ), .Y(new_n2404_));
  INVX1    g02212(.A(new_n2385_), .Y(new_n2405_));
  OAI21X1  g02213(.A0(new_n2361_), .A1(new_n902_), .B0(new_n697_), .Y(new_n2406_));
  OAI21X1  g02214(.A0(new_n2406_), .A1(new_n2403_), .B0(new_n2405_), .Y(new_n2407_));
  NAND3X1  g02215(.A(new_n2407_), .B(new_n2404_), .C(new_n582_), .Y(new_n2408_));
  NAND2X1  g02216(.A(new_n2408_), .B(new_n2399_), .Y(new_n2409_));
  OR4X1    g02217(.A(new_n2263_), .B(new_n2159_), .C(new_n2157_), .D(new_n2186_), .Y(new_n2410_));
  OR2X1    g02218(.A(new_n2159_), .B(new_n2186_), .Y(new_n2411_));
  OAI21X1  g02219(.A0(new_n2411_), .A1(new_n2263_), .B0(new_n2157_), .Y(new_n2412_));
  AND2X1   g02220(.A(new_n2412_), .B(new_n2410_), .Y(new_n2413_));
  AOI21X1  g02221(.A0(new_n2407_), .A1(new_n2404_), .B0(new_n582_), .Y(new_n2414_));
  NOR2X1   g02222(.A(new_n2414_), .B(\asqrt[57] ), .Y(new_n2415_));
  AOI21X1  g02223(.A0(new_n2415_), .A1(new_n2409_), .B0(new_n2413_), .Y(new_n2416_));
  OAI21X1  g02224(.A0(new_n2416_), .A1(new_n2398_), .B0(\asqrt[58] ), .Y(new_n2417_));
  AOI21X1  g02225(.A0(new_n2177_), .A1(new_n2171_), .B0(new_n2206_), .Y(new_n2418_));
  AND2X1   g02226(.A(new_n2418_), .B(new_n2204_), .Y(new_n2419_));
  AOI22X1  g02227(.A0(new_n2177_), .A1(new_n2171_), .B0(new_n2160_), .B1(\asqrt[57] ), .Y(new_n2420_));
  AOI21X1  g02228(.A0(new_n2420_), .A1(\asqrt[46] ), .B0(new_n2176_), .Y(new_n2421_));
  AOI21X1  g02229(.A0(new_n2419_), .A1(\asqrt[46] ), .B0(new_n2421_), .Y(new_n2422_));
  INVX1    g02230(.A(new_n2422_), .Y(new_n2423_));
  AOI21X1  g02231(.A0(new_n2408_), .A1(new_n2399_), .B0(new_n2414_), .Y(new_n2424_));
  OAI21X1  g02232(.A0(new_n2424_), .A1(new_n481_), .B0(new_n399_), .Y(new_n2425_));
  OAI21X1  g02233(.A0(new_n2425_), .A1(new_n2416_), .B0(new_n2423_), .Y(new_n2426_));
  AOI21X1  g02234(.A0(new_n2426_), .A1(new_n2417_), .B0(new_n328_), .Y(new_n2427_));
  AND2X1   g02235(.A(new_n2210_), .B(new_n2208_), .Y(new_n2428_));
  NOR3X1   g02236(.A(new_n2428_), .B(new_n2185_), .C(new_n2209_), .Y(new_n2429_));
  NOR3X1   g02237(.A(new_n2263_), .B(new_n2428_), .C(new_n2209_), .Y(new_n2430_));
  NOR2X1   g02238(.A(new_n2430_), .B(new_n2184_), .Y(new_n2431_));
  AOI21X1  g02239(.A0(new_n2429_), .A1(\asqrt[46] ), .B0(new_n2431_), .Y(new_n2432_));
  INVX1    g02240(.A(new_n2432_), .Y(new_n2433_));
  NAND3X1  g02241(.A(new_n2426_), .B(new_n2417_), .C(new_n328_), .Y(new_n2434_));
  AOI21X1  g02242(.A0(new_n2434_), .A1(new_n2433_), .B0(new_n2427_), .Y(new_n2435_));
  OR2X1    g02243(.A(new_n2435_), .B(new_n292_), .Y(new_n2436_));
  AND2X1   g02244(.A(new_n2434_), .B(new_n2433_), .Y(new_n2437_));
  OR4X1    g02245(.A(new_n2263_), .B(new_n2222_), .C(new_n2193_), .D(new_n2190_), .Y(new_n2438_));
  OR2X1    g02246(.A(new_n2222_), .B(new_n2190_), .Y(new_n2439_));
  OAI21X1  g02247(.A0(new_n2439_), .A1(new_n2263_), .B0(new_n2193_), .Y(new_n2440_));
  AND2X1   g02248(.A(new_n2440_), .B(new_n2438_), .Y(new_n2441_));
  INVX1    g02249(.A(new_n2441_), .Y(new_n2442_));
  OR2X1    g02250(.A(new_n2427_), .B(\asqrt[60] ), .Y(new_n2443_));
  OAI21X1  g02251(.A0(new_n2443_), .A1(new_n2437_), .B0(new_n2442_), .Y(new_n2444_));
  AOI21X1  g02252(.A0(new_n2444_), .A1(new_n2436_), .B0(new_n217_), .Y(new_n2445_));
  AND2X1   g02253(.A(new_n2246_), .B(new_n2245_), .Y(new_n2446_));
  NOR3X1   g02254(.A(new_n2446_), .B(new_n2203_), .C(new_n2244_), .Y(new_n2447_));
  NOR3X1   g02255(.A(new_n2263_), .B(new_n2446_), .C(new_n2244_), .Y(new_n2448_));
  NOR2X1   g02256(.A(new_n2448_), .B(new_n2202_), .Y(new_n2449_));
  AOI21X1  g02257(.A0(new_n2447_), .A1(\asqrt[46] ), .B0(new_n2449_), .Y(new_n2450_));
  OR2X1    g02258(.A(new_n2424_), .B(new_n481_), .Y(new_n2451_));
  AND2X1   g02259(.A(new_n2408_), .B(new_n2399_), .Y(new_n2452_));
  INVX1    g02260(.A(new_n2413_), .Y(new_n2453_));
  OR2X1    g02261(.A(new_n2414_), .B(\asqrt[57] ), .Y(new_n2454_));
  OAI21X1  g02262(.A0(new_n2454_), .A1(new_n2452_), .B0(new_n2453_), .Y(new_n2455_));
  AOI21X1  g02263(.A0(new_n2455_), .A1(new_n2451_), .B0(new_n399_), .Y(new_n2456_));
  AOI21X1  g02264(.A0(new_n2397_), .A1(\asqrt[57] ), .B0(\asqrt[58] ), .Y(new_n2457_));
  AOI21X1  g02265(.A0(new_n2457_), .A1(new_n2455_), .B0(new_n2422_), .Y(new_n2458_));
  OAI21X1  g02266(.A0(new_n2458_), .A1(new_n2456_), .B0(\asqrt[59] ), .Y(new_n2459_));
  NOR3X1   g02267(.A(new_n2458_), .B(new_n2456_), .C(\asqrt[59] ), .Y(new_n2460_));
  OAI21X1  g02268(.A0(new_n2460_), .A1(new_n2432_), .B0(new_n2459_), .Y(new_n2461_));
  AOI21X1  g02269(.A0(new_n2461_), .A1(\asqrt[60] ), .B0(\asqrt[61] ), .Y(new_n2462_));
  AOI21X1  g02270(.A0(new_n2462_), .A1(new_n2444_), .B0(new_n2450_), .Y(new_n2463_));
  OAI21X1  g02271(.A0(new_n2463_), .A1(new_n2445_), .B0(\asqrt[62] ), .Y(new_n2464_));
  AND2X1   g02272(.A(new_n2224_), .B(new_n2214_), .Y(new_n2465_));
  NOR3X1   g02273(.A(new_n2465_), .B(new_n2249_), .C(new_n2215_), .Y(new_n2466_));
  NOR3X1   g02274(.A(new_n2263_), .B(new_n2465_), .C(new_n2215_), .Y(new_n2467_));
  NOR2X1   g02275(.A(new_n2467_), .B(new_n2220_), .Y(new_n2468_));
  AOI21X1  g02276(.A0(new_n2466_), .A1(\asqrt[46] ), .B0(new_n2468_), .Y(new_n2469_));
  NOR3X1   g02277(.A(new_n2463_), .B(new_n2445_), .C(\asqrt[62] ), .Y(new_n2470_));
  OAI21X1  g02278(.A0(new_n2470_), .A1(new_n2469_), .B0(new_n2464_), .Y(new_n2471_));
  NOR4X1   g02279(.A(new_n2263_), .B(new_n2231_), .C(new_n2229_), .D(new_n2269_), .Y(new_n2472_));
  NAND3X1  g02280(.A(\asqrt[46] ), .B(new_n2252_), .C(new_n2226_), .Y(new_n2473_));
  AOI21X1  g02281(.A0(new_n2473_), .A1(new_n2229_), .B0(new_n2472_), .Y(new_n2474_));
  INVX1    g02282(.A(new_n2474_), .Y(new_n2475_));
  NOR2X1   g02283(.A(new_n2237_), .B(new_n2270_), .Y(new_n2476_));
  AOI21X1  g02284(.A0(new_n2476_), .A1(\asqrt[46] ), .B0(new_n2290_), .Y(new_n2477_));
  AND2X1   g02285(.A(new_n2477_), .B(new_n2475_), .Y(new_n2478_));
  AOI21X1  g02286(.A0(new_n2478_), .A1(new_n2471_), .B0(\asqrt[63] ), .Y(new_n2479_));
  INVX1    g02287(.A(new_n2469_), .Y(new_n2480_));
  AND2X1   g02288(.A(new_n2461_), .B(\asqrt[60] ), .Y(new_n2481_));
  NAND2X1  g02289(.A(new_n2434_), .B(new_n2433_), .Y(new_n2482_));
  NOR2X1   g02290(.A(new_n2427_), .B(\asqrt[60] ), .Y(new_n2483_));
  AOI21X1  g02291(.A0(new_n2483_), .A1(new_n2482_), .B0(new_n2441_), .Y(new_n2484_));
  OAI21X1  g02292(.A0(new_n2484_), .A1(new_n2481_), .B0(\asqrt[61] ), .Y(new_n2485_));
  INVX1    g02293(.A(new_n2450_), .Y(new_n2486_));
  OAI21X1  g02294(.A0(new_n2435_), .A1(new_n292_), .B0(new_n217_), .Y(new_n2487_));
  OAI21X1  g02295(.A0(new_n2487_), .A1(new_n2484_), .B0(new_n2486_), .Y(new_n2488_));
  NAND3X1  g02296(.A(new_n2488_), .B(new_n2485_), .C(new_n199_), .Y(new_n2489_));
  AND2X1   g02297(.A(new_n2489_), .B(new_n2480_), .Y(new_n2490_));
  AOI21X1  g02298(.A0(new_n2488_), .A1(new_n2485_), .B0(new_n199_), .Y(new_n2491_));
  OR2X1    g02299(.A(new_n2475_), .B(new_n2491_), .Y(new_n2492_));
  AOI21X1  g02300(.A0(new_n2276_), .A1(new_n2272_), .B0(new_n2237_), .Y(new_n2493_));
  AOI21X1  g02301(.A0(new_n2238_), .A1(new_n2232_), .B0(new_n193_), .Y(new_n2494_));
  OAI21X1  g02302(.A0(new_n2493_), .A1(new_n2232_), .B0(new_n2494_), .Y(new_n2495_));
  NOR4X1   g02303(.A(new_n2260_), .B(new_n2257_), .C(new_n2236_), .D(new_n2234_), .Y(new_n2496_));
  OAI21X1  g02304(.A0(new_n2254_), .A1(new_n2253_), .B0(new_n2496_), .Y(new_n2497_));
  NOR2X1   g02305(.A(new_n2497_), .B(new_n2243_), .Y(new_n2498_));
  INVX1    g02306(.A(new_n2498_), .Y(new_n2499_));
  AND2X1   g02307(.A(new_n2499_), .B(new_n2495_), .Y(new_n2500_));
  OAI21X1  g02308(.A0(new_n2492_), .A1(new_n2490_), .B0(new_n2500_), .Y(new_n2501_));
  OR2X1    g02309(.A(new_n2501_), .B(new_n2479_), .Y(\asqrt[45] ));
  NOR3X1   g02310(.A(\a[90] ), .B(\a[89] ), .C(\a[88] ), .Y(new_n2503_));
  AOI21X1  g02311(.A0(\asqrt[45] ), .A1(\a[90] ), .B0(new_n2503_), .Y(new_n2504_));
  OAI21X1  g02312(.A0(new_n2501_), .A1(new_n2479_), .B0(\a[90] ), .Y(new_n2505_));
  OR2X1    g02313(.A(new_n2503_), .B(new_n2260_), .Y(new_n2506_));
  NOR4X1   g02314(.A(new_n2506_), .B(new_n2257_), .C(new_n2290_), .D(new_n2243_), .Y(new_n2507_));
  AND2X1   g02315(.A(new_n2507_), .B(new_n2505_), .Y(new_n2508_));
  INVX1    g02316(.A(\a[91] ), .Y(new_n2509_));
  AOI21X1  g02317(.A0(new_n2489_), .A1(new_n2480_), .B0(new_n2491_), .Y(new_n2510_));
  INVX1    g02318(.A(new_n2478_), .Y(new_n2511_));
  OAI21X1  g02319(.A0(new_n2511_), .A1(new_n2510_), .B0(new_n193_), .Y(new_n2512_));
  NAND2X1  g02320(.A(new_n2489_), .B(new_n2480_), .Y(new_n2513_));
  NOR2X1   g02321(.A(new_n2475_), .B(new_n2491_), .Y(new_n2514_));
  INVX1    g02322(.A(new_n2500_), .Y(new_n2515_));
  AOI21X1  g02323(.A0(new_n2514_), .A1(new_n2513_), .B0(new_n2515_), .Y(new_n2516_));
  AOI21X1  g02324(.A0(new_n2516_), .A1(new_n2512_), .B0(\a[90] ), .Y(new_n2517_));
  OAI21X1  g02325(.A0(new_n2501_), .A1(new_n2479_), .B0(new_n2266_), .Y(new_n2518_));
  OAI21X1  g02326(.A0(new_n2517_), .A1(new_n2509_), .B0(new_n2518_), .Y(new_n2519_));
  OAI22X1  g02327(.A0(new_n2519_), .A1(new_n2508_), .B0(new_n2504_), .B1(new_n2263_), .Y(new_n2520_));
  AND2X1   g02328(.A(new_n2520_), .B(\asqrt[47] ), .Y(new_n2521_));
  NAND2X1  g02329(.A(new_n2507_), .B(new_n2505_), .Y(new_n2522_));
  INVX1    g02330(.A(\a[90] ), .Y(new_n2523_));
  OAI21X1  g02331(.A0(new_n2501_), .A1(new_n2479_), .B0(new_n2523_), .Y(new_n2524_));
  AOI21X1  g02332(.A0(new_n2516_), .A1(new_n2512_), .B0(new_n2286_), .Y(new_n2525_));
  AOI21X1  g02333(.A0(new_n2524_), .A1(\a[91] ), .B0(new_n2525_), .Y(new_n2526_));
  NAND2X1  g02334(.A(new_n2526_), .B(new_n2522_), .Y(new_n2527_));
  NOR2X1   g02335(.A(\a[89] ), .B(\a[88] ), .Y(new_n2528_));
  MX2X1    g02336(.A(new_n2528_), .B(\asqrt[45] ), .S0(\a[90] ), .Y(new_n2529_));
  AOI21X1  g02337(.A0(new_n2529_), .A1(\asqrt[46] ), .B0(\asqrt[47] ), .Y(new_n2530_));
  INVX1    g02338(.A(new_n2495_), .Y(new_n2531_));
  NOR3X1   g02339(.A(new_n2498_), .B(new_n2531_), .C(new_n2263_), .Y(new_n2532_));
  OAI21X1  g02340(.A0(new_n2492_), .A1(new_n2490_), .B0(new_n2532_), .Y(new_n2533_));
  OR2X1    g02341(.A(new_n2533_), .B(new_n2479_), .Y(new_n2534_));
  AOI21X1  g02342(.A0(new_n2534_), .A1(new_n2518_), .B0(new_n2265_), .Y(new_n2535_));
  OAI21X1  g02343(.A0(new_n2533_), .A1(new_n2479_), .B0(new_n2265_), .Y(new_n2536_));
  NOR2X1   g02344(.A(new_n2536_), .B(new_n2525_), .Y(new_n2537_));
  NOR2X1   g02345(.A(new_n2537_), .B(new_n2535_), .Y(new_n2538_));
  AOI21X1  g02346(.A0(new_n2530_), .A1(new_n2527_), .B0(new_n2538_), .Y(new_n2539_));
  OAI21X1  g02347(.A0(new_n2539_), .A1(new_n2521_), .B0(\asqrt[48] ), .Y(new_n2540_));
  AOI21X1  g02348(.A0(new_n2268_), .A1(\asqrt[47] ), .B0(new_n2305_), .Y(new_n2541_));
  AND2X1   g02349(.A(new_n2541_), .B(new_n2308_), .Y(new_n2542_));
  OAI21X1  g02350(.A0(new_n2501_), .A1(new_n2479_), .B0(new_n2541_), .Y(new_n2543_));
  AOI22X1  g02351(.A0(new_n2543_), .A1(new_n2282_), .B0(new_n2542_), .B1(\asqrt[45] ), .Y(new_n2544_));
  INVX1    g02352(.A(new_n2544_), .Y(new_n2545_));
  AOI22X1  g02353(.A0(new_n2526_), .A1(new_n2522_), .B0(new_n2529_), .B1(\asqrt[46] ), .Y(new_n2546_));
  OAI21X1  g02354(.A0(new_n2546_), .A1(new_n2040_), .B0(new_n1834_), .Y(new_n2547_));
  OAI21X1  g02355(.A0(new_n2547_), .A1(new_n2539_), .B0(new_n2545_), .Y(new_n2548_));
  AOI21X1  g02356(.A0(new_n2548_), .A1(new_n2540_), .B0(new_n1632_), .Y(new_n2549_));
  AOI21X1  g02357(.A0(new_n2326_), .A1(new_n2325_), .B0(new_n2296_), .Y(new_n2550_));
  AND2X1   g02358(.A(new_n2550_), .B(new_n2284_), .Y(new_n2551_));
  AOI22X1  g02359(.A0(new_n2326_), .A1(new_n2325_), .B0(new_n2309_), .B1(\asqrt[48] ), .Y(new_n2552_));
  OAI21X1  g02360(.A0(new_n2501_), .A1(new_n2479_), .B0(new_n2552_), .Y(new_n2553_));
  AOI22X1  g02361(.A0(new_n2553_), .A1(new_n2296_), .B0(new_n2551_), .B1(\asqrt[45] ), .Y(new_n2554_));
  INVX1    g02362(.A(new_n2554_), .Y(new_n2555_));
  NAND3X1  g02363(.A(new_n2548_), .B(new_n2540_), .C(new_n1632_), .Y(new_n2556_));
  AOI21X1  g02364(.A0(new_n2556_), .A1(new_n2555_), .B0(new_n2549_), .Y(new_n2557_));
  OR2X1    g02365(.A(new_n2557_), .B(new_n1469_), .Y(new_n2558_));
  AND2X1   g02366(.A(new_n2556_), .B(new_n2555_), .Y(new_n2559_));
  AND2X1   g02367(.A(new_n2310_), .B(new_n2297_), .Y(new_n2560_));
  NOR3X1   g02368(.A(new_n2560_), .B(new_n2330_), .C(new_n2298_), .Y(new_n2561_));
  NOR2X1   g02369(.A(new_n2560_), .B(new_n2298_), .Y(new_n2562_));
  OAI21X1  g02370(.A0(new_n2501_), .A1(new_n2479_), .B0(new_n2562_), .Y(new_n2563_));
  AOI22X1  g02371(.A0(new_n2563_), .A1(new_n2330_), .B0(new_n2561_), .B1(\asqrt[45] ), .Y(new_n2564_));
  INVX1    g02372(.A(new_n2564_), .Y(new_n2565_));
  OR2X1    g02373(.A(new_n2549_), .B(\asqrt[50] ), .Y(new_n2566_));
  OAI21X1  g02374(.A0(new_n2566_), .A1(new_n2559_), .B0(new_n2565_), .Y(new_n2567_));
  AOI21X1  g02375(.A0(new_n2567_), .A1(new_n2558_), .B0(new_n1277_), .Y(new_n2568_));
  NAND4X1  g02376(.A(\asqrt[45] ), .B(new_n2349_), .C(new_n2319_), .D(new_n2312_), .Y(new_n2569_));
  NOR2X1   g02377(.A(new_n2501_), .B(new_n2479_), .Y(new_n2570_));
  NOR3X1   g02378(.A(new_n2570_), .B(new_n2320_), .C(new_n2333_), .Y(new_n2571_));
  OAI21X1  g02379(.A0(new_n2571_), .A1(new_n2319_), .B0(new_n2569_), .Y(new_n2572_));
  INVX1    g02380(.A(new_n2572_), .Y(new_n2573_));
  OR2X1    g02381(.A(new_n2546_), .B(new_n2040_), .Y(new_n2574_));
  AND2X1   g02382(.A(new_n2526_), .B(new_n2522_), .Y(new_n2575_));
  OAI21X1  g02383(.A0(new_n2504_), .A1(new_n2263_), .B0(new_n2040_), .Y(new_n2576_));
  OR2X1    g02384(.A(new_n2537_), .B(new_n2535_), .Y(new_n2577_));
  OAI21X1  g02385(.A0(new_n2576_), .A1(new_n2575_), .B0(new_n2577_), .Y(new_n2578_));
  AOI21X1  g02386(.A0(new_n2578_), .A1(new_n2574_), .B0(new_n1834_), .Y(new_n2579_));
  AOI21X1  g02387(.A0(new_n2520_), .A1(\asqrt[47] ), .B0(\asqrt[48] ), .Y(new_n2580_));
  AOI21X1  g02388(.A0(new_n2580_), .A1(new_n2578_), .B0(new_n2544_), .Y(new_n2581_));
  OAI21X1  g02389(.A0(new_n2581_), .A1(new_n2579_), .B0(\asqrt[49] ), .Y(new_n2582_));
  NOR3X1   g02390(.A(new_n2581_), .B(new_n2579_), .C(\asqrt[49] ), .Y(new_n2583_));
  OAI21X1  g02391(.A0(new_n2583_), .A1(new_n2554_), .B0(new_n2582_), .Y(new_n2584_));
  AOI21X1  g02392(.A0(new_n2584_), .A1(\asqrt[50] ), .B0(\asqrt[51] ), .Y(new_n2585_));
  AOI21X1  g02393(.A0(new_n2585_), .A1(new_n2567_), .B0(new_n2573_), .Y(new_n2586_));
  OAI21X1  g02394(.A0(new_n2586_), .A1(new_n2568_), .B0(\asqrt[52] ), .Y(new_n2587_));
  NOR3X1   g02395(.A(new_n2586_), .B(new_n2568_), .C(\asqrt[52] ), .Y(new_n2588_));
  AND2X1   g02396(.A(new_n2334_), .B(new_n2323_), .Y(new_n2589_));
  NOR3X1   g02397(.A(new_n2372_), .B(new_n2589_), .C(new_n2322_), .Y(new_n2590_));
  AOI22X1  g02398(.A0(new_n2334_), .A1(new_n2323_), .B0(new_n2321_), .B1(\asqrt[51] ), .Y(new_n2591_));
  AOI21X1  g02399(.A0(new_n2591_), .A1(\asqrt[45] ), .B0(new_n2339_), .Y(new_n2592_));
  AOI21X1  g02400(.A0(new_n2590_), .A1(\asqrt[45] ), .B0(new_n2592_), .Y(new_n2593_));
  OAI21X1  g02401(.A0(new_n2593_), .A1(new_n2588_), .B0(new_n2587_), .Y(new_n2594_));
  AND2X1   g02402(.A(new_n2594_), .B(\asqrt[53] ), .Y(new_n2595_));
  AND2X1   g02403(.A(new_n2584_), .B(\asqrt[50] ), .Y(new_n2596_));
  NAND2X1  g02404(.A(new_n2556_), .B(new_n2555_), .Y(new_n2597_));
  NOR2X1   g02405(.A(new_n2549_), .B(\asqrt[50] ), .Y(new_n2598_));
  AOI21X1  g02406(.A0(new_n2598_), .A1(new_n2597_), .B0(new_n2564_), .Y(new_n2599_));
  OAI21X1  g02407(.A0(new_n2599_), .A1(new_n2596_), .B0(\asqrt[51] ), .Y(new_n2600_));
  OAI21X1  g02408(.A0(new_n2557_), .A1(new_n1469_), .B0(new_n1277_), .Y(new_n2601_));
  OAI21X1  g02409(.A0(new_n2601_), .A1(new_n2599_), .B0(new_n2572_), .Y(new_n2602_));
  NAND3X1  g02410(.A(new_n2602_), .B(new_n2600_), .C(new_n1111_), .Y(new_n2603_));
  INVX1    g02411(.A(new_n2593_), .Y(new_n2604_));
  NAND2X1  g02412(.A(new_n2604_), .B(new_n2603_), .Y(new_n2605_));
  AND2X1   g02413(.A(new_n2375_), .B(new_n2373_), .Y(new_n2606_));
  NOR3X1   g02414(.A(new_n2606_), .B(new_n2347_), .C(new_n2374_), .Y(new_n2607_));
  NOR2X1   g02415(.A(new_n2606_), .B(new_n2374_), .Y(new_n2608_));
  AOI21X1  g02416(.A0(new_n2608_), .A1(\asqrt[45] ), .B0(new_n2346_), .Y(new_n2609_));
  AOI21X1  g02417(.A0(new_n2607_), .A1(\asqrt[45] ), .B0(new_n2609_), .Y(new_n2610_));
  AOI21X1  g02418(.A0(new_n2602_), .A1(new_n2600_), .B0(new_n1111_), .Y(new_n2611_));
  NOR2X1   g02419(.A(new_n2611_), .B(\asqrt[53] ), .Y(new_n2612_));
  AOI21X1  g02420(.A0(new_n2612_), .A1(new_n2605_), .B0(new_n2610_), .Y(new_n2613_));
  OAI21X1  g02421(.A0(new_n2613_), .A1(new_n2595_), .B0(\asqrt[54] ), .Y(new_n2614_));
  OR4X1    g02422(.A(new_n2570_), .B(new_n2386_), .C(new_n2359_), .D(new_n2353_), .Y(new_n2615_));
  OR2X1    g02423(.A(new_n2386_), .B(new_n2353_), .Y(new_n2616_));
  OAI21X1  g02424(.A0(new_n2616_), .A1(new_n2570_), .B0(new_n2359_), .Y(new_n2617_));
  AND2X1   g02425(.A(new_n2617_), .B(new_n2615_), .Y(new_n2618_));
  INVX1    g02426(.A(new_n2618_), .Y(new_n2619_));
  AOI21X1  g02427(.A0(new_n2604_), .A1(new_n2603_), .B0(new_n2611_), .Y(new_n2620_));
  OAI21X1  g02428(.A0(new_n2620_), .A1(new_n968_), .B0(new_n902_), .Y(new_n2621_));
  OAI21X1  g02429(.A0(new_n2621_), .A1(new_n2613_), .B0(new_n2619_), .Y(new_n2622_));
  AOI21X1  g02430(.A0(new_n2622_), .A1(new_n2614_), .B0(new_n697_), .Y(new_n2623_));
  AOI21X1  g02431(.A0(new_n2402_), .A1(new_n2401_), .B0(new_n2368_), .Y(new_n2624_));
  AND2X1   g02432(.A(new_n2624_), .B(new_n2362_), .Y(new_n2625_));
  AOI22X1  g02433(.A0(new_n2402_), .A1(new_n2401_), .B0(new_n2387_), .B1(\asqrt[54] ), .Y(new_n2626_));
  AOI21X1  g02434(.A0(new_n2626_), .A1(\asqrt[45] ), .B0(new_n2367_), .Y(new_n2627_));
  AOI21X1  g02435(.A0(new_n2625_), .A1(\asqrt[45] ), .B0(new_n2627_), .Y(new_n2628_));
  INVX1    g02436(.A(new_n2628_), .Y(new_n2629_));
  NAND3X1  g02437(.A(new_n2622_), .B(new_n2614_), .C(new_n697_), .Y(new_n2630_));
  AOI21X1  g02438(.A0(new_n2630_), .A1(new_n2629_), .B0(new_n2623_), .Y(new_n2631_));
  OR2X1    g02439(.A(new_n2631_), .B(new_n582_), .Y(new_n2632_));
  AND2X1   g02440(.A(new_n2630_), .B(new_n2629_), .Y(new_n2633_));
  AND2X1   g02441(.A(new_n2388_), .B(new_n2379_), .Y(new_n2634_));
  NOR3X1   g02442(.A(new_n2634_), .B(new_n2405_), .C(new_n2380_), .Y(new_n2635_));
  NOR2X1   g02443(.A(new_n2634_), .B(new_n2380_), .Y(new_n2636_));
  AOI21X1  g02444(.A0(new_n2636_), .A1(\asqrt[45] ), .B0(new_n2385_), .Y(new_n2637_));
  AOI21X1  g02445(.A0(new_n2635_), .A1(\asqrt[45] ), .B0(new_n2637_), .Y(new_n2638_));
  INVX1    g02446(.A(new_n2638_), .Y(new_n2639_));
  OR2X1    g02447(.A(new_n2623_), .B(\asqrt[56] ), .Y(new_n2640_));
  OAI21X1  g02448(.A0(new_n2640_), .A1(new_n2633_), .B0(new_n2639_), .Y(new_n2641_));
  AOI21X1  g02449(.A0(new_n2641_), .A1(new_n2632_), .B0(new_n481_), .Y(new_n2642_));
  OR4X1    g02450(.A(new_n2570_), .B(new_n2396_), .C(new_n2399_), .D(new_n2414_), .Y(new_n2643_));
  NAND2X1  g02451(.A(new_n2408_), .B(new_n2390_), .Y(new_n2644_));
  OAI21X1  g02452(.A0(new_n2644_), .A1(new_n2570_), .B0(new_n2399_), .Y(new_n2645_));
  AND2X1   g02453(.A(new_n2645_), .B(new_n2643_), .Y(new_n2646_));
  OR2X1    g02454(.A(new_n2620_), .B(new_n968_), .Y(new_n2647_));
  AND2X1   g02455(.A(new_n2604_), .B(new_n2603_), .Y(new_n2648_));
  INVX1    g02456(.A(new_n2610_), .Y(new_n2649_));
  OR2X1    g02457(.A(new_n2611_), .B(\asqrt[53] ), .Y(new_n2650_));
  OAI21X1  g02458(.A0(new_n2650_), .A1(new_n2648_), .B0(new_n2649_), .Y(new_n2651_));
  AOI21X1  g02459(.A0(new_n2651_), .A1(new_n2647_), .B0(new_n902_), .Y(new_n2652_));
  AOI21X1  g02460(.A0(new_n2594_), .A1(\asqrt[53] ), .B0(\asqrt[54] ), .Y(new_n2653_));
  AOI21X1  g02461(.A0(new_n2653_), .A1(new_n2651_), .B0(new_n2618_), .Y(new_n2654_));
  OAI21X1  g02462(.A0(new_n2654_), .A1(new_n2652_), .B0(\asqrt[55] ), .Y(new_n2655_));
  NOR3X1   g02463(.A(new_n2654_), .B(new_n2652_), .C(\asqrt[55] ), .Y(new_n2656_));
  OAI21X1  g02464(.A0(new_n2656_), .A1(new_n2628_), .B0(new_n2655_), .Y(new_n2657_));
  AOI21X1  g02465(.A0(new_n2657_), .A1(\asqrt[56] ), .B0(\asqrt[57] ), .Y(new_n2658_));
  AOI21X1  g02466(.A0(new_n2658_), .A1(new_n2641_), .B0(new_n2646_), .Y(new_n2659_));
  OAI21X1  g02467(.A0(new_n2659_), .A1(new_n2642_), .B0(\asqrt[58] ), .Y(new_n2660_));
  AND2X1   g02468(.A(new_n2415_), .B(new_n2409_), .Y(new_n2661_));
  NOR3X1   g02469(.A(new_n2661_), .B(new_n2453_), .C(new_n2398_), .Y(new_n2662_));
  AOI22X1  g02470(.A0(new_n2415_), .A1(new_n2409_), .B0(new_n2397_), .B1(\asqrt[57] ), .Y(new_n2663_));
  AOI21X1  g02471(.A0(new_n2663_), .A1(\asqrt[45] ), .B0(new_n2413_), .Y(new_n2664_));
  AOI21X1  g02472(.A0(new_n2662_), .A1(\asqrt[45] ), .B0(new_n2664_), .Y(new_n2665_));
  NOR3X1   g02473(.A(new_n2659_), .B(new_n2642_), .C(\asqrt[58] ), .Y(new_n2666_));
  OAI21X1  g02474(.A0(new_n2666_), .A1(new_n2665_), .B0(new_n2660_), .Y(new_n2667_));
  AND2X1   g02475(.A(new_n2667_), .B(\asqrt[59] ), .Y(new_n2668_));
  INVX1    g02476(.A(new_n2665_), .Y(new_n2669_));
  AND2X1   g02477(.A(new_n2657_), .B(\asqrt[56] ), .Y(new_n2670_));
  NAND2X1  g02478(.A(new_n2630_), .B(new_n2629_), .Y(new_n2671_));
  NOR2X1   g02479(.A(new_n2623_), .B(\asqrt[56] ), .Y(new_n2672_));
  AOI21X1  g02480(.A0(new_n2672_), .A1(new_n2671_), .B0(new_n2638_), .Y(new_n2673_));
  OAI21X1  g02481(.A0(new_n2673_), .A1(new_n2670_), .B0(\asqrt[57] ), .Y(new_n2674_));
  INVX1    g02482(.A(new_n2646_), .Y(new_n2675_));
  OAI21X1  g02483(.A0(new_n2631_), .A1(new_n582_), .B0(new_n481_), .Y(new_n2676_));
  OAI21X1  g02484(.A0(new_n2676_), .A1(new_n2673_), .B0(new_n2675_), .Y(new_n2677_));
  NAND3X1  g02485(.A(new_n2677_), .B(new_n2674_), .C(new_n399_), .Y(new_n2678_));
  NAND2X1  g02486(.A(new_n2678_), .B(new_n2669_), .Y(new_n2679_));
  AND2X1   g02487(.A(new_n2457_), .B(new_n2455_), .Y(new_n2680_));
  NOR3X1   g02488(.A(new_n2680_), .B(new_n2423_), .C(new_n2456_), .Y(new_n2681_));
  NOR2X1   g02489(.A(new_n2680_), .B(new_n2456_), .Y(new_n2682_));
  AOI21X1  g02490(.A0(new_n2682_), .A1(\asqrt[45] ), .B0(new_n2422_), .Y(new_n2683_));
  AOI21X1  g02491(.A0(new_n2681_), .A1(\asqrt[45] ), .B0(new_n2683_), .Y(new_n2684_));
  AOI21X1  g02492(.A0(new_n2677_), .A1(new_n2674_), .B0(new_n399_), .Y(new_n2685_));
  NOR2X1   g02493(.A(new_n2685_), .B(\asqrt[59] ), .Y(new_n2686_));
  AOI21X1  g02494(.A0(new_n2686_), .A1(new_n2679_), .B0(new_n2684_), .Y(new_n2687_));
  OAI21X1  g02495(.A0(new_n2687_), .A1(new_n2668_), .B0(\asqrt[60] ), .Y(new_n2688_));
  OR4X1    g02496(.A(new_n2570_), .B(new_n2460_), .C(new_n2433_), .D(new_n2427_), .Y(new_n2689_));
  NAND2X1  g02497(.A(new_n2434_), .B(new_n2459_), .Y(new_n2690_));
  OAI21X1  g02498(.A0(new_n2690_), .A1(new_n2570_), .B0(new_n2433_), .Y(new_n2691_));
  AND2X1   g02499(.A(new_n2691_), .B(new_n2689_), .Y(new_n2692_));
  INVX1    g02500(.A(new_n2692_), .Y(new_n2693_));
  AOI21X1  g02501(.A0(new_n2678_), .A1(new_n2669_), .B0(new_n2685_), .Y(new_n2694_));
  OAI21X1  g02502(.A0(new_n2694_), .A1(new_n328_), .B0(new_n292_), .Y(new_n2695_));
  OAI21X1  g02503(.A0(new_n2695_), .A1(new_n2687_), .B0(new_n2693_), .Y(new_n2696_));
  AOI21X1  g02504(.A0(new_n2696_), .A1(new_n2688_), .B0(new_n217_), .Y(new_n2697_));
  AOI21X1  g02505(.A0(new_n2483_), .A1(new_n2482_), .B0(new_n2442_), .Y(new_n2698_));
  AND2X1   g02506(.A(new_n2698_), .B(new_n2436_), .Y(new_n2699_));
  AOI22X1  g02507(.A0(new_n2483_), .A1(new_n2482_), .B0(new_n2461_), .B1(\asqrt[60] ), .Y(new_n2700_));
  AOI21X1  g02508(.A0(new_n2700_), .A1(\asqrt[45] ), .B0(new_n2441_), .Y(new_n2701_));
  AOI21X1  g02509(.A0(new_n2699_), .A1(\asqrt[45] ), .B0(new_n2701_), .Y(new_n2702_));
  INVX1    g02510(.A(new_n2702_), .Y(new_n2703_));
  NAND3X1  g02511(.A(new_n2696_), .B(new_n2688_), .C(new_n217_), .Y(new_n2704_));
  AOI21X1  g02512(.A0(new_n2704_), .A1(new_n2703_), .B0(new_n2697_), .Y(new_n2705_));
  OR2X1    g02513(.A(new_n2705_), .B(new_n199_), .Y(new_n2706_));
  AND2X1   g02514(.A(new_n2704_), .B(new_n2703_), .Y(new_n2707_));
  AND2X1   g02515(.A(new_n2462_), .B(new_n2444_), .Y(new_n2708_));
  NOR3X1   g02516(.A(new_n2708_), .B(new_n2486_), .C(new_n2445_), .Y(new_n2709_));
  NOR2X1   g02517(.A(new_n2708_), .B(new_n2445_), .Y(new_n2710_));
  AOI21X1  g02518(.A0(new_n2710_), .A1(\asqrt[45] ), .B0(new_n2450_), .Y(new_n2711_));
  AOI21X1  g02519(.A0(new_n2709_), .A1(\asqrt[45] ), .B0(new_n2711_), .Y(new_n2712_));
  INVX1    g02520(.A(new_n2712_), .Y(new_n2713_));
  OR2X1    g02521(.A(new_n2697_), .B(\asqrt[62] ), .Y(new_n2714_));
  OAI21X1  g02522(.A0(new_n2714_), .A1(new_n2707_), .B0(new_n2713_), .Y(new_n2715_));
  OR4X1    g02523(.A(new_n2570_), .B(new_n2470_), .C(new_n2480_), .D(new_n2491_), .Y(new_n2716_));
  NAND2X1  g02524(.A(new_n2489_), .B(new_n2464_), .Y(new_n2717_));
  OAI21X1  g02525(.A0(new_n2717_), .A1(new_n2570_), .B0(new_n2480_), .Y(new_n2718_));
  AND2X1   g02526(.A(new_n2718_), .B(new_n2716_), .Y(new_n2719_));
  INVX1    g02527(.A(new_n2719_), .Y(new_n2720_));
  NOR2X1   g02528(.A(new_n2474_), .B(new_n2510_), .Y(new_n2721_));
  AOI22X1  g02529(.A0(new_n2721_), .A1(\asqrt[45] ), .B0(new_n2514_), .B1(new_n2513_), .Y(new_n2722_));
  AND2X1   g02530(.A(new_n2722_), .B(new_n2720_), .Y(new_n2723_));
  INVX1    g02531(.A(new_n2723_), .Y(new_n2724_));
  AOI21X1  g02532(.A0(new_n2715_), .A1(new_n2706_), .B0(new_n2724_), .Y(new_n2725_));
  OR2X1    g02533(.A(new_n2694_), .B(new_n328_), .Y(new_n2726_));
  AND2X1   g02534(.A(new_n2678_), .B(new_n2669_), .Y(new_n2727_));
  INVX1    g02535(.A(new_n2684_), .Y(new_n2728_));
  OR2X1    g02536(.A(new_n2685_), .B(\asqrt[59] ), .Y(new_n2729_));
  OAI21X1  g02537(.A0(new_n2729_), .A1(new_n2727_), .B0(new_n2728_), .Y(new_n2730_));
  AOI21X1  g02538(.A0(new_n2730_), .A1(new_n2726_), .B0(new_n292_), .Y(new_n2731_));
  AOI21X1  g02539(.A0(new_n2667_), .A1(\asqrt[59] ), .B0(\asqrt[60] ), .Y(new_n2732_));
  AOI21X1  g02540(.A0(new_n2732_), .A1(new_n2730_), .B0(new_n2692_), .Y(new_n2733_));
  OAI21X1  g02541(.A0(new_n2733_), .A1(new_n2731_), .B0(\asqrt[61] ), .Y(new_n2734_));
  NOR3X1   g02542(.A(new_n2733_), .B(new_n2731_), .C(\asqrt[61] ), .Y(new_n2735_));
  OAI21X1  g02543(.A0(new_n2735_), .A1(new_n2702_), .B0(new_n2734_), .Y(new_n2736_));
  AOI21X1  g02544(.A0(new_n2736_), .A1(\asqrt[62] ), .B0(new_n2720_), .Y(new_n2737_));
  AOI21X1  g02545(.A0(new_n2516_), .A1(new_n2512_), .B0(new_n2474_), .Y(new_n2738_));
  AOI21X1  g02546(.A0(new_n2475_), .A1(new_n2471_), .B0(new_n193_), .Y(new_n2739_));
  OAI21X1  g02547(.A0(new_n2738_), .A1(new_n2471_), .B0(new_n2739_), .Y(new_n2740_));
  OR2X1    g02548(.A(new_n2492_), .B(new_n2490_), .Y(new_n2741_));
  AND2X1   g02549(.A(new_n2473_), .B(new_n2229_), .Y(new_n2742_));
  NOR4X1   g02550(.A(new_n2498_), .B(new_n2531_), .C(new_n2742_), .D(new_n2472_), .Y(new_n2743_));
  NAND3X1  g02551(.A(new_n2743_), .B(new_n2741_), .C(new_n2512_), .Y(new_n2744_));
  AND2X1   g02552(.A(new_n2744_), .B(new_n2740_), .Y(new_n2745_));
  INVX1    g02553(.A(new_n2745_), .Y(new_n2746_));
  AOI21X1  g02554(.A0(new_n2737_), .A1(new_n2715_), .B0(new_n2746_), .Y(new_n2747_));
  OAI21X1  g02555(.A0(new_n2725_), .A1(\asqrt[63] ), .B0(new_n2747_), .Y(\asqrt[44] ));
  NOR2X1   g02556(.A(\a[87] ), .B(\a[86] ), .Y(new_n2749_));
  MX2X1    g02557(.A(new_n2749_), .B(\asqrt[44] ), .S0(\a[88] ), .Y(new_n2750_));
  AND2X1   g02558(.A(new_n2750_), .B(\asqrt[45] ), .Y(new_n2751_));
  NOR3X1   g02559(.A(\a[88] ), .B(\a[87] ), .C(\a[86] ), .Y(new_n2752_));
  NOR3X1   g02560(.A(new_n2752_), .B(new_n2498_), .C(new_n2531_), .Y(new_n2753_));
  NAND3X1  g02561(.A(new_n2753_), .B(new_n2741_), .C(new_n2512_), .Y(new_n2754_));
  AOI21X1  g02562(.A0(\asqrt[44] ), .A1(\a[88] ), .B0(new_n2754_), .Y(new_n2755_));
  INVX1    g02563(.A(\a[88] ), .Y(new_n2756_));
  INVX1    g02564(.A(\a[89] ), .Y(new_n2757_));
  AOI21X1  g02565(.A0(\asqrt[44] ), .A1(new_n2756_), .B0(new_n2757_), .Y(new_n2758_));
  AND2X1   g02566(.A(\asqrt[44] ), .B(new_n2528_), .Y(new_n2759_));
  NOR3X1   g02567(.A(new_n2759_), .B(new_n2758_), .C(new_n2755_), .Y(new_n2760_));
  OAI21X1  g02568(.A0(new_n2760_), .A1(new_n2751_), .B0(\asqrt[46] ), .Y(new_n2761_));
  AND2X1   g02569(.A(new_n2736_), .B(\asqrt[62] ), .Y(new_n2762_));
  NAND2X1  g02570(.A(new_n2704_), .B(new_n2703_), .Y(new_n2763_));
  NOR2X1   g02571(.A(new_n2697_), .B(\asqrt[62] ), .Y(new_n2764_));
  AOI21X1  g02572(.A0(new_n2764_), .A1(new_n2763_), .B0(new_n2712_), .Y(new_n2765_));
  OAI21X1  g02573(.A0(new_n2765_), .A1(new_n2762_), .B0(new_n2723_), .Y(new_n2766_));
  OAI21X1  g02574(.A0(new_n2705_), .A1(new_n199_), .B0(new_n2719_), .Y(new_n2767_));
  OAI21X1  g02575(.A0(new_n2767_), .A1(new_n2765_), .B0(new_n2745_), .Y(new_n2768_));
  AOI21X1  g02576(.A0(new_n2766_), .A1(new_n193_), .B0(new_n2768_), .Y(new_n2769_));
  INVX1    g02577(.A(new_n2749_), .Y(new_n2770_));
  MX2X1    g02578(.A(new_n2770_), .B(new_n2769_), .S0(\a[88] ), .Y(new_n2771_));
  OAI21X1  g02579(.A0(new_n2771_), .A1(new_n2570_), .B0(new_n2263_), .Y(new_n2772_));
  NAND3X1  g02580(.A(new_n2744_), .B(new_n2740_), .C(\asqrt[45] ), .Y(new_n2773_));
  INVX1    g02581(.A(new_n2773_), .Y(new_n2774_));
  OAI21X1  g02582(.A0(new_n2767_), .A1(new_n2765_), .B0(new_n2774_), .Y(new_n2775_));
  AOI21X1  g02583(.A0(new_n2766_), .A1(new_n193_), .B0(new_n2775_), .Y(new_n2776_));
  AOI21X1  g02584(.A0(\asqrt[44] ), .A1(new_n2528_), .B0(new_n2776_), .Y(new_n2777_));
  OR2X1    g02585(.A(new_n2776_), .B(\a[90] ), .Y(new_n2778_));
  OAI22X1  g02586(.A0(new_n2778_), .A1(new_n2759_), .B0(new_n2777_), .B1(new_n2523_), .Y(new_n2779_));
  OAI21X1  g02587(.A0(new_n2772_), .A1(new_n2760_), .B0(new_n2779_), .Y(new_n2780_));
  AOI21X1  g02588(.A0(new_n2780_), .A1(new_n2761_), .B0(new_n2040_), .Y(new_n2781_));
  AOI21X1  g02589(.A0(new_n2529_), .A1(\asqrt[46] ), .B0(new_n2508_), .Y(new_n2782_));
  NAND3X1  g02590(.A(new_n2782_), .B(\asqrt[44] ), .C(new_n2519_), .Y(new_n2783_));
  INVX1    g02591(.A(new_n2782_), .Y(new_n2784_));
  OAI21X1  g02592(.A0(new_n2784_), .A1(new_n2769_), .B0(new_n2526_), .Y(new_n2785_));
  AND2X1   g02593(.A(new_n2785_), .B(new_n2783_), .Y(new_n2786_));
  INVX1    g02594(.A(new_n2786_), .Y(new_n2787_));
  NAND3X1  g02595(.A(new_n2780_), .B(new_n2761_), .C(new_n2040_), .Y(new_n2788_));
  AOI21X1  g02596(.A0(new_n2788_), .A1(new_n2787_), .B0(new_n2781_), .Y(new_n2789_));
  OR2X1    g02597(.A(new_n2789_), .B(new_n1834_), .Y(new_n2790_));
  AND2X1   g02598(.A(new_n2788_), .B(new_n2787_), .Y(new_n2791_));
  OAI21X1  g02599(.A0(new_n2576_), .A1(new_n2575_), .B0(new_n2538_), .Y(new_n2792_));
  NOR3X1   g02600(.A(new_n2792_), .B(new_n2769_), .C(new_n2521_), .Y(new_n2793_));
  OAI22X1  g02601(.A0(new_n2576_), .A1(new_n2575_), .B0(new_n2546_), .B1(new_n2040_), .Y(new_n2794_));
  OR2X1    g02602(.A(new_n2794_), .B(new_n2769_), .Y(new_n2795_));
  AOI21X1  g02603(.A0(new_n2795_), .A1(new_n2577_), .B0(new_n2793_), .Y(new_n2796_));
  INVX1    g02604(.A(new_n2796_), .Y(new_n2797_));
  OR2X1    g02605(.A(new_n2781_), .B(\asqrt[48] ), .Y(new_n2798_));
  OAI21X1  g02606(.A0(new_n2798_), .A1(new_n2791_), .B0(new_n2797_), .Y(new_n2799_));
  AOI21X1  g02607(.A0(new_n2799_), .A1(new_n2790_), .B0(new_n1632_), .Y(new_n2800_));
  AND2X1   g02608(.A(new_n2580_), .B(new_n2578_), .Y(new_n2801_));
  NOR4X1   g02609(.A(new_n2769_), .B(new_n2801_), .C(new_n2545_), .D(new_n2579_), .Y(new_n2802_));
  OR2X1    g02610(.A(new_n2801_), .B(new_n2579_), .Y(new_n2803_));
  OR2X1    g02611(.A(new_n2803_), .B(new_n2769_), .Y(new_n2804_));
  AOI21X1  g02612(.A0(new_n2804_), .A1(new_n2545_), .B0(new_n2802_), .Y(new_n2805_));
  OR2X1    g02613(.A(new_n2771_), .B(new_n2570_), .Y(new_n2806_));
  INVX1    g02614(.A(new_n2754_), .Y(new_n2807_));
  OAI21X1  g02615(.A0(new_n2769_), .A1(new_n2756_), .B0(new_n2807_), .Y(new_n2808_));
  OAI21X1  g02616(.A0(new_n2769_), .A1(\a[88] ), .B0(\a[89] ), .Y(new_n2809_));
  INVX1    g02617(.A(new_n2528_), .Y(new_n2810_));
  OR2X1    g02618(.A(new_n2769_), .B(new_n2810_), .Y(new_n2811_));
  NAND3X1  g02619(.A(new_n2811_), .B(new_n2809_), .C(new_n2808_), .Y(new_n2812_));
  AOI21X1  g02620(.A0(new_n2812_), .A1(new_n2806_), .B0(new_n2263_), .Y(new_n2813_));
  AOI21X1  g02621(.A0(new_n2750_), .A1(\asqrt[45] ), .B0(\asqrt[46] ), .Y(new_n2814_));
  OR2X1    g02622(.A(new_n2777_), .B(new_n2523_), .Y(new_n2815_));
  OR2X1    g02623(.A(new_n2778_), .B(new_n2759_), .Y(new_n2816_));
  AOI22X1  g02624(.A0(new_n2816_), .A1(new_n2815_), .B0(new_n2814_), .B1(new_n2812_), .Y(new_n2817_));
  OAI21X1  g02625(.A0(new_n2817_), .A1(new_n2813_), .B0(\asqrt[47] ), .Y(new_n2818_));
  NOR3X1   g02626(.A(new_n2817_), .B(new_n2813_), .C(\asqrt[47] ), .Y(new_n2819_));
  OAI21X1  g02627(.A0(new_n2819_), .A1(new_n2786_), .B0(new_n2818_), .Y(new_n2820_));
  AOI21X1  g02628(.A0(new_n2820_), .A1(\asqrt[48] ), .B0(\asqrt[49] ), .Y(new_n2821_));
  AOI21X1  g02629(.A0(new_n2821_), .A1(new_n2799_), .B0(new_n2805_), .Y(new_n2822_));
  OAI21X1  g02630(.A0(new_n2822_), .A1(new_n2800_), .B0(\asqrt[50] ), .Y(new_n2823_));
  NAND3X1  g02631(.A(new_n2556_), .B(new_n2554_), .C(new_n2582_), .Y(new_n2824_));
  NOR3X1   g02632(.A(new_n2769_), .B(new_n2583_), .C(new_n2549_), .Y(new_n2825_));
  OAI22X1  g02633(.A0(new_n2825_), .A1(new_n2554_), .B0(new_n2824_), .B1(new_n2769_), .Y(new_n2826_));
  INVX1    g02634(.A(new_n2826_), .Y(new_n2827_));
  NOR3X1   g02635(.A(new_n2822_), .B(new_n2800_), .C(\asqrt[50] ), .Y(new_n2828_));
  OAI21X1  g02636(.A0(new_n2828_), .A1(new_n2827_), .B0(new_n2823_), .Y(new_n2829_));
  AND2X1   g02637(.A(new_n2829_), .B(\asqrt[51] ), .Y(new_n2830_));
  AND2X1   g02638(.A(new_n2820_), .B(\asqrt[48] ), .Y(new_n2831_));
  NAND2X1  g02639(.A(new_n2788_), .B(new_n2787_), .Y(new_n2832_));
  NOR2X1   g02640(.A(new_n2781_), .B(\asqrt[48] ), .Y(new_n2833_));
  AOI21X1  g02641(.A0(new_n2833_), .A1(new_n2832_), .B0(new_n2796_), .Y(new_n2834_));
  OAI21X1  g02642(.A0(new_n2834_), .A1(new_n2831_), .B0(\asqrt[49] ), .Y(new_n2835_));
  INVX1    g02643(.A(new_n2805_), .Y(new_n2836_));
  OAI21X1  g02644(.A0(new_n2789_), .A1(new_n1834_), .B0(new_n1632_), .Y(new_n2837_));
  OAI21X1  g02645(.A0(new_n2837_), .A1(new_n2834_), .B0(new_n2836_), .Y(new_n2838_));
  NAND3X1  g02646(.A(new_n2838_), .B(new_n2835_), .C(new_n1469_), .Y(new_n2839_));
  NAND2X1  g02647(.A(new_n2839_), .B(new_n2826_), .Y(new_n2840_));
  AND2X1   g02648(.A(new_n2598_), .B(new_n2597_), .Y(new_n2841_));
  NOR4X1   g02649(.A(new_n2769_), .B(new_n2841_), .C(new_n2565_), .D(new_n2596_), .Y(new_n2842_));
  AOI22X1  g02650(.A0(new_n2598_), .A1(new_n2597_), .B0(new_n2584_), .B1(\asqrt[50] ), .Y(new_n2843_));
  AOI21X1  g02651(.A0(new_n2843_), .A1(\asqrt[44] ), .B0(new_n2564_), .Y(new_n2844_));
  NOR2X1   g02652(.A(new_n2844_), .B(new_n2842_), .Y(new_n2845_));
  AOI21X1  g02653(.A0(new_n2838_), .A1(new_n2835_), .B0(new_n1469_), .Y(new_n2846_));
  NOR2X1   g02654(.A(new_n2846_), .B(\asqrt[51] ), .Y(new_n2847_));
  AOI21X1  g02655(.A0(new_n2847_), .A1(new_n2840_), .B0(new_n2845_), .Y(new_n2848_));
  OAI21X1  g02656(.A0(new_n2848_), .A1(new_n2830_), .B0(\asqrt[52] ), .Y(new_n2849_));
  AND2X1   g02657(.A(new_n2585_), .B(new_n2567_), .Y(new_n2850_));
  NOR4X1   g02658(.A(new_n2769_), .B(new_n2850_), .C(new_n2572_), .D(new_n2568_), .Y(new_n2851_));
  NOR2X1   g02659(.A(new_n2850_), .B(new_n2568_), .Y(new_n2852_));
  AOI21X1  g02660(.A0(new_n2852_), .A1(\asqrt[44] ), .B0(new_n2573_), .Y(new_n2853_));
  NOR2X1   g02661(.A(new_n2853_), .B(new_n2851_), .Y(new_n2854_));
  INVX1    g02662(.A(new_n2854_), .Y(new_n2855_));
  AOI21X1  g02663(.A0(new_n2839_), .A1(new_n2826_), .B0(new_n2846_), .Y(new_n2856_));
  OAI21X1  g02664(.A0(new_n2856_), .A1(new_n1277_), .B0(new_n1111_), .Y(new_n2857_));
  OAI21X1  g02665(.A0(new_n2857_), .A1(new_n2848_), .B0(new_n2855_), .Y(new_n2858_));
  AOI21X1  g02666(.A0(new_n2858_), .A1(new_n2849_), .B0(new_n968_), .Y(new_n2859_));
  NAND3X1  g02667(.A(new_n2858_), .B(new_n2849_), .C(new_n968_), .Y(new_n2860_));
  OR4X1    g02668(.A(new_n2769_), .B(new_n2604_), .C(new_n2588_), .D(new_n2611_), .Y(new_n2861_));
  OR2X1    g02669(.A(new_n2588_), .B(new_n2611_), .Y(new_n2862_));
  OAI21X1  g02670(.A0(new_n2862_), .A1(new_n2769_), .B0(new_n2604_), .Y(new_n2863_));
  AND2X1   g02671(.A(new_n2863_), .B(new_n2861_), .Y(new_n2864_));
  INVX1    g02672(.A(new_n2864_), .Y(new_n2865_));
  AOI21X1  g02673(.A0(new_n2865_), .A1(new_n2860_), .B0(new_n2859_), .Y(new_n2866_));
  OR2X1    g02674(.A(new_n2866_), .B(new_n902_), .Y(new_n2867_));
  OR2X1    g02675(.A(new_n2856_), .B(new_n1277_), .Y(new_n2868_));
  AND2X1   g02676(.A(new_n2839_), .B(new_n2826_), .Y(new_n2869_));
  INVX1    g02677(.A(new_n2845_), .Y(new_n2870_));
  OR2X1    g02678(.A(new_n2846_), .B(\asqrt[51] ), .Y(new_n2871_));
  OAI21X1  g02679(.A0(new_n2871_), .A1(new_n2869_), .B0(new_n2870_), .Y(new_n2872_));
  AOI21X1  g02680(.A0(new_n2872_), .A1(new_n2868_), .B0(new_n1111_), .Y(new_n2873_));
  AOI21X1  g02681(.A0(new_n2829_), .A1(\asqrt[51] ), .B0(\asqrt[52] ), .Y(new_n2874_));
  AOI21X1  g02682(.A0(new_n2874_), .A1(new_n2872_), .B0(new_n2854_), .Y(new_n2875_));
  NOR3X1   g02683(.A(new_n2875_), .B(new_n2873_), .C(\asqrt[53] ), .Y(new_n2876_));
  NOR2X1   g02684(.A(new_n2864_), .B(new_n2876_), .Y(new_n2877_));
  OAI21X1  g02685(.A0(new_n2650_), .A1(new_n2648_), .B0(new_n2610_), .Y(new_n2878_));
  NOR3X1   g02686(.A(new_n2878_), .B(new_n2769_), .C(new_n2595_), .Y(new_n2879_));
  AOI22X1  g02687(.A0(new_n2612_), .A1(new_n2605_), .B0(new_n2594_), .B1(\asqrt[53] ), .Y(new_n2880_));
  AOI21X1  g02688(.A0(new_n2880_), .A1(\asqrt[44] ), .B0(new_n2610_), .Y(new_n2881_));
  NOR2X1   g02689(.A(new_n2881_), .B(new_n2879_), .Y(new_n2882_));
  INVX1    g02690(.A(new_n2882_), .Y(new_n2883_));
  OAI21X1  g02691(.A0(new_n2875_), .A1(new_n2873_), .B0(\asqrt[53] ), .Y(new_n2884_));
  NAND2X1  g02692(.A(new_n2884_), .B(new_n902_), .Y(new_n2885_));
  OAI21X1  g02693(.A0(new_n2885_), .A1(new_n2877_), .B0(new_n2883_), .Y(new_n2886_));
  AOI21X1  g02694(.A0(new_n2886_), .A1(new_n2867_), .B0(new_n697_), .Y(new_n2887_));
  AND2X1   g02695(.A(new_n2653_), .B(new_n2651_), .Y(new_n2888_));
  OR4X1    g02696(.A(new_n2769_), .B(new_n2888_), .C(new_n2619_), .D(new_n2652_), .Y(new_n2889_));
  OR2X1    g02697(.A(new_n2888_), .B(new_n2652_), .Y(new_n2890_));
  OAI21X1  g02698(.A0(new_n2890_), .A1(new_n2769_), .B0(new_n2619_), .Y(new_n2891_));
  AND2X1   g02699(.A(new_n2891_), .B(new_n2889_), .Y(new_n2892_));
  OAI21X1  g02700(.A0(new_n2864_), .A1(new_n2876_), .B0(new_n2884_), .Y(new_n2893_));
  AOI21X1  g02701(.A0(new_n2893_), .A1(\asqrt[54] ), .B0(\asqrt[55] ), .Y(new_n2894_));
  AOI21X1  g02702(.A0(new_n2894_), .A1(new_n2886_), .B0(new_n2892_), .Y(new_n2895_));
  OAI21X1  g02703(.A0(new_n2895_), .A1(new_n2887_), .B0(\asqrt[56] ), .Y(new_n2896_));
  NAND3X1  g02704(.A(new_n2630_), .B(new_n2628_), .C(new_n2655_), .Y(new_n2897_));
  NOR3X1   g02705(.A(new_n2769_), .B(new_n2656_), .C(new_n2623_), .Y(new_n2898_));
  OAI22X1  g02706(.A0(new_n2898_), .A1(new_n2628_), .B0(new_n2897_), .B1(new_n2769_), .Y(new_n2899_));
  INVX1    g02707(.A(new_n2899_), .Y(new_n2900_));
  NOR3X1   g02708(.A(new_n2895_), .B(new_n2887_), .C(\asqrt[56] ), .Y(new_n2901_));
  OAI21X1  g02709(.A0(new_n2901_), .A1(new_n2900_), .B0(new_n2896_), .Y(new_n2902_));
  AND2X1   g02710(.A(new_n2902_), .B(\asqrt[57] ), .Y(new_n2903_));
  AND2X1   g02711(.A(new_n2893_), .B(\asqrt[54] ), .Y(new_n2904_));
  OR2X1    g02712(.A(new_n2864_), .B(new_n2876_), .Y(new_n2905_));
  AND2X1   g02713(.A(new_n2884_), .B(new_n902_), .Y(new_n2906_));
  AOI21X1  g02714(.A0(new_n2906_), .A1(new_n2905_), .B0(new_n2882_), .Y(new_n2907_));
  OAI21X1  g02715(.A0(new_n2907_), .A1(new_n2904_), .B0(\asqrt[55] ), .Y(new_n2908_));
  INVX1    g02716(.A(new_n2892_), .Y(new_n2909_));
  OAI21X1  g02717(.A0(new_n2866_), .A1(new_n902_), .B0(new_n697_), .Y(new_n2910_));
  OAI21X1  g02718(.A0(new_n2910_), .A1(new_n2907_), .B0(new_n2909_), .Y(new_n2911_));
  NAND3X1  g02719(.A(new_n2911_), .B(new_n2908_), .C(new_n582_), .Y(new_n2912_));
  NAND2X1  g02720(.A(new_n2912_), .B(new_n2899_), .Y(new_n2913_));
  AND2X1   g02721(.A(new_n2672_), .B(new_n2671_), .Y(new_n2914_));
  NOR4X1   g02722(.A(new_n2769_), .B(new_n2914_), .C(new_n2639_), .D(new_n2670_), .Y(new_n2915_));
  AOI22X1  g02723(.A0(new_n2672_), .A1(new_n2671_), .B0(new_n2657_), .B1(\asqrt[56] ), .Y(new_n2916_));
  AOI21X1  g02724(.A0(new_n2916_), .A1(\asqrt[44] ), .B0(new_n2638_), .Y(new_n2917_));
  NOR2X1   g02725(.A(new_n2917_), .B(new_n2915_), .Y(new_n2918_));
  AOI21X1  g02726(.A0(new_n2911_), .A1(new_n2908_), .B0(new_n582_), .Y(new_n2919_));
  NOR2X1   g02727(.A(new_n2919_), .B(\asqrt[57] ), .Y(new_n2920_));
  AOI21X1  g02728(.A0(new_n2920_), .A1(new_n2913_), .B0(new_n2918_), .Y(new_n2921_));
  OAI21X1  g02729(.A0(new_n2921_), .A1(new_n2903_), .B0(\asqrt[58] ), .Y(new_n2922_));
  AND2X1   g02730(.A(new_n2658_), .B(new_n2641_), .Y(new_n2923_));
  OR4X1    g02731(.A(new_n2769_), .B(new_n2923_), .C(new_n2675_), .D(new_n2642_), .Y(new_n2924_));
  OR2X1    g02732(.A(new_n2923_), .B(new_n2642_), .Y(new_n2925_));
  OAI21X1  g02733(.A0(new_n2925_), .A1(new_n2769_), .B0(new_n2675_), .Y(new_n2926_));
  AND2X1   g02734(.A(new_n2926_), .B(new_n2924_), .Y(new_n2927_));
  INVX1    g02735(.A(new_n2927_), .Y(new_n2928_));
  AOI21X1  g02736(.A0(new_n2912_), .A1(new_n2899_), .B0(new_n2919_), .Y(new_n2929_));
  OAI21X1  g02737(.A0(new_n2929_), .A1(new_n481_), .B0(new_n399_), .Y(new_n2930_));
  OAI21X1  g02738(.A0(new_n2930_), .A1(new_n2921_), .B0(new_n2928_), .Y(new_n2931_));
  AOI21X1  g02739(.A0(new_n2931_), .A1(new_n2922_), .B0(new_n328_), .Y(new_n2932_));
  OR4X1    g02740(.A(new_n2769_), .B(new_n2666_), .C(new_n2669_), .D(new_n2685_), .Y(new_n2933_));
  OR2X1    g02741(.A(new_n2666_), .B(new_n2685_), .Y(new_n2934_));
  OAI21X1  g02742(.A0(new_n2934_), .A1(new_n2769_), .B0(new_n2669_), .Y(new_n2935_));
  AND2X1   g02743(.A(new_n2935_), .B(new_n2933_), .Y(new_n2936_));
  INVX1    g02744(.A(new_n2936_), .Y(new_n2937_));
  NAND3X1  g02745(.A(new_n2931_), .B(new_n2922_), .C(new_n328_), .Y(new_n2938_));
  AOI21X1  g02746(.A0(new_n2938_), .A1(new_n2937_), .B0(new_n2932_), .Y(new_n2939_));
  OR2X1    g02747(.A(new_n2939_), .B(new_n292_), .Y(new_n2940_));
  AND2X1   g02748(.A(new_n2938_), .B(new_n2937_), .Y(new_n2941_));
  OAI21X1  g02749(.A0(new_n2729_), .A1(new_n2727_), .B0(new_n2684_), .Y(new_n2942_));
  NOR3X1   g02750(.A(new_n2942_), .B(new_n2769_), .C(new_n2668_), .Y(new_n2943_));
  AOI22X1  g02751(.A0(new_n2686_), .A1(new_n2679_), .B0(new_n2667_), .B1(\asqrt[59] ), .Y(new_n2944_));
  AOI21X1  g02752(.A0(new_n2944_), .A1(\asqrt[44] ), .B0(new_n2684_), .Y(new_n2945_));
  NOR2X1   g02753(.A(new_n2945_), .B(new_n2943_), .Y(new_n2946_));
  INVX1    g02754(.A(new_n2946_), .Y(new_n2947_));
  OR2X1    g02755(.A(new_n2932_), .B(\asqrt[60] ), .Y(new_n2948_));
  OAI21X1  g02756(.A0(new_n2948_), .A1(new_n2941_), .B0(new_n2947_), .Y(new_n2949_));
  AOI21X1  g02757(.A0(new_n2949_), .A1(new_n2940_), .B0(new_n217_), .Y(new_n2950_));
  AND2X1   g02758(.A(new_n2732_), .B(new_n2730_), .Y(new_n2951_));
  NOR4X1   g02759(.A(new_n2769_), .B(new_n2951_), .C(new_n2693_), .D(new_n2731_), .Y(new_n2952_));
  NOR2X1   g02760(.A(new_n2951_), .B(new_n2731_), .Y(new_n2953_));
  AOI21X1  g02761(.A0(new_n2953_), .A1(\asqrt[44] ), .B0(new_n2692_), .Y(new_n2954_));
  NOR2X1   g02762(.A(new_n2954_), .B(new_n2952_), .Y(new_n2955_));
  OR2X1    g02763(.A(new_n2929_), .B(new_n481_), .Y(new_n2956_));
  AND2X1   g02764(.A(new_n2912_), .B(new_n2899_), .Y(new_n2957_));
  INVX1    g02765(.A(new_n2918_), .Y(new_n2958_));
  OR2X1    g02766(.A(new_n2919_), .B(\asqrt[57] ), .Y(new_n2959_));
  OAI21X1  g02767(.A0(new_n2959_), .A1(new_n2957_), .B0(new_n2958_), .Y(new_n2960_));
  AOI21X1  g02768(.A0(new_n2960_), .A1(new_n2956_), .B0(new_n399_), .Y(new_n2961_));
  AOI21X1  g02769(.A0(new_n2902_), .A1(\asqrt[57] ), .B0(\asqrt[58] ), .Y(new_n2962_));
  AOI21X1  g02770(.A0(new_n2962_), .A1(new_n2960_), .B0(new_n2927_), .Y(new_n2963_));
  OAI21X1  g02771(.A0(new_n2963_), .A1(new_n2961_), .B0(\asqrt[59] ), .Y(new_n2964_));
  NOR3X1   g02772(.A(new_n2963_), .B(new_n2961_), .C(\asqrt[59] ), .Y(new_n2965_));
  OAI21X1  g02773(.A0(new_n2965_), .A1(new_n2936_), .B0(new_n2964_), .Y(new_n2966_));
  AOI21X1  g02774(.A0(new_n2966_), .A1(\asqrt[60] ), .B0(\asqrt[61] ), .Y(new_n2967_));
  AOI21X1  g02775(.A0(new_n2967_), .A1(new_n2949_), .B0(new_n2955_), .Y(new_n2968_));
  OAI21X1  g02776(.A0(new_n2968_), .A1(new_n2950_), .B0(\asqrt[62] ), .Y(new_n2969_));
  NAND3X1  g02777(.A(new_n2704_), .B(new_n2702_), .C(new_n2734_), .Y(new_n2970_));
  NOR3X1   g02778(.A(new_n2769_), .B(new_n2735_), .C(new_n2697_), .Y(new_n2971_));
  OAI22X1  g02779(.A0(new_n2971_), .A1(new_n2702_), .B0(new_n2970_), .B1(new_n2769_), .Y(new_n2972_));
  INVX1    g02780(.A(new_n2972_), .Y(new_n2973_));
  NOR3X1   g02781(.A(new_n2968_), .B(new_n2950_), .C(\asqrt[62] ), .Y(new_n2974_));
  OAI21X1  g02782(.A0(new_n2974_), .A1(new_n2973_), .B0(new_n2969_), .Y(new_n2975_));
  AND2X1   g02783(.A(new_n2764_), .B(new_n2763_), .Y(new_n2976_));
  NOR4X1   g02784(.A(new_n2769_), .B(new_n2976_), .C(new_n2713_), .D(new_n2762_), .Y(new_n2977_));
  INVX1    g02785(.A(new_n2977_), .Y(new_n2978_));
  OAI22X1  g02786(.A0(new_n2714_), .A1(new_n2707_), .B0(new_n2705_), .B1(new_n199_), .Y(new_n2979_));
  OAI21X1  g02787(.A0(new_n2979_), .A1(new_n2769_), .B0(new_n2713_), .Y(new_n2980_));
  AND2X1   g02788(.A(new_n2980_), .B(new_n2978_), .Y(new_n2981_));
  INVX1    g02789(.A(new_n2981_), .Y(new_n2982_));
  AND2X1   g02790(.A(new_n2737_), .B(new_n2715_), .Y(new_n2983_));
  AOI21X1  g02791(.A0(new_n2715_), .A1(new_n2706_), .B0(new_n2719_), .Y(new_n2984_));
  AOI21X1  g02792(.A0(new_n2984_), .A1(\asqrt[44] ), .B0(new_n2983_), .Y(new_n2985_));
  AND2X1   g02793(.A(new_n2985_), .B(new_n2982_), .Y(new_n2986_));
  AOI21X1  g02794(.A0(new_n2986_), .A1(new_n2975_), .B0(\asqrt[63] ), .Y(new_n2987_));
  AND2X1   g02795(.A(new_n2966_), .B(\asqrt[60] ), .Y(new_n2988_));
  NAND2X1  g02796(.A(new_n2938_), .B(new_n2937_), .Y(new_n2989_));
  NOR2X1   g02797(.A(new_n2932_), .B(\asqrt[60] ), .Y(new_n2990_));
  AOI21X1  g02798(.A0(new_n2990_), .A1(new_n2989_), .B0(new_n2946_), .Y(new_n2991_));
  OAI21X1  g02799(.A0(new_n2991_), .A1(new_n2988_), .B0(\asqrt[61] ), .Y(new_n2992_));
  INVX1    g02800(.A(new_n2955_), .Y(new_n2993_));
  OAI21X1  g02801(.A0(new_n2939_), .A1(new_n292_), .B0(new_n217_), .Y(new_n2994_));
  OAI21X1  g02802(.A0(new_n2994_), .A1(new_n2991_), .B0(new_n2993_), .Y(new_n2995_));
  NAND3X1  g02803(.A(new_n2995_), .B(new_n2992_), .C(new_n199_), .Y(new_n2996_));
  AND2X1   g02804(.A(new_n2996_), .B(new_n2972_), .Y(new_n2997_));
  NAND2X1  g02805(.A(new_n2981_), .B(new_n2969_), .Y(new_n2998_));
  NAND2X1  g02806(.A(new_n2715_), .B(new_n2706_), .Y(new_n2999_));
  AOI21X1  g02807(.A0(\asqrt[44] ), .A1(new_n2720_), .B0(new_n2999_), .Y(new_n3000_));
  NOR3X1   g02808(.A(new_n3000_), .B(new_n2984_), .C(new_n193_), .Y(new_n3001_));
  AND2X1   g02809(.A(new_n2766_), .B(new_n193_), .Y(new_n3002_));
  NAND4X1  g02810(.A(new_n2744_), .B(new_n2740_), .C(new_n2718_), .D(new_n2716_), .Y(new_n3003_));
  OR2X1    g02811(.A(new_n3003_), .B(new_n2983_), .Y(new_n3004_));
  NOR2X1   g02812(.A(new_n3004_), .B(new_n3002_), .Y(new_n3005_));
  NOR2X1   g02813(.A(new_n3005_), .B(new_n3001_), .Y(new_n3006_));
  OAI21X1  g02814(.A0(new_n2998_), .A1(new_n2997_), .B0(new_n3006_), .Y(new_n3007_));
  NOR2X1   g02815(.A(new_n3007_), .B(new_n2987_), .Y(new_n3008_));
  INVX1    g02816(.A(\a[86] ), .Y(new_n3009_));
  NOR2X1   g02817(.A(\a[85] ), .B(\a[84] ), .Y(new_n3010_));
  NAND2X1  g02818(.A(new_n3010_), .B(new_n3009_), .Y(new_n3011_));
  OAI21X1  g02819(.A0(new_n3008_), .A1(new_n3009_), .B0(new_n3011_), .Y(new_n3012_));
  AOI21X1  g02820(.A0(new_n2995_), .A1(new_n2992_), .B0(new_n199_), .Y(new_n3013_));
  AOI21X1  g02821(.A0(new_n2996_), .A1(new_n2972_), .B0(new_n3013_), .Y(new_n3014_));
  INVX1    g02822(.A(new_n2986_), .Y(new_n3015_));
  OAI21X1  g02823(.A0(new_n3015_), .A1(new_n3014_), .B0(new_n193_), .Y(new_n3016_));
  NAND2X1  g02824(.A(new_n2996_), .B(new_n2972_), .Y(new_n3017_));
  AND2X1   g02825(.A(new_n2981_), .B(new_n2969_), .Y(new_n3018_));
  INVX1    g02826(.A(new_n3006_), .Y(new_n3019_));
  AOI21X1  g02827(.A0(new_n3018_), .A1(new_n3017_), .B0(new_n3019_), .Y(new_n3020_));
  AOI21X1  g02828(.A0(new_n3020_), .A1(new_n3016_), .B0(new_n3009_), .Y(new_n3021_));
  NAND3X1  g02829(.A(new_n3011_), .B(new_n2744_), .C(new_n2740_), .Y(new_n3022_));
  OR4X1    g02830(.A(new_n3022_), .B(new_n3021_), .C(new_n2983_), .D(new_n3002_), .Y(new_n3023_));
  OAI21X1  g02831(.A0(new_n3007_), .A1(new_n2987_), .B0(new_n3009_), .Y(new_n3024_));
  AOI21X1  g02832(.A0(new_n3020_), .A1(new_n3016_), .B0(new_n2770_), .Y(new_n3025_));
  AOI21X1  g02833(.A0(new_n3024_), .A1(\a[87] ), .B0(new_n3025_), .Y(new_n3026_));
  AOI22X1  g02834(.A0(new_n3026_), .A1(new_n3023_), .B0(new_n3012_), .B1(\asqrt[44] ), .Y(new_n3027_));
  OR2X1    g02835(.A(new_n3027_), .B(new_n2570_), .Y(new_n3028_));
  AND2X1   g02836(.A(new_n3026_), .B(new_n3023_), .Y(new_n3029_));
  INVX1    g02837(.A(new_n3010_), .Y(new_n3030_));
  MX2X1    g02838(.A(new_n3030_), .B(new_n3008_), .S0(\a[86] ), .Y(new_n3031_));
  OAI21X1  g02839(.A0(new_n3031_), .A1(new_n2769_), .B0(new_n2570_), .Y(new_n3032_));
  OAI21X1  g02840(.A0(new_n3007_), .A1(new_n2987_), .B0(new_n2749_), .Y(new_n3033_));
  AND2X1   g02841(.A(new_n3018_), .B(new_n3017_), .Y(new_n3034_));
  OAI21X1  g02842(.A0(new_n3004_), .A1(new_n3002_), .B0(\asqrt[44] ), .Y(new_n3035_));
  OR4X1    g02843(.A(new_n3035_), .B(new_n3001_), .C(new_n3034_), .D(new_n2987_), .Y(new_n3036_));
  AOI21X1  g02844(.A0(new_n3036_), .A1(new_n3033_), .B0(new_n2756_), .Y(new_n3037_));
  NOR4X1   g02845(.A(new_n3035_), .B(new_n3001_), .C(new_n3034_), .D(new_n2987_), .Y(new_n3038_));
  NOR3X1   g02846(.A(new_n3038_), .B(new_n3025_), .C(\a[88] ), .Y(new_n3039_));
  OR2X1    g02847(.A(new_n3039_), .B(new_n3037_), .Y(new_n3040_));
  OAI21X1  g02848(.A0(new_n3032_), .A1(new_n3029_), .B0(new_n3040_), .Y(new_n3041_));
  AOI21X1  g02849(.A0(new_n3041_), .A1(new_n3028_), .B0(new_n2263_), .Y(new_n3042_));
  AND2X1   g02850(.A(new_n2811_), .B(new_n2809_), .Y(new_n3043_));
  NOR3X1   g02851(.A(new_n3043_), .B(new_n2755_), .C(new_n2751_), .Y(new_n3044_));
  OAI21X1  g02852(.A0(new_n3007_), .A1(new_n2987_), .B0(new_n3044_), .Y(new_n3045_));
  AOI21X1  g02853(.A0(new_n2750_), .A1(\asqrt[45] ), .B0(new_n2755_), .Y(new_n3046_));
  OAI21X1  g02854(.A0(new_n3007_), .A1(new_n2987_), .B0(new_n3046_), .Y(new_n3047_));
  NAND2X1  g02855(.A(new_n3047_), .B(new_n3043_), .Y(new_n3048_));
  NOR4X1   g02856(.A(new_n3022_), .B(new_n3021_), .C(new_n2983_), .D(new_n3002_), .Y(new_n3049_));
  INVX1    g02857(.A(\a[87] ), .Y(new_n3050_));
  AOI21X1  g02858(.A0(new_n3020_), .A1(new_n3016_), .B0(\a[86] ), .Y(new_n3051_));
  OAI21X1  g02859(.A0(new_n3051_), .A1(new_n3050_), .B0(new_n3033_), .Y(new_n3052_));
  OAI22X1  g02860(.A0(new_n3052_), .A1(new_n3049_), .B0(new_n3031_), .B1(new_n2769_), .Y(new_n3053_));
  AOI21X1  g02861(.A0(new_n3053_), .A1(\asqrt[45] ), .B0(\asqrt[46] ), .Y(new_n3054_));
  AOI22X1  g02862(.A0(new_n3054_), .A1(new_n3041_), .B0(new_n3048_), .B1(new_n3045_), .Y(new_n3055_));
  OAI21X1  g02863(.A0(new_n3055_), .A1(new_n3042_), .B0(\asqrt[47] ), .Y(new_n3056_));
  AND2X1   g02864(.A(new_n2814_), .B(new_n2812_), .Y(new_n3057_));
  NOR3X1   g02865(.A(new_n2779_), .B(new_n3057_), .C(new_n2813_), .Y(new_n3058_));
  OAI21X1  g02866(.A0(new_n3007_), .A1(new_n2987_), .B0(new_n3058_), .Y(new_n3059_));
  NOR2X1   g02867(.A(new_n3057_), .B(new_n2813_), .Y(new_n3060_));
  OAI21X1  g02868(.A0(new_n3007_), .A1(new_n2987_), .B0(new_n3060_), .Y(new_n3061_));
  NAND2X1  g02869(.A(new_n3061_), .B(new_n2779_), .Y(new_n3062_));
  AND2X1   g02870(.A(new_n3062_), .B(new_n3059_), .Y(new_n3063_));
  NOR3X1   g02871(.A(new_n3055_), .B(new_n3042_), .C(\asqrt[47] ), .Y(new_n3064_));
  OAI21X1  g02872(.A0(new_n3064_), .A1(new_n3063_), .B0(new_n3056_), .Y(new_n3065_));
  AND2X1   g02873(.A(new_n3065_), .B(\asqrt[48] ), .Y(new_n3066_));
  OR2X1    g02874(.A(new_n3064_), .B(new_n3063_), .Y(new_n3067_));
  NOR3X1   g02875(.A(new_n2819_), .B(new_n2787_), .C(new_n2781_), .Y(new_n3068_));
  OAI21X1  g02876(.A0(new_n3007_), .A1(new_n2987_), .B0(new_n3068_), .Y(new_n3069_));
  NOR3X1   g02877(.A(new_n3008_), .B(new_n2819_), .C(new_n2781_), .Y(new_n3070_));
  OR2X1    g02878(.A(new_n3070_), .B(new_n2786_), .Y(new_n3071_));
  AND2X1   g02879(.A(new_n3071_), .B(new_n3069_), .Y(new_n3072_));
  AND2X1   g02880(.A(new_n3053_), .B(\asqrt[45] ), .Y(new_n3073_));
  NAND2X1  g02881(.A(new_n3026_), .B(new_n3023_), .Y(new_n3074_));
  AOI21X1  g02882(.A0(new_n3012_), .A1(\asqrt[44] ), .B0(\asqrt[45] ), .Y(new_n3075_));
  NOR2X1   g02883(.A(new_n3039_), .B(new_n3037_), .Y(new_n3076_));
  AOI21X1  g02884(.A0(new_n3075_), .A1(new_n3074_), .B0(new_n3076_), .Y(new_n3077_));
  OAI21X1  g02885(.A0(new_n3077_), .A1(new_n3073_), .B0(\asqrt[46] ), .Y(new_n3078_));
  NAND2X1  g02886(.A(new_n3048_), .B(new_n3045_), .Y(new_n3079_));
  OAI21X1  g02887(.A0(new_n3027_), .A1(new_n2570_), .B0(new_n2263_), .Y(new_n3080_));
  OAI21X1  g02888(.A0(new_n3080_), .A1(new_n3077_), .B0(new_n3079_), .Y(new_n3081_));
  AOI21X1  g02889(.A0(new_n3081_), .A1(new_n3078_), .B0(new_n2040_), .Y(new_n3082_));
  NOR2X1   g02890(.A(new_n3082_), .B(\asqrt[48] ), .Y(new_n3083_));
  AOI21X1  g02891(.A0(new_n3083_), .A1(new_n3067_), .B0(new_n3072_), .Y(new_n3084_));
  OAI21X1  g02892(.A0(new_n3084_), .A1(new_n3066_), .B0(\asqrt[49] ), .Y(new_n3085_));
  INVX1    g02893(.A(new_n3008_), .Y(\asqrt[43] ));
  AOI21X1  g02894(.A0(new_n2833_), .A1(new_n2832_), .B0(new_n2797_), .Y(new_n3087_));
  AND2X1   g02895(.A(new_n3087_), .B(new_n2790_), .Y(new_n3088_));
  AOI22X1  g02896(.A0(new_n2833_), .A1(new_n2832_), .B0(new_n2820_), .B1(\asqrt[48] ), .Y(new_n3089_));
  AOI21X1  g02897(.A0(new_n3089_), .A1(\asqrt[43] ), .B0(new_n2796_), .Y(new_n3090_));
  AOI21X1  g02898(.A0(new_n3088_), .A1(\asqrt[43] ), .B0(new_n3090_), .Y(new_n3091_));
  INVX1    g02899(.A(new_n3091_), .Y(new_n3092_));
  INVX1    g02900(.A(new_n3063_), .Y(new_n3093_));
  NAND3X1  g02901(.A(new_n3081_), .B(new_n3078_), .C(new_n2040_), .Y(new_n3094_));
  AOI21X1  g02902(.A0(new_n3094_), .A1(new_n3093_), .B0(new_n3082_), .Y(new_n3095_));
  OAI21X1  g02903(.A0(new_n3095_), .A1(new_n1834_), .B0(new_n1632_), .Y(new_n3096_));
  OAI21X1  g02904(.A0(new_n3096_), .A1(new_n3084_), .B0(new_n3092_), .Y(new_n3097_));
  AOI21X1  g02905(.A0(new_n3097_), .A1(new_n3085_), .B0(new_n1469_), .Y(new_n3098_));
  AND2X1   g02906(.A(new_n2821_), .B(new_n2799_), .Y(new_n3099_));
  NOR3X1   g02907(.A(new_n3099_), .B(new_n2836_), .C(new_n2800_), .Y(new_n3100_));
  NOR3X1   g02908(.A(new_n3008_), .B(new_n3099_), .C(new_n2800_), .Y(new_n3101_));
  NOR2X1   g02909(.A(new_n3101_), .B(new_n2805_), .Y(new_n3102_));
  AOI21X1  g02910(.A0(new_n3100_), .A1(\asqrt[43] ), .B0(new_n3102_), .Y(new_n3103_));
  INVX1    g02911(.A(new_n3103_), .Y(new_n3104_));
  NAND3X1  g02912(.A(new_n3097_), .B(new_n3085_), .C(new_n1469_), .Y(new_n3105_));
  AOI21X1  g02913(.A0(new_n3105_), .A1(new_n3104_), .B0(new_n3098_), .Y(new_n3106_));
  OR2X1    g02914(.A(new_n3106_), .B(new_n1277_), .Y(new_n3107_));
  OR2X1    g02915(.A(new_n3095_), .B(new_n1834_), .Y(new_n3108_));
  NOR2X1   g02916(.A(new_n3064_), .B(new_n3063_), .Y(new_n3109_));
  INVX1    g02917(.A(new_n3072_), .Y(new_n3110_));
  OR2X1    g02918(.A(new_n3082_), .B(\asqrt[48] ), .Y(new_n3111_));
  OAI21X1  g02919(.A0(new_n3111_), .A1(new_n3109_), .B0(new_n3110_), .Y(new_n3112_));
  AOI21X1  g02920(.A0(new_n3112_), .A1(new_n3108_), .B0(new_n1632_), .Y(new_n3113_));
  AOI21X1  g02921(.A0(new_n3065_), .A1(\asqrt[48] ), .B0(\asqrt[49] ), .Y(new_n3114_));
  AOI21X1  g02922(.A0(new_n3114_), .A1(new_n3112_), .B0(new_n3091_), .Y(new_n3115_));
  NOR3X1   g02923(.A(new_n3115_), .B(new_n3113_), .C(\asqrt[50] ), .Y(new_n3116_));
  NOR2X1   g02924(.A(new_n3116_), .B(new_n3103_), .Y(new_n3117_));
  OR4X1    g02925(.A(new_n3008_), .B(new_n2828_), .C(new_n2826_), .D(new_n2846_), .Y(new_n3118_));
  NAND2X1  g02926(.A(new_n2839_), .B(new_n2823_), .Y(new_n3119_));
  OAI21X1  g02927(.A0(new_n3119_), .A1(new_n3008_), .B0(new_n2826_), .Y(new_n3120_));
  AND2X1   g02928(.A(new_n3120_), .B(new_n3118_), .Y(new_n3121_));
  INVX1    g02929(.A(new_n3121_), .Y(new_n3122_));
  OAI21X1  g02930(.A0(new_n3115_), .A1(new_n3113_), .B0(\asqrt[50] ), .Y(new_n3123_));
  NAND2X1  g02931(.A(new_n3123_), .B(new_n1277_), .Y(new_n3124_));
  OAI21X1  g02932(.A0(new_n3124_), .A1(new_n3117_), .B0(new_n3122_), .Y(new_n3125_));
  AOI21X1  g02933(.A0(new_n3125_), .A1(new_n3107_), .B0(new_n1111_), .Y(new_n3126_));
  AND2X1   g02934(.A(new_n2847_), .B(new_n2840_), .Y(new_n3127_));
  NOR3X1   g02935(.A(new_n3127_), .B(new_n2870_), .C(new_n2830_), .Y(new_n3128_));
  NOR3X1   g02936(.A(new_n3008_), .B(new_n3127_), .C(new_n2830_), .Y(new_n3129_));
  NOR2X1   g02937(.A(new_n3129_), .B(new_n2845_), .Y(new_n3130_));
  AOI21X1  g02938(.A0(new_n3128_), .A1(\asqrt[43] ), .B0(new_n3130_), .Y(new_n3131_));
  OAI21X1  g02939(.A0(new_n3116_), .A1(new_n3103_), .B0(new_n3123_), .Y(new_n3132_));
  AOI21X1  g02940(.A0(new_n3132_), .A1(\asqrt[51] ), .B0(\asqrt[52] ), .Y(new_n3133_));
  AOI21X1  g02941(.A0(new_n3133_), .A1(new_n3125_), .B0(new_n3131_), .Y(new_n3134_));
  OAI21X1  g02942(.A0(new_n3134_), .A1(new_n3126_), .B0(\asqrt[53] ), .Y(new_n3135_));
  AND2X1   g02943(.A(new_n2874_), .B(new_n2872_), .Y(new_n3136_));
  NOR3X1   g02944(.A(new_n3136_), .B(new_n2855_), .C(new_n2873_), .Y(new_n3137_));
  NOR3X1   g02945(.A(new_n3008_), .B(new_n3136_), .C(new_n2873_), .Y(new_n3138_));
  NOR2X1   g02946(.A(new_n3138_), .B(new_n2854_), .Y(new_n3139_));
  AOI21X1  g02947(.A0(new_n3137_), .A1(\asqrt[43] ), .B0(new_n3139_), .Y(new_n3140_));
  NOR3X1   g02948(.A(new_n3134_), .B(new_n3126_), .C(\asqrt[53] ), .Y(new_n3141_));
  OAI21X1  g02949(.A0(new_n3141_), .A1(new_n3140_), .B0(new_n3135_), .Y(new_n3142_));
  AND2X1   g02950(.A(new_n3142_), .B(\asqrt[54] ), .Y(new_n3143_));
  INVX1    g02951(.A(new_n3140_), .Y(new_n3144_));
  AND2X1   g02952(.A(new_n3132_), .B(\asqrt[51] ), .Y(new_n3145_));
  OR2X1    g02953(.A(new_n3116_), .B(new_n3103_), .Y(new_n3146_));
  AND2X1   g02954(.A(new_n3123_), .B(new_n1277_), .Y(new_n3147_));
  AOI21X1  g02955(.A0(new_n3147_), .A1(new_n3146_), .B0(new_n3121_), .Y(new_n3148_));
  OAI21X1  g02956(.A0(new_n3148_), .A1(new_n3145_), .B0(\asqrt[52] ), .Y(new_n3149_));
  INVX1    g02957(.A(new_n3131_), .Y(new_n3150_));
  OAI21X1  g02958(.A0(new_n3106_), .A1(new_n1277_), .B0(new_n1111_), .Y(new_n3151_));
  OAI21X1  g02959(.A0(new_n3151_), .A1(new_n3148_), .B0(new_n3150_), .Y(new_n3152_));
  NAND3X1  g02960(.A(new_n3152_), .B(new_n3149_), .C(new_n968_), .Y(new_n3153_));
  NAND2X1  g02961(.A(new_n3153_), .B(new_n3144_), .Y(new_n3154_));
  AOI21X1  g02962(.A0(new_n3152_), .A1(new_n3149_), .B0(new_n968_), .Y(new_n3155_));
  NOR2X1   g02963(.A(new_n3155_), .B(\asqrt[54] ), .Y(new_n3156_));
  OR4X1    g02964(.A(new_n3008_), .B(new_n2865_), .C(new_n2876_), .D(new_n2859_), .Y(new_n3157_));
  OR2X1    g02965(.A(new_n2876_), .B(new_n2859_), .Y(new_n3158_));
  OAI21X1  g02966(.A0(new_n3158_), .A1(new_n3008_), .B0(new_n2865_), .Y(new_n3159_));
  AND2X1   g02967(.A(new_n3159_), .B(new_n3157_), .Y(new_n3160_));
  AOI21X1  g02968(.A0(new_n3156_), .A1(new_n3154_), .B0(new_n3160_), .Y(new_n3161_));
  OAI21X1  g02969(.A0(new_n3161_), .A1(new_n3143_), .B0(\asqrt[55] ), .Y(new_n3162_));
  AOI21X1  g02970(.A0(new_n2906_), .A1(new_n2905_), .B0(new_n2883_), .Y(new_n3163_));
  AND2X1   g02971(.A(new_n3163_), .B(new_n2867_), .Y(new_n3164_));
  AOI22X1  g02972(.A0(new_n2906_), .A1(new_n2905_), .B0(new_n2893_), .B1(\asqrt[54] ), .Y(new_n3165_));
  AOI21X1  g02973(.A0(new_n3165_), .A1(\asqrt[43] ), .B0(new_n2882_), .Y(new_n3166_));
  AOI21X1  g02974(.A0(new_n3164_), .A1(\asqrt[43] ), .B0(new_n3166_), .Y(new_n3167_));
  INVX1    g02975(.A(new_n3167_), .Y(new_n3168_));
  AOI21X1  g02976(.A0(new_n3153_), .A1(new_n3144_), .B0(new_n3155_), .Y(new_n3169_));
  OAI21X1  g02977(.A0(new_n3169_), .A1(new_n902_), .B0(new_n697_), .Y(new_n3170_));
  OAI21X1  g02978(.A0(new_n3170_), .A1(new_n3161_), .B0(new_n3168_), .Y(new_n3171_));
  AOI21X1  g02979(.A0(new_n3171_), .A1(new_n3162_), .B0(new_n582_), .Y(new_n3172_));
  AND2X1   g02980(.A(new_n2894_), .B(new_n2886_), .Y(new_n3173_));
  NOR3X1   g02981(.A(new_n3173_), .B(new_n2909_), .C(new_n2887_), .Y(new_n3174_));
  NOR3X1   g02982(.A(new_n3008_), .B(new_n3173_), .C(new_n2887_), .Y(new_n3175_));
  NOR2X1   g02983(.A(new_n3175_), .B(new_n2892_), .Y(new_n3176_));
  AOI21X1  g02984(.A0(new_n3174_), .A1(\asqrt[43] ), .B0(new_n3176_), .Y(new_n3177_));
  INVX1    g02985(.A(new_n3177_), .Y(new_n3178_));
  NAND3X1  g02986(.A(new_n3171_), .B(new_n3162_), .C(new_n582_), .Y(new_n3179_));
  AOI21X1  g02987(.A0(new_n3179_), .A1(new_n3178_), .B0(new_n3172_), .Y(new_n3180_));
  OR2X1    g02988(.A(new_n3180_), .B(new_n481_), .Y(new_n3181_));
  AND2X1   g02989(.A(new_n3179_), .B(new_n3178_), .Y(new_n3182_));
  OR4X1    g02990(.A(new_n3008_), .B(new_n2901_), .C(new_n2899_), .D(new_n2919_), .Y(new_n3183_));
  NAND2X1  g02991(.A(new_n2912_), .B(new_n2896_), .Y(new_n3184_));
  OAI21X1  g02992(.A0(new_n3184_), .A1(new_n3008_), .B0(new_n2899_), .Y(new_n3185_));
  AND2X1   g02993(.A(new_n3185_), .B(new_n3183_), .Y(new_n3186_));
  INVX1    g02994(.A(new_n3186_), .Y(new_n3187_));
  OR2X1    g02995(.A(new_n3172_), .B(\asqrt[57] ), .Y(new_n3188_));
  OAI21X1  g02996(.A0(new_n3188_), .A1(new_n3182_), .B0(new_n3187_), .Y(new_n3189_));
  AOI21X1  g02997(.A0(new_n3189_), .A1(new_n3181_), .B0(new_n399_), .Y(new_n3190_));
  AND2X1   g02998(.A(new_n2920_), .B(new_n2913_), .Y(new_n3191_));
  NOR3X1   g02999(.A(new_n3191_), .B(new_n2958_), .C(new_n2903_), .Y(new_n3192_));
  NOR3X1   g03000(.A(new_n3008_), .B(new_n3191_), .C(new_n2903_), .Y(new_n3193_));
  NOR2X1   g03001(.A(new_n3193_), .B(new_n2918_), .Y(new_n3194_));
  AOI21X1  g03002(.A0(new_n3192_), .A1(\asqrt[43] ), .B0(new_n3194_), .Y(new_n3195_));
  OR2X1    g03003(.A(new_n3169_), .B(new_n902_), .Y(new_n3196_));
  AND2X1   g03004(.A(new_n3153_), .B(new_n3144_), .Y(new_n3197_));
  OR2X1    g03005(.A(new_n3155_), .B(\asqrt[54] ), .Y(new_n3198_));
  INVX1    g03006(.A(new_n3160_), .Y(new_n3199_));
  OAI21X1  g03007(.A0(new_n3198_), .A1(new_n3197_), .B0(new_n3199_), .Y(new_n3200_));
  AOI21X1  g03008(.A0(new_n3200_), .A1(new_n3196_), .B0(new_n697_), .Y(new_n3201_));
  AOI21X1  g03009(.A0(new_n3142_), .A1(\asqrt[54] ), .B0(\asqrt[55] ), .Y(new_n3202_));
  AOI21X1  g03010(.A0(new_n3202_), .A1(new_n3200_), .B0(new_n3167_), .Y(new_n3203_));
  OAI21X1  g03011(.A0(new_n3203_), .A1(new_n3201_), .B0(\asqrt[56] ), .Y(new_n3204_));
  NOR3X1   g03012(.A(new_n3203_), .B(new_n3201_), .C(\asqrt[56] ), .Y(new_n3205_));
  OAI21X1  g03013(.A0(new_n3205_), .A1(new_n3177_), .B0(new_n3204_), .Y(new_n3206_));
  AOI21X1  g03014(.A0(new_n3206_), .A1(\asqrt[57] ), .B0(\asqrt[58] ), .Y(new_n3207_));
  AOI21X1  g03015(.A0(new_n3207_), .A1(new_n3189_), .B0(new_n3195_), .Y(new_n3208_));
  OAI21X1  g03016(.A0(new_n3208_), .A1(new_n3190_), .B0(\asqrt[59] ), .Y(new_n3209_));
  AND2X1   g03017(.A(new_n2962_), .B(new_n2960_), .Y(new_n3210_));
  NOR3X1   g03018(.A(new_n3210_), .B(new_n2928_), .C(new_n2961_), .Y(new_n3211_));
  NOR3X1   g03019(.A(new_n3008_), .B(new_n3210_), .C(new_n2961_), .Y(new_n3212_));
  NOR2X1   g03020(.A(new_n3212_), .B(new_n2927_), .Y(new_n3213_));
  AOI21X1  g03021(.A0(new_n3211_), .A1(\asqrt[43] ), .B0(new_n3213_), .Y(new_n3214_));
  NOR3X1   g03022(.A(new_n3208_), .B(new_n3190_), .C(\asqrt[59] ), .Y(new_n3215_));
  OAI21X1  g03023(.A0(new_n3215_), .A1(new_n3214_), .B0(new_n3209_), .Y(new_n3216_));
  AND2X1   g03024(.A(new_n3216_), .B(\asqrt[60] ), .Y(new_n3217_));
  INVX1    g03025(.A(new_n3214_), .Y(new_n3218_));
  AND2X1   g03026(.A(new_n3206_), .B(\asqrt[57] ), .Y(new_n3219_));
  NAND2X1  g03027(.A(new_n3179_), .B(new_n3178_), .Y(new_n3220_));
  NOR2X1   g03028(.A(new_n3172_), .B(\asqrt[57] ), .Y(new_n3221_));
  AOI21X1  g03029(.A0(new_n3221_), .A1(new_n3220_), .B0(new_n3186_), .Y(new_n3222_));
  OAI21X1  g03030(.A0(new_n3222_), .A1(new_n3219_), .B0(\asqrt[58] ), .Y(new_n3223_));
  INVX1    g03031(.A(new_n3195_), .Y(new_n3224_));
  OAI21X1  g03032(.A0(new_n3180_), .A1(new_n481_), .B0(new_n399_), .Y(new_n3225_));
  OAI21X1  g03033(.A0(new_n3225_), .A1(new_n3222_), .B0(new_n3224_), .Y(new_n3226_));
  NAND3X1  g03034(.A(new_n3226_), .B(new_n3223_), .C(new_n328_), .Y(new_n3227_));
  NAND2X1  g03035(.A(new_n3227_), .B(new_n3218_), .Y(new_n3228_));
  NAND4X1  g03036(.A(\asqrt[43] ), .B(new_n2938_), .C(new_n2936_), .D(new_n2964_), .Y(new_n3229_));
  NAND2X1  g03037(.A(new_n2938_), .B(new_n2964_), .Y(new_n3230_));
  OAI21X1  g03038(.A0(new_n3230_), .A1(new_n3008_), .B0(new_n2937_), .Y(new_n3231_));
  AND2X1   g03039(.A(new_n3231_), .B(new_n3229_), .Y(new_n3232_));
  AOI21X1  g03040(.A0(new_n3226_), .A1(new_n3223_), .B0(new_n328_), .Y(new_n3233_));
  NOR2X1   g03041(.A(new_n3233_), .B(\asqrt[60] ), .Y(new_n3234_));
  AOI21X1  g03042(.A0(new_n3234_), .A1(new_n3228_), .B0(new_n3232_), .Y(new_n3235_));
  OAI21X1  g03043(.A0(new_n3235_), .A1(new_n3217_), .B0(\asqrt[61] ), .Y(new_n3236_));
  AOI21X1  g03044(.A0(new_n2990_), .A1(new_n2989_), .B0(new_n2947_), .Y(new_n3237_));
  AND2X1   g03045(.A(new_n3237_), .B(new_n2940_), .Y(new_n3238_));
  AOI22X1  g03046(.A0(new_n2990_), .A1(new_n2989_), .B0(new_n2966_), .B1(\asqrt[60] ), .Y(new_n3239_));
  AOI21X1  g03047(.A0(new_n3239_), .A1(\asqrt[43] ), .B0(new_n2946_), .Y(new_n3240_));
  AOI21X1  g03048(.A0(new_n3238_), .A1(\asqrt[43] ), .B0(new_n3240_), .Y(new_n3241_));
  INVX1    g03049(.A(new_n3241_), .Y(new_n3242_));
  AOI21X1  g03050(.A0(new_n3227_), .A1(new_n3218_), .B0(new_n3233_), .Y(new_n3243_));
  OAI21X1  g03051(.A0(new_n3243_), .A1(new_n292_), .B0(new_n217_), .Y(new_n3244_));
  OAI21X1  g03052(.A0(new_n3244_), .A1(new_n3235_), .B0(new_n3242_), .Y(new_n3245_));
  AOI21X1  g03053(.A0(new_n3245_), .A1(new_n3236_), .B0(new_n199_), .Y(new_n3246_));
  AND2X1   g03054(.A(new_n2967_), .B(new_n2949_), .Y(new_n3247_));
  NOR3X1   g03055(.A(new_n3247_), .B(new_n2993_), .C(new_n2950_), .Y(new_n3248_));
  NOR3X1   g03056(.A(new_n3008_), .B(new_n3247_), .C(new_n2950_), .Y(new_n3249_));
  NOR2X1   g03057(.A(new_n3249_), .B(new_n2955_), .Y(new_n3250_));
  AOI21X1  g03058(.A0(new_n3248_), .A1(\asqrt[43] ), .B0(new_n3250_), .Y(new_n3251_));
  INVX1    g03059(.A(new_n3251_), .Y(new_n3252_));
  NAND3X1  g03060(.A(new_n3245_), .B(new_n3236_), .C(new_n199_), .Y(new_n3253_));
  AOI21X1  g03061(.A0(new_n3253_), .A1(new_n3252_), .B0(new_n3246_), .Y(new_n3254_));
  NOR4X1   g03062(.A(new_n3008_), .B(new_n2974_), .C(new_n2972_), .D(new_n3013_), .Y(new_n3255_));
  NAND3X1  g03063(.A(\asqrt[43] ), .B(new_n2996_), .C(new_n2969_), .Y(new_n3256_));
  AOI21X1  g03064(.A0(new_n3256_), .A1(new_n2972_), .B0(new_n3255_), .Y(new_n3257_));
  NOR3X1   g03065(.A(new_n3008_), .B(new_n2981_), .C(new_n3014_), .Y(new_n3258_));
  NOR3X1   g03066(.A(new_n3258_), .B(new_n3257_), .C(new_n3034_), .Y(new_n3259_));
  INVX1    g03067(.A(new_n3259_), .Y(new_n3260_));
  OAI21X1  g03068(.A0(new_n3260_), .A1(new_n3254_), .B0(new_n193_), .Y(new_n3261_));
  NAND2X1  g03069(.A(new_n3253_), .B(new_n3252_), .Y(new_n3262_));
  INVX1    g03070(.A(new_n3257_), .Y(new_n3263_));
  NOR2X1   g03071(.A(new_n3263_), .B(new_n3246_), .Y(new_n3264_));
  AOI21X1  g03072(.A0(new_n3020_), .A1(new_n3016_), .B0(new_n2981_), .Y(new_n3265_));
  AOI21X1  g03073(.A0(new_n2982_), .A1(new_n2975_), .B0(new_n193_), .Y(new_n3266_));
  OAI21X1  g03074(.A0(new_n3265_), .A1(new_n2975_), .B0(new_n3266_), .Y(new_n3267_));
  INVX1    g03075(.A(new_n2980_), .Y(new_n3268_));
  OR4X1    g03076(.A(new_n3005_), .B(new_n3001_), .C(new_n3268_), .D(new_n2977_), .Y(new_n3269_));
  AOI21X1  g03077(.A0(new_n3018_), .A1(new_n3017_), .B0(new_n3269_), .Y(new_n3270_));
  AND2X1   g03078(.A(new_n3270_), .B(new_n3016_), .Y(new_n3271_));
  INVX1    g03079(.A(new_n3271_), .Y(new_n3272_));
  AND2X1   g03080(.A(new_n3272_), .B(new_n3267_), .Y(new_n3273_));
  INVX1    g03081(.A(new_n3273_), .Y(new_n3274_));
  AOI21X1  g03082(.A0(new_n3264_), .A1(new_n3262_), .B0(new_n3274_), .Y(new_n3275_));
  AND2X1   g03083(.A(new_n3275_), .B(new_n3261_), .Y(new_n3276_));
  NOR2X1   g03084(.A(\a[83] ), .B(\a[82] ), .Y(new_n3277_));
  INVX1    g03085(.A(new_n3277_), .Y(new_n3278_));
  MX2X1    g03086(.A(new_n3278_), .B(new_n3276_), .S0(\a[84] ), .Y(new_n3279_));
  OR2X1    g03087(.A(new_n3243_), .B(new_n292_), .Y(new_n3280_));
  AND2X1   g03088(.A(new_n3227_), .B(new_n3218_), .Y(new_n3281_));
  INVX1    g03089(.A(new_n3232_), .Y(new_n3282_));
  OR2X1    g03090(.A(new_n3233_), .B(\asqrt[60] ), .Y(new_n3283_));
  OAI21X1  g03091(.A0(new_n3283_), .A1(new_n3281_), .B0(new_n3282_), .Y(new_n3284_));
  AOI21X1  g03092(.A0(new_n3284_), .A1(new_n3280_), .B0(new_n217_), .Y(new_n3285_));
  AOI21X1  g03093(.A0(new_n3216_), .A1(\asqrt[60] ), .B0(\asqrt[61] ), .Y(new_n3286_));
  AOI21X1  g03094(.A0(new_n3286_), .A1(new_n3284_), .B0(new_n3241_), .Y(new_n3287_));
  OAI21X1  g03095(.A0(new_n3287_), .A1(new_n3285_), .B0(\asqrt[62] ), .Y(new_n3288_));
  NOR3X1   g03096(.A(new_n3287_), .B(new_n3285_), .C(\asqrt[62] ), .Y(new_n3289_));
  OAI21X1  g03097(.A0(new_n3289_), .A1(new_n3251_), .B0(new_n3288_), .Y(new_n3290_));
  AOI21X1  g03098(.A0(new_n3259_), .A1(new_n3290_), .B0(\asqrt[63] ), .Y(new_n3291_));
  AND2X1   g03099(.A(new_n3253_), .B(new_n3252_), .Y(new_n3292_));
  OR2X1    g03100(.A(new_n3263_), .B(new_n3246_), .Y(new_n3293_));
  OAI21X1  g03101(.A0(new_n3293_), .A1(new_n3292_), .B0(new_n3273_), .Y(new_n3294_));
  OAI21X1  g03102(.A0(new_n3294_), .A1(new_n3291_), .B0(\a[84] ), .Y(new_n3295_));
  OAI22X1  g03103(.A0(new_n3278_), .A1(\a[84] ), .B0(new_n3004_), .B1(new_n3002_), .Y(new_n3296_));
  NOR4X1   g03104(.A(new_n3296_), .B(new_n3001_), .C(new_n3034_), .D(new_n2987_), .Y(new_n3297_));
  AND2X1   g03105(.A(new_n3297_), .B(new_n3295_), .Y(new_n3298_));
  INVX1    g03106(.A(\a[85] ), .Y(new_n3299_));
  AOI21X1  g03107(.A0(new_n3275_), .A1(new_n3261_), .B0(\a[84] ), .Y(new_n3300_));
  OAI21X1  g03108(.A0(new_n3294_), .A1(new_n3291_), .B0(new_n3010_), .Y(new_n3301_));
  OAI21X1  g03109(.A0(new_n3300_), .A1(new_n3299_), .B0(new_n3301_), .Y(new_n3302_));
  OAI22X1  g03110(.A0(new_n3302_), .A1(new_n3298_), .B0(new_n3279_), .B1(new_n3008_), .Y(new_n3303_));
  AND2X1   g03111(.A(new_n3303_), .B(\asqrt[44] ), .Y(new_n3304_));
  OR2X1    g03112(.A(new_n3302_), .B(new_n3298_), .Y(new_n3305_));
  NAND2X1  g03113(.A(new_n3275_), .B(new_n3261_), .Y(\asqrt[42] ));
  MX2X1    g03114(.A(new_n3277_), .B(\asqrt[42] ), .S0(\a[84] ), .Y(new_n3307_));
  AOI21X1  g03115(.A0(new_n3307_), .A1(\asqrt[43] ), .B0(\asqrt[44] ), .Y(new_n3308_));
  INVX1    g03116(.A(new_n3267_), .Y(new_n3309_));
  NOR3X1   g03117(.A(new_n3271_), .B(new_n3309_), .C(new_n3008_), .Y(new_n3310_));
  OAI21X1  g03118(.A0(new_n3293_), .A1(new_n3292_), .B0(new_n3310_), .Y(new_n3311_));
  OR2X1    g03119(.A(new_n3311_), .B(new_n3291_), .Y(new_n3312_));
  AOI21X1  g03120(.A0(new_n3312_), .A1(new_n3301_), .B0(new_n3009_), .Y(new_n3313_));
  AOI21X1  g03121(.A0(new_n3275_), .A1(new_n3261_), .B0(new_n3030_), .Y(new_n3314_));
  OAI21X1  g03122(.A0(new_n3311_), .A1(new_n3291_), .B0(new_n3009_), .Y(new_n3315_));
  NOR2X1   g03123(.A(new_n3315_), .B(new_n3314_), .Y(new_n3316_));
  NOR2X1   g03124(.A(new_n3316_), .B(new_n3313_), .Y(new_n3317_));
  AOI21X1  g03125(.A0(new_n3308_), .A1(new_n3305_), .B0(new_n3317_), .Y(new_n3318_));
  OAI21X1  g03126(.A0(new_n3318_), .A1(new_n3304_), .B0(\asqrt[45] ), .Y(new_n3319_));
  AOI21X1  g03127(.A0(new_n3012_), .A1(\asqrt[44] ), .B0(new_n3049_), .Y(new_n3320_));
  NAND3X1  g03128(.A(new_n3320_), .B(\asqrt[42] ), .C(new_n3052_), .Y(new_n3321_));
  OAI21X1  g03129(.A0(new_n3294_), .A1(new_n3291_), .B0(new_n3320_), .Y(new_n3322_));
  NAND2X1  g03130(.A(new_n3322_), .B(new_n3026_), .Y(new_n3323_));
  NAND2X1  g03131(.A(new_n3323_), .B(new_n3321_), .Y(new_n3324_));
  NAND2X1  g03132(.A(new_n3297_), .B(new_n3295_), .Y(new_n3325_));
  INVX1    g03133(.A(\a[84] ), .Y(new_n3326_));
  OAI21X1  g03134(.A0(new_n3294_), .A1(new_n3291_), .B0(new_n3326_), .Y(new_n3327_));
  AOI21X1  g03135(.A0(new_n3327_), .A1(\a[85] ), .B0(new_n3314_), .Y(new_n3328_));
  AOI22X1  g03136(.A0(new_n3328_), .A1(new_n3325_), .B0(new_n3307_), .B1(\asqrt[43] ), .Y(new_n3329_));
  OAI21X1  g03137(.A0(new_n3329_), .A1(new_n2769_), .B0(new_n2570_), .Y(new_n3330_));
  OAI21X1  g03138(.A0(new_n3330_), .A1(new_n3318_), .B0(new_n3324_), .Y(new_n3331_));
  AOI21X1  g03139(.A0(new_n3331_), .A1(new_n3319_), .B0(new_n2263_), .Y(new_n3332_));
  AOI21X1  g03140(.A0(new_n3075_), .A1(new_n3074_), .B0(new_n3040_), .Y(new_n3333_));
  AND2X1   g03141(.A(new_n3333_), .B(new_n3028_), .Y(new_n3334_));
  AOI22X1  g03142(.A0(new_n3075_), .A1(new_n3074_), .B0(new_n3053_), .B1(\asqrt[45] ), .Y(new_n3335_));
  OAI21X1  g03143(.A0(new_n3294_), .A1(new_n3291_), .B0(new_n3335_), .Y(new_n3336_));
  AOI22X1  g03144(.A0(new_n3336_), .A1(new_n3040_), .B0(new_n3334_), .B1(\asqrt[42] ), .Y(new_n3337_));
  INVX1    g03145(.A(new_n3337_), .Y(new_n3338_));
  NAND3X1  g03146(.A(new_n3331_), .B(new_n3319_), .C(new_n2263_), .Y(new_n3339_));
  AOI21X1  g03147(.A0(new_n3339_), .A1(new_n3338_), .B0(new_n3332_), .Y(new_n3340_));
  OR2X1    g03148(.A(new_n3340_), .B(new_n2040_), .Y(new_n3341_));
  OR2X1    g03149(.A(new_n3329_), .B(new_n2769_), .Y(new_n3342_));
  NOR2X1   g03150(.A(new_n3302_), .B(new_n3298_), .Y(new_n3343_));
  OAI21X1  g03151(.A0(new_n3279_), .A1(new_n3008_), .B0(new_n2769_), .Y(new_n3344_));
  OR2X1    g03152(.A(new_n3316_), .B(new_n3313_), .Y(new_n3345_));
  OAI21X1  g03153(.A0(new_n3344_), .A1(new_n3343_), .B0(new_n3345_), .Y(new_n3346_));
  AOI21X1  g03154(.A0(new_n3346_), .A1(new_n3342_), .B0(new_n2570_), .Y(new_n3347_));
  AOI21X1  g03155(.A0(new_n3303_), .A1(\asqrt[44] ), .B0(\asqrt[45] ), .Y(new_n3348_));
  AOI22X1  g03156(.A0(new_n3348_), .A1(new_n3346_), .B0(new_n3323_), .B1(new_n3321_), .Y(new_n3349_));
  NOR3X1   g03157(.A(new_n3349_), .B(new_n3347_), .C(\asqrt[46] ), .Y(new_n3350_));
  NOR2X1   g03158(.A(new_n3350_), .B(new_n3337_), .Y(new_n3351_));
  AND2X1   g03159(.A(new_n3054_), .B(new_n3041_), .Y(new_n3352_));
  NOR3X1   g03160(.A(new_n3352_), .B(new_n3079_), .C(new_n3042_), .Y(new_n3353_));
  NOR2X1   g03161(.A(new_n3352_), .B(new_n3042_), .Y(new_n3354_));
  OAI21X1  g03162(.A0(new_n3294_), .A1(new_n3291_), .B0(new_n3354_), .Y(new_n3355_));
  AOI22X1  g03163(.A0(new_n3355_), .A1(new_n3079_), .B0(new_n3353_), .B1(\asqrt[42] ), .Y(new_n3356_));
  INVX1    g03164(.A(new_n3356_), .Y(new_n3357_));
  OAI21X1  g03165(.A0(new_n3349_), .A1(new_n3347_), .B0(\asqrt[46] ), .Y(new_n3358_));
  NAND2X1  g03166(.A(new_n3358_), .B(new_n2040_), .Y(new_n3359_));
  OAI21X1  g03167(.A0(new_n3359_), .A1(new_n3351_), .B0(new_n3357_), .Y(new_n3360_));
  AOI21X1  g03168(.A0(new_n3360_), .A1(new_n3341_), .B0(new_n1834_), .Y(new_n3361_));
  NAND4X1  g03169(.A(\asqrt[42] ), .B(new_n3094_), .C(new_n3063_), .D(new_n3056_), .Y(new_n3362_));
  NOR3X1   g03170(.A(new_n3276_), .B(new_n3064_), .C(new_n3082_), .Y(new_n3363_));
  OAI21X1  g03171(.A0(new_n3363_), .A1(new_n3063_), .B0(new_n3362_), .Y(new_n3364_));
  INVX1    g03172(.A(new_n3364_), .Y(new_n3365_));
  OAI21X1  g03173(.A0(new_n3350_), .A1(new_n3337_), .B0(new_n3358_), .Y(new_n3366_));
  AOI21X1  g03174(.A0(new_n3366_), .A1(\asqrt[47] ), .B0(\asqrt[48] ), .Y(new_n3367_));
  AOI21X1  g03175(.A0(new_n3367_), .A1(new_n3360_), .B0(new_n3365_), .Y(new_n3368_));
  OAI21X1  g03176(.A0(new_n3368_), .A1(new_n3361_), .B0(\asqrt[49] ), .Y(new_n3369_));
  AND2X1   g03177(.A(new_n3083_), .B(new_n3067_), .Y(new_n3370_));
  NOR3X1   g03178(.A(new_n3370_), .B(new_n3110_), .C(new_n3066_), .Y(new_n3371_));
  AOI22X1  g03179(.A0(new_n3083_), .A1(new_n3067_), .B0(new_n3065_), .B1(\asqrt[48] ), .Y(new_n3372_));
  AOI21X1  g03180(.A0(new_n3372_), .A1(\asqrt[42] ), .B0(new_n3072_), .Y(new_n3373_));
  AOI21X1  g03181(.A0(new_n3371_), .A1(\asqrt[42] ), .B0(new_n3373_), .Y(new_n3374_));
  NOR3X1   g03182(.A(new_n3368_), .B(new_n3361_), .C(\asqrt[49] ), .Y(new_n3375_));
  OAI21X1  g03183(.A0(new_n3375_), .A1(new_n3374_), .B0(new_n3369_), .Y(new_n3376_));
  AND2X1   g03184(.A(new_n3376_), .B(\asqrt[50] ), .Y(new_n3377_));
  INVX1    g03185(.A(new_n3374_), .Y(new_n3378_));
  AND2X1   g03186(.A(new_n3366_), .B(\asqrt[47] ), .Y(new_n3379_));
  OR2X1    g03187(.A(new_n3350_), .B(new_n3337_), .Y(new_n3380_));
  AND2X1   g03188(.A(new_n3358_), .B(new_n2040_), .Y(new_n3381_));
  AOI21X1  g03189(.A0(new_n3381_), .A1(new_n3380_), .B0(new_n3356_), .Y(new_n3382_));
  OAI21X1  g03190(.A0(new_n3382_), .A1(new_n3379_), .B0(\asqrt[48] ), .Y(new_n3383_));
  OAI21X1  g03191(.A0(new_n3340_), .A1(new_n2040_), .B0(new_n1834_), .Y(new_n3384_));
  OAI21X1  g03192(.A0(new_n3384_), .A1(new_n3382_), .B0(new_n3364_), .Y(new_n3385_));
  NAND3X1  g03193(.A(new_n3385_), .B(new_n3383_), .C(new_n1632_), .Y(new_n3386_));
  NAND2X1  g03194(.A(new_n3386_), .B(new_n3378_), .Y(new_n3387_));
  AND2X1   g03195(.A(new_n3114_), .B(new_n3112_), .Y(new_n3388_));
  NOR3X1   g03196(.A(new_n3388_), .B(new_n3092_), .C(new_n3113_), .Y(new_n3389_));
  NOR2X1   g03197(.A(new_n3388_), .B(new_n3113_), .Y(new_n3390_));
  AOI21X1  g03198(.A0(new_n3390_), .A1(\asqrt[42] ), .B0(new_n3091_), .Y(new_n3391_));
  AOI21X1  g03199(.A0(new_n3389_), .A1(\asqrt[42] ), .B0(new_n3391_), .Y(new_n3392_));
  AND2X1   g03200(.A(new_n3369_), .B(new_n1469_), .Y(new_n3393_));
  AOI21X1  g03201(.A0(new_n3393_), .A1(new_n3387_), .B0(new_n3392_), .Y(new_n3394_));
  OAI21X1  g03202(.A0(new_n3394_), .A1(new_n3377_), .B0(\asqrt[51] ), .Y(new_n3395_));
  OR4X1    g03203(.A(new_n3276_), .B(new_n3116_), .C(new_n3104_), .D(new_n3098_), .Y(new_n3396_));
  OR2X1    g03204(.A(new_n3116_), .B(new_n3098_), .Y(new_n3397_));
  OAI21X1  g03205(.A0(new_n3397_), .A1(new_n3276_), .B0(new_n3104_), .Y(new_n3398_));
  AND2X1   g03206(.A(new_n3398_), .B(new_n3396_), .Y(new_n3399_));
  INVX1    g03207(.A(new_n3399_), .Y(new_n3400_));
  AOI21X1  g03208(.A0(new_n3385_), .A1(new_n3383_), .B0(new_n1632_), .Y(new_n3401_));
  AOI21X1  g03209(.A0(new_n3386_), .A1(new_n3378_), .B0(new_n3401_), .Y(new_n3402_));
  OAI21X1  g03210(.A0(new_n3402_), .A1(new_n1469_), .B0(new_n1277_), .Y(new_n3403_));
  OAI21X1  g03211(.A0(new_n3403_), .A1(new_n3394_), .B0(new_n3400_), .Y(new_n3404_));
  AOI21X1  g03212(.A0(new_n3404_), .A1(new_n3395_), .B0(new_n1111_), .Y(new_n3405_));
  AOI21X1  g03213(.A0(new_n3147_), .A1(new_n3146_), .B0(new_n3122_), .Y(new_n3406_));
  AND2X1   g03214(.A(new_n3406_), .B(new_n3107_), .Y(new_n3407_));
  AOI22X1  g03215(.A0(new_n3147_), .A1(new_n3146_), .B0(new_n3132_), .B1(\asqrt[51] ), .Y(new_n3408_));
  AOI21X1  g03216(.A0(new_n3408_), .A1(\asqrt[42] ), .B0(new_n3121_), .Y(new_n3409_));
  AOI21X1  g03217(.A0(new_n3407_), .A1(\asqrt[42] ), .B0(new_n3409_), .Y(new_n3410_));
  INVX1    g03218(.A(new_n3410_), .Y(new_n3411_));
  NAND3X1  g03219(.A(new_n3404_), .B(new_n3395_), .C(new_n1111_), .Y(new_n3412_));
  AOI21X1  g03220(.A0(new_n3412_), .A1(new_n3411_), .B0(new_n3405_), .Y(new_n3413_));
  OR2X1    g03221(.A(new_n3413_), .B(new_n968_), .Y(new_n3414_));
  AND2X1   g03222(.A(new_n3412_), .B(new_n3411_), .Y(new_n3415_));
  AND2X1   g03223(.A(new_n3133_), .B(new_n3125_), .Y(new_n3416_));
  NOR3X1   g03224(.A(new_n3416_), .B(new_n3150_), .C(new_n3126_), .Y(new_n3417_));
  NOR2X1   g03225(.A(new_n3416_), .B(new_n3126_), .Y(new_n3418_));
  AOI21X1  g03226(.A0(new_n3418_), .A1(\asqrt[42] ), .B0(new_n3131_), .Y(new_n3419_));
  AOI21X1  g03227(.A0(new_n3417_), .A1(\asqrt[42] ), .B0(new_n3419_), .Y(new_n3420_));
  INVX1    g03228(.A(new_n3420_), .Y(new_n3421_));
  OR2X1    g03229(.A(new_n3402_), .B(new_n1469_), .Y(new_n3422_));
  AND2X1   g03230(.A(new_n3386_), .B(new_n3378_), .Y(new_n3423_));
  INVX1    g03231(.A(new_n3392_), .Y(new_n3424_));
  NAND2X1  g03232(.A(new_n3369_), .B(new_n1469_), .Y(new_n3425_));
  OAI21X1  g03233(.A0(new_n3425_), .A1(new_n3423_), .B0(new_n3424_), .Y(new_n3426_));
  AOI21X1  g03234(.A0(new_n3426_), .A1(new_n3422_), .B0(new_n1277_), .Y(new_n3427_));
  AOI21X1  g03235(.A0(new_n3376_), .A1(\asqrt[50] ), .B0(\asqrt[51] ), .Y(new_n3428_));
  AOI21X1  g03236(.A0(new_n3428_), .A1(new_n3426_), .B0(new_n3399_), .Y(new_n3429_));
  OAI21X1  g03237(.A0(new_n3429_), .A1(new_n3427_), .B0(\asqrt[52] ), .Y(new_n3430_));
  NAND2X1  g03238(.A(new_n3430_), .B(new_n968_), .Y(new_n3431_));
  OAI21X1  g03239(.A0(new_n3431_), .A1(new_n3415_), .B0(new_n3421_), .Y(new_n3432_));
  AOI21X1  g03240(.A0(new_n3432_), .A1(new_n3414_), .B0(new_n902_), .Y(new_n3433_));
  OR4X1    g03241(.A(new_n3276_), .B(new_n3141_), .C(new_n3144_), .D(new_n3155_), .Y(new_n3434_));
  NAND2X1  g03242(.A(new_n3153_), .B(new_n3135_), .Y(new_n3435_));
  OAI21X1  g03243(.A0(new_n3435_), .A1(new_n3276_), .B0(new_n3144_), .Y(new_n3436_));
  AND2X1   g03244(.A(new_n3436_), .B(new_n3434_), .Y(new_n3437_));
  NOR3X1   g03245(.A(new_n3429_), .B(new_n3427_), .C(\asqrt[52] ), .Y(new_n3438_));
  OAI21X1  g03246(.A0(new_n3438_), .A1(new_n3410_), .B0(new_n3430_), .Y(new_n3439_));
  AOI21X1  g03247(.A0(new_n3439_), .A1(\asqrt[53] ), .B0(\asqrt[54] ), .Y(new_n3440_));
  AOI21X1  g03248(.A0(new_n3440_), .A1(new_n3432_), .B0(new_n3437_), .Y(new_n3441_));
  OAI21X1  g03249(.A0(new_n3441_), .A1(new_n3433_), .B0(\asqrt[55] ), .Y(new_n3442_));
  NOR3X1   g03250(.A(new_n3441_), .B(new_n3433_), .C(\asqrt[55] ), .Y(new_n3443_));
  AND2X1   g03251(.A(new_n3156_), .B(new_n3154_), .Y(new_n3444_));
  NOR3X1   g03252(.A(new_n3199_), .B(new_n3444_), .C(new_n3143_), .Y(new_n3445_));
  AOI22X1  g03253(.A0(new_n3156_), .A1(new_n3154_), .B0(new_n3142_), .B1(\asqrt[54] ), .Y(new_n3446_));
  AOI21X1  g03254(.A0(new_n3446_), .A1(\asqrt[42] ), .B0(new_n3160_), .Y(new_n3447_));
  AOI21X1  g03255(.A0(new_n3445_), .A1(\asqrt[42] ), .B0(new_n3447_), .Y(new_n3448_));
  OAI21X1  g03256(.A0(new_n3448_), .A1(new_n3443_), .B0(new_n3442_), .Y(new_n3449_));
  AND2X1   g03257(.A(new_n3449_), .B(\asqrt[56] ), .Y(new_n3450_));
  OR2X1    g03258(.A(new_n3448_), .B(new_n3443_), .Y(new_n3451_));
  AND2X1   g03259(.A(new_n3202_), .B(new_n3200_), .Y(new_n3452_));
  NOR3X1   g03260(.A(new_n3452_), .B(new_n3168_), .C(new_n3201_), .Y(new_n3453_));
  NOR2X1   g03261(.A(new_n3452_), .B(new_n3201_), .Y(new_n3454_));
  AOI21X1  g03262(.A0(new_n3454_), .A1(\asqrt[42] ), .B0(new_n3167_), .Y(new_n3455_));
  AOI21X1  g03263(.A0(new_n3453_), .A1(\asqrt[42] ), .B0(new_n3455_), .Y(new_n3456_));
  AND2X1   g03264(.A(new_n3442_), .B(new_n582_), .Y(new_n3457_));
  AOI21X1  g03265(.A0(new_n3457_), .A1(new_n3451_), .B0(new_n3456_), .Y(new_n3458_));
  OAI21X1  g03266(.A0(new_n3458_), .A1(new_n3450_), .B0(\asqrt[57] ), .Y(new_n3459_));
  NAND4X1  g03267(.A(\asqrt[42] ), .B(new_n3179_), .C(new_n3177_), .D(new_n3204_), .Y(new_n3460_));
  NAND2X1  g03268(.A(new_n3179_), .B(new_n3204_), .Y(new_n3461_));
  OAI21X1  g03269(.A0(new_n3461_), .A1(new_n3276_), .B0(new_n3178_), .Y(new_n3462_));
  AND2X1   g03270(.A(new_n3462_), .B(new_n3460_), .Y(new_n3463_));
  INVX1    g03271(.A(new_n3463_), .Y(new_n3464_));
  AND2X1   g03272(.A(new_n3439_), .B(\asqrt[53] ), .Y(new_n3465_));
  NAND2X1  g03273(.A(new_n3412_), .B(new_n3411_), .Y(new_n3466_));
  AND2X1   g03274(.A(new_n3430_), .B(new_n968_), .Y(new_n3467_));
  AOI21X1  g03275(.A0(new_n3467_), .A1(new_n3466_), .B0(new_n3420_), .Y(new_n3468_));
  OAI21X1  g03276(.A0(new_n3468_), .A1(new_n3465_), .B0(\asqrt[54] ), .Y(new_n3469_));
  INVX1    g03277(.A(new_n3437_), .Y(new_n3470_));
  OAI21X1  g03278(.A0(new_n3413_), .A1(new_n968_), .B0(new_n902_), .Y(new_n3471_));
  OAI21X1  g03279(.A0(new_n3471_), .A1(new_n3468_), .B0(new_n3470_), .Y(new_n3472_));
  AOI21X1  g03280(.A0(new_n3472_), .A1(new_n3469_), .B0(new_n697_), .Y(new_n3473_));
  NAND3X1  g03281(.A(new_n3472_), .B(new_n3469_), .C(new_n697_), .Y(new_n3474_));
  INVX1    g03282(.A(new_n3448_), .Y(new_n3475_));
  AOI21X1  g03283(.A0(new_n3475_), .A1(new_n3474_), .B0(new_n3473_), .Y(new_n3476_));
  OAI21X1  g03284(.A0(new_n3476_), .A1(new_n582_), .B0(new_n481_), .Y(new_n3477_));
  OAI21X1  g03285(.A0(new_n3477_), .A1(new_n3458_), .B0(new_n3464_), .Y(new_n3478_));
  AOI21X1  g03286(.A0(new_n3478_), .A1(new_n3459_), .B0(new_n399_), .Y(new_n3479_));
  AOI21X1  g03287(.A0(new_n3221_), .A1(new_n3220_), .B0(new_n3187_), .Y(new_n3480_));
  AND2X1   g03288(.A(new_n3480_), .B(new_n3181_), .Y(new_n3481_));
  AOI22X1  g03289(.A0(new_n3221_), .A1(new_n3220_), .B0(new_n3206_), .B1(\asqrt[57] ), .Y(new_n3482_));
  AOI21X1  g03290(.A0(new_n3482_), .A1(\asqrt[42] ), .B0(new_n3186_), .Y(new_n3483_));
  AOI21X1  g03291(.A0(new_n3481_), .A1(\asqrt[42] ), .B0(new_n3483_), .Y(new_n3484_));
  INVX1    g03292(.A(new_n3484_), .Y(new_n3485_));
  NAND3X1  g03293(.A(new_n3478_), .B(new_n3459_), .C(new_n399_), .Y(new_n3486_));
  AOI21X1  g03294(.A0(new_n3486_), .A1(new_n3485_), .B0(new_n3479_), .Y(new_n3487_));
  OR2X1    g03295(.A(new_n3487_), .B(new_n328_), .Y(new_n3488_));
  AND2X1   g03296(.A(new_n3486_), .B(new_n3485_), .Y(new_n3489_));
  AND2X1   g03297(.A(new_n3207_), .B(new_n3189_), .Y(new_n3490_));
  NOR3X1   g03298(.A(new_n3490_), .B(new_n3224_), .C(new_n3190_), .Y(new_n3491_));
  NOR2X1   g03299(.A(new_n3490_), .B(new_n3190_), .Y(new_n3492_));
  AOI21X1  g03300(.A0(new_n3492_), .A1(\asqrt[42] ), .B0(new_n3195_), .Y(new_n3493_));
  AOI21X1  g03301(.A0(new_n3491_), .A1(\asqrt[42] ), .B0(new_n3493_), .Y(new_n3494_));
  INVX1    g03302(.A(new_n3494_), .Y(new_n3495_));
  OR2X1    g03303(.A(new_n3476_), .B(new_n582_), .Y(new_n3496_));
  NOR2X1   g03304(.A(new_n3448_), .B(new_n3443_), .Y(new_n3497_));
  INVX1    g03305(.A(new_n3456_), .Y(new_n3498_));
  NAND2X1  g03306(.A(new_n3442_), .B(new_n582_), .Y(new_n3499_));
  OAI21X1  g03307(.A0(new_n3499_), .A1(new_n3497_), .B0(new_n3498_), .Y(new_n3500_));
  AOI21X1  g03308(.A0(new_n3500_), .A1(new_n3496_), .B0(new_n481_), .Y(new_n3501_));
  AOI21X1  g03309(.A0(new_n3449_), .A1(\asqrt[56] ), .B0(\asqrt[57] ), .Y(new_n3502_));
  AOI21X1  g03310(.A0(new_n3502_), .A1(new_n3500_), .B0(new_n3463_), .Y(new_n3503_));
  OAI21X1  g03311(.A0(new_n3503_), .A1(new_n3501_), .B0(\asqrt[58] ), .Y(new_n3504_));
  NAND2X1  g03312(.A(new_n3504_), .B(new_n328_), .Y(new_n3505_));
  OAI21X1  g03313(.A0(new_n3505_), .A1(new_n3489_), .B0(new_n3495_), .Y(new_n3506_));
  AOI21X1  g03314(.A0(new_n3506_), .A1(new_n3488_), .B0(new_n292_), .Y(new_n3507_));
  NAND4X1  g03315(.A(\asqrt[42] ), .B(new_n3227_), .C(new_n3214_), .D(new_n3209_), .Y(new_n3508_));
  NAND2X1  g03316(.A(new_n3227_), .B(new_n3209_), .Y(new_n3509_));
  OAI21X1  g03317(.A0(new_n3509_), .A1(new_n3276_), .B0(new_n3218_), .Y(new_n3510_));
  AND2X1   g03318(.A(new_n3510_), .B(new_n3508_), .Y(new_n3511_));
  NOR3X1   g03319(.A(new_n3503_), .B(new_n3501_), .C(\asqrt[58] ), .Y(new_n3512_));
  OAI21X1  g03320(.A0(new_n3512_), .A1(new_n3484_), .B0(new_n3504_), .Y(new_n3513_));
  AOI21X1  g03321(.A0(new_n3513_), .A1(\asqrt[59] ), .B0(\asqrt[60] ), .Y(new_n3514_));
  AOI21X1  g03322(.A0(new_n3514_), .A1(new_n3506_), .B0(new_n3511_), .Y(new_n3515_));
  OAI21X1  g03323(.A0(new_n3515_), .A1(new_n3507_), .B0(\asqrt[61] ), .Y(new_n3516_));
  AND2X1   g03324(.A(new_n3234_), .B(new_n3228_), .Y(new_n3517_));
  NOR3X1   g03325(.A(new_n3517_), .B(new_n3282_), .C(new_n3217_), .Y(new_n3518_));
  AOI22X1  g03326(.A0(new_n3234_), .A1(new_n3228_), .B0(new_n3216_), .B1(\asqrt[60] ), .Y(new_n3519_));
  AOI21X1  g03327(.A0(new_n3519_), .A1(\asqrt[42] ), .B0(new_n3232_), .Y(new_n3520_));
  AOI21X1  g03328(.A0(new_n3518_), .A1(\asqrt[42] ), .B0(new_n3520_), .Y(new_n3521_));
  NOR3X1   g03329(.A(new_n3515_), .B(new_n3507_), .C(\asqrt[61] ), .Y(new_n3522_));
  OAI21X1  g03330(.A0(new_n3522_), .A1(new_n3521_), .B0(new_n3516_), .Y(new_n3523_));
  AND2X1   g03331(.A(new_n3523_), .B(\asqrt[62] ), .Y(new_n3524_));
  INVX1    g03332(.A(new_n3521_), .Y(new_n3525_));
  AND2X1   g03333(.A(new_n3513_), .B(\asqrt[59] ), .Y(new_n3526_));
  NAND2X1  g03334(.A(new_n3486_), .B(new_n3485_), .Y(new_n3527_));
  AND2X1   g03335(.A(new_n3504_), .B(new_n328_), .Y(new_n3528_));
  AOI21X1  g03336(.A0(new_n3528_), .A1(new_n3527_), .B0(new_n3494_), .Y(new_n3529_));
  OAI21X1  g03337(.A0(new_n3529_), .A1(new_n3526_), .B0(\asqrt[60] ), .Y(new_n3530_));
  INVX1    g03338(.A(new_n3511_), .Y(new_n3531_));
  OAI21X1  g03339(.A0(new_n3487_), .A1(new_n328_), .B0(new_n292_), .Y(new_n3532_));
  OAI21X1  g03340(.A0(new_n3532_), .A1(new_n3529_), .B0(new_n3531_), .Y(new_n3533_));
  NAND3X1  g03341(.A(new_n3533_), .B(new_n3530_), .C(new_n217_), .Y(new_n3534_));
  NAND2X1  g03342(.A(new_n3534_), .B(new_n3525_), .Y(new_n3535_));
  AND2X1   g03343(.A(new_n3286_), .B(new_n3284_), .Y(new_n3536_));
  NOR3X1   g03344(.A(new_n3536_), .B(new_n3242_), .C(new_n3285_), .Y(new_n3537_));
  NOR2X1   g03345(.A(new_n3536_), .B(new_n3285_), .Y(new_n3538_));
  AOI21X1  g03346(.A0(new_n3538_), .A1(\asqrt[42] ), .B0(new_n3241_), .Y(new_n3539_));
  AOI21X1  g03347(.A0(new_n3537_), .A1(\asqrt[42] ), .B0(new_n3539_), .Y(new_n3540_));
  AOI21X1  g03348(.A0(new_n3533_), .A1(new_n3530_), .B0(new_n217_), .Y(new_n3541_));
  NOR2X1   g03349(.A(new_n3541_), .B(\asqrt[62] ), .Y(new_n3542_));
  AOI21X1  g03350(.A0(new_n3542_), .A1(new_n3535_), .B0(new_n3540_), .Y(new_n3543_));
  OR4X1    g03351(.A(new_n3276_), .B(new_n3289_), .C(new_n3252_), .D(new_n3246_), .Y(new_n3544_));
  NAND2X1  g03352(.A(new_n3253_), .B(new_n3288_), .Y(new_n3545_));
  OAI21X1  g03353(.A0(new_n3545_), .A1(new_n3276_), .B0(new_n3252_), .Y(new_n3546_));
  AND2X1   g03354(.A(new_n3546_), .B(new_n3544_), .Y(new_n3547_));
  INVX1    g03355(.A(new_n3547_), .Y(new_n3548_));
  NOR2X1   g03356(.A(new_n3257_), .B(new_n3254_), .Y(new_n3549_));
  AOI22X1  g03357(.A0(new_n3549_), .A1(\asqrt[42] ), .B0(new_n3264_), .B1(new_n3262_), .Y(new_n3550_));
  AND2X1   g03358(.A(new_n3550_), .B(new_n3548_), .Y(new_n3551_));
  OAI21X1  g03359(.A0(new_n3543_), .A1(new_n3524_), .B0(new_n3551_), .Y(new_n3552_));
  AOI21X1  g03360(.A0(new_n3534_), .A1(new_n3525_), .B0(new_n3541_), .Y(new_n3553_));
  OAI21X1  g03361(.A0(new_n3553_), .A1(new_n199_), .B0(new_n3547_), .Y(new_n3554_));
  AOI21X1  g03362(.A0(new_n3275_), .A1(new_n3261_), .B0(new_n3257_), .Y(new_n3555_));
  AOI21X1  g03363(.A0(new_n3263_), .A1(new_n3290_), .B0(new_n193_), .Y(new_n3556_));
  OAI21X1  g03364(.A0(new_n3555_), .A1(new_n3290_), .B0(new_n3556_), .Y(new_n3557_));
  OR2X1    g03365(.A(new_n3293_), .B(new_n3292_), .Y(new_n3558_));
  AND2X1   g03366(.A(new_n3256_), .B(new_n2972_), .Y(new_n3559_));
  NOR4X1   g03367(.A(new_n3271_), .B(new_n3309_), .C(new_n3559_), .D(new_n3255_), .Y(new_n3560_));
  NAND3X1  g03368(.A(new_n3560_), .B(new_n3558_), .C(new_n3261_), .Y(new_n3561_));
  AND2X1   g03369(.A(new_n3561_), .B(new_n3557_), .Y(new_n3562_));
  OAI21X1  g03370(.A0(new_n3554_), .A1(new_n3543_), .B0(new_n3562_), .Y(new_n3563_));
  AOI21X1  g03371(.A0(new_n3552_), .A1(new_n193_), .B0(new_n3563_), .Y(new_n3564_));
  NOR2X1   g03372(.A(\a[81] ), .B(\a[80] ), .Y(new_n3565_));
  INVX1    g03373(.A(new_n3565_), .Y(new_n3566_));
  MX2X1    g03374(.A(new_n3566_), .B(new_n3564_), .S0(\a[82] ), .Y(new_n3567_));
  OR2X1    g03375(.A(new_n3567_), .B(new_n3276_), .Y(new_n3568_));
  INVX1    g03376(.A(\a[82] ), .Y(new_n3569_));
  NOR3X1   g03377(.A(\a[82] ), .B(\a[81] ), .C(\a[80] ), .Y(new_n3570_));
  NOR3X1   g03378(.A(new_n3570_), .B(new_n3271_), .C(new_n3309_), .Y(new_n3571_));
  NAND3X1  g03379(.A(new_n3571_), .B(new_n3558_), .C(new_n3261_), .Y(new_n3572_));
  INVX1    g03380(.A(new_n3572_), .Y(new_n3573_));
  OAI21X1  g03381(.A0(new_n3564_), .A1(new_n3569_), .B0(new_n3573_), .Y(new_n3574_));
  OAI21X1  g03382(.A0(new_n3564_), .A1(\a[82] ), .B0(\a[83] ), .Y(new_n3575_));
  OR2X1    g03383(.A(new_n3564_), .B(new_n3278_), .Y(new_n3576_));
  NAND3X1  g03384(.A(new_n3576_), .B(new_n3575_), .C(new_n3574_), .Y(new_n3577_));
  AOI21X1  g03385(.A0(new_n3577_), .A1(new_n3568_), .B0(new_n3008_), .Y(new_n3578_));
  OR2X1    g03386(.A(new_n3553_), .B(new_n199_), .Y(new_n3579_));
  AND2X1   g03387(.A(new_n3534_), .B(new_n3525_), .Y(new_n3580_));
  INVX1    g03388(.A(new_n3540_), .Y(new_n3581_));
  OR2X1    g03389(.A(new_n3541_), .B(\asqrt[62] ), .Y(new_n3582_));
  OAI21X1  g03390(.A0(new_n3582_), .A1(new_n3580_), .B0(new_n3581_), .Y(new_n3583_));
  INVX1    g03391(.A(new_n3551_), .Y(new_n3584_));
  AOI21X1  g03392(.A0(new_n3583_), .A1(new_n3579_), .B0(new_n3584_), .Y(new_n3585_));
  AOI21X1  g03393(.A0(new_n3523_), .A1(\asqrt[62] ), .B0(new_n3548_), .Y(new_n3586_));
  INVX1    g03394(.A(new_n3562_), .Y(new_n3587_));
  AOI21X1  g03395(.A0(new_n3586_), .A1(new_n3583_), .B0(new_n3587_), .Y(new_n3588_));
  OAI21X1  g03396(.A0(new_n3585_), .A1(\asqrt[63] ), .B0(new_n3588_), .Y(\asqrt[41] ));
  MX2X1    g03397(.A(new_n3565_), .B(\asqrt[41] ), .S0(\a[82] ), .Y(new_n3590_));
  AOI21X1  g03398(.A0(new_n3590_), .A1(\asqrt[42] ), .B0(\asqrt[43] ), .Y(new_n3591_));
  NAND3X1  g03399(.A(new_n3561_), .B(new_n3557_), .C(\asqrt[42] ), .Y(new_n3592_));
  INVX1    g03400(.A(new_n3592_), .Y(new_n3593_));
  OAI21X1  g03401(.A0(new_n3554_), .A1(new_n3543_), .B0(new_n3593_), .Y(new_n3594_));
  AOI21X1  g03402(.A0(new_n3552_), .A1(new_n193_), .B0(new_n3594_), .Y(new_n3595_));
  AOI21X1  g03403(.A0(\asqrt[41] ), .A1(new_n3277_), .B0(new_n3595_), .Y(new_n3596_));
  OR2X1    g03404(.A(new_n3596_), .B(new_n3326_), .Y(new_n3597_));
  AND2X1   g03405(.A(\asqrt[41] ), .B(new_n3277_), .Y(new_n3598_));
  OR2X1    g03406(.A(new_n3595_), .B(\a[84] ), .Y(new_n3599_));
  OR2X1    g03407(.A(new_n3599_), .B(new_n3598_), .Y(new_n3600_));
  AOI22X1  g03408(.A0(new_n3600_), .A1(new_n3597_), .B0(new_n3591_), .B1(new_n3577_), .Y(new_n3601_));
  OAI21X1  g03409(.A0(new_n3601_), .A1(new_n3578_), .B0(\asqrt[44] ), .Y(new_n3602_));
  AOI21X1  g03410(.A0(new_n3307_), .A1(\asqrt[43] ), .B0(new_n3298_), .Y(new_n3603_));
  NAND3X1  g03411(.A(new_n3603_), .B(\asqrt[41] ), .C(new_n3302_), .Y(new_n3604_));
  INVX1    g03412(.A(new_n3603_), .Y(new_n3605_));
  OAI21X1  g03413(.A0(new_n3605_), .A1(new_n3564_), .B0(new_n3328_), .Y(new_n3606_));
  AND2X1   g03414(.A(new_n3606_), .B(new_n3604_), .Y(new_n3607_));
  NOR3X1   g03415(.A(new_n3601_), .B(new_n3578_), .C(\asqrt[44] ), .Y(new_n3608_));
  OAI21X1  g03416(.A0(new_n3608_), .A1(new_n3607_), .B0(new_n3602_), .Y(new_n3609_));
  AND2X1   g03417(.A(new_n3609_), .B(\asqrt[45] ), .Y(new_n3610_));
  INVX1    g03418(.A(new_n3607_), .Y(new_n3611_));
  AND2X1   g03419(.A(new_n3590_), .B(\asqrt[42] ), .Y(new_n3612_));
  AOI21X1  g03420(.A0(\asqrt[41] ), .A1(\a[82] ), .B0(new_n3572_), .Y(new_n3613_));
  INVX1    g03421(.A(\a[83] ), .Y(new_n3614_));
  AOI21X1  g03422(.A0(\asqrt[41] ), .A1(new_n3569_), .B0(new_n3614_), .Y(new_n3615_));
  NOR3X1   g03423(.A(new_n3598_), .B(new_n3615_), .C(new_n3613_), .Y(new_n3616_));
  OAI21X1  g03424(.A0(new_n3616_), .A1(new_n3612_), .B0(\asqrt[43] ), .Y(new_n3617_));
  OAI21X1  g03425(.A0(new_n3567_), .A1(new_n3276_), .B0(new_n3008_), .Y(new_n3618_));
  OAI22X1  g03426(.A0(new_n3599_), .A1(new_n3598_), .B0(new_n3596_), .B1(new_n3326_), .Y(new_n3619_));
  OAI21X1  g03427(.A0(new_n3618_), .A1(new_n3616_), .B0(new_n3619_), .Y(new_n3620_));
  NAND3X1  g03428(.A(new_n3620_), .B(new_n3617_), .C(new_n2769_), .Y(new_n3621_));
  NAND2X1  g03429(.A(new_n3621_), .B(new_n3611_), .Y(new_n3622_));
  OAI21X1  g03430(.A0(new_n3344_), .A1(new_n3343_), .B0(new_n3317_), .Y(new_n3623_));
  NOR3X1   g03431(.A(new_n3623_), .B(new_n3564_), .C(new_n3304_), .Y(new_n3624_));
  OAI22X1  g03432(.A0(new_n3344_), .A1(new_n3343_), .B0(new_n3329_), .B1(new_n2769_), .Y(new_n3625_));
  OR2X1    g03433(.A(new_n3625_), .B(new_n3564_), .Y(new_n3626_));
  AOI21X1  g03434(.A0(new_n3626_), .A1(new_n3345_), .B0(new_n3624_), .Y(new_n3627_));
  AOI21X1  g03435(.A0(new_n3620_), .A1(new_n3617_), .B0(new_n2769_), .Y(new_n3628_));
  NOR2X1   g03436(.A(new_n3628_), .B(\asqrt[45] ), .Y(new_n3629_));
  AOI21X1  g03437(.A0(new_n3629_), .A1(new_n3622_), .B0(new_n3627_), .Y(new_n3630_));
  OAI21X1  g03438(.A0(new_n3630_), .A1(new_n3610_), .B0(\asqrt[46] ), .Y(new_n3631_));
  AND2X1   g03439(.A(new_n3348_), .B(new_n3346_), .Y(new_n3632_));
  OR4X1    g03440(.A(new_n3564_), .B(new_n3632_), .C(new_n3324_), .D(new_n3347_), .Y(new_n3633_));
  OR2X1    g03441(.A(new_n3632_), .B(new_n3347_), .Y(new_n3634_));
  OAI21X1  g03442(.A0(new_n3634_), .A1(new_n3564_), .B0(new_n3324_), .Y(new_n3635_));
  AND2X1   g03443(.A(new_n3635_), .B(new_n3633_), .Y(new_n3636_));
  INVX1    g03444(.A(new_n3636_), .Y(new_n3637_));
  AOI21X1  g03445(.A0(new_n3621_), .A1(new_n3611_), .B0(new_n3628_), .Y(new_n3638_));
  OAI21X1  g03446(.A0(new_n3638_), .A1(new_n2570_), .B0(new_n2263_), .Y(new_n3639_));
  OAI21X1  g03447(.A0(new_n3639_), .A1(new_n3630_), .B0(new_n3637_), .Y(new_n3640_));
  AOI21X1  g03448(.A0(new_n3640_), .A1(new_n3631_), .B0(new_n2040_), .Y(new_n3641_));
  NAND3X1  g03449(.A(new_n3339_), .B(new_n3337_), .C(new_n3358_), .Y(new_n3642_));
  NOR3X1   g03450(.A(new_n3564_), .B(new_n3350_), .C(new_n3332_), .Y(new_n3643_));
  OAI22X1  g03451(.A0(new_n3643_), .A1(new_n3337_), .B0(new_n3642_), .B1(new_n3564_), .Y(new_n3644_));
  NAND3X1  g03452(.A(new_n3640_), .B(new_n3631_), .C(new_n2040_), .Y(new_n3645_));
  AOI21X1  g03453(.A0(new_n3645_), .A1(new_n3644_), .B0(new_n3641_), .Y(new_n3646_));
  OR2X1    g03454(.A(new_n3646_), .B(new_n1834_), .Y(new_n3647_));
  AND2X1   g03455(.A(new_n3645_), .B(new_n3644_), .Y(new_n3648_));
  AND2X1   g03456(.A(new_n3381_), .B(new_n3380_), .Y(new_n3649_));
  NOR4X1   g03457(.A(new_n3564_), .B(new_n3649_), .C(new_n3357_), .D(new_n3379_), .Y(new_n3650_));
  AOI22X1  g03458(.A0(new_n3381_), .A1(new_n3380_), .B0(new_n3366_), .B1(\asqrt[47] ), .Y(new_n3651_));
  AOI21X1  g03459(.A0(new_n3651_), .A1(\asqrt[41] ), .B0(new_n3356_), .Y(new_n3652_));
  NOR2X1   g03460(.A(new_n3652_), .B(new_n3650_), .Y(new_n3653_));
  INVX1    g03461(.A(new_n3653_), .Y(new_n3654_));
  OR2X1    g03462(.A(new_n3641_), .B(\asqrt[48] ), .Y(new_n3655_));
  OAI21X1  g03463(.A0(new_n3655_), .A1(new_n3648_), .B0(new_n3654_), .Y(new_n3656_));
  AOI21X1  g03464(.A0(new_n3656_), .A1(new_n3647_), .B0(new_n1632_), .Y(new_n3657_));
  AND2X1   g03465(.A(new_n3367_), .B(new_n3360_), .Y(new_n3658_));
  OR4X1    g03466(.A(new_n3564_), .B(new_n3658_), .C(new_n3364_), .D(new_n3361_), .Y(new_n3659_));
  OR2X1    g03467(.A(new_n3658_), .B(new_n3361_), .Y(new_n3660_));
  OAI21X1  g03468(.A0(new_n3660_), .A1(new_n3564_), .B0(new_n3364_), .Y(new_n3661_));
  AND2X1   g03469(.A(new_n3661_), .B(new_n3659_), .Y(new_n3662_));
  OR2X1    g03470(.A(new_n3638_), .B(new_n2570_), .Y(new_n3663_));
  AND2X1   g03471(.A(new_n3621_), .B(new_n3611_), .Y(new_n3664_));
  INVX1    g03472(.A(new_n3627_), .Y(new_n3665_));
  OR2X1    g03473(.A(new_n3628_), .B(\asqrt[45] ), .Y(new_n3666_));
  OAI21X1  g03474(.A0(new_n3666_), .A1(new_n3664_), .B0(new_n3665_), .Y(new_n3667_));
  AOI21X1  g03475(.A0(new_n3667_), .A1(new_n3663_), .B0(new_n2263_), .Y(new_n3668_));
  AOI21X1  g03476(.A0(new_n3609_), .A1(\asqrt[45] ), .B0(\asqrt[46] ), .Y(new_n3669_));
  AOI21X1  g03477(.A0(new_n3669_), .A1(new_n3667_), .B0(new_n3636_), .Y(new_n3670_));
  OAI21X1  g03478(.A0(new_n3670_), .A1(new_n3668_), .B0(\asqrt[47] ), .Y(new_n3671_));
  INVX1    g03479(.A(new_n3644_), .Y(new_n3672_));
  NOR3X1   g03480(.A(new_n3670_), .B(new_n3668_), .C(\asqrt[47] ), .Y(new_n3673_));
  OAI21X1  g03481(.A0(new_n3673_), .A1(new_n3672_), .B0(new_n3671_), .Y(new_n3674_));
  AOI21X1  g03482(.A0(new_n3674_), .A1(\asqrt[48] ), .B0(\asqrt[49] ), .Y(new_n3675_));
  AOI21X1  g03483(.A0(new_n3675_), .A1(new_n3656_), .B0(new_n3662_), .Y(new_n3676_));
  OAI21X1  g03484(.A0(new_n3676_), .A1(new_n3657_), .B0(\asqrt[50] ), .Y(new_n3677_));
  OR4X1    g03485(.A(new_n3564_), .B(new_n3375_), .C(new_n3378_), .D(new_n3401_), .Y(new_n3678_));
  NAND2X1  g03486(.A(new_n3386_), .B(new_n3369_), .Y(new_n3679_));
  OAI21X1  g03487(.A0(new_n3679_), .A1(new_n3564_), .B0(new_n3378_), .Y(new_n3680_));
  AND2X1   g03488(.A(new_n3680_), .B(new_n3678_), .Y(new_n3681_));
  NOR3X1   g03489(.A(new_n3676_), .B(new_n3657_), .C(\asqrt[50] ), .Y(new_n3682_));
  OAI21X1  g03490(.A0(new_n3682_), .A1(new_n3681_), .B0(new_n3677_), .Y(new_n3683_));
  AND2X1   g03491(.A(new_n3683_), .B(\asqrt[51] ), .Y(new_n3684_));
  INVX1    g03492(.A(new_n3681_), .Y(new_n3685_));
  AND2X1   g03493(.A(new_n3674_), .B(\asqrt[48] ), .Y(new_n3686_));
  NAND2X1  g03494(.A(new_n3645_), .B(new_n3644_), .Y(new_n3687_));
  NOR2X1   g03495(.A(new_n3641_), .B(\asqrt[48] ), .Y(new_n3688_));
  AOI21X1  g03496(.A0(new_n3688_), .A1(new_n3687_), .B0(new_n3653_), .Y(new_n3689_));
  OAI21X1  g03497(.A0(new_n3689_), .A1(new_n3686_), .B0(\asqrt[49] ), .Y(new_n3690_));
  INVX1    g03498(.A(new_n3662_), .Y(new_n3691_));
  OAI21X1  g03499(.A0(new_n3646_), .A1(new_n1834_), .B0(new_n1632_), .Y(new_n3692_));
  OAI21X1  g03500(.A0(new_n3692_), .A1(new_n3689_), .B0(new_n3691_), .Y(new_n3693_));
  NAND3X1  g03501(.A(new_n3693_), .B(new_n3690_), .C(new_n1469_), .Y(new_n3694_));
  NAND2X1  g03502(.A(new_n3694_), .B(new_n3685_), .Y(new_n3695_));
  OAI21X1  g03503(.A0(new_n3425_), .A1(new_n3423_), .B0(new_n3392_), .Y(new_n3696_));
  OR2X1    g03504(.A(new_n3696_), .B(new_n3377_), .Y(new_n3697_));
  AOI22X1  g03505(.A0(new_n3393_), .A1(new_n3387_), .B0(new_n3376_), .B1(\asqrt[50] ), .Y(new_n3698_));
  AND2X1   g03506(.A(new_n3698_), .B(\asqrt[41] ), .Y(new_n3699_));
  OAI22X1  g03507(.A0(new_n3699_), .A1(new_n3392_), .B0(new_n3697_), .B1(new_n3564_), .Y(new_n3700_));
  INVX1    g03508(.A(new_n3700_), .Y(new_n3701_));
  AOI21X1  g03509(.A0(new_n3693_), .A1(new_n3690_), .B0(new_n1469_), .Y(new_n3702_));
  NOR2X1   g03510(.A(new_n3702_), .B(\asqrt[51] ), .Y(new_n3703_));
  AOI21X1  g03511(.A0(new_n3703_), .A1(new_n3695_), .B0(new_n3701_), .Y(new_n3704_));
  OAI21X1  g03512(.A0(new_n3704_), .A1(new_n3684_), .B0(\asqrt[52] ), .Y(new_n3705_));
  AND2X1   g03513(.A(new_n3428_), .B(new_n3426_), .Y(new_n3706_));
  OR4X1    g03514(.A(new_n3564_), .B(new_n3706_), .C(new_n3400_), .D(new_n3427_), .Y(new_n3707_));
  OR2X1    g03515(.A(new_n3706_), .B(new_n3427_), .Y(new_n3708_));
  OAI21X1  g03516(.A0(new_n3708_), .A1(new_n3564_), .B0(new_n3400_), .Y(new_n3709_));
  AND2X1   g03517(.A(new_n3709_), .B(new_n3707_), .Y(new_n3710_));
  INVX1    g03518(.A(new_n3710_), .Y(new_n3711_));
  AOI21X1  g03519(.A0(new_n3694_), .A1(new_n3685_), .B0(new_n3702_), .Y(new_n3712_));
  OAI21X1  g03520(.A0(new_n3712_), .A1(new_n1277_), .B0(new_n1111_), .Y(new_n3713_));
  OAI21X1  g03521(.A0(new_n3713_), .A1(new_n3704_), .B0(new_n3711_), .Y(new_n3714_));
  AOI21X1  g03522(.A0(new_n3714_), .A1(new_n3705_), .B0(new_n968_), .Y(new_n3715_));
  OR4X1    g03523(.A(new_n3564_), .B(new_n3438_), .C(new_n3411_), .D(new_n3405_), .Y(new_n3716_));
  NAND2X1  g03524(.A(new_n3412_), .B(new_n3430_), .Y(new_n3717_));
  OAI21X1  g03525(.A0(new_n3717_), .A1(new_n3564_), .B0(new_n3411_), .Y(new_n3718_));
  AND2X1   g03526(.A(new_n3718_), .B(new_n3716_), .Y(new_n3719_));
  INVX1    g03527(.A(new_n3719_), .Y(new_n3720_));
  NAND3X1  g03528(.A(new_n3714_), .B(new_n3705_), .C(new_n968_), .Y(new_n3721_));
  AOI21X1  g03529(.A0(new_n3721_), .A1(new_n3720_), .B0(new_n3715_), .Y(new_n3722_));
  OR2X1    g03530(.A(new_n3722_), .B(new_n902_), .Y(new_n3723_));
  AND2X1   g03531(.A(new_n3721_), .B(new_n3720_), .Y(new_n3724_));
  AND2X1   g03532(.A(new_n3467_), .B(new_n3466_), .Y(new_n3725_));
  NOR3X1   g03533(.A(new_n3725_), .B(new_n3421_), .C(new_n3465_), .Y(new_n3726_));
  AOI22X1  g03534(.A0(new_n3467_), .A1(new_n3466_), .B0(new_n3439_), .B1(\asqrt[53] ), .Y(new_n3727_));
  AOI21X1  g03535(.A0(new_n3727_), .A1(\asqrt[41] ), .B0(new_n3420_), .Y(new_n3728_));
  AOI21X1  g03536(.A0(new_n3726_), .A1(\asqrt[41] ), .B0(new_n3728_), .Y(new_n3729_));
  INVX1    g03537(.A(new_n3729_), .Y(new_n3730_));
  OR2X1    g03538(.A(new_n3715_), .B(\asqrt[54] ), .Y(new_n3731_));
  OAI21X1  g03539(.A0(new_n3731_), .A1(new_n3724_), .B0(new_n3730_), .Y(new_n3732_));
  AOI21X1  g03540(.A0(new_n3732_), .A1(new_n3723_), .B0(new_n697_), .Y(new_n3733_));
  AOI21X1  g03541(.A0(new_n3440_), .A1(new_n3432_), .B0(new_n3470_), .Y(new_n3734_));
  NAND3X1  g03542(.A(new_n3734_), .B(\asqrt[41] ), .C(new_n3469_), .Y(new_n3735_));
  OAI21X1  g03543(.A0(new_n3471_), .A1(new_n3468_), .B0(new_n3469_), .Y(new_n3736_));
  OAI21X1  g03544(.A0(new_n3736_), .A1(new_n3564_), .B0(new_n3470_), .Y(new_n3737_));
  AND2X1   g03545(.A(new_n3737_), .B(new_n3735_), .Y(new_n3738_));
  OR2X1    g03546(.A(new_n3712_), .B(new_n1277_), .Y(new_n3739_));
  AND2X1   g03547(.A(new_n3694_), .B(new_n3685_), .Y(new_n3740_));
  OR2X1    g03548(.A(new_n3702_), .B(\asqrt[51] ), .Y(new_n3741_));
  OAI21X1  g03549(.A0(new_n3741_), .A1(new_n3740_), .B0(new_n3700_), .Y(new_n3742_));
  AOI21X1  g03550(.A0(new_n3742_), .A1(new_n3739_), .B0(new_n1111_), .Y(new_n3743_));
  AOI21X1  g03551(.A0(new_n3683_), .A1(\asqrt[51] ), .B0(\asqrt[52] ), .Y(new_n3744_));
  AOI21X1  g03552(.A0(new_n3744_), .A1(new_n3742_), .B0(new_n3710_), .Y(new_n3745_));
  OAI21X1  g03553(.A0(new_n3745_), .A1(new_n3743_), .B0(\asqrt[53] ), .Y(new_n3746_));
  NOR3X1   g03554(.A(new_n3745_), .B(new_n3743_), .C(\asqrt[53] ), .Y(new_n3747_));
  OAI21X1  g03555(.A0(new_n3747_), .A1(new_n3719_), .B0(new_n3746_), .Y(new_n3748_));
  AOI21X1  g03556(.A0(new_n3748_), .A1(\asqrt[54] ), .B0(\asqrt[55] ), .Y(new_n3749_));
  AOI21X1  g03557(.A0(new_n3749_), .A1(new_n3732_), .B0(new_n3738_), .Y(new_n3750_));
  OAI21X1  g03558(.A0(new_n3750_), .A1(new_n3733_), .B0(\asqrt[56] ), .Y(new_n3751_));
  NOR3X1   g03559(.A(new_n3750_), .B(new_n3733_), .C(\asqrt[56] ), .Y(new_n3752_));
  OR4X1    g03560(.A(new_n3564_), .B(new_n3475_), .C(new_n3443_), .D(new_n3473_), .Y(new_n3753_));
  OR2X1    g03561(.A(new_n3443_), .B(new_n3473_), .Y(new_n3754_));
  OAI21X1  g03562(.A0(new_n3754_), .A1(new_n3564_), .B0(new_n3475_), .Y(new_n3755_));
  AND2X1   g03563(.A(new_n3755_), .B(new_n3753_), .Y(new_n3756_));
  OAI21X1  g03564(.A0(new_n3756_), .A1(new_n3752_), .B0(new_n3751_), .Y(new_n3757_));
  AND2X1   g03565(.A(new_n3757_), .B(\asqrt[57] ), .Y(new_n3758_));
  AND2X1   g03566(.A(new_n3748_), .B(\asqrt[54] ), .Y(new_n3759_));
  NAND2X1  g03567(.A(new_n3721_), .B(new_n3720_), .Y(new_n3760_));
  NOR2X1   g03568(.A(new_n3715_), .B(\asqrt[54] ), .Y(new_n3761_));
  AOI21X1  g03569(.A0(new_n3761_), .A1(new_n3760_), .B0(new_n3729_), .Y(new_n3762_));
  OAI21X1  g03570(.A0(new_n3762_), .A1(new_n3759_), .B0(\asqrt[55] ), .Y(new_n3763_));
  INVX1    g03571(.A(new_n3738_), .Y(new_n3764_));
  OAI21X1  g03572(.A0(new_n3722_), .A1(new_n902_), .B0(new_n697_), .Y(new_n3765_));
  OAI21X1  g03573(.A0(new_n3765_), .A1(new_n3762_), .B0(new_n3764_), .Y(new_n3766_));
  NAND3X1  g03574(.A(new_n3766_), .B(new_n3763_), .C(new_n582_), .Y(new_n3767_));
  INVX1    g03575(.A(new_n3756_), .Y(new_n3768_));
  NAND2X1  g03576(.A(new_n3768_), .B(new_n3767_), .Y(new_n3769_));
  OAI21X1  g03577(.A0(new_n3499_), .A1(new_n3497_), .B0(new_n3456_), .Y(new_n3770_));
  OR2X1    g03578(.A(new_n3770_), .B(new_n3450_), .Y(new_n3771_));
  AOI22X1  g03579(.A0(new_n3457_), .A1(new_n3451_), .B0(new_n3449_), .B1(\asqrt[56] ), .Y(new_n3772_));
  AND2X1   g03580(.A(new_n3772_), .B(\asqrt[41] ), .Y(new_n3773_));
  OAI22X1  g03581(.A0(new_n3773_), .A1(new_n3456_), .B0(new_n3771_), .B1(new_n3564_), .Y(new_n3774_));
  INVX1    g03582(.A(new_n3774_), .Y(new_n3775_));
  AOI21X1  g03583(.A0(new_n3766_), .A1(new_n3763_), .B0(new_n582_), .Y(new_n3776_));
  NOR2X1   g03584(.A(new_n3776_), .B(\asqrt[57] ), .Y(new_n3777_));
  AOI21X1  g03585(.A0(new_n3777_), .A1(new_n3769_), .B0(new_n3775_), .Y(new_n3778_));
  OAI21X1  g03586(.A0(new_n3778_), .A1(new_n3758_), .B0(\asqrt[58] ), .Y(new_n3779_));
  AND2X1   g03587(.A(new_n3502_), .B(new_n3500_), .Y(new_n3780_));
  OR4X1    g03588(.A(new_n3564_), .B(new_n3780_), .C(new_n3464_), .D(new_n3501_), .Y(new_n3781_));
  OR2X1    g03589(.A(new_n3780_), .B(new_n3501_), .Y(new_n3782_));
  OAI21X1  g03590(.A0(new_n3782_), .A1(new_n3564_), .B0(new_n3464_), .Y(new_n3783_));
  AND2X1   g03591(.A(new_n3783_), .B(new_n3781_), .Y(new_n3784_));
  INVX1    g03592(.A(new_n3784_), .Y(new_n3785_));
  AOI21X1  g03593(.A0(new_n3768_), .A1(new_n3767_), .B0(new_n3776_), .Y(new_n3786_));
  OAI21X1  g03594(.A0(new_n3786_), .A1(new_n481_), .B0(new_n399_), .Y(new_n3787_));
  OAI21X1  g03595(.A0(new_n3787_), .A1(new_n3778_), .B0(new_n3785_), .Y(new_n3788_));
  AOI21X1  g03596(.A0(new_n3788_), .A1(new_n3779_), .B0(new_n328_), .Y(new_n3789_));
  OR4X1    g03597(.A(new_n3564_), .B(new_n3512_), .C(new_n3485_), .D(new_n3479_), .Y(new_n3790_));
  NAND2X1  g03598(.A(new_n3486_), .B(new_n3504_), .Y(new_n3791_));
  OAI21X1  g03599(.A0(new_n3791_), .A1(new_n3564_), .B0(new_n3485_), .Y(new_n3792_));
  AND2X1   g03600(.A(new_n3792_), .B(new_n3790_), .Y(new_n3793_));
  INVX1    g03601(.A(new_n3793_), .Y(new_n3794_));
  NAND3X1  g03602(.A(new_n3788_), .B(new_n3779_), .C(new_n328_), .Y(new_n3795_));
  AOI21X1  g03603(.A0(new_n3795_), .A1(new_n3794_), .B0(new_n3789_), .Y(new_n3796_));
  OR2X1    g03604(.A(new_n3796_), .B(new_n292_), .Y(new_n3797_));
  OR2X1    g03605(.A(new_n3786_), .B(new_n481_), .Y(new_n3798_));
  AND2X1   g03606(.A(new_n3768_), .B(new_n3767_), .Y(new_n3799_));
  OR2X1    g03607(.A(new_n3776_), .B(\asqrt[57] ), .Y(new_n3800_));
  OAI21X1  g03608(.A0(new_n3800_), .A1(new_n3799_), .B0(new_n3774_), .Y(new_n3801_));
  AOI21X1  g03609(.A0(new_n3801_), .A1(new_n3798_), .B0(new_n399_), .Y(new_n3802_));
  AOI21X1  g03610(.A0(new_n3757_), .A1(\asqrt[57] ), .B0(\asqrt[58] ), .Y(new_n3803_));
  AOI21X1  g03611(.A0(new_n3803_), .A1(new_n3801_), .B0(new_n3784_), .Y(new_n3804_));
  NOR3X1   g03612(.A(new_n3804_), .B(new_n3802_), .C(\asqrt[59] ), .Y(new_n3805_));
  NOR2X1   g03613(.A(new_n3805_), .B(new_n3793_), .Y(new_n3806_));
  AND2X1   g03614(.A(new_n3528_), .B(new_n3527_), .Y(new_n3807_));
  OAI21X1  g03615(.A0(new_n3487_), .A1(new_n328_), .B0(new_n3494_), .Y(new_n3808_));
  OR2X1    g03616(.A(new_n3808_), .B(new_n3807_), .Y(new_n3809_));
  NOR3X1   g03617(.A(new_n3564_), .B(new_n3807_), .C(new_n3526_), .Y(new_n3810_));
  OAI22X1  g03618(.A0(new_n3810_), .A1(new_n3494_), .B0(new_n3809_), .B1(new_n3564_), .Y(new_n3811_));
  OAI21X1  g03619(.A0(new_n3804_), .A1(new_n3802_), .B0(\asqrt[59] ), .Y(new_n3812_));
  NAND2X1  g03620(.A(new_n3812_), .B(new_n292_), .Y(new_n3813_));
  OAI21X1  g03621(.A0(new_n3813_), .A1(new_n3806_), .B0(new_n3811_), .Y(new_n3814_));
  AOI21X1  g03622(.A0(new_n3814_), .A1(new_n3797_), .B0(new_n217_), .Y(new_n3815_));
  AND2X1   g03623(.A(new_n3514_), .B(new_n3506_), .Y(new_n3816_));
  NOR4X1   g03624(.A(new_n3564_), .B(new_n3816_), .C(new_n3531_), .D(new_n3507_), .Y(new_n3817_));
  NOR2X1   g03625(.A(new_n3816_), .B(new_n3507_), .Y(new_n3818_));
  AOI21X1  g03626(.A0(new_n3818_), .A1(\asqrt[41] ), .B0(new_n3511_), .Y(new_n3819_));
  NOR2X1   g03627(.A(new_n3819_), .B(new_n3817_), .Y(new_n3820_));
  OAI21X1  g03628(.A0(new_n3805_), .A1(new_n3793_), .B0(new_n3812_), .Y(new_n3821_));
  AOI21X1  g03629(.A0(new_n3821_), .A1(\asqrt[60] ), .B0(\asqrt[61] ), .Y(new_n3822_));
  AOI21X1  g03630(.A0(new_n3822_), .A1(new_n3814_), .B0(new_n3820_), .Y(new_n3823_));
  OAI21X1  g03631(.A0(new_n3823_), .A1(new_n3815_), .B0(\asqrt[62] ), .Y(new_n3824_));
  OR4X1    g03632(.A(new_n3564_), .B(new_n3522_), .C(new_n3525_), .D(new_n3541_), .Y(new_n3825_));
  NAND2X1  g03633(.A(new_n3534_), .B(new_n3516_), .Y(new_n3826_));
  OAI21X1  g03634(.A0(new_n3826_), .A1(new_n3564_), .B0(new_n3525_), .Y(new_n3827_));
  AND2X1   g03635(.A(new_n3827_), .B(new_n3825_), .Y(new_n3828_));
  NOR3X1   g03636(.A(new_n3823_), .B(new_n3815_), .C(\asqrt[62] ), .Y(new_n3829_));
  OAI21X1  g03637(.A0(new_n3829_), .A1(new_n3828_), .B0(new_n3824_), .Y(new_n3830_));
  AND2X1   g03638(.A(new_n3542_), .B(new_n3535_), .Y(new_n3831_));
  NOR4X1   g03639(.A(new_n3564_), .B(new_n3831_), .C(new_n3581_), .D(new_n3524_), .Y(new_n3832_));
  AOI22X1  g03640(.A0(new_n3542_), .A1(new_n3535_), .B0(new_n3523_), .B1(\asqrt[62] ), .Y(new_n3833_));
  AOI21X1  g03641(.A0(new_n3833_), .A1(\asqrt[41] ), .B0(new_n3540_), .Y(new_n3834_));
  NOR2X1   g03642(.A(new_n3834_), .B(new_n3832_), .Y(new_n3835_));
  INVX1    g03643(.A(new_n3835_), .Y(new_n3836_));
  AND2X1   g03644(.A(new_n3586_), .B(new_n3583_), .Y(new_n3837_));
  AOI21X1  g03645(.A0(new_n3583_), .A1(new_n3579_), .B0(new_n3547_), .Y(new_n3838_));
  AOI21X1  g03646(.A0(new_n3838_), .A1(\asqrt[41] ), .B0(new_n3837_), .Y(new_n3839_));
  AND2X1   g03647(.A(new_n3839_), .B(new_n3836_), .Y(new_n3840_));
  AOI21X1  g03648(.A0(new_n3840_), .A1(new_n3830_), .B0(\asqrt[63] ), .Y(new_n3841_));
  INVX1    g03649(.A(new_n3828_), .Y(new_n3842_));
  AND2X1   g03650(.A(new_n3821_), .B(\asqrt[60] ), .Y(new_n3843_));
  OR2X1    g03651(.A(new_n3805_), .B(new_n3793_), .Y(new_n3844_));
  INVX1    g03652(.A(new_n3811_), .Y(new_n3845_));
  AND2X1   g03653(.A(new_n3812_), .B(new_n292_), .Y(new_n3846_));
  AOI21X1  g03654(.A0(new_n3846_), .A1(new_n3844_), .B0(new_n3845_), .Y(new_n3847_));
  OAI21X1  g03655(.A0(new_n3847_), .A1(new_n3843_), .B0(\asqrt[61] ), .Y(new_n3848_));
  INVX1    g03656(.A(new_n3820_), .Y(new_n3849_));
  OAI21X1  g03657(.A0(new_n3796_), .A1(new_n292_), .B0(new_n217_), .Y(new_n3850_));
  OAI21X1  g03658(.A0(new_n3850_), .A1(new_n3847_), .B0(new_n3849_), .Y(new_n3851_));
  NAND3X1  g03659(.A(new_n3851_), .B(new_n3848_), .C(new_n199_), .Y(new_n3852_));
  AND2X1   g03660(.A(new_n3852_), .B(new_n3842_), .Y(new_n3853_));
  NAND2X1  g03661(.A(new_n3835_), .B(new_n3824_), .Y(new_n3854_));
  OR2X1    g03662(.A(new_n3543_), .B(new_n3524_), .Y(new_n3855_));
  AOI21X1  g03663(.A0(\asqrt[41] ), .A1(new_n3548_), .B0(new_n3855_), .Y(new_n3856_));
  NOR3X1   g03664(.A(new_n3856_), .B(new_n3838_), .C(new_n193_), .Y(new_n3857_));
  AND2X1   g03665(.A(new_n3552_), .B(new_n193_), .Y(new_n3858_));
  NAND4X1  g03666(.A(new_n3561_), .B(new_n3557_), .C(new_n3546_), .D(new_n3544_), .Y(new_n3859_));
  NOR3X1   g03667(.A(new_n3859_), .B(new_n3837_), .C(new_n3858_), .Y(new_n3860_));
  NOR2X1   g03668(.A(new_n3860_), .B(new_n3857_), .Y(new_n3861_));
  OAI21X1  g03669(.A0(new_n3854_), .A1(new_n3853_), .B0(new_n3861_), .Y(new_n3862_));
  NOR2X1   g03670(.A(new_n3862_), .B(new_n3841_), .Y(new_n3863_));
  INVX1    g03671(.A(new_n3863_), .Y(\asqrt[40] ));
  INVX1    g03672(.A(\a[80] ), .Y(new_n3865_));
  NOR2X1   g03673(.A(\a[79] ), .B(\a[78] ), .Y(new_n3866_));
  NAND2X1  g03674(.A(new_n3866_), .B(new_n3865_), .Y(new_n3867_));
  OAI21X1  g03675(.A0(new_n3863_), .A1(new_n3865_), .B0(new_n3867_), .Y(new_n3868_));
  AOI21X1  g03676(.A0(new_n3851_), .A1(new_n3848_), .B0(new_n199_), .Y(new_n3869_));
  AOI21X1  g03677(.A0(new_n3852_), .A1(new_n3842_), .B0(new_n3869_), .Y(new_n3870_));
  INVX1    g03678(.A(new_n3840_), .Y(new_n3871_));
  OAI21X1  g03679(.A0(new_n3871_), .A1(new_n3870_), .B0(new_n193_), .Y(new_n3872_));
  OR2X1    g03680(.A(new_n3829_), .B(new_n3828_), .Y(new_n3873_));
  AND2X1   g03681(.A(new_n3835_), .B(new_n3824_), .Y(new_n3874_));
  INVX1    g03682(.A(new_n3861_), .Y(new_n3875_));
  AOI21X1  g03683(.A0(new_n3874_), .A1(new_n3873_), .B0(new_n3875_), .Y(new_n3876_));
  AOI21X1  g03684(.A0(new_n3876_), .A1(new_n3872_), .B0(new_n3865_), .Y(new_n3877_));
  NAND3X1  g03685(.A(new_n3867_), .B(new_n3561_), .C(new_n3557_), .Y(new_n3878_));
  OR4X1    g03686(.A(new_n3878_), .B(new_n3877_), .C(new_n3837_), .D(new_n3858_), .Y(new_n3879_));
  OAI21X1  g03687(.A0(new_n3862_), .A1(new_n3841_), .B0(new_n3865_), .Y(new_n3880_));
  AOI21X1  g03688(.A0(new_n3876_), .A1(new_n3872_), .B0(new_n3566_), .Y(new_n3881_));
  AOI21X1  g03689(.A0(new_n3880_), .A1(\a[81] ), .B0(new_n3881_), .Y(new_n3882_));
  AOI22X1  g03690(.A0(new_n3882_), .A1(new_n3879_), .B0(new_n3868_), .B1(\asqrt[41] ), .Y(new_n3883_));
  OR2X1    g03691(.A(new_n3883_), .B(new_n3276_), .Y(new_n3884_));
  AND2X1   g03692(.A(new_n3882_), .B(new_n3879_), .Y(new_n3885_));
  INVX1    g03693(.A(new_n3866_), .Y(new_n3886_));
  MX2X1    g03694(.A(new_n3886_), .B(new_n3863_), .S0(\a[80] ), .Y(new_n3887_));
  OAI21X1  g03695(.A0(new_n3887_), .A1(new_n3564_), .B0(new_n3276_), .Y(new_n3888_));
  OAI21X1  g03696(.A0(new_n3862_), .A1(new_n3841_), .B0(new_n3565_), .Y(new_n3889_));
  AND2X1   g03697(.A(new_n3874_), .B(new_n3873_), .Y(new_n3890_));
  OR2X1    g03698(.A(new_n3860_), .B(new_n3564_), .Y(new_n3891_));
  OR4X1    g03699(.A(new_n3891_), .B(new_n3857_), .C(new_n3890_), .D(new_n3841_), .Y(new_n3892_));
  AOI21X1  g03700(.A0(new_n3892_), .A1(new_n3889_), .B0(new_n3569_), .Y(new_n3893_));
  NOR4X1   g03701(.A(new_n3891_), .B(new_n3857_), .C(new_n3890_), .D(new_n3841_), .Y(new_n3894_));
  NOR3X1   g03702(.A(new_n3894_), .B(new_n3881_), .C(\a[82] ), .Y(new_n3895_));
  OR2X1    g03703(.A(new_n3895_), .B(new_n3893_), .Y(new_n3896_));
  OAI21X1  g03704(.A0(new_n3888_), .A1(new_n3885_), .B0(new_n3896_), .Y(new_n3897_));
  AOI21X1  g03705(.A0(new_n3897_), .A1(new_n3884_), .B0(new_n3008_), .Y(new_n3898_));
  AND2X1   g03706(.A(new_n3576_), .B(new_n3575_), .Y(new_n3899_));
  NOR3X1   g03707(.A(new_n3899_), .B(new_n3613_), .C(new_n3612_), .Y(new_n3900_));
  OAI21X1  g03708(.A0(new_n3862_), .A1(new_n3841_), .B0(new_n3900_), .Y(new_n3901_));
  AOI21X1  g03709(.A0(new_n3590_), .A1(\asqrt[42] ), .B0(new_n3613_), .Y(new_n3902_));
  OAI21X1  g03710(.A0(new_n3862_), .A1(new_n3841_), .B0(new_n3902_), .Y(new_n3903_));
  NAND2X1  g03711(.A(new_n3903_), .B(new_n3899_), .Y(new_n3904_));
  NOR4X1   g03712(.A(new_n3878_), .B(new_n3877_), .C(new_n3837_), .D(new_n3858_), .Y(new_n3905_));
  INVX1    g03713(.A(\a[81] ), .Y(new_n3906_));
  AOI21X1  g03714(.A0(new_n3876_), .A1(new_n3872_), .B0(\a[80] ), .Y(new_n3907_));
  OAI21X1  g03715(.A0(new_n3907_), .A1(new_n3906_), .B0(new_n3889_), .Y(new_n3908_));
  OAI22X1  g03716(.A0(new_n3908_), .A1(new_n3905_), .B0(new_n3887_), .B1(new_n3564_), .Y(new_n3909_));
  AOI21X1  g03717(.A0(new_n3909_), .A1(\asqrt[42] ), .B0(\asqrt[43] ), .Y(new_n3910_));
  AOI22X1  g03718(.A0(new_n3910_), .A1(new_n3897_), .B0(new_n3904_), .B1(new_n3901_), .Y(new_n3911_));
  OAI21X1  g03719(.A0(new_n3911_), .A1(new_n3898_), .B0(\asqrt[44] ), .Y(new_n3912_));
  AND2X1   g03720(.A(new_n3591_), .B(new_n3577_), .Y(new_n3913_));
  NOR3X1   g03721(.A(new_n3619_), .B(new_n3913_), .C(new_n3578_), .Y(new_n3914_));
  OAI21X1  g03722(.A0(new_n3862_), .A1(new_n3841_), .B0(new_n3914_), .Y(new_n3915_));
  NOR2X1   g03723(.A(new_n3913_), .B(new_n3578_), .Y(new_n3916_));
  OAI21X1  g03724(.A0(new_n3862_), .A1(new_n3841_), .B0(new_n3916_), .Y(new_n3917_));
  NAND2X1  g03725(.A(new_n3917_), .B(new_n3619_), .Y(new_n3918_));
  AND2X1   g03726(.A(new_n3918_), .B(new_n3915_), .Y(new_n3919_));
  NOR3X1   g03727(.A(new_n3911_), .B(new_n3898_), .C(\asqrt[44] ), .Y(new_n3920_));
  OAI21X1  g03728(.A0(new_n3920_), .A1(new_n3919_), .B0(new_n3912_), .Y(new_n3921_));
  AND2X1   g03729(.A(new_n3921_), .B(\asqrt[45] ), .Y(new_n3922_));
  OR2X1    g03730(.A(new_n3920_), .B(new_n3919_), .Y(new_n3923_));
  NOR3X1   g03731(.A(new_n3608_), .B(new_n3611_), .C(new_n3628_), .Y(new_n3924_));
  OAI21X1  g03732(.A0(new_n3862_), .A1(new_n3841_), .B0(new_n3924_), .Y(new_n3925_));
  NOR3X1   g03733(.A(new_n3863_), .B(new_n3608_), .C(new_n3628_), .Y(new_n3926_));
  OR2X1    g03734(.A(new_n3926_), .B(new_n3607_), .Y(new_n3927_));
  AND2X1   g03735(.A(new_n3927_), .B(new_n3925_), .Y(new_n3928_));
  AND2X1   g03736(.A(new_n3909_), .B(\asqrt[42] ), .Y(new_n3929_));
  NAND2X1  g03737(.A(new_n3882_), .B(new_n3879_), .Y(new_n3930_));
  AOI21X1  g03738(.A0(new_n3868_), .A1(\asqrt[41] ), .B0(\asqrt[42] ), .Y(new_n3931_));
  NOR2X1   g03739(.A(new_n3895_), .B(new_n3893_), .Y(new_n3932_));
  AOI21X1  g03740(.A0(new_n3931_), .A1(new_n3930_), .B0(new_n3932_), .Y(new_n3933_));
  OAI21X1  g03741(.A0(new_n3933_), .A1(new_n3929_), .B0(\asqrt[43] ), .Y(new_n3934_));
  NAND2X1  g03742(.A(new_n3904_), .B(new_n3901_), .Y(new_n3935_));
  OAI21X1  g03743(.A0(new_n3883_), .A1(new_n3276_), .B0(new_n3008_), .Y(new_n3936_));
  OAI21X1  g03744(.A0(new_n3936_), .A1(new_n3933_), .B0(new_n3935_), .Y(new_n3937_));
  AOI21X1  g03745(.A0(new_n3937_), .A1(new_n3934_), .B0(new_n2769_), .Y(new_n3938_));
  NOR2X1   g03746(.A(new_n3938_), .B(\asqrt[45] ), .Y(new_n3939_));
  AOI21X1  g03747(.A0(new_n3939_), .A1(new_n3923_), .B0(new_n3928_), .Y(new_n3940_));
  OAI21X1  g03748(.A0(new_n3940_), .A1(new_n3922_), .B0(\asqrt[46] ), .Y(new_n3941_));
  AOI21X1  g03749(.A0(new_n3629_), .A1(new_n3622_), .B0(new_n3665_), .Y(new_n3942_));
  AND2X1   g03750(.A(new_n3942_), .B(new_n3663_), .Y(new_n3943_));
  AOI22X1  g03751(.A0(new_n3629_), .A1(new_n3622_), .B0(new_n3609_), .B1(\asqrt[45] ), .Y(new_n3944_));
  AOI21X1  g03752(.A0(new_n3944_), .A1(\asqrt[40] ), .B0(new_n3627_), .Y(new_n3945_));
  AOI21X1  g03753(.A0(new_n3943_), .A1(\asqrt[40] ), .B0(new_n3945_), .Y(new_n3946_));
  INVX1    g03754(.A(new_n3946_), .Y(new_n3947_));
  INVX1    g03755(.A(new_n3919_), .Y(new_n3948_));
  NAND3X1  g03756(.A(new_n3937_), .B(new_n3934_), .C(new_n2769_), .Y(new_n3949_));
  AOI21X1  g03757(.A0(new_n3949_), .A1(new_n3948_), .B0(new_n3938_), .Y(new_n3950_));
  OAI21X1  g03758(.A0(new_n3950_), .A1(new_n2570_), .B0(new_n2263_), .Y(new_n3951_));
  OAI21X1  g03759(.A0(new_n3951_), .A1(new_n3940_), .B0(new_n3947_), .Y(new_n3952_));
  AOI21X1  g03760(.A0(new_n3952_), .A1(new_n3941_), .B0(new_n2040_), .Y(new_n3953_));
  AND2X1   g03761(.A(new_n3669_), .B(new_n3667_), .Y(new_n3954_));
  NOR3X1   g03762(.A(new_n3954_), .B(new_n3637_), .C(new_n3668_), .Y(new_n3955_));
  NOR3X1   g03763(.A(new_n3863_), .B(new_n3954_), .C(new_n3668_), .Y(new_n3956_));
  NOR2X1   g03764(.A(new_n3956_), .B(new_n3636_), .Y(new_n3957_));
  AOI21X1  g03765(.A0(new_n3955_), .A1(\asqrt[40] ), .B0(new_n3957_), .Y(new_n3958_));
  INVX1    g03766(.A(new_n3958_), .Y(new_n3959_));
  NAND3X1  g03767(.A(new_n3952_), .B(new_n3941_), .C(new_n2040_), .Y(new_n3960_));
  AOI21X1  g03768(.A0(new_n3960_), .A1(new_n3959_), .B0(new_n3953_), .Y(new_n3961_));
  OR2X1    g03769(.A(new_n3961_), .B(new_n1834_), .Y(new_n3962_));
  AND2X1   g03770(.A(new_n3960_), .B(new_n3959_), .Y(new_n3963_));
  OR4X1    g03771(.A(new_n3863_), .B(new_n3673_), .C(new_n3644_), .D(new_n3641_), .Y(new_n3964_));
  NAND2X1  g03772(.A(new_n3645_), .B(new_n3671_), .Y(new_n3965_));
  OAI21X1  g03773(.A0(new_n3965_), .A1(new_n3863_), .B0(new_n3644_), .Y(new_n3966_));
  AND2X1   g03774(.A(new_n3966_), .B(new_n3964_), .Y(new_n3967_));
  INVX1    g03775(.A(new_n3967_), .Y(new_n3968_));
  OR2X1    g03776(.A(new_n3953_), .B(\asqrt[48] ), .Y(new_n3969_));
  OAI21X1  g03777(.A0(new_n3969_), .A1(new_n3963_), .B0(new_n3968_), .Y(new_n3970_));
  AOI21X1  g03778(.A0(new_n3970_), .A1(new_n3962_), .B0(new_n1632_), .Y(new_n3971_));
  AND2X1   g03779(.A(new_n3688_), .B(new_n3687_), .Y(new_n3972_));
  NOR3X1   g03780(.A(new_n3972_), .B(new_n3654_), .C(new_n3686_), .Y(new_n3973_));
  NOR3X1   g03781(.A(new_n3863_), .B(new_n3972_), .C(new_n3686_), .Y(new_n3974_));
  NOR2X1   g03782(.A(new_n3974_), .B(new_n3653_), .Y(new_n3975_));
  AOI21X1  g03783(.A0(new_n3973_), .A1(\asqrt[40] ), .B0(new_n3975_), .Y(new_n3976_));
  OR2X1    g03784(.A(new_n3950_), .B(new_n2570_), .Y(new_n3977_));
  NOR2X1   g03785(.A(new_n3920_), .B(new_n3919_), .Y(new_n3978_));
  INVX1    g03786(.A(new_n3928_), .Y(new_n3979_));
  OR2X1    g03787(.A(new_n3938_), .B(\asqrt[45] ), .Y(new_n3980_));
  OAI21X1  g03788(.A0(new_n3980_), .A1(new_n3978_), .B0(new_n3979_), .Y(new_n3981_));
  AOI21X1  g03789(.A0(new_n3981_), .A1(new_n3977_), .B0(new_n2263_), .Y(new_n3982_));
  AOI21X1  g03790(.A0(new_n3921_), .A1(\asqrt[45] ), .B0(\asqrt[46] ), .Y(new_n3983_));
  AOI21X1  g03791(.A0(new_n3983_), .A1(new_n3981_), .B0(new_n3946_), .Y(new_n3984_));
  OAI21X1  g03792(.A0(new_n3984_), .A1(new_n3982_), .B0(\asqrt[47] ), .Y(new_n3985_));
  NOR3X1   g03793(.A(new_n3984_), .B(new_n3982_), .C(\asqrt[47] ), .Y(new_n3986_));
  OAI21X1  g03794(.A0(new_n3986_), .A1(new_n3958_), .B0(new_n3985_), .Y(new_n3987_));
  AOI21X1  g03795(.A0(new_n3987_), .A1(\asqrt[48] ), .B0(\asqrt[49] ), .Y(new_n3988_));
  AOI21X1  g03796(.A0(new_n3988_), .A1(new_n3970_), .B0(new_n3976_), .Y(new_n3989_));
  OAI21X1  g03797(.A0(new_n3989_), .A1(new_n3971_), .B0(\asqrt[50] ), .Y(new_n3990_));
  AND2X1   g03798(.A(new_n3675_), .B(new_n3656_), .Y(new_n3991_));
  NOR3X1   g03799(.A(new_n3991_), .B(new_n3691_), .C(new_n3657_), .Y(new_n3992_));
  NOR3X1   g03800(.A(new_n3863_), .B(new_n3991_), .C(new_n3657_), .Y(new_n3993_));
  NOR2X1   g03801(.A(new_n3993_), .B(new_n3662_), .Y(new_n3994_));
  AOI21X1  g03802(.A0(new_n3992_), .A1(\asqrt[40] ), .B0(new_n3994_), .Y(new_n3995_));
  NOR3X1   g03803(.A(new_n3989_), .B(new_n3971_), .C(\asqrt[50] ), .Y(new_n3996_));
  OAI21X1  g03804(.A0(new_n3996_), .A1(new_n3995_), .B0(new_n3990_), .Y(new_n3997_));
  AND2X1   g03805(.A(new_n3997_), .B(\asqrt[51] ), .Y(new_n3998_));
  INVX1    g03806(.A(new_n3995_), .Y(new_n3999_));
  AND2X1   g03807(.A(new_n3987_), .B(\asqrt[48] ), .Y(new_n4000_));
  OR2X1    g03808(.A(new_n3986_), .B(new_n3958_), .Y(new_n4001_));
  NOR2X1   g03809(.A(new_n3953_), .B(\asqrt[48] ), .Y(new_n4002_));
  AOI21X1  g03810(.A0(new_n4002_), .A1(new_n4001_), .B0(new_n3967_), .Y(new_n4003_));
  OAI21X1  g03811(.A0(new_n4003_), .A1(new_n4000_), .B0(\asqrt[49] ), .Y(new_n4004_));
  INVX1    g03812(.A(new_n3976_), .Y(new_n4005_));
  OAI21X1  g03813(.A0(new_n3961_), .A1(new_n1834_), .B0(new_n1632_), .Y(new_n4006_));
  OAI21X1  g03814(.A0(new_n4006_), .A1(new_n4003_), .B0(new_n4005_), .Y(new_n4007_));
  NAND3X1  g03815(.A(new_n4007_), .B(new_n4004_), .C(new_n1469_), .Y(new_n4008_));
  NAND2X1  g03816(.A(new_n4008_), .B(new_n3999_), .Y(new_n4009_));
  NAND4X1  g03817(.A(\asqrt[40] ), .B(new_n3694_), .C(new_n3681_), .D(new_n3677_), .Y(new_n4010_));
  NAND2X1  g03818(.A(new_n3694_), .B(new_n3677_), .Y(new_n4011_));
  OAI21X1  g03819(.A0(new_n4011_), .A1(new_n3863_), .B0(new_n3685_), .Y(new_n4012_));
  AND2X1   g03820(.A(new_n4012_), .B(new_n4010_), .Y(new_n4013_));
  AOI21X1  g03821(.A0(new_n4007_), .A1(new_n4004_), .B0(new_n1469_), .Y(new_n4014_));
  NOR2X1   g03822(.A(new_n4014_), .B(\asqrt[51] ), .Y(new_n4015_));
  AOI21X1  g03823(.A0(new_n4015_), .A1(new_n4009_), .B0(new_n4013_), .Y(new_n4016_));
  OAI21X1  g03824(.A0(new_n4016_), .A1(new_n3998_), .B0(\asqrt[52] ), .Y(new_n4017_));
  AOI21X1  g03825(.A0(new_n3703_), .A1(new_n3695_), .B0(new_n3700_), .Y(new_n4018_));
  AND2X1   g03826(.A(new_n4018_), .B(new_n3739_), .Y(new_n4019_));
  AOI22X1  g03827(.A0(new_n3703_), .A1(new_n3695_), .B0(new_n3683_), .B1(\asqrt[51] ), .Y(new_n4020_));
  AOI21X1  g03828(.A0(new_n4020_), .A1(\asqrt[40] ), .B0(new_n3701_), .Y(new_n4021_));
  AOI21X1  g03829(.A0(new_n4019_), .A1(\asqrt[40] ), .B0(new_n4021_), .Y(new_n4022_));
  INVX1    g03830(.A(new_n4022_), .Y(new_n4023_));
  AOI21X1  g03831(.A0(new_n4008_), .A1(new_n3999_), .B0(new_n4014_), .Y(new_n4024_));
  OAI21X1  g03832(.A0(new_n4024_), .A1(new_n1277_), .B0(new_n1111_), .Y(new_n4025_));
  OAI21X1  g03833(.A0(new_n4025_), .A1(new_n4016_), .B0(new_n4023_), .Y(new_n4026_));
  AOI21X1  g03834(.A0(new_n4026_), .A1(new_n4017_), .B0(new_n968_), .Y(new_n4027_));
  AND2X1   g03835(.A(new_n3744_), .B(new_n3742_), .Y(new_n4028_));
  NOR3X1   g03836(.A(new_n4028_), .B(new_n3711_), .C(new_n3743_), .Y(new_n4029_));
  NOR3X1   g03837(.A(new_n3863_), .B(new_n4028_), .C(new_n3743_), .Y(new_n4030_));
  NOR2X1   g03838(.A(new_n4030_), .B(new_n3710_), .Y(new_n4031_));
  AOI21X1  g03839(.A0(new_n4029_), .A1(\asqrt[40] ), .B0(new_n4031_), .Y(new_n4032_));
  INVX1    g03840(.A(new_n4032_), .Y(new_n4033_));
  NAND3X1  g03841(.A(new_n4026_), .B(new_n4017_), .C(new_n968_), .Y(new_n4034_));
  AOI21X1  g03842(.A0(new_n4034_), .A1(new_n4033_), .B0(new_n4027_), .Y(new_n4035_));
  OR2X1    g03843(.A(new_n4035_), .B(new_n902_), .Y(new_n4036_));
  AND2X1   g03844(.A(new_n4034_), .B(new_n4033_), .Y(new_n4037_));
  NAND4X1  g03845(.A(\asqrt[40] ), .B(new_n3721_), .C(new_n3719_), .D(new_n3746_), .Y(new_n4038_));
  NAND2X1  g03846(.A(new_n3721_), .B(new_n3746_), .Y(new_n4039_));
  OAI21X1  g03847(.A0(new_n4039_), .A1(new_n3863_), .B0(new_n3720_), .Y(new_n4040_));
  AND2X1   g03848(.A(new_n4040_), .B(new_n4038_), .Y(new_n4041_));
  INVX1    g03849(.A(new_n4041_), .Y(new_n4042_));
  OR2X1    g03850(.A(new_n4027_), .B(\asqrt[54] ), .Y(new_n4043_));
  OAI21X1  g03851(.A0(new_n4043_), .A1(new_n4037_), .B0(new_n4042_), .Y(new_n4044_));
  AOI21X1  g03852(.A0(new_n4044_), .A1(new_n4036_), .B0(new_n697_), .Y(new_n4045_));
  AND2X1   g03853(.A(new_n3761_), .B(new_n3760_), .Y(new_n4046_));
  NOR3X1   g03854(.A(new_n4046_), .B(new_n3730_), .C(new_n3759_), .Y(new_n4047_));
  NOR3X1   g03855(.A(new_n3863_), .B(new_n4046_), .C(new_n3759_), .Y(new_n4048_));
  NOR2X1   g03856(.A(new_n4048_), .B(new_n3729_), .Y(new_n4049_));
  AOI21X1  g03857(.A0(new_n4047_), .A1(\asqrt[40] ), .B0(new_n4049_), .Y(new_n4050_));
  OR2X1    g03858(.A(new_n4024_), .B(new_n1277_), .Y(new_n4051_));
  AND2X1   g03859(.A(new_n4008_), .B(new_n3999_), .Y(new_n4052_));
  INVX1    g03860(.A(new_n4013_), .Y(new_n4053_));
  OR2X1    g03861(.A(new_n4014_), .B(\asqrt[51] ), .Y(new_n4054_));
  OAI21X1  g03862(.A0(new_n4054_), .A1(new_n4052_), .B0(new_n4053_), .Y(new_n4055_));
  AOI21X1  g03863(.A0(new_n4055_), .A1(new_n4051_), .B0(new_n1111_), .Y(new_n4056_));
  AOI21X1  g03864(.A0(new_n3997_), .A1(\asqrt[51] ), .B0(\asqrt[52] ), .Y(new_n4057_));
  AOI21X1  g03865(.A0(new_n4057_), .A1(new_n4055_), .B0(new_n4022_), .Y(new_n4058_));
  OAI21X1  g03866(.A0(new_n4058_), .A1(new_n4056_), .B0(\asqrt[53] ), .Y(new_n4059_));
  NOR3X1   g03867(.A(new_n4058_), .B(new_n4056_), .C(\asqrt[53] ), .Y(new_n4060_));
  OAI21X1  g03868(.A0(new_n4060_), .A1(new_n4032_), .B0(new_n4059_), .Y(new_n4061_));
  AOI21X1  g03869(.A0(new_n4061_), .A1(\asqrt[54] ), .B0(\asqrt[55] ), .Y(new_n4062_));
  AOI21X1  g03870(.A0(new_n4062_), .A1(new_n4044_), .B0(new_n4050_), .Y(new_n4063_));
  OAI21X1  g03871(.A0(new_n4063_), .A1(new_n4045_), .B0(\asqrt[56] ), .Y(new_n4064_));
  AND2X1   g03872(.A(new_n3749_), .B(new_n3732_), .Y(new_n4065_));
  NOR3X1   g03873(.A(new_n4065_), .B(new_n3764_), .C(new_n3733_), .Y(new_n4066_));
  NOR3X1   g03874(.A(new_n3863_), .B(new_n4065_), .C(new_n3733_), .Y(new_n4067_));
  NOR2X1   g03875(.A(new_n4067_), .B(new_n3738_), .Y(new_n4068_));
  AOI21X1  g03876(.A0(new_n4066_), .A1(\asqrt[40] ), .B0(new_n4068_), .Y(new_n4069_));
  NOR3X1   g03877(.A(new_n4063_), .B(new_n4045_), .C(\asqrt[56] ), .Y(new_n4070_));
  OAI21X1  g03878(.A0(new_n4070_), .A1(new_n4069_), .B0(new_n4064_), .Y(new_n4071_));
  AND2X1   g03879(.A(new_n4071_), .B(\asqrt[57] ), .Y(new_n4072_));
  OR2X1    g03880(.A(new_n4070_), .B(new_n4069_), .Y(new_n4073_));
  AND2X1   g03881(.A(new_n4064_), .B(new_n481_), .Y(new_n4074_));
  NAND4X1  g03882(.A(\asqrt[40] ), .B(new_n3756_), .C(new_n3767_), .D(new_n3751_), .Y(new_n4075_));
  NAND2X1  g03883(.A(new_n3767_), .B(new_n3751_), .Y(new_n4076_));
  OAI21X1  g03884(.A0(new_n4076_), .A1(new_n3863_), .B0(new_n3768_), .Y(new_n4077_));
  AND2X1   g03885(.A(new_n4077_), .B(new_n4075_), .Y(new_n4078_));
  AOI21X1  g03886(.A0(new_n4074_), .A1(new_n4073_), .B0(new_n4078_), .Y(new_n4079_));
  OAI21X1  g03887(.A0(new_n4079_), .A1(new_n4072_), .B0(\asqrt[58] ), .Y(new_n4080_));
  AOI21X1  g03888(.A0(new_n3777_), .A1(new_n3769_), .B0(new_n3774_), .Y(new_n4081_));
  AND2X1   g03889(.A(new_n4081_), .B(new_n3798_), .Y(new_n4082_));
  AOI22X1  g03890(.A0(new_n3777_), .A1(new_n3769_), .B0(new_n3757_), .B1(\asqrt[57] ), .Y(new_n4083_));
  AOI21X1  g03891(.A0(new_n4083_), .A1(\asqrt[40] ), .B0(new_n3775_), .Y(new_n4084_));
  AOI21X1  g03892(.A0(new_n4082_), .A1(\asqrt[40] ), .B0(new_n4084_), .Y(new_n4085_));
  INVX1    g03893(.A(new_n4085_), .Y(new_n4086_));
  AND2X1   g03894(.A(new_n4061_), .B(\asqrt[54] ), .Y(new_n4087_));
  NAND2X1  g03895(.A(new_n4034_), .B(new_n4033_), .Y(new_n4088_));
  NOR2X1   g03896(.A(new_n4027_), .B(\asqrt[54] ), .Y(new_n4089_));
  AOI21X1  g03897(.A0(new_n4089_), .A1(new_n4088_), .B0(new_n4041_), .Y(new_n4090_));
  OAI21X1  g03898(.A0(new_n4090_), .A1(new_n4087_), .B0(\asqrt[55] ), .Y(new_n4091_));
  INVX1    g03899(.A(new_n4050_), .Y(new_n4092_));
  OAI21X1  g03900(.A0(new_n4035_), .A1(new_n902_), .B0(new_n697_), .Y(new_n4093_));
  OAI21X1  g03901(.A0(new_n4093_), .A1(new_n4090_), .B0(new_n4092_), .Y(new_n4094_));
  AOI21X1  g03902(.A0(new_n4094_), .A1(new_n4091_), .B0(new_n582_), .Y(new_n4095_));
  INVX1    g03903(.A(new_n4069_), .Y(new_n4096_));
  NAND3X1  g03904(.A(new_n4094_), .B(new_n4091_), .C(new_n582_), .Y(new_n4097_));
  AOI21X1  g03905(.A0(new_n4097_), .A1(new_n4096_), .B0(new_n4095_), .Y(new_n4098_));
  OAI21X1  g03906(.A0(new_n4098_), .A1(new_n481_), .B0(new_n399_), .Y(new_n4099_));
  OAI21X1  g03907(.A0(new_n4099_), .A1(new_n4079_), .B0(new_n4086_), .Y(new_n4100_));
  AOI21X1  g03908(.A0(new_n4100_), .A1(new_n4080_), .B0(new_n328_), .Y(new_n4101_));
  AND2X1   g03909(.A(new_n3803_), .B(new_n3801_), .Y(new_n4102_));
  NOR3X1   g03910(.A(new_n4102_), .B(new_n3785_), .C(new_n3802_), .Y(new_n4103_));
  NOR3X1   g03911(.A(new_n3863_), .B(new_n4102_), .C(new_n3802_), .Y(new_n4104_));
  NOR2X1   g03912(.A(new_n4104_), .B(new_n3784_), .Y(new_n4105_));
  AOI21X1  g03913(.A0(new_n4103_), .A1(\asqrt[40] ), .B0(new_n4105_), .Y(new_n4106_));
  INVX1    g03914(.A(new_n4106_), .Y(new_n4107_));
  NAND3X1  g03915(.A(new_n4100_), .B(new_n4080_), .C(new_n328_), .Y(new_n4108_));
  AOI21X1  g03916(.A0(new_n4108_), .A1(new_n4107_), .B0(new_n4101_), .Y(new_n4109_));
  OR2X1    g03917(.A(new_n4109_), .B(new_n292_), .Y(new_n4110_));
  OR2X1    g03918(.A(new_n4098_), .B(new_n481_), .Y(new_n4111_));
  NOR2X1   g03919(.A(new_n4070_), .B(new_n4069_), .Y(new_n4112_));
  NAND2X1  g03920(.A(new_n4064_), .B(new_n481_), .Y(new_n4113_));
  INVX1    g03921(.A(new_n4078_), .Y(new_n4114_));
  OAI21X1  g03922(.A0(new_n4113_), .A1(new_n4112_), .B0(new_n4114_), .Y(new_n4115_));
  AOI21X1  g03923(.A0(new_n4115_), .A1(new_n4111_), .B0(new_n399_), .Y(new_n4116_));
  AOI21X1  g03924(.A0(new_n4071_), .A1(\asqrt[57] ), .B0(\asqrt[58] ), .Y(new_n4117_));
  AOI21X1  g03925(.A0(new_n4117_), .A1(new_n4115_), .B0(new_n4085_), .Y(new_n4118_));
  NOR3X1   g03926(.A(new_n4118_), .B(new_n4116_), .C(\asqrt[59] ), .Y(new_n4119_));
  NOR2X1   g03927(.A(new_n4119_), .B(new_n4106_), .Y(new_n4120_));
  OR4X1    g03928(.A(new_n3863_), .B(new_n3805_), .C(new_n3794_), .D(new_n3789_), .Y(new_n4121_));
  OR2X1    g03929(.A(new_n3805_), .B(new_n3789_), .Y(new_n4122_));
  OAI21X1  g03930(.A0(new_n4122_), .A1(new_n3863_), .B0(new_n3794_), .Y(new_n4123_));
  AND2X1   g03931(.A(new_n4123_), .B(new_n4121_), .Y(new_n4124_));
  INVX1    g03932(.A(new_n4124_), .Y(new_n4125_));
  OAI21X1  g03933(.A0(new_n4118_), .A1(new_n4116_), .B0(\asqrt[59] ), .Y(new_n4126_));
  NAND2X1  g03934(.A(new_n4126_), .B(new_n292_), .Y(new_n4127_));
  OAI21X1  g03935(.A0(new_n4127_), .A1(new_n4120_), .B0(new_n4125_), .Y(new_n4128_));
  AOI21X1  g03936(.A0(new_n4128_), .A1(new_n4110_), .B0(new_n217_), .Y(new_n4129_));
  AND2X1   g03937(.A(new_n3846_), .B(new_n3844_), .Y(new_n4130_));
  NOR3X1   g03938(.A(new_n4130_), .B(new_n3811_), .C(new_n3843_), .Y(new_n4131_));
  NOR3X1   g03939(.A(new_n3863_), .B(new_n4130_), .C(new_n3843_), .Y(new_n4132_));
  NOR2X1   g03940(.A(new_n4132_), .B(new_n3845_), .Y(new_n4133_));
  AOI21X1  g03941(.A0(new_n4131_), .A1(\asqrt[40] ), .B0(new_n4133_), .Y(new_n4134_));
  OAI21X1  g03942(.A0(new_n4119_), .A1(new_n4106_), .B0(new_n4126_), .Y(new_n4135_));
  AOI21X1  g03943(.A0(new_n4135_), .A1(\asqrt[60] ), .B0(\asqrt[61] ), .Y(new_n4136_));
  AOI21X1  g03944(.A0(new_n4136_), .A1(new_n4128_), .B0(new_n4134_), .Y(new_n4137_));
  OAI21X1  g03945(.A0(new_n4137_), .A1(new_n4129_), .B0(\asqrt[62] ), .Y(new_n4138_));
  AND2X1   g03946(.A(new_n3822_), .B(new_n3814_), .Y(new_n4139_));
  NOR3X1   g03947(.A(new_n4139_), .B(new_n3849_), .C(new_n3815_), .Y(new_n4140_));
  NOR3X1   g03948(.A(new_n3863_), .B(new_n4139_), .C(new_n3815_), .Y(new_n4141_));
  NOR2X1   g03949(.A(new_n4141_), .B(new_n3820_), .Y(new_n4142_));
  AOI21X1  g03950(.A0(new_n4140_), .A1(\asqrt[40] ), .B0(new_n4142_), .Y(new_n4143_));
  NOR3X1   g03951(.A(new_n4137_), .B(new_n4129_), .C(\asqrt[62] ), .Y(new_n4144_));
  OAI21X1  g03952(.A0(new_n4144_), .A1(new_n4143_), .B0(new_n4138_), .Y(new_n4145_));
  NOR4X1   g03953(.A(new_n3863_), .B(new_n3829_), .C(new_n3842_), .D(new_n3869_), .Y(new_n4146_));
  NAND3X1  g03954(.A(\asqrt[40] ), .B(new_n3852_), .C(new_n3824_), .Y(new_n4147_));
  AOI21X1  g03955(.A0(new_n4147_), .A1(new_n3842_), .B0(new_n4146_), .Y(new_n4148_));
  INVX1    g03956(.A(new_n4148_), .Y(new_n4149_));
  AND2X1   g03957(.A(new_n3836_), .B(new_n3830_), .Y(new_n4150_));
  AOI21X1  g03958(.A0(new_n4150_), .A1(\asqrt[40] ), .B0(new_n3890_), .Y(new_n4151_));
  AND2X1   g03959(.A(new_n4151_), .B(new_n4149_), .Y(new_n4152_));
  AOI21X1  g03960(.A0(new_n4152_), .A1(new_n4145_), .B0(\asqrt[63] ), .Y(new_n4153_));
  NOR2X1   g03961(.A(new_n4144_), .B(new_n4143_), .Y(new_n4154_));
  NAND2X1  g03962(.A(new_n4148_), .B(new_n4138_), .Y(new_n4155_));
  AOI21X1  g03963(.A0(new_n3876_), .A1(new_n3872_), .B0(new_n3835_), .Y(new_n4156_));
  AOI21X1  g03964(.A0(new_n3836_), .A1(new_n3830_), .B0(new_n193_), .Y(new_n4157_));
  OAI21X1  g03965(.A0(new_n4156_), .A1(new_n3830_), .B0(new_n4157_), .Y(new_n4158_));
  NOR4X1   g03966(.A(new_n3860_), .B(new_n3857_), .C(new_n3834_), .D(new_n3832_), .Y(new_n4159_));
  OAI21X1  g03967(.A0(new_n3854_), .A1(new_n3853_), .B0(new_n4159_), .Y(new_n4160_));
  NOR2X1   g03968(.A(new_n4160_), .B(new_n3841_), .Y(new_n4161_));
  INVX1    g03969(.A(new_n4161_), .Y(new_n4162_));
  AND2X1   g03970(.A(new_n4162_), .B(new_n4158_), .Y(new_n4163_));
  OAI21X1  g03971(.A0(new_n4155_), .A1(new_n4154_), .B0(new_n4163_), .Y(new_n4164_));
  NOR2X1   g03972(.A(new_n4164_), .B(new_n4153_), .Y(new_n4165_));
  OR2X1    g03973(.A(new_n4164_), .B(new_n4153_), .Y(\asqrt[39] ));
  NOR2X1   g03974(.A(\a[77] ), .B(\a[76] ), .Y(new_n4167_));
  MX2X1    g03975(.A(new_n4167_), .B(\asqrt[39] ), .S0(\a[78] ), .Y(new_n4168_));
  OAI21X1  g03976(.A0(new_n4164_), .A1(new_n4153_), .B0(\a[78] ), .Y(new_n4169_));
  NOR3X1   g03977(.A(\a[78] ), .B(\a[77] ), .C(\a[76] ), .Y(new_n4170_));
  OR2X1    g03978(.A(new_n4170_), .B(new_n3860_), .Y(new_n4171_));
  NOR4X1   g03979(.A(new_n4171_), .B(new_n3857_), .C(new_n3890_), .D(new_n3841_), .Y(new_n4172_));
  NAND2X1  g03980(.A(new_n4172_), .B(new_n4169_), .Y(new_n4173_));
  INVX1    g03981(.A(\a[78] ), .Y(new_n4174_));
  OAI21X1  g03982(.A0(new_n4164_), .A1(new_n4153_), .B0(new_n4174_), .Y(new_n4175_));
  AND2X1   g03983(.A(new_n4135_), .B(\asqrt[60] ), .Y(new_n4176_));
  OR2X1    g03984(.A(new_n4119_), .B(new_n4106_), .Y(new_n4177_));
  AND2X1   g03985(.A(new_n4126_), .B(new_n292_), .Y(new_n4178_));
  AOI21X1  g03986(.A0(new_n4178_), .A1(new_n4177_), .B0(new_n4124_), .Y(new_n4179_));
  OAI21X1  g03987(.A0(new_n4179_), .A1(new_n4176_), .B0(\asqrt[61] ), .Y(new_n4180_));
  INVX1    g03988(.A(new_n4134_), .Y(new_n4181_));
  OAI21X1  g03989(.A0(new_n4109_), .A1(new_n292_), .B0(new_n217_), .Y(new_n4182_));
  OAI21X1  g03990(.A0(new_n4182_), .A1(new_n4179_), .B0(new_n4181_), .Y(new_n4183_));
  AOI21X1  g03991(.A0(new_n4183_), .A1(new_n4180_), .B0(new_n199_), .Y(new_n4184_));
  INVX1    g03992(.A(new_n4143_), .Y(new_n4185_));
  NAND3X1  g03993(.A(new_n4183_), .B(new_n4180_), .C(new_n199_), .Y(new_n4186_));
  AOI21X1  g03994(.A0(new_n4186_), .A1(new_n4185_), .B0(new_n4184_), .Y(new_n4187_));
  INVX1    g03995(.A(new_n4152_), .Y(new_n4188_));
  OAI21X1  g03996(.A0(new_n4188_), .A1(new_n4187_), .B0(new_n193_), .Y(new_n4189_));
  OR2X1    g03997(.A(new_n4144_), .B(new_n4143_), .Y(new_n4190_));
  AND2X1   g03998(.A(new_n4148_), .B(new_n4138_), .Y(new_n4191_));
  INVX1    g03999(.A(new_n4163_), .Y(new_n4192_));
  AOI21X1  g04000(.A0(new_n4191_), .A1(new_n4190_), .B0(new_n4192_), .Y(new_n4193_));
  AOI21X1  g04001(.A0(new_n4193_), .A1(new_n4189_), .B0(new_n3886_), .Y(new_n4194_));
  AOI21X1  g04002(.A0(new_n4175_), .A1(\a[79] ), .B0(new_n4194_), .Y(new_n4195_));
  AOI22X1  g04003(.A0(new_n4195_), .A1(new_n4173_), .B0(new_n4168_), .B1(\asqrt[40] ), .Y(new_n4196_));
  OR2X1    g04004(.A(new_n4196_), .B(new_n3564_), .Y(new_n4197_));
  AND2X1   g04005(.A(new_n4195_), .B(new_n4173_), .Y(new_n4198_));
  AOI21X1  g04006(.A0(\asqrt[39] ), .A1(\a[78] ), .B0(new_n4170_), .Y(new_n4199_));
  OAI21X1  g04007(.A0(new_n4199_), .A1(new_n3863_), .B0(new_n3564_), .Y(new_n4200_));
  OAI21X1  g04008(.A0(new_n4164_), .A1(new_n4153_), .B0(new_n3866_), .Y(new_n4201_));
  INVX1    g04009(.A(new_n4158_), .Y(new_n4202_));
  NOR3X1   g04010(.A(new_n4161_), .B(new_n4202_), .C(new_n3863_), .Y(new_n4203_));
  OAI21X1  g04011(.A0(new_n4155_), .A1(new_n4154_), .B0(new_n4203_), .Y(new_n4204_));
  OR2X1    g04012(.A(new_n4204_), .B(new_n4153_), .Y(new_n4205_));
  AOI21X1  g04013(.A0(new_n4205_), .A1(new_n4201_), .B0(new_n3865_), .Y(new_n4206_));
  OAI21X1  g04014(.A0(new_n4204_), .A1(new_n4153_), .B0(new_n3865_), .Y(new_n4207_));
  NOR2X1   g04015(.A(new_n4207_), .B(new_n4194_), .Y(new_n4208_));
  OR2X1    g04016(.A(new_n4208_), .B(new_n4206_), .Y(new_n4209_));
  OAI21X1  g04017(.A0(new_n4200_), .A1(new_n4198_), .B0(new_n4209_), .Y(new_n4210_));
  AOI21X1  g04018(.A0(new_n4210_), .A1(new_n4197_), .B0(new_n3276_), .Y(new_n4211_));
  AOI21X1  g04019(.A0(new_n3868_), .A1(\asqrt[41] ), .B0(new_n3905_), .Y(new_n4212_));
  AND2X1   g04020(.A(new_n4212_), .B(new_n3908_), .Y(new_n4213_));
  OAI21X1  g04021(.A0(new_n4164_), .A1(new_n4153_), .B0(new_n4212_), .Y(new_n4214_));
  AOI22X1  g04022(.A0(new_n4214_), .A1(new_n3882_), .B0(new_n4213_), .B1(\asqrt[39] ), .Y(new_n4215_));
  AND2X1   g04023(.A(new_n4172_), .B(new_n4169_), .Y(new_n4216_));
  INVX1    g04024(.A(\a[79] ), .Y(new_n4217_));
  AOI21X1  g04025(.A0(new_n4193_), .A1(new_n4189_), .B0(\a[78] ), .Y(new_n4218_));
  OAI21X1  g04026(.A0(new_n4218_), .A1(new_n4217_), .B0(new_n4201_), .Y(new_n4219_));
  OAI22X1  g04027(.A0(new_n4219_), .A1(new_n4216_), .B0(new_n4199_), .B1(new_n3863_), .Y(new_n4220_));
  AOI21X1  g04028(.A0(new_n4220_), .A1(\asqrt[41] ), .B0(\asqrt[42] ), .Y(new_n4221_));
  AOI21X1  g04029(.A0(new_n4221_), .A1(new_n4210_), .B0(new_n4215_), .Y(new_n4222_));
  OAI21X1  g04030(.A0(new_n4222_), .A1(new_n4211_), .B0(\asqrt[43] ), .Y(new_n4223_));
  AOI21X1  g04031(.A0(new_n3931_), .A1(new_n3930_), .B0(new_n3896_), .Y(new_n4224_));
  AND2X1   g04032(.A(new_n4224_), .B(new_n3884_), .Y(new_n4225_));
  AOI22X1  g04033(.A0(new_n3931_), .A1(new_n3930_), .B0(new_n3909_), .B1(\asqrt[42] ), .Y(new_n4226_));
  OAI21X1  g04034(.A0(new_n4164_), .A1(new_n4153_), .B0(new_n4226_), .Y(new_n4227_));
  AOI22X1  g04035(.A0(new_n4227_), .A1(new_n3896_), .B0(new_n4225_), .B1(\asqrt[39] ), .Y(new_n4228_));
  NOR3X1   g04036(.A(new_n4222_), .B(new_n4211_), .C(\asqrt[43] ), .Y(new_n4229_));
  OAI21X1  g04037(.A0(new_n4229_), .A1(new_n4228_), .B0(new_n4223_), .Y(new_n4230_));
  AND2X1   g04038(.A(new_n4230_), .B(\asqrt[44] ), .Y(new_n4231_));
  OR2X1    g04039(.A(new_n4229_), .B(new_n4228_), .Y(new_n4232_));
  AND2X1   g04040(.A(new_n3910_), .B(new_n3897_), .Y(new_n4233_));
  NOR3X1   g04041(.A(new_n4233_), .B(new_n3935_), .C(new_n3898_), .Y(new_n4234_));
  NOR2X1   g04042(.A(new_n4233_), .B(new_n3898_), .Y(new_n4235_));
  OAI21X1  g04043(.A0(new_n4164_), .A1(new_n4153_), .B0(new_n4235_), .Y(new_n4236_));
  AOI22X1  g04044(.A0(new_n4236_), .A1(new_n3935_), .B0(new_n4234_), .B1(\asqrt[39] ), .Y(new_n4237_));
  AND2X1   g04045(.A(new_n4223_), .B(new_n2769_), .Y(new_n4238_));
  AOI21X1  g04046(.A0(new_n4238_), .A1(new_n4232_), .B0(new_n4237_), .Y(new_n4239_));
  OAI21X1  g04047(.A0(new_n4239_), .A1(new_n4231_), .B0(\asqrt[45] ), .Y(new_n4240_));
  NAND4X1  g04048(.A(\asqrt[39] ), .B(new_n3949_), .C(new_n3919_), .D(new_n3912_), .Y(new_n4241_));
  NOR3X1   g04049(.A(new_n4165_), .B(new_n3920_), .C(new_n3938_), .Y(new_n4242_));
  OAI21X1  g04050(.A0(new_n4242_), .A1(new_n3919_), .B0(new_n4241_), .Y(new_n4243_));
  AND2X1   g04051(.A(new_n4220_), .B(\asqrt[41] ), .Y(new_n4244_));
  NAND2X1  g04052(.A(new_n4195_), .B(new_n4173_), .Y(new_n4245_));
  AOI21X1  g04053(.A0(new_n4168_), .A1(\asqrt[40] ), .B0(\asqrt[41] ), .Y(new_n4246_));
  NOR2X1   g04054(.A(new_n4208_), .B(new_n4206_), .Y(new_n4247_));
  AOI21X1  g04055(.A0(new_n4246_), .A1(new_n4245_), .B0(new_n4247_), .Y(new_n4248_));
  OAI21X1  g04056(.A0(new_n4248_), .A1(new_n4244_), .B0(\asqrt[42] ), .Y(new_n4249_));
  INVX1    g04057(.A(new_n4215_), .Y(new_n4250_));
  OAI21X1  g04058(.A0(new_n4196_), .A1(new_n3564_), .B0(new_n3276_), .Y(new_n4251_));
  OAI21X1  g04059(.A0(new_n4251_), .A1(new_n4248_), .B0(new_n4250_), .Y(new_n4252_));
  AOI21X1  g04060(.A0(new_n4252_), .A1(new_n4249_), .B0(new_n3008_), .Y(new_n4253_));
  INVX1    g04061(.A(new_n4228_), .Y(new_n4254_));
  NAND3X1  g04062(.A(new_n4252_), .B(new_n4249_), .C(new_n3008_), .Y(new_n4255_));
  AOI21X1  g04063(.A0(new_n4255_), .A1(new_n4254_), .B0(new_n4253_), .Y(new_n4256_));
  OAI21X1  g04064(.A0(new_n4256_), .A1(new_n2769_), .B0(new_n2570_), .Y(new_n4257_));
  OAI21X1  g04065(.A0(new_n4257_), .A1(new_n4239_), .B0(new_n4243_), .Y(new_n4258_));
  AOI21X1  g04066(.A0(new_n4258_), .A1(new_n4240_), .B0(new_n2263_), .Y(new_n4259_));
  AND2X1   g04067(.A(new_n3939_), .B(new_n3923_), .Y(new_n4260_));
  NOR3X1   g04068(.A(new_n4260_), .B(new_n3979_), .C(new_n3922_), .Y(new_n4261_));
  AOI22X1  g04069(.A0(new_n3939_), .A1(new_n3923_), .B0(new_n3921_), .B1(\asqrt[45] ), .Y(new_n4262_));
  AOI21X1  g04070(.A0(new_n4262_), .A1(\asqrt[39] ), .B0(new_n3928_), .Y(new_n4263_));
  AOI21X1  g04071(.A0(new_n4261_), .A1(\asqrt[39] ), .B0(new_n4263_), .Y(new_n4264_));
  INVX1    g04072(.A(new_n4264_), .Y(new_n4265_));
  NAND3X1  g04073(.A(new_n4258_), .B(new_n4240_), .C(new_n2263_), .Y(new_n4266_));
  AOI21X1  g04074(.A0(new_n4266_), .A1(new_n4265_), .B0(new_n4259_), .Y(new_n4267_));
  OR2X1    g04075(.A(new_n4267_), .B(new_n2040_), .Y(new_n4268_));
  AND2X1   g04076(.A(new_n4266_), .B(new_n4265_), .Y(new_n4269_));
  AND2X1   g04077(.A(new_n3983_), .B(new_n3981_), .Y(new_n4270_));
  NOR3X1   g04078(.A(new_n4270_), .B(new_n3947_), .C(new_n3982_), .Y(new_n4271_));
  NOR2X1   g04079(.A(new_n4270_), .B(new_n3982_), .Y(new_n4272_));
  AOI21X1  g04080(.A0(new_n4272_), .A1(\asqrt[39] ), .B0(new_n3946_), .Y(new_n4273_));
  AOI21X1  g04081(.A0(new_n4271_), .A1(\asqrt[39] ), .B0(new_n4273_), .Y(new_n4274_));
  INVX1    g04082(.A(new_n4274_), .Y(new_n4275_));
  OR2X1    g04083(.A(new_n4256_), .B(new_n2769_), .Y(new_n4276_));
  NOR2X1   g04084(.A(new_n4229_), .B(new_n4228_), .Y(new_n4277_));
  INVX1    g04085(.A(new_n4237_), .Y(new_n4278_));
  NAND2X1  g04086(.A(new_n4223_), .B(new_n2769_), .Y(new_n4279_));
  OAI21X1  g04087(.A0(new_n4279_), .A1(new_n4277_), .B0(new_n4278_), .Y(new_n4280_));
  AOI21X1  g04088(.A0(new_n4280_), .A1(new_n4276_), .B0(new_n2570_), .Y(new_n4281_));
  INVX1    g04089(.A(new_n4243_), .Y(new_n4282_));
  AOI21X1  g04090(.A0(new_n4230_), .A1(\asqrt[44] ), .B0(\asqrt[45] ), .Y(new_n4283_));
  AOI21X1  g04091(.A0(new_n4283_), .A1(new_n4280_), .B0(new_n4282_), .Y(new_n4284_));
  OAI21X1  g04092(.A0(new_n4284_), .A1(new_n4281_), .B0(\asqrt[46] ), .Y(new_n4285_));
  NAND2X1  g04093(.A(new_n4285_), .B(new_n2040_), .Y(new_n4286_));
  OAI21X1  g04094(.A0(new_n4286_), .A1(new_n4269_), .B0(new_n4275_), .Y(new_n4287_));
  AOI21X1  g04095(.A0(new_n4287_), .A1(new_n4268_), .B0(new_n1834_), .Y(new_n4288_));
  NAND4X1  g04096(.A(\asqrt[39] ), .B(new_n3960_), .C(new_n3958_), .D(new_n3985_), .Y(new_n4289_));
  OR2X1    g04097(.A(new_n3986_), .B(new_n3953_), .Y(new_n4290_));
  OAI21X1  g04098(.A0(new_n4290_), .A1(new_n4165_), .B0(new_n3959_), .Y(new_n4291_));
  AND2X1   g04099(.A(new_n4291_), .B(new_n4289_), .Y(new_n4292_));
  NOR3X1   g04100(.A(new_n4284_), .B(new_n4281_), .C(\asqrt[46] ), .Y(new_n4293_));
  OAI21X1  g04101(.A0(new_n4293_), .A1(new_n4264_), .B0(new_n4285_), .Y(new_n4294_));
  AOI21X1  g04102(.A0(new_n4294_), .A1(\asqrt[47] ), .B0(\asqrt[48] ), .Y(new_n4295_));
  AOI21X1  g04103(.A0(new_n4295_), .A1(new_n4287_), .B0(new_n4292_), .Y(new_n4296_));
  OAI21X1  g04104(.A0(new_n4296_), .A1(new_n4288_), .B0(\asqrt[49] ), .Y(new_n4297_));
  AOI21X1  g04105(.A0(new_n4002_), .A1(new_n4001_), .B0(new_n3968_), .Y(new_n4298_));
  AND2X1   g04106(.A(new_n4298_), .B(new_n3962_), .Y(new_n4299_));
  AOI22X1  g04107(.A0(new_n4002_), .A1(new_n4001_), .B0(new_n3987_), .B1(\asqrt[48] ), .Y(new_n4300_));
  AOI21X1  g04108(.A0(new_n4300_), .A1(\asqrt[39] ), .B0(new_n3967_), .Y(new_n4301_));
  AOI21X1  g04109(.A0(new_n4299_), .A1(\asqrt[39] ), .B0(new_n4301_), .Y(new_n4302_));
  NOR3X1   g04110(.A(new_n4296_), .B(new_n4288_), .C(\asqrt[49] ), .Y(new_n4303_));
  OAI21X1  g04111(.A0(new_n4303_), .A1(new_n4302_), .B0(new_n4297_), .Y(new_n4304_));
  AND2X1   g04112(.A(new_n4304_), .B(\asqrt[50] ), .Y(new_n4305_));
  INVX1    g04113(.A(new_n4302_), .Y(new_n4306_));
  AND2X1   g04114(.A(new_n4294_), .B(\asqrt[47] ), .Y(new_n4307_));
  NAND2X1  g04115(.A(new_n4266_), .B(new_n4265_), .Y(new_n4308_));
  AND2X1   g04116(.A(new_n4285_), .B(new_n2040_), .Y(new_n4309_));
  AOI21X1  g04117(.A0(new_n4309_), .A1(new_n4308_), .B0(new_n4274_), .Y(new_n4310_));
  OAI21X1  g04118(.A0(new_n4310_), .A1(new_n4307_), .B0(\asqrt[48] ), .Y(new_n4311_));
  INVX1    g04119(.A(new_n4292_), .Y(new_n4312_));
  OAI21X1  g04120(.A0(new_n4267_), .A1(new_n2040_), .B0(new_n1834_), .Y(new_n4313_));
  OAI21X1  g04121(.A0(new_n4313_), .A1(new_n4310_), .B0(new_n4312_), .Y(new_n4314_));
  NAND3X1  g04122(.A(new_n4314_), .B(new_n4311_), .C(new_n1632_), .Y(new_n4315_));
  NAND2X1  g04123(.A(new_n4315_), .B(new_n4306_), .Y(new_n4316_));
  AND2X1   g04124(.A(new_n3988_), .B(new_n3970_), .Y(new_n4317_));
  NOR3X1   g04125(.A(new_n4317_), .B(new_n4005_), .C(new_n3971_), .Y(new_n4318_));
  NOR2X1   g04126(.A(new_n4317_), .B(new_n3971_), .Y(new_n4319_));
  AOI21X1  g04127(.A0(new_n4319_), .A1(\asqrt[39] ), .B0(new_n3976_), .Y(new_n4320_));
  AOI21X1  g04128(.A0(new_n4318_), .A1(\asqrt[39] ), .B0(new_n4320_), .Y(new_n4321_));
  AND2X1   g04129(.A(new_n4297_), .B(new_n1469_), .Y(new_n4322_));
  AOI21X1  g04130(.A0(new_n4322_), .A1(new_n4316_), .B0(new_n4321_), .Y(new_n4323_));
  OAI21X1  g04131(.A0(new_n4323_), .A1(new_n4305_), .B0(\asqrt[51] ), .Y(new_n4324_));
  NAND4X1  g04132(.A(\asqrt[39] ), .B(new_n4008_), .C(new_n3995_), .D(new_n3990_), .Y(new_n4325_));
  NAND2X1  g04133(.A(new_n4008_), .B(new_n3990_), .Y(new_n4326_));
  OAI21X1  g04134(.A0(new_n4326_), .A1(new_n4165_), .B0(new_n3999_), .Y(new_n4327_));
  AND2X1   g04135(.A(new_n4327_), .B(new_n4325_), .Y(new_n4328_));
  INVX1    g04136(.A(new_n4328_), .Y(new_n4329_));
  AOI21X1  g04137(.A0(new_n4314_), .A1(new_n4311_), .B0(new_n1632_), .Y(new_n4330_));
  AOI21X1  g04138(.A0(new_n4315_), .A1(new_n4306_), .B0(new_n4330_), .Y(new_n4331_));
  OAI21X1  g04139(.A0(new_n4331_), .A1(new_n1469_), .B0(new_n1277_), .Y(new_n4332_));
  OAI21X1  g04140(.A0(new_n4332_), .A1(new_n4323_), .B0(new_n4329_), .Y(new_n4333_));
  AOI21X1  g04141(.A0(new_n4333_), .A1(new_n4324_), .B0(new_n1111_), .Y(new_n4334_));
  AND2X1   g04142(.A(new_n4015_), .B(new_n4009_), .Y(new_n4335_));
  NOR3X1   g04143(.A(new_n4335_), .B(new_n4053_), .C(new_n3998_), .Y(new_n4336_));
  AOI22X1  g04144(.A0(new_n4015_), .A1(new_n4009_), .B0(new_n3997_), .B1(\asqrt[51] ), .Y(new_n4337_));
  AOI21X1  g04145(.A0(new_n4337_), .A1(\asqrt[39] ), .B0(new_n4013_), .Y(new_n4338_));
  AOI21X1  g04146(.A0(new_n4336_), .A1(\asqrt[39] ), .B0(new_n4338_), .Y(new_n4339_));
  INVX1    g04147(.A(new_n4339_), .Y(new_n4340_));
  NAND3X1  g04148(.A(new_n4333_), .B(new_n4324_), .C(new_n1111_), .Y(new_n4341_));
  AOI21X1  g04149(.A0(new_n4341_), .A1(new_n4340_), .B0(new_n4334_), .Y(new_n4342_));
  OR2X1    g04150(.A(new_n4342_), .B(new_n968_), .Y(new_n4343_));
  AND2X1   g04151(.A(new_n4341_), .B(new_n4340_), .Y(new_n4344_));
  AND2X1   g04152(.A(new_n4057_), .B(new_n4055_), .Y(new_n4345_));
  NOR3X1   g04153(.A(new_n4345_), .B(new_n4023_), .C(new_n4056_), .Y(new_n4346_));
  NOR2X1   g04154(.A(new_n4345_), .B(new_n4056_), .Y(new_n4347_));
  AOI21X1  g04155(.A0(new_n4347_), .A1(\asqrt[39] ), .B0(new_n4022_), .Y(new_n4348_));
  AOI21X1  g04156(.A0(new_n4346_), .A1(\asqrt[39] ), .B0(new_n4348_), .Y(new_n4349_));
  INVX1    g04157(.A(new_n4349_), .Y(new_n4350_));
  OR2X1    g04158(.A(new_n4331_), .B(new_n1469_), .Y(new_n4351_));
  AND2X1   g04159(.A(new_n4315_), .B(new_n4306_), .Y(new_n4352_));
  INVX1    g04160(.A(new_n4321_), .Y(new_n4353_));
  NAND2X1  g04161(.A(new_n4297_), .B(new_n1469_), .Y(new_n4354_));
  OAI21X1  g04162(.A0(new_n4354_), .A1(new_n4352_), .B0(new_n4353_), .Y(new_n4355_));
  AOI21X1  g04163(.A0(new_n4355_), .A1(new_n4351_), .B0(new_n1277_), .Y(new_n4356_));
  AOI21X1  g04164(.A0(new_n4304_), .A1(\asqrt[50] ), .B0(\asqrt[51] ), .Y(new_n4357_));
  AOI21X1  g04165(.A0(new_n4357_), .A1(new_n4355_), .B0(new_n4328_), .Y(new_n4358_));
  OAI21X1  g04166(.A0(new_n4358_), .A1(new_n4356_), .B0(\asqrt[52] ), .Y(new_n4359_));
  NAND2X1  g04167(.A(new_n4359_), .B(new_n968_), .Y(new_n4360_));
  OAI21X1  g04168(.A0(new_n4360_), .A1(new_n4344_), .B0(new_n4350_), .Y(new_n4361_));
  AOI21X1  g04169(.A0(new_n4361_), .A1(new_n4343_), .B0(new_n902_), .Y(new_n4362_));
  NAND4X1  g04170(.A(\asqrt[39] ), .B(new_n4034_), .C(new_n4032_), .D(new_n4059_), .Y(new_n4363_));
  NAND2X1  g04171(.A(new_n4034_), .B(new_n4059_), .Y(new_n4364_));
  OAI21X1  g04172(.A0(new_n4364_), .A1(new_n4165_), .B0(new_n4033_), .Y(new_n4365_));
  AND2X1   g04173(.A(new_n4365_), .B(new_n4363_), .Y(new_n4366_));
  NOR3X1   g04174(.A(new_n4358_), .B(new_n4356_), .C(\asqrt[52] ), .Y(new_n4367_));
  OAI21X1  g04175(.A0(new_n4367_), .A1(new_n4339_), .B0(new_n4359_), .Y(new_n4368_));
  AOI21X1  g04176(.A0(new_n4368_), .A1(\asqrt[53] ), .B0(\asqrt[54] ), .Y(new_n4369_));
  AOI21X1  g04177(.A0(new_n4369_), .A1(new_n4361_), .B0(new_n4366_), .Y(new_n4370_));
  OAI21X1  g04178(.A0(new_n4370_), .A1(new_n4362_), .B0(\asqrt[55] ), .Y(new_n4371_));
  AOI21X1  g04179(.A0(new_n4089_), .A1(new_n4088_), .B0(new_n4042_), .Y(new_n4372_));
  AND2X1   g04180(.A(new_n4372_), .B(new_n4036_), .Y(new_n4373_));
  AOI22X1  g04181(.A0(new_n4089_), .A1(new_n4088_), .B0(new_n4061_), .B1(\asqrt[54] ), .Y(new_n4374_));
  AOI21X1  g04182(.A0(new_n4374_), .A1(\asqrt[39] ), .B0(new_n4041_), .Y(new_n4375_));
  AOI21X1  g04183(.A0(new_n4373_), .A1(\asqrt[39] ), .B0(new_n4375_), .Y(new_n4376_));
  NOR3X1   g04184(.A(new_n4370_), .B(new_n4362_), .C(\asqrt[55] ), .Y(new_n4377_));
  OAI21X1  g04185(.A0(new_n4377_), .A1(new_n4376_), .B0(new_n4371_), .Y(new_n4378_));
  AND2X1   g04186(.A(new_n4378_), .B(\asqrt[56] ), .Y(new_n4379_));
  INVX1    g04187(.A(new_n4376_), .Y(new_n4380_));
  AND2X1   g04188(.A(new_n4368_), .B(\asqrt[53] ), .Y(new_n4381_));
  NAND2X1  g04189(.A(new_n4341_), .B(new_n4340_), .Y(new_n4382_));
  AND2X1   g04190(.A(new_n4359_), .B(new_n968_), .Y(new_n4383_));
  AOI21X1  g04191(.A0(new_n4383_), .A1(new_n4382_), .B0(new_n4349_), .Y(new_n4384_));
  OAI21X1  g04192(.A0(new_n4384_), .A1(new_n4381_), .B0(\asqrt[54] ), .Y(new_n4385_));
  INVX1    g04193(.A(new_n4366_), .Y(new_n4386_));
  OAI21X1  g04194(.A0(new_n4342_), .A1(new_n968_), .B0(new_n902_), .Y(new_n4387_));
  OAI21X1  g04195(.A0(new_n4387_), .A1(new_n4384_), .B0(new_n4386_), .Y(new_n4388_));
  NAND3X1  g04196(.A(new_n4388_), .B(new_n4385_), .C(new_n697_), .Y(new_n4389_));
  NAND2X1  g04197(.A(new_n4389_), .B(new_n4380_), .Y(new_n4390_));
  AND2X1   g04198(.A(new_n4062_), .B(new_n4044_), .Y(new_n4391_));
  NOR3X1   g04199(.A(new_n4391_), .B(new_n4092_), .C(new_n4045_), .Y(new_n4392_));
  NOR2X1   g04200(.A(new_n4391_), .B(new_n4045_), .Y(new_n4393_));
  AOI21X1  g04201(.A0(new_n4393_), .A1(\asqrt[39] ), .B0(new_n4050_), .Y(new_n4394_));
  AOI21X1  g04202(.A0(new_n4392_), .A1(\asqrt[39] ), .B0(new_n4394_), .Y(new_n4395_));
  AND2X1   g04203(.A(new_n4371_), .B(new_n582_), .Y(new_n4396_));
  AOI21X1  g04204(.A0(new_n4396_), .A1(new_n4390_), .B0(new_n4395_), .Y(new_n4397_));
  OAI21X1  g04205(.A0(new_n4397_), .A1(new_n4379_), .B0(\asqrt[57] ), .Y(new_n4398_));
  NAND4X1  g04206(.A(\asqrt[39] ), .B(new_n4097_), .C(new_n4069_), .D(new_n4064_), .Y(new_n4399_));
  OR2X1    g04207(.A(new_n4070_), .B(new_n4095_), .Y(new_n4400_));
  OAI21X1  g04208(.A0(new_n4400_), .A1(new_n4165_), .B0(new_n4096_), .Y(new_n4401_));
  AND2X1   g04209(.A(new_n4401_), .B(new_n4399_), .Y(new_n4402_));
  INVX1    g04210(.A(new_n4402_), .Y(new_n4403_));
  AOI21X1  g04211(.A0(new_n4388_), .A1(new_n4385_), .B0(new_n697_), .Y(new_n4404_));
  AOI21X1  g04212(.A0(new_n4389_), .A1(new_n4380_), .B0(new_n4404_), .Y(new_n4405_));
  OAI21X1  g04213(.A0(new_n4405_), .A1(new_n582_), .B0(new_n481_), .Y(new_n4406_));
  OAI21X1  g04214(.A0(new_n4406_), .A1(new_n4397_), .B0(new_n4403_), .Y(new_n4407_));
  AOI21X1  g04215(.A0(new_n4407_), .A1(new_n4398_), .B0(new_n399_), .Y(new_n4408_));
  NAND3X1  g04216(.A(new_n4407_), .B(new_n4398_), .C(new_n399_), .Y(new_n4409_));
  AND2X1   g04217(.A(new_n4074_), .B(new_n4073_), .Y(new_n4410_));
  NOR3X1   g04218(.A(new_n4114_), .B(new_n4410_), .C(new_n4072_), .Y(new_n4411_));
  AOI22X1  g04219(.A0(new_n4074_), .A1(new_n4073_), .B0(new_n4071_), .B1(\asqrt[57] ), .Y(new_n4412_));
  AOI21X1  g04220(.A0(new_n4412_), .A1(\asqrt[39] ), .B0(new_n4078_), .Y(new_n4413_));
  AOI21X1  g04221(.A0(new_n4411_), .A1(\asqrt[39] ), .B0(new_n4413_), .Y(new_n4414_));
  INVX1    g04222(.A(new_n4414_), .Y(new_n4415_));
  AOI21X1  g04223(.A0(new_n4415_), .A1(new_n4409_), .B0(new_n4408_), .Y(new_n4416_));
  OR2X1    g04224(.A(new_n4416_), .B(new_n328_), .Y(new_n4417_));
  AND2X1   g04225(.A(new_n4415_), .B(new_n4409_), .Y(new_n4418_));
  AND2X1   g04226(.A(new_n4117_), .B(new_n4115_), .Y(new_n4419_));
  NOR3X1   g04227(.A(new_n4419_), .B(new_n4086_), .C(new_n4116_), .Y(new_n4420_));
  NOR2X1   g04228(.A(new_n4419_), .B(new_n4116_), .Y(new_n4421_));
  AOI21X1  g04229(.A0(new_n4421_), .A1(\asqrt[39] ), .B0(new_n4085_), .Y(new_n4422_));
  AOI21X1  g04230(.A0(new_n4420_), .A1(\asqrt[39] ), .B0(new_n4422_), .Y(new_n4423_));
  INVX1    g04231(.A(new_n4423_), .Y(new_n4424_));
  OR2X1    g04232(.A(new_n4405_), .B(new_n582_), .Y(new_n4425_));
  AND2X1   g04233(.A(new_n4389_), .B(new_n4380_), .Y(new_n4426_));
  INVX1    g04234(.A(new_n4395_), .Y(new_n4427_));
  NAND2X1  g04235(.A(new_n4371_), .B(new_n582_), .Y(new_n4428_));
  OAI21X1  g04236(.A0(new_n4428_), .A1(new_n4426_), .B0(new_n4427_), .Y(new_n4429_));
  AOI21X1  g04237(.A0(new_n4429_), .A1(new_n4425_), .B0(new_n481_), .Y(new_n4430_));
  AOI21X1  g04238(.A0(new_n4378_), .A1(\asqrt[56] ), .B0(\asqrt[57] ), .Y(new_n4431_));
  AOI21X1  g04239(.A0(new_n4431_), .A1(new_n4429_), .B0(new_n4402_), .Y(new_n4432_));
  OAI21X1  g04240(.A0(new_n4432_), .A1(new_n4430_), .B0(\asqrt[58] ), .Y(new_n4433_));
  NAND2X1  g04241(.A(new_n4433_), .B(new_n328_), .Y(new_n4434_));
  OAI21X1  g04242(.A0(new_n4434_), .A1(new_n4418_), .B0(new_n4424_), .Y(new_n4435_));
  AOI21X1  g04243(.A0(new_n4435_), .A1(new_n4417_), .B0(new_n292_), .Y(new_n4436_));
  OR4X1    g04244(.A(new_n4165_), .B(new_n4119_), .C(new_n4107_), .D(new_n4101_), .Y(new_n4437_));
  OR2X1    g04245(.A(new_n4119_), .B(new_n4101_), .Y(new_n4438_));
  OAI21X1  g04246(.A0(new_n4438_), .A1(new_n4165_), .B0(new_n4107_), .Y(new_n4439_));
  AND2X1   g04247(.A(new_n4439_), .B(new_n4437_), .Y(new_n4440_));
  NOR3X1   g04248(.A(new_n4432_), .B(new_n4430_), .C(\asqrt[58] ), .Y(new_n4441_));
  OAI21X1  g04249(.A0(new_n4414_), .A1(new_n4441_), .B0(new_n4433_), .Y(new_n4442_));
  AOI21X1  g04250(.A0(new_n4442_), .A1(\asqrt[59] ), .B0(\asqrt[60] ), .Y(new_n4443_));
  AOI21X1  g04251(.A0(new_n4443_), .A1(new_n4435_), .B0(new_n4440_), .Y(new_n4444_));
  OAI21X1  g04252(.A0(new_n4444_), .A1(new_n4436_), .B0(\asqrt[61] ), .Y(new_n4445_));
  AOI21X1  g04253(.A0(new_n4178_), .A1(new_n4177_), .B0(new_n4125_), .Y(new_n4446_));
  AND2X1   g04254(.A(new_n4446_), .B(new_n4110_), .Y(new_n4447_));
  AOI22X1  g04255(.A0(new_n4178_), .A1(new_n4177_), .B0(new_n4135_), .B1(\asqrt[60] ), .Y(new_n4448_));
  AOI21X1  g04256(.A0(new_n4448_), .A1(\asqrt[39] ), .B0(new_n4124_), .Y(new_n4449_));
  AOI21X1  g04257(.A0(new_n4447_), .A1(\asqrt[39] ), .B0(new_n4449_), .Y(new_n4450_));
  NOR3X1   g04258(.A(new_n4444_), .B(new_n4436_), .C(\asqrt[61] ), .Y(new_n4451_));
  OAI21X1  g04259(.A0(new_n4451_), .A1(new_n4450_), .B0(new_n4445_), .Y(new_n4452_));
  AND2X1   g04260(.A(new_n4452_), .B(\asqrt[62] ), .Y(new_n4453_));
  OR2X1    g04261(.A(new_n4451_), .B(new_n4450_), .Y(new_n4454_));
  AND2X1   g04262(.A(new_n4136_), .B(new_n4128_), .Y(new_n4455_));
  NOR3X1   g04263(.A(new_n4455_), .B(new_n4181_), .C(new_n4129_), .Y(new_n4456_));
  NOR2X1   g04264(.A(new_n4455_), .B(new_n4129_), .Y(new_n4457_));
  AOI21X1  g04265(.A0(new_n4457_), .A1(\asqrt[39] ), .B0(new_n4134_), .Y(new_n4458_));
  AOI21X1  g04266(.A0(new_n4456_), .A1(\asqrt[39] ), .B0(new_n4458_), .Y(new_n4459_));
  AND2X1   g04267(.A(new_n4445_), .B(new_n199_), .Y(new_n4460_));
  AOI21X1  g04268(.A0(new_n4460_), .A1(new_n4454_), .B0(new_n4459_), .Y(new_n4461_));
  NAND3X1  g04269(.A(new_n4186_), .B(new_n4143_), .C(new_n4138_), .Y(new_n4462_));
  AOI21X1  g04270(.A0(new_n4193_), .A1(new_n4189_), .B0(new_n4462_), .Y(new_n4463_));
  NAND3X1  g04271(.A(\asqrt[39] ), .B(new_n4186_), .C(new_n4138_), .Y(new_n4464_));
  AOI21X1  g04272(.A0(new_n4464_), .A1(new_n4185_), .B0(new_n4463_), .Y(new_n4465_));
  INVX1    g04273(.A(new_n4465_), .Y(new_n4466_));
  AND2X1   g04274(.A(new_n4149_), .B(new_n4145_), .Y(new_n4467_));
  AOI22X1  g04275(.A0(new_n4467_), .A1(\asqrt[39] ), .B0(new_n4191_), .B1(new_n4190_), .Y(new_n4468_));
  AND2X1   g04276(.A(new_n4468_), .B(new_n4466_), .Y(new_n4469_));
  OAI21X1  g04277(.A0(new_n4461_), .A1(new_n4453_), .B0(new_n4469_), .Y(new_n4470_));
  AND2X1   g04278(.A(new_n4442_), .B(\asqrt[59] ), .Y(new_n4471_));
  NAND2X1  g04279(.A(new_n4415_), .B(new_n4409_), .Y(new_n4472_));
  AND2X1   g04280(.A(new_n4433_), .B(new_n328_), .Y(new_n4473_));
  AOI21X1  g04281(.A0(new_n4473_), .A1(new_n4472_), .B0(new_n4423_), .Y(new_n4474_));
  OAI21X1  g04282(.A0(new_n4474_), .A1(new_n4471_), .B0(\asqrt[60] ), .Y(new_n4475_));
  INVX1    g04283(.A(new_n4440_), .Y(new_n4476_));
  OAI21X1  g04284(.A0(new_n4416_), .A1(new_n328_), .B0(new_n292_), .Y(new_n4477_));
  OAI21X1  g04285(.A0(new_n4477_), .A1(new_n4474_), .B0(new_n4476_), .Y(new_n4478_));
  AOI21X1  g04286(.A0(new_n4478_), .A1(new_n4475_), .B0(new_n217_), .Y(new_n4479_));
  INVX1    g04287(.A(new_n4450_), .Y(new_n4480_));
  NAND3X1  g04288(.A(new_n4478_), .B(new_n4475_), .C(new_n217_), .Y(new_n4481_));
  AOI21X1  g04289(.A0(new_n4481_), .A1(new_n4480_), .B0(new_n4479_), .Y(new_n4482_));
  OAI21X1  g04290(.A0(new_n4482_), .A1(new_n199_), .B0(new_n4465_), .Y(new_n4483_));
  AOI21X1  g04291(.A0(new_n4193_), .A1(new_n4189_), .B0(new_n4148_), .Y(new_n4484_));
  AOI21X1  g04292(.A0(new_n4149_), .A1(new_n4145_), .B0(new_n193_), .Y(new_n4485_));
  OAI21X1  g04293(.A0(new_n4484_), .A1(new_n4145_), .B0(new_n4485_), .Y(new_n4486_));
  OR2X1    g04294(.A(new_n4155_), .B(new_n4154_), .Y(new_n4487_));
  AND2X1   g04295(.A(new_n4147_), .B(new_n3842_), .Y(new_n4488_));
  NOR4X1   g04296(.A(new_n4161_), .B(new_n4202_), .C(new_n4488_), .D(new_n4146_), .Y(new_n4489_));
  NAND3X1  g04297(.A(new_n4489_), .B(new_n4487_), .C(new_n4189_), .Y(new_n4490_));
  AND2X1   g04298(.A(new_n4490_), .B(new_n4486_), .Y(new_n4491_));
  OAI21X1  g04299(.A0(new_n4483_), .A1(new_n4461_), .B0(new_n4491_), .Y(new_n4492_));
  AOI21X1  g04300(.A0(new_n4470_), .A1(new_n193_), .B0(new_n4492_), .Y(new_n4493_));
  OR2X1    g04301(.A(new_n4482_), .B(new_n199_), .Y(new_n4494_));
  NOR2X1   g04302(.A(new_n4451_), .B(new_n4450_), .Y(new_n4495_));
  INVX1    g04303(.A(new_n4459_), .Y(new_n4496_));
  NAND2X1  g04304(.A(new_n4445_), .B(new_n199_), .Y(new_n4497_));
  OAI21X1  g04305(.A0(new_n4497_), .A1(new_n4495_), .B0(new_n4496_), .Y(new_n4498_));
  INVX1    g04306(.A(new_n4469_), .Y(new_n4499_));
  AOI21X1  g04307(.A0(new_n4498_), .A1(new_n4494_), .B0(new_n4499_), .Y(new_n4500_));
  AOI21X1  g04308(.A0(new_n4452_), .A1(\asqrt[62] ), .B0(new_n4466_), .Y(new_n4501_));
  INVX1    g04309(.A(new_n4491_), .Y(new_n4502_));
  AOI21X1  g04310(.A0(new_n4501_), .A1(new_n4498_), .B0(new_n4502_), .Y(new_n4503_));
  OAI21X1  g04311(.A0(new_n4500_), .A1(\asqrt[63] ), .B0(new_n4503_), .Y(\asqrt[38] ));
  NOR2X1   g04312(.A(\a[75] ), .B(\a[74] ), .Y(new_n4505_));
  MX2X1    g04313(.A(new_n4505_), .B(\asqrt[38] ), .S0(\a[76] ), .Y(new_n4506_));
  AND2X1   g04314(.A(new_n4506_), .B(\asqrt[39] ), .Y(new_n4507_));
  NOR3X1   g04315(.A(\a[76] ), .B(\a[75] ), .C(\a[74] ), .Y(new_n4508_));
  NOR3X1   g04316(.A(new_n4508_), .B(new_n4161_), .C(new_n4202_), .Y(new_n4509_));
  NAND3X1  g04317(.A(new_n4509_), .B(new_n4487_), .C(new_n4189_), .Y(new_n4510_));
  AOI21X1  g04318(.A0(\asqrt[38] ), .A1(\a[76] ), .B0(new_n4510_), .Y(new_n4511_));
  INVX1    g04319(.A(\a[76] ), .Y(new_n4512_));
  INVX1    g04320(.A(\a[77] ), .Y(new_n4513_));
  AOI21X1  g04321(.A0(\asqrt[38] ), .A1(new_n4512_), .B0(new_n4513_), .Y(new_n4514_));
  AND2X1   g04322(.A(\asqrt[38] ), .B(new_n4167_), .Y(new_n4515_));
  NOR3X1   g04323(.A(new_n4515_), .B(new_n4514_), .C(new_n4511_), .Y(new_n4516_));
  OAI21X1  g04324(.A0(new_n4516_), .A1(new_n4507_), .B0(\asqrt[40] ), .Y(new_n4517_));
  INVX1    g04325(.A(new_n4505_), .Y(new_n4518_));
  MX2X1    g04326(.A(new_n4518_), .B(new_n4493_), .S0(\a[76] ), .Y(new_n4519_));
  OAI21X1  g04327(.A0(new_n4519_), .A1(new_n4165_), .B0(new_n3863_), .Y(new_n4520_));
  NAND3X1  g04328(.A(new_n4490_), .B(new_n4486_), .C(\asqrt[39] ), .Y(new_n4521_));
  INVX1    g04329(.A(new_n4521_), .Y(new_n4522_));
  OAI21X1  g04330(.A0(new_n4483_), .A1(new_n4461_), .B0(new_n4522_), .Y(new_n4523_));
  AOI21X1  g04331(.A0(new_n4470_), .A1(new_n193_), .B0(new_n4523_), .Y(new_n4524_));
  AOI21X1  g04332(.A0(\asqrt[38] ), .A1(new_n4167_), .B0(new_n4524_), .Y(new_n4525_));
  OR2X1    g04333(.A(new_n4524_), .B(\a[78] ), .Y(new_n4526_));
  OAI22X1  g04334(.A0(new_n4526_), .A1(new_n4515_), .B0(new_n4525_), .B1(new_n4174_), .Y(new_n4527_));
  OAI21X1  g04335(.A0(new_n4520_), .A1(new_n4516_), .B0(new_n4527_), .Y(new_n4528_));
  AOI21X1  g04336(.A0(new_n4528_), .A1(new_n4517_), .B0(new_n3564_), .Y(new_n4529_));
  AOI21X1  g04337(.A0(new_n4168_), .A1(\asqrt[40] ), .B0(new_n4216_), .Y(new_n4530_));
  NAND3X1  g04338(.A(new_n4530_), .B(\asqrt[38] ), .C(new_n4219_), .Y(new_n4531_));
  INVX1    g04339(.A(new_n4530_), .Y(new_n4532_));
  OAI21X1  g04340(.A0(new_n4532_), .A1(new_n4493_), .B0(new_n4195_), .Y(new_n4533_));
  AND2X1   g04341(.A(new_n4533_), .B(new_n4531_), .Y(new_n4534_));
  INVX1    g04342(.A(new_n4534_), .Y(new_n4535_));
  NAND3X1  g04343(.A(new_n4528_), .B(new_n4517_), .C(new_n3564_), .Y(new_n4536_));
  AOI21X1  g04344(.A0(new_n4536_), .A1(new_n4535_), .B0(new_n4529_), .Y(new_n4537_));
  OR2X1    g04345(.A(new_n4537_), .B(new_n3276_), .Y(new_n4538_));
  AND2X1   g04346(.A(new_n4536_), .B(new_n4535_), .Y(new_n4539_));
  OAI21X1  g04347(.A0(new_n4200_), .A1(new_n4198_), .B0(new_n4247_), .Y(new_n4540_));
  OR2X1    g04348(.A(new_n4540_), .B(new_n4244_), .Y(new_n4541_));
  OR2X1    g04349(.A(new_n4541_), .B(new_n4493_), .Y(new_n4542_));
  OAI22X1  g04350(.A0(new_n4200_), .A1(new_n4198_), .B0(new_n4196_), .B1(new_n3564_), .Y(new_n4543_));
  OAI21X1  g04351(.A0(new_n4543_), .A1(new_n4493_), .B0(new_n4209_), .Y(new_n4544_));
  AND2X1   g04352(.A(new_n4544_), .B(new_n4542_), .Y(new_n4545_));
  INVX1    g04353(.A(new_n4545_), .Y(new_n4546_));
  OR2X1    g04354(.A(new_n4529_), .B(\asqrt[42] ), .Y(new_n4547_));
  OAI21X1  g04355(.A0(new_n4547_), .A1(new_n4539_), .B0(new_n4546_), .Y(new_n4548_));
  AOI21X1  g04356(.A0(new_n4548_), .A1(new_n4538_), .B0(new_n3008_), .Y(new_n4549_));
  AND2X1   g04357(.A(new_n4221_), .B(new_n4210_), .Y(new_n4550_));
  OR4X1    g04358(.A(new_n4493_), .B(new_n4550_), .C(new_n4250_), .D(new_n4211_), .Y(new_n4551_));
  OR2X1    g04359(.A(new_n4550_), .B(new_n4211_), .Y(new_n4552_));
  OAI21X1  g04360(.A0(new_n4552_), .A1(new_n4493_), .B0(new_n4250_), .Y(new_n4553_));
  AND2X1   g04361(.A(new_n4553_), .B(new_n4551_), .Y(new_n4554_));
  OR2X1    g04362(.A(new_n4519_), .B(new_n4165_), .Y(new_n4555_));
  INVX1    g04363(.A(new_n4510_), .Y(new_n4556_));
  OAI21X1  g04364(.A0(new_n4493_), .A1(new_n4512_), .B0(new_n4556_), .Y(new_n4557_));
  OAI21X1  g04365(.A0(new_n4493_), .A1(\a[76] ), .B0(\a[77] ), .Y(new_n4558_));
  INVX1    g04366(.A(new_n4167_), .Y(new_n4559_));
  OR2X1    g04367(.A(new_n4493_), .B(new_n4559_), .Y(new_n4560_));
  NAND3X1  g04368(.A(new_n4560_), .B(new_n4558_), .C(new_n4557_), .Y(new_n4561_));
  AOI21X1  g04369(.A0(new_n4561_), .A1(new_n4555_), .B0(new_n3863_), .Y(new_n4562_));
  AOI21X1  g04370(.A0(new_n4506_), .A1(\asqrt[39] ), .B0(\asqrt[40] ), .Y(new_n4563_));
  OR2X1    g04371(.A(new_n4525_), .B(new_n4174_), .Y(new_n4564_));
  OR2X1    g04372(.A(new_n4526_), .B(new_n4515_), .Y(new_n4565_));
  AOI22X1  g04373(.A0(new_n4565_), .A1(new_n4564_), .B0(new_n4563_), .B1(new_n4561_), .Y(new_n4566_));
  OAI21X1  g04374(.A0(new_n4566_), .A1(new_n4562_), .B0(\asqrt[41] ), .Y(new_n4567_));
  NOR3X1   g04375(.A(new_n4566_), .B(new_n4562_), .C(\asqrt[41] ), .Y(new_n4568_));
  OAI21X1  g04376(.A0(new_n4568_), .A1(new_n4534_), .B0(new_n4567_), .Y(new_n4569_));
  AOI21X1  g04377(.A0(new_n4569_), .A1(\asqrt[42] ), .B0(\asqrt[43] ), .Y(new_n4570_));
  AOI21X1  g04378(.A0(new_n4570_), .A1(new_n4548_), .B0(new_n4554_), .Y(new_n4571_));
  OAI21X1  g04379(.A0(new_n4571_), .A1(new_n4549_), .B0(\asqrt[44] ), .Y(new_n4572_));
  OR4X1    g04380(.A(new_n4493_), .B(new_n4229_), .C(new_n4254_), .D(new_n4253_), .Y(new_n4573_));
  NAND2X1  g04381(.A(new_n4255_), .B(new_n4223_), .Y(new_n4574_));
  OAI21X1  g04382(.A0(new_n4574_), .A1(new_n4493_), .B0(new_n4254_), .Y(new_n4575_));
  AND2X1   g04383(.A(new_n4575_), .B(new_n4573_), .Y(new_n4576_));
  NOR3X1   g04384(.A(new_n4571_), .B(new_n4549_), .C(\asqrt[44] ), .Y(new_n4577_));
  OAI21X1  g04385(.A0(new_n4577_), .A1(new_n4576_), .B0(new_n4572_), .Y(new_n4578_));
  AND2X1   g04386(.A(new_n4578_), .B(\asqrt[45] ), .Y(new_n4579_));
  INVX1    g04387(.A(new_n4576_), .Y(new_n4580_));
  AND2X1   g04388(.A(new_n4569_), .B(\asqrt[42] ), .Y(new_n4581_));
  NAND2X1  g04389(.A(new_n4536_), .B(new_n4535_), .Y(new_n4582_));
  NOR2X1   g04390(.A(new_n4529_), .B(\asqrt[42] ), .Y(new_n4583_));
  AOI21X1  g04391(.A0(new_n4583_), .A1(new_n4582_), .B0(new_n4545_), .Y(new_n4584_));
  OAI21X1  g04392(.A0(new_n4584_), .A1(new_n4581_), .B0(\asqrt[43] ), .Y(new_n4585_));
  INVX1    g04393(.A(new_n4554_), .Y(new_n4586_));
  OAI21X1  g04394(.A0(new_n4537_), .A1(new_n3276_), .B0(new_n3008_), .Y(new_n4587_));
  OAI21X1  g04395(.A0(new_n4587_), .A1(new_n4584_), .B0(new_n4586_), .Y(new_n4588_));
  NAND3X1  g04396(.A(new_n4588_), .B(new_n4585_), .C(new_n2769_), .Y(new_n4589_));
  NAND2X1  g04397(.A(new_n4589_), .B(new_n4580_), .Y(new_n4590_));
  AND2X1   g04398(.A(new_n4238_), .B(new_n4232_), .Y(new_n4591_));
  NOR4X1   g04399(.A(new_n4493_), .B(new_n4591_), .C(new_n4278_), .D(new_n4231_), .Y(new_n4592_));
  AOI22X1  g04400(.A0(new_n4238_), .A1(new_n4232_), .B0(new_n4230_), .B1(\asqrt[44] ), .Y(new_n4593_));
  AOI21X1  g04401(.A0(new_n4593_), .A1(\asqrt[38] ), .B0(new_n4237_), .Y(new_n4594_));
  NOR2X1   g04402(.A(new_n4594_), .B(new_n4592_), .Y(new_n4595_));
  AOI21X1  g04403(.A0(new_n4588_), .A1(new_n4585_), .B0(new_n2769_), .Y(new_n4596_));
  NOR2X1   g04404(.A(new_n4596_), .B(\asqrt[45] ), .Y(new_n4597_));
  AOI21X1  g04405(.A0(new_n4597_), .A1(new_n4590_), .B0(new_n4595_), .Y(new_n4598_));
  OAI21X1  g04406(.A0(new_n4598_), .A1(new_n4579_), .B0(\asqrt[46] ), .Y(new_n4599_));
  AND2X1   g04407(.A(new_n4283_), .B(new_n4280_), .Y(new_n4600_));
  OR4X1    g04408(.A(new_n4493_), .B(new_n4600_), .C(new_n4243_), .D(new_n4281_), .Y(new_n4601_));
  OR2X1    g04409(.A(new_n4600_), .B(new_n4281_), .Y(new_n4602_));
  OAI21X1  g04410(.A0(new_n4602_), .A1(new_n4493_), .B0(new_n4243_), .Y(new_n4603_));
  AND2X1   g04411(.A(new_n4603_), .B(new_n4601_), .Y(new_n4604_));
  INVX1    g04412(.A(new_n4604_), .Y(new_n4605_));
  AOI21X1  g04413(.A0(new_n4589_), .A1(new_n4580_), .B0(new_n4596_), .Y(new_n4606_));
  OAI21X1  g04414(.A0(new_n4606_), .A1(new_n2570_), .B0(new_n2263_), .Y(new_n4607_));
  OAI21X1  g04415(.A0(new_n4607_), .A1(new_n4598_), .B0(new_n4605_), .Y(new_n4608_));
  AOI21X1  g04416(.A0(new_n4608_), .A1(new_n4599_), .B0(new_n2040_), .Y(new_n4609_));
  NOR3X1   g04417(.A(new_n4293_), .B(new_n4265_), .C(new_n4259_), .Y(new_n4610_));
  AND2X1   g04418(.A(new_n4266_), .B(new_n4285_), .Y(new_n4611_));
  AOI21X1  g04419(.A0(new_n4611_), .A1(\asqrt[38] ), .B0(new_n4264_), .Y(new_n4612_));
  AOI21X1  g04420(.A0(new_n4610_), .A1(\asqrt[38] ), .B0(new_n4612_), .Y(new_n4613_));
  INVX1    g04421(.A(new_n4613_), .Y(new_n4614_));
  NAND3X1  g04422(.A(new_n4608_), .B(new_n4599_), .C(new_n2040_), .Y(new_n4615_));
  AOI21X1  g04423(.A0(new_n4615_), .A1(new_n4614_), .B0(new_n4609_), .Y(new_n4616_));
  OR2X1    g04424(.A(new_n4616_), .B(new_n1834_), .Y(new_n4617_));
  AND2X1   g04425(.A(new_n4615_), .B(new_n4614_), .Y(new_n4618_));
  OAI21X1  g04426(.A0(new_n4286_), .A1(new_n4269_), .B0(new_n4274_), .Y(new_n4619_));
  OR2X1    g04427(.A(new_n4619_), .B(new_n4307_), .Y(new_n4620_));
  AOI22X1  g04428(.A0(new_n4309_), .A1(new_n4308_), .B0(new_n4294_), .B1(\asqrt[47] ), .Y(new_n4621_));
  AND2X1   g04429(.A(new_n4621_), .B(\asqrt[38] ), .Y(new_n4622_));
  OAI22X1  g04430(.A0(new_n4622_), .A1(new_n4274_), .B0(new_n4620_), .B1(new_n4493_), .Y(new_n4623_));
  OR2X1    g04431(.A(new_n4609_), .B(\asqrt[48] ), .Y(new_n4624_));
  OAI21X1  g04432(.A0(new_n4624_), .A1(new_n4618_), .B0(new_n4623_), .Y(new_n4625_));
  AOI21X1  g04433(.A0(new_n4625_), .A1(new_n4617_), .B0(new_n1632_), .Y(new_n4626_));
  AND2X1   g04434(.A(new_n4295_), .B(new_n4287_), .Y(new_n4627_));
  OR4X1    g04435(.A(new_n4493_), .B(new_n4627_), .C(new_n4312_), .D(new_n4288_), .Y(new_n4628_));
  OR2X1    g04436(.A(new_n4627_), .B(new_n4288_), .Y(new_n4629_));
  OAI21X1  g04437(.A0(new_n4629_), .A1(new_n4493_), .B0(new_n4312_), .Y(new_n4630_));
  AND2X1   g04438(.A(new_n4630_), .B(new_n4628_), .Y(new_n4631_));
  OR2X1    g04439(.A(new_n4606_), .B(new_n2570_), .Y(new_n4632_));
  AND2X1   g04440(.A(new_n4589_), .B(new_n4580_), .Y(new_n4633_));
  INVX1    g04441(.A(new_n4595_), .Y(new_n4634_));
  OR2X1    g04442(.A(new_n4596_), .B(\asqrt[45] ), .Y(new_n4635_));
  OAI21X1  g04443(.A0(new_n4635_), .A1(new_n4633_), .B0(new_n4634_), .Y(new_n4636_));
  AOI21X1  g04444(.A0(new_n4636_), .A1(new_n4632_), .B0(new_n2263_), .Y(new_n4637_));
  AOI21X1  g04445(.A0(new_n4578_), .A1(\asqrt[45] ), .B0(\asqrt[46] ), .Y(new_n4638_));
  AOI21X1  g04446(.A0(new_n4638_), .A1(new_n4636_), .B0(new_n4604_), .Y(new_n4639_));
  OAI21X1  g04447(.A0(new_n4639_), .A1(new_n4637_), .B0(\asqrt[47] ), .Y(new_n4640_));
  NOR3X1   g04448(.A(new_n4639_), .B(new_n4637_), .C(\asqrt[47] ), .Y(new_n4641_));
  OAI21X1  g04449(.A0(new_n4641_), .A1(new_n4613_), .B0(new_n4640_), .Y(new_n4642_));
  AOI21X1  g04450(.A0(new_n4642_), .A1(\asqrt[48] ), .B0(\asqrt[49] ), .Y(new_n4643_));
  AOI21X1  g04451(.A0(new_n4643_), .A1(new_n4625_), .B0(new_n4631_), .Y(new_n4644_));
  OAI21X1  g04452(.A0(new_n4644_), .A1(new_n4626_), .B0(\asqrt[50] ), .Y(new_n4645_));
  OR4X1    g04453(.A(new_n4493_), .B(new_n4303_), .C(new_n4306_), .D(new_n4330_), .Y(new_n4646_));
  NAND2X1  g04454(.A(new_n4315_), .B(new_n4297_), .Y(new_n4647_));
  OAI21X1  g04455(.A0(new_n4647_), .A1(new_n4493_), .B0(new_n4306_), .Y(new_n4648_));
  AND2X1   g04456(.A(new_n4648_), .B(new_n4646_), .Y(new_n4649_));
  NOR3X1   g04457(.A(new_n4644_), .B(new_n4626_), .C(\asqrt[50] ), .Y(new_n4650_));
  OAI21X1  g04458(.A0(new_n4650_), .A1(new_n4649_), .B0(new_n4645_), .Y(new_n4651_));
  AND2X1   g04459(.A(new_n4651_), .B(\asqrt[51] ), .Y(new_n4652_));
  INVX1    g04460(.A(new_n4649_), .Y(new_n4653_));
  AND2X1   g04461(.A(new_n4642_), .B(\asqrt[48] ), .Y(new_n4654_));
  NAND2X1  g04462(.A(new_n4615_), .B(new_n4614_), .Y(new_n4655_));
  INVX1    g04463(.A(new_n4623_), .Y(new_n4656_));
  NOR2X1   g04464(.A(new_n4609_), .B(\asqrt[48] ), .Y(new_n4657_));
  AOI21X1  g04465(.A0(new_n4657_), .A1(new_n4655_), .B0(new_n4656_), .Y(new_n4658_));
  OAI21X1  g04466(.A0(new_n4658_), .A1(new_n4654_), .B0(\asqrt[49] ), .Y(new_n4659_));
  INVX1    g04467(.A(new_n4631_), .Y(new_n4660_));
  OAI21X1  g04468(.A0(new_n4616_), .A1(new_n1834_), .B0(new_n1632_), .Y(new_n4661_));
  OAI21X1  g04469(.A0(new_n4661_), .A1(new_n4658_), .B0(new_n4660_), .Y(new_n4662_));
  NAND3X1  g04470(.A(new_n4662_), .B(new_n4659_), .C(new_n1469_), .Y(new_n4663_));
  NAND2X1  g04471(.A(new_n4663_), .B(new_n4653_), .Y(new_n4664_));
  AND2X1   g04472(.A(new_n4322_), .B(new_n4316_), .Y(new_n4665_));
  NOR3X1   g04473(.A(new_n4665_), .B(new_n4353_), .C(new_n4305_), .Y(new_n4666_));
  AOI22X1  g04474(.A0(new_n4322_), .A1(new_n4316_), .B0(new_n4304_), .B1(\asqrt[50] ), .Y(new_n4667_));
  AOI21X1  g04475(.A0(new_n4667_), .A1(\asqrt[38] ), .B0(new_n4321_), .Y(new_n4668_));
  AOI21X1  g04476(.A0(new_n4666_), .A1(\asqrt[38] ), .B0(new_n4668_), .Y(new_n4669_));
  AOI21X1  g04477(.A0(new_n4662_), .A1(new_n4659_), .B0(new_n1469_), .Y(new_n4670_));
  NOR2X1   g04478(.A(new_n4670_), .B(\asqrt[51] ), .Y(new_n4671_));
  AOI21X1  g04479(.A0(new_n4671_), .A1(new_n4664_), .B0(new_n4669_), .Y(new_n4672_));
  OAI21X1  g04480(.A0(new_n4672_), .A1(new_n4652_), .B0(\asqrt[52] ), .Y(new_n4673_));
  AND2X1   g04481(.A(new_n4357_), .B(new_n4355_), .Y(new_n4674_));
  OR4X1    g04482(.A(new_n4493_), .B(new_n4674_), .C(new_n4329_), .D(new_n4356_), .Y(new_n4675_));
  OR2X1    g04483(.A(new_n4674_), .B(new_n4356_), .Y(new_n4676_));
  OAI21X1  g04484(.A0(new_n4676_), .A1(new_n4493_), .B0(new_n4329_), .Y(new_n4677_));
  AND2X1   g04485(.A(new_n4677_), .B(new_n4675_), .Y(new_n4678_));
  INVX1    g04486(.A(new_n4678_), .Y(new_n4679_));
  AOI21X1  g04487(.A0(new_n4663_), .A1(new_n4653_), .B0(new_n4670_), .Y(new_n4680_));
  OAI21X1  g04488(.A0(new_n4680_), .A1(new_n1277_), .B0(new_n1111_), .Y(new_n4681_));
  OAI21X1  g04489(.A0(new_n4681_), .A1(new_n4672_), .B0(new_n4679_), .Y(new_n4682_));
  AOI21X1  g04490(.A0(new_n4682_), .A1(new_n4673_), .B0(new_n968_), .Y(new_n4683_));
  OR4X1    g04491(.A(new_n4493_), .B(new_n4367_), .C(new_n4340_), .D(new_n4334_), .Y(new_n4684_));
  NAND2X1  g04492(.A(new_n4341_), .B(new_n4359_), .Y(new_n4685_));
  OAI21X1  g04493(.A0(new_n4685_), .A1(new_n4493_), .B0(new_n4340_), .Y(new_n4686_));
  AND2X1   g04494(.A(new_n4686_), .B(new_n4684_), .Y(new_n4687_));
  INVX1    g04495(.A(new_n4687_), .Y(new_n4688_));
  NAND3X1  g04496(.A(new_n4682_), .B(new_n4673_), .C(new_n968_), .Y(new_n4689_));
  AOI21X1  g04497(.A0(new_n4689_), .A1(new_n4688_), .B0(new_n4683_), .Y(new_n4690_));
  OR2X1    g04498(.A(new_n4690_), .B(new_n902_), .Y(new_n4691_));
  AND2X1   g04499(.A(new_n4689_), .B(new_n4688_), .Y(new_n4692_));
  AOI21X1  g04500(.A0(new_n4383_), .A1(new_n4382_), .B0(new_n4350_), .Y(new_n4693_));
  AND2X1   g04501(.A(new_n4693_), .B(new_n4343_), .Y(new_n4694_));
  AOI22X1  g04502(.A0(new_n4383_), .A1(new_n4382_), .B0(new_n4368_), .B1(\asqrt[53] ), .Y(new_n4695_));
  AOI21X1  g04503(.A0(new_n4695_), .A1(\asqrt[38] ), .B0(new_n4349_), .Y(new_n4696_));
  AOI21X1  g04504(.A0(new_n4694_), .A1(\asqrt[38] ), .B0(new_n4696_), .Y(new_n4697_));
  INVX1    g04505(.A(new_n4697_), .Y(new_n4698_));
  OR2X1    g04506(.A(new_n4683_), .B(\asqrt[54] ), .Y(new_n4699_));
  OAI21X1  g04507(.A0(new_n4699_), .A1(new_n4692_), .B0(new_n4698_), .Y(new_n4700_));
  AOI21X1  g04508(.A0(new_n4700_), .A1(new_n4691_), .B0(new_n697_), .Y(new_n4701_));
  AND2X1   g04509(.A(new_n4369_), .B(new_n4361_), .Y(new_n4702_));
  OR4X1    g04510(.A(new_n4493_), .B(new_n4702_), .C(new_n4386_), .D(new_n4362_), .Y(new_n4703_));
  OR2X1    g04511(.A(new_n4702_), .B(new_n4362_), .Y(new_n4704_));
  OAI21X1  g04512(.A0(new_n4704_), .A1(new_n4493_), .B0(new_n4386_), .Y(new_n4705_));
  AND2X1   g04513(.A(new_n4705_), .B(new_n4703_), .Y(new_n4706_));
  OR2X1    g04514(.A(new_n4680_), .B(new_n1277_), .Y(new_n4707_));
  AND2X1   g04515(.A(new_n4663_), .B(new_n4653_), .Y(new_n4708_));
  INVX1    g04516(.A(new_n4669_), .Y(new_n4709_));
  OR2X1    g04517(.A(new_n4670_), .B(\asqrt[51] ), .Y(new_n4710_));
  OAI21X1  g04518(.A0(new_n4710_), .A1(new_n4708_), .B0(new_n4709_), .Y(new_n4711_));
  AOI21X1  g04519(.A0(new_n4711_), .A1(new_n4707_), .B0(new_n1111_), .Y(new_n4712_));
  AOI21X1  g04520(.A0(new_n4651_), .A1(\asqrt[51] ), .B0(\asqrt[52] ), .Y(new_n4713_));
  AOI21X1  g04521(.A0(new_n4713_), .A1(new_n4711_), .B0(new_n4678_), .Y(new_n4714_));
  OAI21X1  g04522(.A0(new_n4714_), .A1(new_n4712_), .B0(\asqrt[53] ), .Y(new_n4715_));
  NOR3X1   g04523(.A(new_n4714_), .B(new_n4712_), .C(\asqrt[53] ), .Y(new_n4716_));
  OAI21X1  g04524(.A0(new_n4716_), .A1(new_n4687_), .B0(new_n4715_), .Y(new_n4717_));
  AOI21X1  g04525(.A0(new_n4717_), .A1(\asqrt[54] ), .B0(\asqrt[55] ), .Y(new_n4718_));
  AOI21X1  g04526(.A0(new_n4718_), .A1(new_n4700_), .B0(new_n4706_), .Y(new_n4719_));
  OAI21X1  g04527(.A0(new_n4719_), .A1(new_n4701_), .B0(\asqrt[56] ), .Y(new_n4720_));
  OR4X1    g04528(.A(new_n4493_), .B(new_n4377_), .C(new_n4380_), .D(new_n4404_), .Y(new_n4721_));
  NAND2X1  g04529(.A(new_n4389_), .B(new_n4371_), .Y(new_n4722_));
  OAI21X1  g04530(.A0(new_n4722_), .A1(new_n4493_), .B0(new_n4380_), .Y(new_n4723_));
  AND2X1   g04531(.A(new_n4723_), .B(new_n4721_), .Y(new_n4724_));
  NOR3X1   g04532(.A(new_n4719_), .B(new_n4701_), .C(\asqrt[56] ), .Y(new_n4725_));
  OAI21X1  g04533(.A0(new_n4725_), .A1(new_n4724_), .B0(new_n4720_), .Y(new_n4726_));
  AND2X1   g04534(.A(new_n4726_), .B(\asqrt[57] ), .Y(new_n4727_));
  OR2X1    g04535(.A(new_n4725_), .B(new_n4724_), .Y(new_n4728_));
  AND2X1   g04536(.A(new_n4396_), .B(new_n4390_), .Y(new_n4729_));
  NOR4X1   g04537(.A(new_n4493_), .B(new_n4729_), .C(new_n4427_), .D(new_n4379_), .Y(new_n4730_));
  AOI22X1  g04538(.A0(new_n4396_), .A1(new_n4390_), .B0(new_n4378_), .B1(\asqrt[56] ), .Y(new_n4731_));
  AOI21X1  g04539(.A0(new_n4731_), .A1(\asqrt[38] ), .B0(new_n4395_), .Y(new_n4732_));
  NOR2X1   g04540(.A(new_n4732_), .B(new_n4730_), .Y(new_n4733_));
  AND2X1   g04541(.A(new_n4720_), .B(new_n481_), .Y(new_n4734_));
  AOI21X1  g04542(.A0(new_n4734_), .A1(new_n4728_), .B0(new_n4733_), .Y(new_n4735_));
  OAI21X1  g04543(.A0(new_n4735_), .A1(new_n4727_), .B0(\asqrt[58] ), .Y(new_n4736_));
  AND2X1   g04544(.A(new_n4431_), .B(new_n4429_), .Y(new_n4737_));
  OR4X1    g04545(.A(new_n4493_), .B(new_n4737_), .C(new_n4403_), .D(new_n4430_), .Y(new_n4738_));
  OR2X1    g04546(.A(new_n4737_), .B(new_n4430_), .Y(new_n4739_));
  OAI21X1  g04547(.A0(new_n4739_), .A1(new_n4493_), .B0(new_n4403_), .Y(new_n4740_));
  AND2X1   g04548(.A(new_n4740_), .B(new_n4738_), .Y(new_n4741_));
  INVX1    g04549(.A(new_n4741_), .Y(new_n4742_));
  AND2X1   g04550(.A(new_n4717_), .B(\asqrt[54] ), .Y(new_n4743_));
  NAND2X1  g04551(.A(new_n4689_), .B(new_n4688_), .Y(new_n4744_));
  NOR2X1   g04552(.A(new_n4683_), .B(\asqrt[54] ), .Y(new_n4745_));
  AOI21X1  g04553(.A0(new_n4745_), .A1(new_n4744_), .B0(new_n4697_), .Y(new_n4746_));
  OAI21X1  g04554(.A0(new_n4746_), .A1(new_n4743_), .B0(\asqrt[55] ), .Y(new_n4747_));
  INVX1    g04555(.A(new_n4706_), .Y(new_n4748_));
  OAI21X1  g04556(.A0(new_n4690_), .A1(new_n902_), .B0(new_n697_), .Y(new_n4749_));
  OAI21X1  g04557(.A0(new_n4749_), .A1(new_n4746_), .B0(new_n4748_), .Y(new_n4750_));
  AOI21X1  g04558(.A0(new_n4750_), .A1(new_n4747_), .B0(new_n582_), .Y(new_n4751_));
  INVX1    g04559(.A(new_n4724_), .Y(new_n4752_));
  NAND3X1  g04560(.A(new_n4750_), .B(new_n4747_), .C(new_n582_), .Y(new_n4753_));
  AOI21X1  g04561(.A0(new_n4753_), .A1(new_n4752_), .B0(new_n4751_), .Y(new_n4754_));
  OAI21X1  g04562(.A0(new_n4754_), .A1(new_n481_), .B0(new_n399_), .Y(new_n4755_));
  OAI21X1  g04563(.A0(new_n4755_), .A1(new_n4735_), .B0(new_n4742_), .Y(new_n4756_));
  AOI21X1  g04564(.A0(new_n4756_), .A1(new_n4736_), .B0(new_n328_), .Y(new_n4757_));
  NAND3X1  g04565(.A(new_n4756_), .B(new_n4736_), .C(new_n328_), .Y(new_n4758_));
  OR4X1    g04566(.A(new_n4493_), .B(new_n4415_), .C(new_n4441_), .D(new_n4408_), .Y(new_n4759_));
  NAND2X1  g04567(.A(new_n4409_), .B(new_n4433_), .Y(new_n4760_));
  OAI21X1  g04568(.A0(new_n4760_), .A1(new_n4493_), .B0(new_n4415_), .Y(new_n4761_));
  AND2X1   g04569(.A(new_n4761_), .B(new_n4759_), .Y(new_n4762_));
  INVX1    g04570(.A(new_n4762_), .Y(new_n4763_));
  AOI21X1  g04571(.A0(new_n4763_), .A1(new_n4758_), .B0(new_n4757_), .Y(new_n4764_));
  OR2X1    g04572(.A(new_n4764_), .B(new_n292_), .Y(new_n4765_));
  OR2X1    g04573(.A(new_n4754_), .B(new_n481_), .Y(new_n4766_));
  NOR2X1   g04574(.A(new_n4725_), .B(new_n4724_), .Y(new_n4767_));
  INVX1    g04575(.A(new_n4733_), .Y(new_n4768_));
  NAND2X1  g04576(.A(new_n4720_), .B(new_n481_), .Y(new_n4769_));
  OAI21X1  g04577(.A0(new_n4769_), .A1(new_n4767_), .B0(new_n4768_), .Y(new_n4770_));
  AOI21X1  g04578(.A0(new_n4770_), .A1(new_n4766_), .B0(new_n399_), .Y(new_n4771_));
  AOI21X1  g04579(.A0(new_n4726_), .A1(\asqrt[57] ), .B0(\asqrt[58] ), .Y(new_n4772_));
  AOI21X1  g04580(.A0(new_n4772_), .A1(new_n4770_), .B0(new_n4741_), .Y(new_n4773_));
  NOR3X1   g04581(.A(new_n4773_), .B(new_n4771_), .C(\asqrt[59] ), .Y(new_n4774_));
  NOR2X1   g04582(.A(new_n4762_), .B(new_n4774_), .Y(new_n4775_));
  OAI21X1  g04583(.A0(new_n4434_), .A1(new_n4418_), .B0(new_n4423_), .Y(new_n4776_));
  NOR3X1   g04584(.A(new_n4776_), .B(new_n4493_), .C(new_n4471_), .Y(new_n4777_));
  AOI22X1  g04585(.A0(new_n4473_), .A1(new_n4472_), .B0(new_n4442_), .B1(\asqrt[59] ), .Y(new_n4778_));
  AOI21X1  g04586(.A0(new_n4778_), .A1(\asqrt[38] ), .B0(new_n4423_), .Y(new_n4779_));
  NOR2X1   g04587(.A(new_n4779_), .B(new_n4777_), .Y(new_n4780_));
  INVX1    g04588(.A(new_n4780_), .Y(new_n4781_));
  OAI21X1  g04589(.A0(new_n4773_), .A1(new_n4771_), .B0(\asqrt[59] ), .Y(new_n4782_));
  NAND2X1  g04590(.A(new_n4782_), .B(new_n292_), .Y(new_n4783_));
  OAI21X1  g04591(.A0(new_n4783_), .A1(new_n4775_), .B0(new_n4781_), .Y(new_n4784_));
  AOI21X1  g04592(.A0(new_n4784_), .A1(new_n4765_), .B0(new_n217_), .Y(new_n4785_));
  AND2X1   g04593(.A(new_n4443_), .B(new_n4435_), .Y(new_n4786_));
  OR4X1    g04594(.A(new_n4493_), .B(new_n4786_), .C(new_n4476_), .D(new_n4436_), .Y(new_n4787_));
  OR2X1    g04595(.A(new_n4786_), .B(new_n4436_), .Y(new_n4788_));
  OAI21X1  g04596(.A0(new_n4788_), .A1(new_n4493_), .B0(new_n4476_), .Y(new_n4789_));
  AND2X1   g04597(.A(new_n4789_), .B(new_n4787_), .Y(new_n4790_));
  OAI21X1  g04598(.A0(new_n4762_), .A1(new_n4774_), .B0(new_n4782_), .Y(new_n4791_));
  AOI21X1  g04599(.A0(new_n4791_), .A1(\asqrt[60] ), .B0(\asqrt[61] ), .Y(new_n4792_));
  AOI21X1  g04600(.A0(new_n4792_), .A1(new_n4784_), .B0(new_n4790_), .Y(new_n4793_));
  OAI21X1  g04601(.A0(new_n4793_), .A1(new_n4785_), .B0(\asqrt[62] ), .Y(new_n4794_));
  OR4X1    g04602(.A(new_n4493_), .B(new_n4451_), .C(new_n4480_), .D(new_n4479_), .Y(new_n4795_));
  OR2X1    g04603(.A(new_n4451_), .B(new_n4479_), .Y(new_n4796_));
  OAI21X1  g04604(.A0(new_n4796_), .A1(new_n4493_), .B0(new_n4480_), .Y(new_n4797_));
  AND2X1   g04605(.A(new_n4797_), .B(new_n4795_), .Y(new_n4798_));
  NOR3X1   g04606(.A(new_n4793_), .B(new_n4785_), .C(\asqrt[62] ), .Y(new_n4799_));
  OAI21X1  g04607(.A0(new_n4799_), .A1(new_n4798_), .B0(new_n4794_), .Y(new_n4800_));
  AND2X1   g04608(.A(new_n4460_), .B(new_n4454_), .Y(new_n4801_));
  NOR4X1   g04609(.A(new_n4493_), .B(new_n4801_), .C(new_n4496_), .D(new_n4453_), .Y(new_n4802_));
  INVX1    g04610(.A(new_n4802_), .Y(new_n4803_));
  OAI22X1  g04611(.A0(new_n4497_), .A1(new_n4495_), .B0(new_n4482_), .B1(new_n199_), .Y(new_n4804_));
  OAI21X1  g04612(.A0(new_n4804_), .A1(new_n4493_), .B0(new_n4496_), .Y(new_n4805_));
  AND2X1   g04613(.A(new_n4805_), .B(new_n4803_), .Y(new_n4806_));
  INVX1    g04614(.A(new_n4806_), .Y(new_n4807_));
  AND2X1   g04615(.A(new_n4501_), .B(new_n4498_), .Y(new_n4808_));
  AOI21X1  g04616(.A0(new_n4498_), .A1(new_n4494_), .B0(new_n4465_), .Y(new_n4809_));
  AOI21X1  g04617(.A0(new_n4809_), .A1(\asqrt[38] ), .B0(new_n4808_), .Y(new_n4810_));
  AND2X1   g04618(.A(new_n4810_), .B(new_n4807_), .Y(new_n4811_));
  AOI21X1  g04619(.A0(new_n4811_), .A1(new_n4800_), .B0(\asqrt[63] ), .Y(new_n4812_));
  NOR2X1   g04620(.A(new_n4799_), .B(new_n4798_), .Y(new_n4813_));
  NAND2X1  g04621(.A(new_n4806_), .B(new_n4794_), .Y(new_n4814_));
  NAND2X1  g04622(.A(new_n4498_), .B(new_n4494_), .Y(new_n4815_));
  AOI21X1  g04623(.A0(\asqrt[38] ), .A1(new_n4466_), .B0(new_n4815_), .Y(new_n4816_));
  NOR3X1   g04624(.A(new_n4816_), .B(new_n4809_), .C(new_n193_), .Y(new_n4817_));
  AND2X1   g04625(.A(new_n4470_), .B(new_n193_), .Y(new_n4818_));
  OAI21X1  g04626(.A0(new_n4462_), .A1(new_n4165_), .B0(new_n4490_), .Y(new_n4819_));
  AOI21X1  g04627(.A0(new_n4464_), .A1(new_n4185_), .B0(new_n4819_), .Y(new_n4820_));
  NAND2X1  g04628(.A(new_n4820_), .B(new_n4486_), .Y(new_n4821_));
  OR2X1    g04629(.A(new_n4821_), .B(new_n4808_), .Y(new_n4822_));
  NOR2X1   g04630(.A(new_n4822_), .B(new_n4818_), .Y(new_n4823_));
  NOR2X1   g04631(.A(new_n4823_), .B(new_n4817_), .Y(new_n4824_));
  OAI21X1  g04632(.A0(new_n4814_), .A1(new_n4813_), .B0(new_n4824_), .Y(new_n4825_));
  NOR2X1   g04633(.A(new_n4825_), .B(new_n4812_), .Y(new_n4826_));
  INVX1    g04634(.A(new_n4826_), .Y(\asqrt[37] ));
  NOR2X1   g04635(.A(\a[73] ), .B(\a[72] ), .Y(new_n4828_));
  INVX1    g04636(.A(new_n4828_), .Y(new_n4829_));
  MX2X1    g04637(.A(new_n4829_), .B(new_n4826_), .S0(\a[74] ), .Y(new_n4830_));
  INVX1    g04638(.A(\a[74] ), .Y(new_n4831_));
  AND2X1   g04639(.A(new_n4791_), .B(\asqrt[60] ), .Y(new_n4832_));
  OR2X1    g04640(.A(new_n4762_), .B(new_n4774_), .Y(new_n4833_));
  AND2X1   g04641(.A(new_n4782_), .B(new_n292_), .Y(new_n4834_));
  AOI21X1  g04642(.A0(new_n4834_), .A1(new_n4833_), .B0(new_n4780_), .Y(new_n4835_));
  OAI21X1  g04643(.A0(new_n4835_), .A1(new_n4832_), .B0(\asqrt[61] ), .Y(new_n4836_));
  INVX1    g04644(.A(new_n4790_), .Y(new_n4837_));
  OAI21X1  g04645(.A0(new_n4764_), .A1(new_n292_), .B0(new_n217_), .Y(new_n4838_));
  OAI21X1  g04646(.A0(new_n4838_), .A1(new_n4835_), .B0(new_n4837_), .Y(new_n4839_));
  AOI21X1  g04647(.A0(new_n4839_), .A1(new_n4836_), .B0(new_n199_), .Y(new_n4840_));
  INVX1    g04648(.A(new_n4798_), .Y(new_n4841_));
  NAND3X1  g04649(.A(new_n4839_), .B(new_n4836_), .C(new_n199_), .Y(new_n4842_));
  AOI21X1  g04650(.A0(new_n4842_), .A1(new_n4841_), .B0(new_n4840_), .Y(new_n4843_));
  INVX1    g04651(.A(new_n4811_), .Y(new_n4844_));
  OAI21X1  g04652(.A0(new_n4844_), .A1(new_n4843_), .B0(new_n193_), .Y(new_n4845_));
  OR2X1    g04653(.A(new_n4799_), .B(new_n4798_), .Y(new_n4846_));
  AND2X1   g04654(.A(new_n4806_), .B(new_n4794_), .Y(new_n4847_));
  INVX1    g04655(.A(new_n4824_), .Y(new_n4848_));
  AOI21X1  g04656(.A0(new_n4847_), .A1(new_n4846_), .B0(new_n4848_), .Y(new_n4849_));
  AOI21X1  g04657(.A0(new_n4849_), .A1(new_n4845_), .B0(new_n4831_), .Y(new_n4850_));
  NAND2X1  g04658(.A(new_n4828_), .B(new_n4831_), .Y(new_n4851_));
  NAND3X1  g04659(.A(new_n4851_), .B(new_n4490_), .C(new_n4486_), .Y(new_n4852_));
  NOR4X1   g04660(.A(new_n4852_), .B(new_n4850_), .C(new_n4808_), .D(new_n4818_), .Y(new_n4853_));
  INVX1    g04661(.A(\a[75] ), .Y(new_n4854_));
  AOI21X1  g04662(.A0(new_n4849_), .A1(new_n4845_), .B0(\a[74] ), .Y(new_n4855_));
  OAI21X1  g04663(.A0(new_n4825_), .A1(new_n4812_), .B0(new_n4505_), .Y(new_n4856_));
  OAI21X1  g04664(.A0(new_n4855_), .A1(new_n4854_), .B0(new_n4856_), .Y(new_n4857_));
  OAI22X1  g04665(.A0(new_n4857_), .A1(new_n4853_), .B0(new_n4830_), .B1(new_n4493_), .Y(new_n4858_));
  AND2X1   g04666(.A(new_n4858_), .B(\asqrt[39] ), .Y(new_n4859_));
  OR4X1    g04667(.A(new_n4852_), .B(new_n4850_), .C(new_n4808_), .D(new_n4818_), .Y(new_n4860_));
  OAI21X1  g04668(.A0(new_n4825_), .A1(new_n4812_), .B0(new_n4831_), .Y(new_n4861_));
  AOI21X1  g04669(.A0(new_n4849_), .A1(new_n4845_), .B0(new_n4518_), .Y(new_n4862_));
  AOI21X1  g04670(.A0(new_n4861_), .A1(\a[75] ), .B0(new_n4862_), .Y(new_n4863_));
  NAND2X1  g04671(.A(new_n4863_), .B(new_n4860_), .Y(new_n4864_));
  OAI21X1  g04672(.A0(new_n4826_), .A1(new_n4831_), .B0(new_n4851_), .Y(new_n4865_));
  AOI21X1  g04673(.A0(new_n4865_), .A1(\asqrt[38] ), .B0(\asqrt[39] ), .Y(new_n4866_));
  AND2X1   g04674(.A(new_n4847_), .B(new_n4846_), .Y(new_n4867_));
  OAI21X1  g04675(.A0(new_n4822_), .A1(new_n4818_), .B0(\asqrt[38] ), .Y(new_n4868_));
  OR4X1    g04676(.A(new_n4868_), .B(new_n4817_), .C(new_n4867_), .D(new_n4812_), .Y(new_n4869_));
  AOI21X1  g04677(.A0(new_n4869_), .A1(new_n4856_), .B0(new_n4512_), .Y(new_n4870_));
  NOR4X1   g04678(.A(new_n4868_), .B(new_n4817_), .C(new_n4867_), .D(new_n4812_), .Y(new_n4871_));
  NOR3X1   g04679(.A(new_n4871_), .B(new_n4862_), .C(\a[76] ), .Y(new_n4872_));
  NOR2X1   g04680(.A(new_n4872_), .B(new_n4870_), .Y(new_n4873_));
  AOI21X1  g04681(.A0(new_n4866_), .A1(new_n4864_), .B0(new_n4873_), .Y(new_n4874_));
  OAI21X1  g04682(.A0(new_n4874_), .A1(new_n4859_), .B0(\asqrt[40] ), .Y(new_n4875_));
  AND2X1   g04683(.A(new_n4560_), .B(new_n4558_), .Y(new_n4876_));
  NOR3X1   g04684(.A(new_n4876_), .B(new_n4511_), .C(new_n4507_), .Y(new_n4877_));
  OAI21X1  g04685(.A0(new_n4825_), .A1(new_n4812_), .B0(new_n4877_), .Y(new_n4878_));
  AOI21X1  g04686(.A0(new_n4506_), .A1(\asqrt[39] ), .B0(new_n4511_), .Y(new_n4879_));
  OAI21X1  g04687(.A0(new_n4825_), .A1(new_n4812_), .B0(new_n4879_), .Y(new_n4880_));
  NAND2X1  g04688(.A(new_n4880_), .B(new_n4876_), .Y(new_n4881_));
  NAND2X1  g04689(.A(new_n4881_), .B(new_n4878_), .Y(new_n4882_));
  AOI22X1  g04690(.A0(new_n4863_), .A1(new_n4860_), .B0(new_n4865_), .B1(\asqrt[38] ), .Y(new_n4883_));
  OAI21X1  g04691(.A0(new_n4883_), .A1(new_n4165_), .B0(new_n3863_), .Y(new_n4884_));
  OAI21X1  g04692(.A0(new_n4884_), .A1(new_n4874_), .B0(new_n4882_), .Y(new_n4885_));
  AOI21X1  g04693(.A0(new_n4885_), .A1(new_n4875_), .B0(new_n3564_), .Y(new_n4886_));
  AND2X1   g04694(.A(new_n4563_), .B(new_n4561_), .Y(new_n4887_));
  NOR3X1   g04695(.A(new_n4527_), .B(new_n4887_), .C(new_n4562_), .Y(new_n4888_));
  OAI21X1  g04696(.A0(new_n4825_), .A1(new_n4812_), .B0(new_n4888_), .Y(new_n4889_));
  NOR2X1   g04697(.A(new_n4887_), .B(new_n4562_), .Y(new_n4890_));
  OAI21X1  g04698(.A0(new_n4825_), .A1(new_n4812_), .B0(new_n4890_), .Y(new_n4891_));
  NAND2X1  g04699(.A(new_n4891_), .B(new_n4527_), .Y(new_n4892_));
  AND2X1   g04700(.A(new_n4892_), .B(new_n4889_), .Y(new_n4893_));
  INVX1    g04701(.A(new_n4893_), .Y(new_n4894_));
  NAND3X1  g04702(.A(new_n4885_), .B(new_n4875_), .C(new_n3564_), .Y(new_n4895_));
  AOI21X1  g04703(.A0(new_n4895_), .A1(new_n4894_), .B0(new_n4886_), .Y(new_n4896_));
  OR2X1    g04704(.A(new_n4896_), .B(new_n3276_), .Y(new_n4897_));
  OR2X1    g04705(.A(new_n4883_), .B(new_n4165_), .Y(new_n4898_));
  AND2X1   g04706(.A(new_n4863_), .B(new_n4860_), .Y(new_n4899_));
  OAI21X1  g04707(.A0(new_n4830_), .A1(new_n4493_), .B0(new_n4165_), .Y(new_n4900_));
  OR2X1    g04708(.A(new_n4872_), .B(new_n4870_), .Y(new_n4901_));
  OAI21X1  g04709(.A0(new_n4900_), .A1(new_n4899_), .B0(new_n4901_), .Y(new_n4902_));
  AOI21X1  g04710(.A0(new_n4902_), .A1(new_n4898_), .B0(new_n3863_), .Y(new_n4903_));
  AOI21X1  g04711(.A0(new_n4858_), .A1(\asqrt[39] ), .B0(\asqrt[40] ), .Y(new_n4904_));
  AOI22X1  g04712(.A0(new_n4904_), .A1(new_n4902_), .B0(new_n4881_), .B1(new_n4878_), .Y(new_n4905_));
  NOR3X1   g04713(.A(new_n4905_), .B(new_n4903_), .C(\asqrt[41] ), .Y(new_n4906_));
  NOR2X1   g04714(.A(new_n4906_), .B(new_n4893_), .Y(new_n4907_));
  NOR3X1   g04715(.A(new_n4568_), .B(new_n4535_), .C(new_n4529_), .Y(new_n4908_));
  OAI21X1  g04716(.A0(new_n4825_), .A1(new_n4812_), .B0(new_n4908_), .Y(new_n4909_));
  NOR3X1   g04717(.A(new_n4826_), .B(new_n4568_), .C(new_n4529_), .Y(new_n4910_));
  OR2X1    g04718(.A(new_n4910_), .B(new_n4534_), .Y(new_n4911_));
  AND2X1   g04719(.A(new_n4911_), .B(new_n4909_), .Y(new_n4912_));
  INVX1    g04720(.A(new_n4912_), .Y(new_n4913_));
  OR2X1    g04721(.A(new_n4886_), .B(\asqrt[42] ), .Y(new_n4914_));
  OAI21X1  g04722(.A0(new_n4914_), .A1(new_n4907_), .B0(new_n4913_), .Y(new_n4915_));
  AOI21X1  g04723(.A0(new_n4915_), .A1(new_n4897_), .B0(new_n3008_), .Y(new_n4916_));
  AOI21X1  g04724(.A0(new_n4583_), .A1(new_n4582_), .B0(new_n4546_), .Y(new_n4917_));
  AND2X1   g04725(.A(new_n4917_), .B(new_n4538_), .Y(new_n4918_));
  AOI22X1  g04726(.A0(new_n4583_), .A1(new_n4582_), .B0(new_n4569_), .B1(\asqrt[42] ), .Y(new_n4919_));
  AOI21X1  g04727(.A0(new_n4919_), .A1(\asqrt[37] ), .B0(new_n4545_), .Y(new_n4920_));
  AOI21X1  g04728(.A0(new_n4918_), .A1(\asqrt[37] ), .B0(new_n4920_), .Y(new_n4921_));
  OAI21X1  g04729(.A0(new_n4905_), .A1(new_n4903_), .B0(\asqrt[41] ), .Y(new_n4922_));
  OAI21X1  g04730(.A0(new_n4906_), .A1(new_n4893_), .B0(new_n4922_), .Y(new_n4923_));
  AOI21X1  g04731(.A0(new_n4923_), .A1(\asqrt[42] ), .B0(\asqrt[43] ), .Y(new_n4924_));
  AOI21X1  g04732(.A0(new_n4924_), .A1(new_n4915_), .B0(new_n4921_), .Y(new_n4925_));
  OAI21X1  g04733(.A0(new_n4925_), .A1(new_n4916_), .B0(\asqrt[44] ), .Y(new_n4926_));
  AND2X1   g04734(.A(new_n4570_), .B(new_n4548_), .Y(new_n4927_));
  NOR3X1   g04735(.A(new_n4927_), .B(new_n4586_), .C(new_n4549_), .Y(new_n4928_));
  NOR3X1   g04736(.A(new_n4826_), .B(new_n4927_), .C(new_n4549_), .Y(new_n4929_));
  NOR2X1   g04737(.A(new_n4929_), .B(new_n4554_), .Y(new_n4930_));
  AOI21X1  g04738(.A0(new_n4928_), .A1(\asqrt[37] ), .B0(new_n4930_), .Y(new_n4931_));
  NOR3X1   g04739(.A(new_n4925_), .B(new_n4916_), .C(\asqrt[44] ), .Y(new_n4932_));
  OAI21X1  g04740(.A0(new_n4932_), .A1(new_n4931_), .B0(new_n4926_), .Y(new_n4933_));
  AND2X1   g04741(.A(new_n4933_), .B(\asqrt[45] ), .Y(new_n4934_));
  OR2X1    g04742(.A(new_n4932_), .B(new_n4931_), .Y(new_n4935_));
  NAND4X1  g04743(.A(\asqrt[37] ), .B(new_n4589_), .C(new_n4576_), .D(new_n4572_), .Y(new_n4936_));
  NAND2X1  g04744(.A(new_n4589_), .B(new_n4572_), .Y(new_n4937_));
  OAI21X1  g04745(.A0(new_n4937_), .A1(new_n4826_), .B0(new_n4580_), .Y(new_n4938_));
  AND2X1   g04746(.A(new_n4938_), .B(new_n4936_), .Y(new_n4939_));
  AND2X1   g04747(.A(new_n4926_), .B(new_n2570_), .Y(new_n4940_));
  AOI21X1  g04748(.A0(new_n4940_), .A1(new_n4935_), .B0(new_n4939_), .Y(new_n4941_));
  OAI21X1  g04749(.A0(new_n4941_), .A1(new_n4934_), .B0(\asqrt[46] ), .Y(new_n4942_));
  AND2X1   g04750(.A(new_n4597_), .B(new_n4590_), .Y(new_n4943_));
  NOR3X1   g04751(.A(new_n4943_), .B(new_n4634_), .C(new_n4579_), .Y(new_n4944_));
  NOR3X1   g04752(.A(new_n4826_), .B(new_n4943_), .C(new_n4579_), .Y(new_n4945_));
  NOR2X1   g04753(.A(new_n4945_), .B(new_n4595_), .Y(new_n4946_));
  AOI21X1  g04754(.A0(new_n4944_), .A1(\asqrt[37] ), .B0(new_n4946_), .Y(new_n4947_));
  INVX1    g04755(.A(new_n4947_), .Y(new_n4948_));
  AND2X1   g04756(.A(new_n4923_), .B(\asqrt[42] ), .Y(new_n4949_));
  OR2X1    g04757(.A(new_n4906_), .B(new_n4893_), .Y(new_n4950_));
  NOR2X1   g04758(.A(new_n4886_), .B(\asqrt[42] ), .Y(new_n4951_));
  AOI21X1  g04759(.A0(new_n4951_), .A1(new_n4950_), .B0(new_n4912_), .Y(new_n4952_));
  OAI21X1  g04760(.A0(new_n4952_), .A1(new_n4949_), .B0(\asqrt[43] ), .Y(new_n4953_));
  INVX1    g04761(.A(new_n4921_), .Y(new_n4954_));
  OAI21X1  g04762(.A0(new_n4896_), .A1(new_n3276_), .B0(new_n3008_), .Y(new_n4955_));
  OAI21X1  g04763(.A0(new_n4955_), .A1(new_n4952_), .B0(new_n4954_), .Y(new_n4956_));
  AOI21X1  g04764(.A0(new_n4956_), .A1(new_n4953_), .B0(new_n2769_), .Y(new_n4957_));
  INVX1    g04765(.A(new_n4931_), .Y(new_n4958_));
  NAND3X1  g04766(.A(new_n4956_), .B(new_n4953_), .C(new_n2769_), .Y(new_n4959_));
  AOI21X1  g04767(.A0(new_n4959_), .A1(new_n4958_), .B0(new_n4957_), .Y(new_n4960_));
  OAI21X1  g04768(.A0(new_n4960_), .A1(new_n2570_), .B0(new_n2263_), .Y(new_n4961_));
  OAI21X1  g04769(.A0(new_n4961_), .A1(new_n4941_), .B0(new_n4948_), .Y(new_n4962_));
  AOI21X1  g04770(.A0(new_n4962_), .A1(new_n4942_), .B0(new_n2040_), .Y(new_n4963_));
  AND2X1   g04771(.A(new_n4638_), .B(new_n4636_), .Y(new_n4964_));
  NOR3X1   g04772(.A(new_n4964_), .B(new_n4605_), .C(new_n4637_), .Y(new_n4965_));
  NOR3X1   g04773(.A(new_n4826_), .B(new_n4964_), .C(new_n4637_), .Y(new_n4966_));
  NOR2X1   g04774(.A(new_n4966_), .B(new_n4604_), .Y(new_n4967_));
  AOI21X1  g04775(.A0(new_n4965_), .A1(\asqrt[37] ), .B0(new_n4967_), .Y(new_n4968_));
  INVX1    g04776(.A(new_n4968_), .Y(new_n4969_));
  NAND3X1  g04777(.A(new_n4962_), .B(new_n4942_), .C(new_n2040_), .Y(new_n4970_));
  AOI21X1  g04778(.A0(new_n4970_), .A1(new_n4969_), .B0(new_n4963_), .Y(new_n4971_));
  OR2X1    g04779(.A(new_n4971_), .B(new_n1834_), .Y(new_n4972_));
  AND2X1   g04780(.A(new_n4970_), .B(new_n4969_), .Y(new_n4973_));
  OR4X1    g04781(.A(new_n4826_), .B(new_n4641_), .C(new_n4614_), .D(new_n4609_), .Y(new_n4974_));
  NAND2X1  g04782(.A(new_n4615_), .B(new_n4640_), .Y(new_n4975_));
  OAI21X1  g04783(.A0(new_n4975_), .A1(new_n4826_), .B0(new_n4614_), .Y(new_n4976_));
  AND2X1   g04784(.A(new_n4976_), .B(new_n4974_), .Y(new_n4977_));
  INVX1    g04785(.A(new_n4977_), .Y(new_n4978_));
  OR2X1    g04786(.A(new_n4963_), .B(\asqrt[48] ), .Y(new_n4979_));
  OAI21X1  g04787(.A0(new_n4979_), .A1(new_n4973_), .B0(new_n4978_), .Y(new_n4980_));
  AOI21X1  g04788(.A0(new_n4980_), .A1(new_n4972_), .B0(new_n1632_), .Y(new_n4981_));
  AOI21X1  g04789(.A0(new_n4657_), .A1(new_n4655_), .B0(new_n4623_), .Y(new_n4982_));
  AND2X1   g04790(.A(new_n4982_), .B(new_n4617_), .Y(new_n4983_));
  AOI22X1  g04791(.A0(new_n4657_), .A1(new_n4655_), .B0(new_n4642_), .B1(\asqrt[48] ), .Y(new_n4984_));
  AOI21X1  g04792(.A0(new_n4984_), .A1(\asqrt[37] ), .B0(new_n4656_), .Y(new_n4985_));
  AOI21X1  g04793(.A0(new_n4983_), .A1(\asqrt[37] ), .B0(new_n4985_), .Y(new_n4986_));
  OR2X1    g04794(.A(new_n4960_), .B(new_n2570_), .Y(new_n4987_));
  NOR2X1   g04795(.A(new_n4932_), .B(new_n4931_), .Y(new_n4988_));
  INVX1    g04796(.A(new_n4939_), .Y(new_n4989_));
  NAND2X1  g04797(.A(new_n4926_), .B(new_n2570_), .Y(new_n4990_));
  OAI21X1  g04798(.A0(new_n4990_), .A1(new_n4988_), .B0(new_n4989_), .Y(new_n4991_));
  AOI21X1  g04799(.A0(new_n4991_), .A1(new_n4987_), .B0(new_n2263_), .Y(new_n4992_));
  AOI21X1  g04800(.A0(new_n4933_), .A1(\asqrt[45] ), .B0(\asqrt[46] ), .Y(new_n4993_));
  AOI21X1  g04801(.A0(new_n4993_), .A1(new_n4991_), .B0(new_n4947_), .Y(new_n4994_));
  OAI21X1  g04802(.A0(new_n4994_), .A1(new_n4992_), .B0(\asqrt[47] ), .Y(new_n4995_));
  NOR3X1   g04803(.A(new_n4994_), .B(new_n4992_), .C(\asqrt[47] ), .Y(new_n4996_));
  OAI21X1  g04804(.A0(new_n4996_), .A1(new_n4968_), .B0(new_n4995_), .Y(new_n4997_));
  AOI21X1  g04805(.A0(new_n4997_), .A1(\asqrt[48] ), .B0(\asqrt[49] ), .Y(new_n4998_));
  AOI21X1  g04806(.A0(new_n4998_), .A1(new_n4980_), .B0(new_n4986_), .Y(new_n4999_));
  OAI21X1  g04807(.A0(new_n4999_), .A1(new_n4981_), .B0(\asqrt[50] ), .Y(new_n5000_));
  AND2X1   g04808(.A(new_n4643_), .B(new_n4625_), .Y(new_n5001_));
  NOR3X1   g04809(.A(new_n5001_), .B(new_n4660_), .C(new_n4626_), .Y(new_n5002_));
  NOR3X1   g04810(.A(new_n4826_), .B(new_n5001_), .C(new_n4626_), .Y(new_n5003_));
  NOR2X1   g04811(.A(new_n5003_), .B(new_n4631_), .Y(new_n5004_));
  AOI21X1  g04812(.A0(new_n5002_), .A1(\asqrt[37] ), .B0(new_n5004_), .Y(new_n5005_));
  NOR3X1   g04813(.A(new_n4999_), .B(new_n4981_), .C(\asqrt[50] ), .Y(new_n5006_));
  OAI21X1  g04814(.A0(new_n5006_), .A1(new_n5005_), .B0(new_n5000_), .Y(new_n5007_));
  AND2X1   g04815(.A(new_n5007_), .B(\asqrt[51] ), .Y(new_n5008_));
  INVX1    g04816(.A(new_n5005_), .Y(new_n5009_));
  AND2X1   g04817(.A(new_n4997_), .B(\asqrt[48] ), .Y(new_n5010_));
  NAND2X1  g04818(.A(new_n4970_), .B(new_n4969_), .Y(new_n5011_));
  NOR2X1   g04819(.A(new_n4963_), .B(\asqrt[48] ), .Y(new_n5012_));
  AOI21X1  g04820(.A0(new_n5012_), .A1(new_n5011_), .B0(new_n4977_), .Y(new_n5013_));
  OAI21X1  g04821(.A0(new_n5013_), .A1(new_n5010_), .B0(\asqrt[49] ), .Y(new_n5014_));
  INVX1    g04822(.A(new_n4986_), .Y(new_n5015_));
  OAI21X1  g04823(.A0(new_n4971_), .A1(new_n1834_), .B0(new_n1632_), .Y(new_n5016_));
  OAI21X1  g04824(.A0(new_n5016_), .A1(new_n5013_), .B0(new_n5015_), .Y(new_n5017_));
  NAND3X1  g04825(.A(new_n5017_), .B(new_n5014_), .C(new_n1469_), .Y(new_n5018_));
  NAND2X1  g04826(.A(new_n5018_), .B(new_n5009_), .Y(new_n5019_));
  NAND4X1  g04827(.A(\asqrt[37] ), .B(new_n4663_), .C(new_n4649_), .D(new_n4645_), .Y(new_n5020_));
  NAND2X1  g04828(.A(new_n4663_), .B(new_n4645_), .Y(new_n5021_));
  OAI21X1  g04829(.A0(new_n5021_), .A1(new_n4826_), .B0(new_n4653_), .Y(new_n5022_));
  AND2X1   g04830(.A(new_n5022_), .B(new_n5020_), .Y(new_n5023_));
  AOI21X1  g04831(.A0(new_n5017_), .A1(new_n5014_), .B0(new_n1469_), .Y(new_n5024_));
  NOR2X1   g04832(.A(new_n5024_), .B(\asqrt[51] ), .Y(new_n5025_));
  AOI21X1  g04833(.A0(new_n5025_), .A1(new_n5019_), .B0(new_n5023_), .Y(new_n5026_));
  OAI21X1  g04834(.A0(new_n5026_), .A1(new_n5008_), .B0(\asqrt[52] ), .Y(new_n5027_));
  AND2X1   g04835(.A(new_n4671_), .B(new_n4664_), .Y(new_n5028_));
  NOR3X1   g04836(.A(new_n5028_), .B(new_n4709_), .C(new_n4652_), .Y(new_n5029_));
  NOR3X1   g04837(.A(new_n4826_), .B(new_n5028_), .C(new_n4652_), .Y(new_n5030_));
  NOR2X1   g04838(.A(new_n5030_), .B(new_n4669_), .Y(new_n5031_));
  AOI21X1  g04839(.A0(new_n5029_), .A1(\asqrt[37] ), .B0(new_n5031_), .Y(new_n5032_));
  INVX1    g04840(.A(new_n5032_), .Y(new_n5033_));
  AOI21X1  g04841(.A0(new_n5018_), .A1(new_n5009_), .B0(new_n5024_), .Y(new_n5034_));
  OAI21X1  g04842(.A0(new_n5034_), .A1(new_n1277_), .B0(new_n1111_), .Y(new_n5035_));
  OAI21X1  g04843(.A0(new_n5035_), .A1(new_n5026_), .B0(new_n5033_), .Y(new_n5036_));
  AOI21X1  g04844(.A0(new_n5036_), .A1(new_n5027_), .B0(new_n968_), .Y(new_n5037_));
  AND2X1   g04845(.A(new_n4713_), .B(new_n4711_), .Y(new_n5038_));
  NOR3X1   g04846(.A(new_n5038_), .B(new_n4679_), .C(new_n4712_), .Y(new_n5039_));
  NOR3X1   g04847(.A(new_n4826_), .B(new_n5038_), .C(new_n4712_), .Y(new_n5040_));
  NOR2X1   g04848(.A(new_n5040_), .B(new_n4678_), .Y(new_n5041_));
  AOI21X1  g04849(.A0(new_n5039_), .A1(\asqrt[37] ), .B0(new_n5041_), .Y(new_n5042_));
  INVX1    g04850(.A(new_n5042_), .Y(new_n5043_));
  NAND3X1  g04851(.A(new_n5036_), .B(new_n5027_), .C(new_n968_), .Y(new_n5044_));
  AOI21X1  g04852(.A0(new_n5044_), .A1(new_n5043_), .B0(new_n5037_), .Y(new_n5045_));
  OR2X1    g04853(.A(new_n5045_), .B(new_n902_), .Y(new_n5046_));
  AND2X1   g04854(.A(new_n5044_), .B(new_n5043_), .Y(new_n5047_));
  NAND4X1  g04855(.A(\asqrt[37] ), .B(new_n4689_), .C(new_n4687_), .D(new_n4715_), .Y(new_n5048_));
  NAND2X1  g04856(.A(new_n4689_), .B(new_n4715_), .Y(new_n5049_));
  OAI21X1  g04857(.A0(new_n5049_), .A1(new_n4826_), .B0(new_n4688_), .Y(new_n5050_));
  AND2X1   g04858(.A(new_n5050_), .B(new_n5048_), .Y(new_n5051_));
  INVX1    g04859(.A(new_n5051_), .Y(new_n5052_));
  OR2X1    g04860(.A(new_n5037_), .B(\asqrt[54] ), .Y(new_n5053_));
  OAI21X1  g04861(.A0(new_n5053_), .A1(new_n5047_), .B0(new_n5052_), .Y(new_n5054_));
  AOI21X1  g04862(.A0(new_n5054_), .A1(new_n5046_), .B0(new_n697_), .Y(new_n5055_));
  AOI21X1  g04863(.A0(new_n4745_), .A1(new_n4744_), .B0(new_n4698_), .Y(new_n5056_));
  AND2X1   g04864(.A(new_n5056_), .B(new_n4691_), .Y(new_n5057_));
  AOI22X1  g04865(.A0(new_n4745_), .A1(new_n4744_), .B0(new_n4717_), .B1(\asqrt[54] ), .Y(new_n5058_));
  AOI21X1  g04866(.A0(new_n5058_), .A1(\asqrt[37] ), .B0(new_n4697_), .Y(new_n5059_));
  AOI21X1  g04867(.A0(new_n5057_), .A1(\asqrt[37] ), .B0(new_n5059_), .Y(new_n5060_));
  OR2X1    g04868(.A(new_n5034_), .B(new_n1277_), .Y(new_n5061_));
  AND2X1   g04869(.A(new_n5018_), .B(new_n5009_), .Y(new_n5062_));
  INVX1    g04870(.A(new_n5023_), .Y(new_n5063_));
  OR2X1    g04871(.A(new_n5024_), .B(\asqrt[51] ), .Y(new_n5064_));
  OAI21X1  g04872(.A0(new_n5064_), .A1(new_n5062_), .B0(new_n5063_), .Y(new_n5065_));
  AOI21X1  g04873(.A0(new_n5065_), .A1(new_n5061_), .B0(new_n1111_), .Y(new_n5066_));
  AOI21X1  g04874(.A0(new_n5007_), .A1(\asqrt[51] ), .B0(\asqrt[52] ), .Y(new_n5067_));
  AOI21X1  g04875(.A0(new_n5067_), .A1(new_n5065_), .B0(new_n5032_), .Y(new_n5068_));
  OAI21X1  g04876(.A0(new_n5068_), .A1(new_n5066_), .B0(\asqrt[53] ), .Y(new_n5069_));
  NOR3X1   g04877(.A(new_n5068_), .B(new_n5066_), .C(\asqrt[53] ), .Y(new_n5070_));
  OAI21X1  g04878(.A0(new_n5070_), .A1(new_n5042_), .B0(new_n5069_), .Y(new_n5071_));
  AOI21X1  g04879(.A0(new_n5071_), .A1(\asqrt[54] ), .B0(\asqrt[55] ), .Y(new_n5072_));
  AOI21X1  g04880(.A0(new_n5072_), .A1(new_n5054_), .B0(new_n5060_), .Y(new_n5073_));
  OAI21X1  g04881(.A0(new_n5073_), .A1(new_n5055_), .B0(\asqrt[56] ), .Y(new_n5074_));
  AND2X1   g04882(.A(new_n4718_), .B(new_n4700_), .Y(new_n5075_));
  NOR3X1   g04883(.A(new_n5075_), .B(new_n4748_), .C(new_n4701_), .Y(new_n5076_));
  NOR3X1   g04884(.A(new_n4826_), .B(new_n5075_), .C(new_n4701_), .Y(new_n5077_));
  NOR2X1   g04885(.A(new_n5077_), .B(new_n4706_), .Y(new_n5078_));
  AOI21X1  g04886(.A0(new_n5076_), .A1(\asqrt[37] ), .B0(new_n5078_), .Y(new_n5079_));
  NOR3X1   g04887(.A(new_n5073_), .B(new_n5055_), .C(\asqrt[56] ), .Y(new_n5080_));
  OAI21X1  g04888(.A0(new_n5080_), .A1(new_n5079_), .B0(new_n5074_), .Y(new_n5081_));
  AND2X1   g04889(.A(new_n5081_), .B(\asqrt[57] ), .Y(new_n5082_));
  OR2X1    g04890(.A(new_n5080_), .B(new_n5079_), .Y(new_n5083_));
  OR4X1    g04891(.A(new_n4826_), .B(new_n4725_), .C(new_n4752_), .D(new_n4751_), .Y(new_n5084_));
  OR2X1    g04892(.A(new_n4725_), .B(new_n4751_), .Y(new_n5085_));
  OAI21X1  g04893(.A0(new_n5085_), .A1(new_n4826_), .B0(new_n4752_), .Y(new_n5086_));
  AND2X1   g04894(.A(new_n5086_), .B(new_n5084_), .Y(new_n5087_));
  AND2X1   g04895(.A(new_n5074_), .B(new_n481_), .Y(new_n5088_));
  AOI21X1  g04896(.A0(new_n5088_), .A1(new_n5083_), .B0(new_n5087_), .Y(new_n5089_));
  OAI21X1  g04897(.A0(new_n5089_), .A1(new_n5082_), .B0(\asqrt[58] ), .Y(new_n5090_));
  AND2X1   g04898(.A(new_n4734_), .B(new_n4728_), .Y(new_n5091_));
  NOR3X1   g04899(.A(new_n5091_), .B(new_n4768_), .C(new_n4727_), .Y(new_n5092_));
  NOR3X1   g04900(.A(new_n4826_), .B(new_n5091_), .C(new_n4727_), .Y(new_n5093_));
  NOR2X1   g04901(.A(new_n5093_), .B(new_n4733_), .Y(new_n5094_));
  AOI21X1  g04902(.A0(new_n5092_), .A1(\asqrt[37] ), .B0(new_n5094_), .Y(new_n5095_));
  INVX1    g04903(.A(new_n5095_), .Y(new_n5096_));
  AND2X1   g04904(.A(new_n5071_), .B(\asqrt[54] ), .Y(new_n5097_));
  NAND2X1  g04905(.A(new_n5044_), .B(new_n5043_), .Y(new_n5098_));
  NOR2X1   g04906(.A(new_n5037_), .B(\asqrt[54] ), .Y(new_n5099_));
  AOI21X1  g04907(.A0(new_n5099_), .A1(new_n5098_), .B0(new_n5051_), .Y(new_n5100_));
  OAI21X1  g04908(.A0(new_n5100_), .A1(new_n5097_), .B0(\asqrt[55] ), .Y(new_n5101_));
  INVX1    g04909(.A(new_n5060_), .Y(new_n5102_));
  OAI21X1  g04910(.A0(new_n5045_), .A1(new_n902_), .B0(new_n697_), .Y(new_n5103_));
  OAI21X1  g04911(.A0(new_n5103_), .A1(new_n5100_), .B0(new_n5102_), .Y(new_n5104_));
  AOI21X1  g04912(.A0(new_n5104_), .A1(new_n5101_), .B0(new_n582_), .Y(new_n5105_));
  INVX1    g04913(.A(new_n5079_), .Y(new_n5106_));
  NAND3X1  g04914(.A(new_n5104_), .B(new_n5101_), .C(new_n582_), .Y(new_n5107_));
  AOI21X1  g04915(.A0(new_n5107_), .A1(new_n5106_), .B0(new_n5105_), .Y(new_n5108_));
  OAI21X1  g04916(.A0(new_n5108_), .A1(new_n481_), .B0(new_n399_), .Y(new_n5109_));
  OAI21X1  g04917(.A0(new_n5109_), .A1(new_n5089_), .B0(new_n5096_), .Y(new_n5110_));
  AOI21X1  g04918(.A0(new_n5110_), .A1(new_n5090_), .B0(new_n328_), .Y(new_n5111_));
  AND2X1   g04919(.A(new_n4772_), .B(new_n4770_), .Y(new_n5112_));
  NOR3X1   g04920(.A(new_n5112_), .B(new_n4742_), .C(new_n4771_), .Y(new_n5113_));
  NOR3X1   g04921(.A(new_n4826_), .B(new_n5112_), .C(new_n4771_), .Y(new_n5114_));
  NOR2X1   g04922(.A(new_n5114_), .B(new_n4741_), .Y(new_n5115_));
  AOI21X1  g04923(.A0(new_n5113_), .A1(\asqrt[37] ), .B0(new_n5115_), .Y(new_n5116_));
  INVX1    g04924(.A(new_n5116_), .Y(new_n5117_));
  NAND3X1  g04925(.A(new_n5110_), .B(new_n5090_), .C(new_n328_), .Y(new_n5118_));
  AOI21X1  g04926(.A0(new_n5118_), .A1(new_n5117_), .B0(new_n5111_), .Y(new_n5119_));
  OR2X1    g04927(.A(new_n5119_), .B(new_n292_), .Y(new_n5120_));
  OR2X1    g04928(.A(new_n5108_), .B(new_n481_), .Y(new_n5121_));
  NOR2X1   g04929(.A(new_n5080_), .B(new_n5079_), .Y(new_n5122_));
  INVX1    g04930(.A(new_n5087_), .Y(new_n5123_));
  NAND2X1  g04931(.A(new_n5074_), .B(new_n481_), .Y(new_n5124_));
  OAI21X1  g04932(.A0(new_n5124_), .A1(new_n5122_), .B0(new_n5123_), .Y(new_n5125_));
  AOI21X1  g04933(.A0(new_n5125_), .A1(new_n5121_), .B0(new_n399_), .Y(new_n5126_));
  AOI21X1  g04934(.A0(new_n5081_), .A1(\asqrt[57] ), .B0(\asqrt[58] ), .Y(new_n5127_));
  AOI21X1  g04935(.A0(new_n5127_), .A1(new_n5125_), .B0(new_n5095_), .Y(new_n5128_));
  NOR3X1   g04936(.A(new_n5128_), .B(new_n5126_), .C(\asqrt[59] ), .Y(new_n5129_));
  NOR2X1   g04937(.A(new_n5129_), .B(new_n5116_), .Y(new_n5130_));
  OAI21X1  g04938(.A0(new_n5128_), .A1(new_n5126_), .B0(\asqrt[59] ), .Y(new_n5131_));
  NAND2X1  g04939(.A(new_n5131_), .B(new_n292_), .Y(new_n5132_));
  OR4X1    g04940(.A(new_n4826_), .B(new_n4763_), .C(new_n4774_), .D(new_n4757_), .Y(new_n5133_));
  OR2X1    g04941(.A(new_n4774_), .B(new_n4757_), .Y(new_n5134_));
  OAI21X1  g04942(.A0(new_n5134_), .A1(new_n4826_), .B0(new_n4763_), .Y(new_n5135_));
  AND2X1   g04943(.A(new_n5135_), .B(new_n5133_), .Y(new_n5136_));
  INVX1    g04944(.A(new_n5136_), .Y(new_n5137_));
  OAI21X1  g04945(.A0(new_n5132_), .A1(new_n5130_), .B0(new_n5137_), .Y(new_n5138_));
  AOI21X1  g04946(.A0(new_n5138_), .A1(new_n5120_), .B0(new_n217_), .Y(new_n5139_));
  AOI21X1  g04947(.A0(new_n4834_), .A1(new_n4833_), .B0(new_n4781_), .Y(new_n5140_));
  AND2X1   g04948(.A(new_n5140_), .B(new_n4765_), .Y(new_n5141_));
  AOI22X1  g04949(.A0(new_n4834_), .A1(new_n4833_), .B0(new_n4791_), .B1(\asqrt[60] ), .Y(new_n5142_));
  AOI21X1  g04950(.A0(new_n5142_), .A1(\asqrt[37] ), .B0(new_n4780_), .Y(new_n5143_));
  AOI21X1  g04951(.A0(new_n5141_), .A1(\asqrt[37] ), .B0(new_n5143_), .Y(new_n5144_));
  OAI21X1  g04952(.A0(new_n5129_), .A1(new_n5116_), .B0(new_n5131_), .Y(new_n5145_));
  AOI21X1  g04953(.A0(new_n5145_), .A1(\asqrt[60] ), .B0(\asqrt[61] ), .Y(new_n5146_));
  AOI21X1  g04954(.A0(new_n5146_), .A1(new_n5138_), .B0(new_n5144_), .Y(new_n5147_));
  OAI21X1  g04955(.A0(new_n5147_), .A1(new_n5139_), .B0(\asqrt[62] ), .Y(new_n5148_));
  AND2X1   g04956(.A(new_n4792_), .B(new_n4784_), .Y(new_n5149_));
  NOR3X1   g04957(.A(new_n5149_), .B(new_n4837_), .C(new_n4785_), .Y(new_n5150_));
  NOR3X1   g04958(.A(new_n4826_), .B(new_n5149_), .C(new_n4785_), .Y(new_n5151_));
  NOR2X1   g04959(.A(new_n5151_), .B(new_n4790_), .Y(new_n5152_));
  AOI21X1  g04960(.A0(new_n5150_), .A1(\asqrt[37] ), .B0(new_n5152_), .Y(new_n5153_));
  NOR3X1   g04961(.A(new_n5147_), .B(new_n5139_), .C(\asqrt[62] ), .Y(new_n5154_));
  OAI21X1  g04962(.A0(new_n5154_), .A1(new_n5153_), .B0(new_n5148_), .Y(new_n5155_));
  NOR4X1   g04963(.A(new_n4826_), .B(new_n4799_), .C(new_n4841_), .D(new_n4840_), .Y(new_n5156_));
  NAND3X1  g04964(.A(\asqrt[37] ), .B(new_n4842_), .C(new_n4794_), .Y(new_n5157_));
  AOI21X1  g04965(.A0(new_n5157_), .A1(new_n4841_), .B0(new_n5156_), .Y(new_n5158_));
  INVX1    g04966(.A(new_n5158_), .Y(new_n5159_));
  AND2X1   g04967(.A(new_n4807_), .B(new_n4800_), .Y(new_n5160_));
  AOI21X1  g04968(.A0(new_n5160_), .A1(\asqrt[37] ), .B0(new_n4867_), .Y(new_n5161_));
  AND2X1   g04969(.A(new_n5161_), .B(new_n5159_), .Y(new_n5162_));
  AOI21X1  g04970(.A0(new_n5162_), .A1(new_n5155_), .B0(\asqrt[63] ), .Y(new_n5163_));
  NOR2X1   g04971(.A(new_n5154_), .B(new_n5153_), .Y(new_n5164_));
  NAND2X1  g04972(.A(new_n5158_), .B(new_n5148_), .Y(new_n5165_));
  AOI21X1  g04973(.A0(new_n4849_), .A1(new_n4845_), .B0(new_n4806_), .Y(new_n5166_));
  AOI21X1  g04974(.A0(new_n4807_), .A1(new_n4800_), .B0(new_n193_), .Y(new_n5167_));
  OAI21X1  g04975(.A0(new_n5166_), .A1(new_n4800_), .B0(new_n5167_), .Y(new_n5168_));
  INVX1    g04976(.A(new_n4805_), .Y(new_n5169_));
  NOR4X1   g04977(.A(new_n4823_), .B(new_n4817_), .C(new_n5169_), .D(new_n4802_), .Y(new_n5170_));
  OAI21X1  g04978(.A0(new_n4814_), .A1(new_n4813_), .B0(new_n5170_), .Y(new_n5171_));
  NOR2X1   g04979(.A(new_n5171_), .B(new_n4812_), .Y(new_n5172_));
  INVX1    g04980(.A(new_n5172_), .Y(new_n5173_));
  AND2X1   g04981(.A(new_n5173_), .B(new_n5168_), .Y(new_n5174_));
  OAI21X1  g04982(.A0(new_n5165_), .A1(new_n5164_), .B0(new_n5174_), .Y(new_n5175_));
  NOR2X1   g04983(.A(new_n5175_), .B(new_n5163_), .Y(new_n5176_));
  NOR2X1   g04984(.A(\a[71] ), .B(\a[70] ), .Y(new_n5177_));
  INVX1    g04985(.A(new_n5177_), .Y(new_n5178_));
  MX2X1    g04986(.A(new_n5178_), .B(new_n5176_), .S0(\a[72] ), .Y(new_n5179_));
  OAI21X1  g04987(.A0(new_n5175_), .A1(new_n5163_), .B0(\a[72] ), .Y(new_n5180_));
  OAI22X1  g04988(.A0(new_n5178_), .A1(\a[72] ), .B0(new_n4822_), .B1(new_n4818_), .Y(new_n5181_));
  NOR4X1   g04989(.A(new_n5181_), .B(new_n4817_), .C(new_n4867_), .D(new_n4812_), .Y(new_n5182_));
  AND2X1   g04990(.A(new_n5182_), .B(new_n5180_), .Y(new_n5183_));
  INVX1    g04991(.A(\a[73] ), .Y(new_n5184_));
  AND2X1   g04992(.A(new_n5145_), .B(\asqrt[60] ), .Y(new_n5185_));
  OR2X1    g04993(.A(new_n5129_), .B(new_n5116_), .Y(new_n5186_));
  AND2X1   g04994(.A(new_n5131_), .B(new_n292_), .Y(new_n5187_));
  AOI21X1  g04995(.A0(new_n5187_), .A1(new_n5186_), .B0(new_n5136_), .Y(new_n5188_));
  OAI21X1  g04996(.A0(new_n5188_), .A1(new_n5185_), .B0(\asqrt[61] ), .Y(new_n5189_));
  INVX1    g04997(.A(new_n5144_), .Y(new_n5190_));
  OAI21X1  g04998(.A0(new_n5119_), .A1(new_n292_), .B0(new_n217_), .Y(new_n5191_));
  OAI21X1  g04999(.A0(new_n5191_), .A1(new_n5188_), .B0(new_n5190_), .Y(new_n5192_));
  AOI21X1  g05000(.A0(new_n5192_), .A1(new_n5189_), .B0(new_n199_), .Y(new_n5193_));
  INVX1    g05001(.A(new_n5153_), .Y(new_n5194_));
  NAND3X1  g05002(.A(new_n5192_), .B(new_n5189_), .C(new_n199_), .Y(new_n5195_));
  AOI21X1  g05003(.A0(new_n5195_), .A1(new_n5194_), .B0(new_n5193_), .Y(new_n5196_));
  INVX1    g05004(.A(new_n5162_), .Y(new_n5197_));
  OAI21X1  g05005(.A0(new_n5197_), .A1(new_n5196_), .B0(new_n193_), .Y(new_n5198_));
  OR2X1    g05006(.A(new_n5154_), .B(new_n5153_), .Y(new_n5199_));
  AND2X1   g05007(.A(new_n5158_), .B(new_n5148_), .Y(new_n5200_));
  INVX1    g05008(.A(new_n5174_), .Y(new_n5201_));
  AOI21X1  g05009(.A0(new_n5200_), .A1(new_n5199_), .B0(new_n5201_), .Y(new_n5202_));
  AOI21X1  g05010(.A0(new_n5202_), .A1(new_n5198_), .B0(\a[72] ), .Y(new_n5203_));
  OAI21X1  g05011(.A0(new_n5175_), .A1(new_n5163_), .B0(new_n4828_), .Y(new_n5204_));
  OAI21X1  g05012(.A0(new_n5203_), .A1(new_n5184_), .B0(new_n5204_), .Y(new_n5205_));
  OAI22X1  g05013(.A0(new_n5205_), .A1(new_n5183_), .B0(new_n5179_), .B1(new_n4826_), .Y(new_n5206_));
  AND2X1   g05014(.A(new_n5206_), .B(\asqrt[38] ), .Y(new_n5207_));
  OR2X1    g05015(.A(new_n5205_), .B(new_n5183_), .Y(new_n5208_));
  OR2X1    g05016(.A(new_n5175_), .B(new_n5163_), .Y(\asqrt[36] ));
  MX2X1    g05017(.A(new_n5177_), .B(\asqrt[36] ), .S0(\a[72] ), .Y(new_n5210_));
  AOI21X1  g05018(.A0(new_n5210_), .A1(\asqrt[37] ), .B0(\asqrt[38] ), .Y(new_n5211_));
  INVX1    g05019(.A(new_n5168_), .Y(new_n5212_));
  NOR3X1   g05020(.A(new_n5172_), .B(new_n5212_), .C(new_n4826_), .Y(new_n5213_));
  OAI21X1  g05021(.A0(new_n5165_), .A1(new_n5164_), .B0(new_n5213_), .Y(new_n5214_));
  OR2X1    g05022(.A(new_n5214_), .B(new_n5163_), .Y(new_n5215_));
  AOI21X1  g05023(.A0(new_n5215_), .A1(new_n5204_), .B0(new_n4831_), .Y(new_n5216_));
  AOI21X1  g05024(.A0(new_n5202_), .A1(new_n5198_), .B0(new_n4829_), .Y(new_n5217_));
  OAI21X1  g05025(.A0(new_n5214_), .A1(new_n5163_), .B0(new_n4831_), .Y(new_n5218_));
  NOR2X1   g05026(.A(new_n5218_), .B(new_n5217_), .Y(new_n5219_));
  NOR2X1   g05027(.A(new_n5219_), .B(new_n5216_), .Y(new_n5220_));
  AOI21X1  g05028(.A0(new_n5211_), .A1(new_n5208_), .B0(new_n5220_), .Y(new_n5221_));
  OAI21X1  g05029(.A0(new_n5221_), .A1(new_n5207_), .B0(\asqrt[39] ), .Y(new_n5222_));
  AOI21X1  g05030(.A0(new_n4865_), .A1(\asqrt[38] ), .B0(new_n4853_), .Y(new_n5223_));
  AND2X1   g05031(.A(new_n5223_), .B(new_n4857_), .Y(new_n5224_));
  OAI21X1  g05032(.A0(new_n5175_), .A1(new_n5163_), .B0(new_n5223_), .Y(new_n5225_));
  AOI22X1  g05033(.A0(new_n5225_), .A1(new_n4863_), .B0(new_n5224_), .B1(\asqrt[36] ), .Y(new_n5226_));
  INVX1    g05034(.A(new_n5226_), .Y(new_n5227_));
  NAND2X1  g05035(.A(new_n5182_), .B(new_n5180_), .Y(new_n5228_));
  INVX1    g05036(.A(\a[72] ), .Y(new_n5229_));
  OAI21X1  g05037(.A0(new_n5175_), .A1(new_n5163_), .B0(new_n5229_), .Y(new_n5230_));
  AOI21X1  g05038(.A0(new_n5230_), .A1(\a[73] ), .B0(new_n5217_), .Y(new_n5231_));
  AOI22X1  g05039(.A0(new_n5231_), .A1(new_n5228_), .B0(new_n5210_), .B1(\asqrt[37] ), .Y(new_n5232_));
  OAI21X1  g05040(.A0(new_n5232_), .A1(new_n4493_), .B0(new_n4165_), .Y(new_n5233_));
  OAI21X1  g05041(.A0(new_n5233_), .A1(new_n5221_), .B0(new_n5227_), .Y(new_n5234_));
  AOI21X1  g05042(.A0(new_n5234_), .A1(new_n5222_), .B0(new_n3863_), .Y(new_n5235_));
  AOI21X1  g05043(.A0(new_n4866_), .A1(new_n4864_), .B0(new_n4901_), .Y(new_n5236_));
  AND2X1   g05044(.A(new_n5236_), .B(new_n4898_), .Y(new_n5237_));
  AOI22X1  g05045(.A0(new_n4866_), .A1(new_n4864_), .B0(new_n4858_), .B1(\asqrt[39] ), .Y(new_n5238_));
  OAI21X1  g05046(.A0(new_n5175_), .A1(new_n5163_), .B0(new_n5238_), .Y(new_n5239_));
  AOI22X1  g05047(.A0(new_n5239_), .A1(new_n4901_), .B0(new_n5237_), .B1(\asqrt[36] ), .Y(new_n5240_));
  INVX1    g05048(.A(new_n5240_), .Y(new_n5241_));
  NAND3X1  g05049(.A(new_n5234_), .B(new_n5222_), .C(new_n3863_), .Y(new_n5242_));
  AOI21X1  g05050(.A0(new_n5242_), .A1(new_n5241_), .B0(new_n5235_), .Y(new_n5243_));
  OR2X1    g05051(.A(new_n5243_), .B(new_n3564_), .Y(new_n5244_));
  OR2X1    g05052(.A(new_n5232_), .B(new_n4493_), .Y(new_n5245_));
  AND2X1   g05053(.A(new_n5231_), .B(new_n5228_), .Y(new_n5246_));
  OAI21X1  g05054(.A0(new_n5179_), .A1(new_n4826_), .B0(new_n4493_), .Y(new_n5247_));
  OR2X1    g05055(.A(new_n5219_), .B(new_n5216_), .Y(new_n5248_));
  OAI21X1  g05056(.A0(new_n5247_), .A1(new_n5246_), .B0(new_n5248_), .Y(new_n5249_));
  AOI21X1  g05057(.A0(new_n5249_), .A1(new_n5245_), .B0(new_n4165_), .Y(new_n5250_));
  AOI21X1  g05058(.A0(new_n5206_), .A1(\asqrt[38] ), .B0(\asqrt[39] ), .Y(new_n5251_));
  AOI21X1  g05059(.A0(new_n5251_), .A1(new_n5249_), .B0(new_n5226_), .Y(new_n5252_));
  NOR3X1   g05060(.A(new_n5252_), .B(new_n5250_), .C(\asqrt[40] ), .Y(new_n5253_));
  NOR2X1   g05061(.A(new_n5253_), .B(new_n5240_), .Y(new_n5254_));
  AND2X1   g05062(.A(new_n4904_), .B(new_n4902_), .Y(new_n5255_));
  NOR3X1   g05063(.A(new_n5255_), .B(new_n4882_), .C(new_n4903_), .Y(new_n5256_));
  NOR2X1   g05064(.A(new_n5255_), .B(new_n4903_), .Y(new_n5257_));
  OAI21X1  g05065(.A0(new_n5175_), .A1(new_n5163_), .B0(new_n5257_), .Y(new_n5258_));
  AOI22X1  g05066(.A0(new_n5258_), .A1(new_n4882_), .B0(new_n5256_), .B1(\asqrt[36] ), .Y(new_n5259_));
  INVX1    g05067(.A(new_n5259_), .Y(new_n5260_));
  OAI21X1  g05068(.A0(new_n5252_), .A1(new_n5250_), .B0(\asqrt[40] ), .Y(new_n5261_));
  NAND2X1  g05069(.A(new_n5261_), .B(new_n3564_), .Y(new_n5262_));
  OAI21X1  g05070(.A0(new_n5262_), .A1(new_n5254_), .B0(new_n5260_), .Y(new_n5263_));
  AOI21X1  g05071(.A0(new_n5263_), .A1(new_n5244_), .B0(new_n3276_), .Y(new_n5264_));
  NAND4X1  g05072(.A(\asqrt[36] ), .B(new_n4895_), .C(new_n4893_), .D(new_n4922_), .Y(new_n5265_));
  NOR3X1   g05073(.A(new_n5176_), .B(new_n4906_), .C(new_n4886_), .Y(new_n5266_));
  OAI21X1  g05074(.A0(new_n5266_), .A1(new_n4893_), .B0(new_n5265_), .Y(new_n5267_));
  INVX1    g05075(.A(new_n5267_), .Y(new_n5268_));
  OAI21X1  g05076(.A0(new_n5253_), .A1(new_n5240_), .B0(new_n5261_), .Y(new_n5269_));
  AOI21X1  g05077(.A0(new_n5269_), .A1(\asqrt[41] ), .B0(\asqrt[42] ), .Y(new_n5270_));
  AOI21X1  g05078(.A0(new_n5270_), .A1(new_n5263_), .B0(new_n5268_), .Y(new_n5271_));
  OAI21X1  g05079(.A0(new_n5271_), .A1(new_n5264_), .B0(\asqrt[43] ), .Y(new_n5272_));
  AND2X1   g05080(.A(new_n4951_), .B(new_n4950_), .Y(new_n5273_));
  NOR3X1   g05081(.A(new_n5273_), .B(new_n4913_), .C(new_n4949_), .Y(new_n5274_));
  AOI22X1  g05082(.A0(new_n4951_), .A1(new_n4950_), .B0(new_n4923_), .B1(\asqrt[42] ), .Y(new_n5275_));
  AOI21X1  g05083(.A0(new_n5275_), .A1(\asqrt[36] ), .B0(new_n4912_), .Y(new_n5276_));
  AOI21X1  g05084(.A0(new_n5274_), .A1(\asqrt[36] ), .B0(new_n5276_), .Y(new_n5277_));
  NOR3X1   g05085(.A(new_n5271_), .B(new_n5264_), .C(\asqrt[43] ), .Y(new_n5278_));
  OAI21X1  g05086(.A0(new_n5278_), .A1(new_n5277_), .B0(new_n5272_), .Y(new_n5279_));
  AND2X1   g05087(.A(new_n5279_), .B(\asqrt[44] ), .Y(new_n5280_));
  INVX1    g05088(.A(new_n5277_), .Y(new_n5281_));
  AND2X1   g05089(.A(new_n5269_), .B(\asqrt[41] ), .Y(new_n5282_));
  OR2X1    g05090(.A(new_n5253_), .B(new_n5240_), .Y(new_n5283_));
  AND2X1   g05091(.A(new_n5261_), .B(new_n3564_), .Y(new_n5284_));
  AOI21X1  g05092(.A0(new_n5284_), .A1(new_n5283_), .B0(new_n5259_), .Y(new_n5285_));
  OAI21X1  g05093(.A0(new_n5285_), .A1(new_n5282_), .B0(\asqrt[42] ), .Y(new_n5286_));
  OAI21X1  g05094(.A0(new_n5243_), .A1(new_n3564_), .B0(new_n3276_), .Y(new_n5287_));
  OAI21X1  g05095(.A0(new_n5287_), .A1(new_n5285_), .B0(new_n5267_), .Y(new_n5288_));
  NAND3X1  g05096(.A(new_n5288_), .B(new_n5286_), .C(new_n3008_), .Y(new_n5289_));
  NAND2X1  g05097(.A(new_n5289_), .B(new_n5281_), .Y(new_n5290_));
  AND2X1   g05098(.A(new_n4924_), .B(new_n4915_), .Y(new_n5291_));
  NOR3X1   g05099(.A(new_n5291_), .B(new_n4954_), .C(new_n4916_), .Y(new_n5292_));
  NOR2X1   g05100(.A(new_n5291_), .B(new_n4916_), .Y(new_n5293_));
  AOI21X1  g05101(.A0(new_n5293_), .A1(\asqrt[36] ), .B0(new_n4921_), .Y(new_n5294_));
  AOI21X1  g05102(.A0(new_n5292_), .A1(\asqrt[36] ), .B0(new_n5294_), .Y(new_n5295_));
  AND2X1   g05103(.A(new_n5272_), .B(new_n2769_), .Y(new_n5296_));
  AOI21X1  g05104(.A0(new_n5296_), .A1(new_n5290_), .B0(new_n5295_), .Y(new_n5297_));
  OAI21X1  g05105(.A0(new_n5297_), .A1(new_n5280_), .B0(\asqrt[45] ), .Y(new_n5298_));
  OR4X1    g05106(.A(new_n5176_), .B(new_n4932_), .C(new_n4958_), .D(new_n4957_), .Y(new_n5299_));
  OR2X1    g05107(.A(new_n4932_), .B(new_n4957_), .Y(new_n5300_));
  OAI21X1  g05108(.A0(new_n5300_), .A1(new_n5176_), .B0(new_n4958_), .Y(new_n5301_));
  AND2X1   g05109(.A(new_n5301_), .B(new_n5299_), .Y(new_n5302_));
  INVX1    g05110(.A(new_n5302_), .Y(new_n5303_));
  AOI21X1  g05111(.A0(new_n5288_), .A1(new_n5286_), .B0(new_n3008_), .Y(new_n5304_));
  AOI21X1  g05112(.A0(new_n5289_), .A1(new_n5281_), .B0(new_n5304_), .Y(new_n5305_));
  OAI21X1  g05113(.A0(new_n5305_), .A1(new_n2769_), .B0(new_n2570_), .Y(new_n5306_));
  OAI21X1  g05114(.A0(new_n5306_), .A1(new_n5297_), .B0(new_n5303_), .Y(new_n5307_));
  AOI21X1  g05115(.A0(new_n5307_), .A1(new_n5298_), .B0(new_n2263_), .Y(new_n5308_));
  AOI21X1  g05116(.A0(new_n4940_), .A1(new_n4935_), .B0(new_n4989_), .Y(new_n5309_));
  AND2X1   g05117(.A(new_n5309_), .B(new_n4987_), .Y(new_n5310_));
  AOI22X1  g05118(.A0(new_n4940_), .A1(new_n4935_), .B0(new_n4933_), .B1(\asqrt[45] ), .Y(new_n5311_));
  AOI21X1  g05119(.A0(new_n5311_), .A1(\asqrt[36] ), .B0(new_n4939_), .Y(new_n5312_));
  AOI21X1  g05120(.A0(new_n5310_), .A1(\asqrt[36] ), .B0(new_n5312_), .Y(new_n5313_));
  INVX1    g05121(.A(new_n5313_), .Y(new_n5314_));
  NAND3X1  g05122(.A(new_n5307_), .B(new_n5298_), .C(new_n2263_), .Y(new_n5315_));
  AOI21X1  g05123(.A0(new_n5315_), .A1(new_n5314_), .B0(new_n5308_), .Y(new_n5316_));
  OR2X1    g05124(.A(new_n5316_), .B(new_n2040_), .Y(new_n5317_));
  AND2X1   g05125(.A(new_n5315_), .B(new_n5314_), .Y(new_n5318_));
  AND2X1   g05126(.A(new_n4993_), .B(new_n4991_), .Y(new_n5319_));
  NOR3X1   g05127(.A(new_n5319_), .B(new_n4948_), .C(new_n4992_), .Y(new_n5320_));
  NOR2X1   g05128(.A(new_n5319_), .B(new_n4992_), .Y(new_n5321_));
  AOI21X1  g05129(.A0(new_n5321_), .A1(\asqrt[36] ), .B0(new_n4947_), .Y(new_n5322_));
  AOI21X1  g05130(.A0(new_n5320_), .A1(\asqrt[36] ), .B0(new_n5322_), .Y(new_n5323_));
  INVX1    g05131(.A(new_n5323_), .Y(new_n5324_));
  OR2X1    g05132(.A(new_n5305_), .B(new_n2769_), .Y(new_n5325_));
  AND2X1   g05133(.A(new_n5289_), .B(new_n5281_), .Y(new_n5326_));
  INVX1    g05134(.A(new_n5295_), .Y(new_n5327_));
  NAND2X1  g05135(.A(new_n5272_), .B(new_n2769_), .Y(new_n5328_));
  OAI21X1  g05136(.A0(new_n5328_), .A1(new_n5326_), .B0(new_n5327_), .Y(new_n5329_));
  AOI21X1  g05137(.A0(new_n5329_), .A1(new_n5325_), .B0(new_n2570_), .Y(new_n5330_));
  AOI21X1  g05138(.A0(new_n5279_), .A1(\asqrt[44] ), .B0(\asqrt[45] ), .Y(new_n5331_));
  AOI21X1  g05139(.A0(new_n5331_), .A1(new_n5329_), .B0(new_n5302_), .Y(new_n5332_));
  OAI21X1  g05140(.A0(new_n5332_), .A1(new_n5330_), .B0(\asqrt[46] ), .Y(new_n5333_));
  NAND2X1  g05141(.A(new_n5333_), .B(new_n2040_), .Y(new_n5334_));
  OAI21X1  g05142(.A0(new_n5334_), .A1(new_n5318_), .B0(new_n5324_), .Y(new_n5335_));
  AOI21X1  g05143(.A0(new_n5335_), .A1(new_n5317_), .B0(new_n1834_), .Y(new_n5336_));
  NAND4X1  g05144(.A(\asqrt[36] ), .B(new_n4970_), .C(new_n4968_), .D(new_n4995_), .Y(new_n5337_));
  NAND2X1  g05145(.A(new_n4970_), .B(new_n4995_), .Y(new_n5338_));
  OAI21X1  g05146(.A0(new_n5338_), .A1(new_n5176_), .B0(new_n4969_), .Y(new_n5339_));
  AND2X1   g05147(.A(new_n5339_), .B(new_n5337_), .Y(new_n5340_));
  NOR3X1   g05148(.A(new_n5332_), .B(new_n5330_), .C(\asqrt[46] ), .Y(new_n5341_));
  OAI21X1  g05149(.A0(new_n5341_), .A1(new_n5313_), .B0(new_n5333_), .Y(new_n5342_));
  AOI21X1  g05150(.A0(new_n5342_), .A1(\asqrt[47] ), .B0(\asqrt[48] ), .Y(new_n5343_));
  AOI21X1  g05151(.A0(new_n5343_), .A1(new_n5335_), .B0(new_n5340_), .Y(new_n5344_));
  OAI21X1  g05152(.A0(new_n5344_), .A1(new_n5336_), .B0(\asqrt[49] ), .Y(new_n5345_));
  AND2X1   g05153(.A(new_n5012_), .B(new_n5011_), .Y(new_n5346_));
  NOR3X1   g05154(.A(new_n5346_), .B(new_n4978_), .C(new_n5010_), .Y(new_n5347_));
  AOI22X1  g05155(.A0(new_n5012_), .A1(new_n5011_), .B0(new_n4997_), .B1(\asqrt[48] ), .Y(new_n5348_));
  AOI21X1  g05156(.A0(new_n5348_), .A1(\asqrt[36] ), .B0(new_n4977_), .Y(new_n5349_));
  AOI21X1  g05157(.A0(new_n5347_), .A1(\asqrt[36] ), .B0(new_n5349_), .Y(new_n5350_));
  NOR3X1   g05158(.A(new_n5344_), .B(new_n5336_), .C(\asqrt[49] ), .Y(new_n5351_));
  OAI21X1  g05159(.A0(new_n5351_), .A1(new_n5350_), .B0(new_n5345_), .Y(new_n5352_));
  AND2X1   g05160(.A(new_n5352_), .B(\asqrt[50] ), .Y(new_n5353_));
  INVX1    g05161(.A(new_n5350_), .Y(new_n5354_));
  AND2X1   g05162(.A(new_n5342_), .B(\asqrt[47] ), .Y(new_n5355_));
  NAND2X1  g05163(.A(new_n5315_), .B(new_n5314_), .Y(new_n5356_));
  AND2X1   g05164(.A(new_n5333_), .B(new_n2040_), .Y(new_n5357_));
  AOI21X1  g05165(.A0(new_n5357_), .A1(new_n5356_), .B0(new_n5323_), .Y(new_n5358_));
  OAI21X1  g05166(.A0(new_n5358_), .A1(new_n5355_), .B0(\asqrt[48] ), .Y(new_n5359_));
  INVX1    g05167(.A(new_n5340_), .Y(new_n5360_));
  OAI21X1  g05168(.A0(new_n5316_), .A1(new_n2040_), .B0(new_n1834_), .Y(new_n5361_));
  OAI21X1  g05169(.A0(new_n5361_), .A1(new_n5358_), .B0(new_n5360_), .Y(new_n5362_));
  NAND3X1  g05170(.A(new_n5362_), .B(new_n5359_), .C(new_n1632_), .Y(new_n5363_));
  NAND2X1  g05171(.A(new_n5363_), .B(new_n5354_), .Y(new_n5364_));
  AND2X1   g05172(.A(new_n4998_), .B(new_n4980_), .Y(new_n5365_));
  NOR3X1   g05173(.A(new_n5365_), .B(new_n5015_), .C(new_n4981_), .Y(new_n5366_));
  NOR2X1   g05174(.A(new_n5365_), .B(new_n4981_), .Y(new_n5367_));
  AOI21X1  g05175(.A0(new_n5367_), .A1(\asqrt[36] ), .B0(new_n4986_), .Y(new_n5368_));
  AOI21X1  g05176(.A0(new_n5366_), .A1(\asqrt[36] ), .B0(new_n5368_), .Y(new_n5369_));
  AND2X1   g05177(.A(new_n5345_), .B(new_n1469_), .Y(new_n5370_));
  AOI21X1  g05178(.A0(new_n5370_), .A1(new_n5364_), .B0(new_n5369_), .Y(new_n5371_));
  OAI21X1  g05179(.A0(new_n5371_), .A1(new_n5353_), .B0(\asqrt[51] ), .Y(new_n5372_));
  NAND4X1  g05180(.A(\asqrt[36] ), .B(new_n5018_), .C(new_n5005_), .D(new_n5000_), .Y(new_n5373_));
  NAND2X1  g05181(.A(new_n5018_), .B(new_n5000_), .Y(new_n5374_));
  OAI21X1  g05182(.A0(new_n5374_), .A1(new_n5176_), .B0(new_n5009_), .Y(new_n5375_));
  AND2X1   g05183(.A(new_n5375_), .B(new_n5373_), .Y(new_n5376_));
  INVX1    g05184(.A(new_n5376_), .Y(new_n5377_));
  AOI21X1  g05185(.A0(new_n5362_), .A1(new_n5359_), .B0(new_n1632_), .Y(new_n5378_));
  AOI21X1  g05186(.A0(new_n5363_), .A1(new_n5354_), .B0(new_n5378_), .Y(new_n5379_));
  OAI21X1  g05187(.A0(new_n5379_), .A1(new_n1469_), .B0(new_n1277_), .Y(new_n5380_));
  OAI21X1  g05188(.A0(new_n5380_), .A1(new_n5371_), .B0(new_n5377_), .Y(new_n5381_));
  AOI21X1  g05189(.A0(new_n5381_), .A1(new_n5372_), .B0(new_n1111_), .Y(new_n5382_));
  AOI21X1  g05190(.A0(new_n5025_), .A1(new_n5019_), .B0(new_n5063_), .Y(new_n5383_));
  AND2X1   g05191(.A(new_n5383_), .B(new_n5061_), .Y(new_n5384_));
  AOI22X1  g05192(.A0(new_n5025_), .A1(new_n5019_), .B0(new_n5007_), .B1(\asqrt[51] ), .Y(new_n5385_));
  AOI21X1  g05193(.A0(new_n5385_), .A1(\asqrt[36] ), .B0(new_n5023_), .Y(new_n5386_));
  AOI21X1  g05194(.A0(new_n5384_), .A1(\asqrt[36] ), .B0(new_n5386_), .Y(new_n5387_));
  INVX1    g05195(.A(new_n5387_), .Y(new_n5388_));
  NAND3X1  g05196(.A(new_n5381_), .B(new_n5372_), .C(new_n1111_), .Y(new_n5389_));
  AOI21X1  g05197(.A0(new_n5389_), .A1(new_n5388_), .B0(new_n5382_), .Y(new_n5390_));
  OR2X1    g05198(.A(new_n5390_), .B(new_n968_), .Y(new_n5391_));
  AND2X1   g05199(.A(new_n5389_), .B(new_n5388_), .Y(new_n5392_));
  AND2X1   g05200(.A(new_n5067_), .B(new_n5065_), .Y(new_n5393_));
  NOR3X1   g05201(.A(new_n5393_), .B(new_n5033_), .C(new_n5066_), .Y(new_n5394_));
  NOR2X1   g05202(.A(new_n5393_), .B(new_n5066_), .Y(new_n5395_));
  AOI21X1  g05203(.A0(new_n5395_), .A1(\asqrt[36] ), .B0(new_n5032_), .Y(new_n5396_));
  AOI21X1  g05204(.A0(new_n5394_), .A1(\asqrt[36] ), .B0(new_n5396_), .Y(new_n5397_));
  INVX1    g05205(.A(new_n5397_), .Y(new_n5398_));
  OR2X1    g05206(.A(new_n5379_), .B(new_n1469_), .Y(new_n5399_));
  AND2X1   g05207(.A(new_n5363_), .B(new_n5354_), .Y(new_n5400_));
  INVX1    g05208(.A(new_n5369_), .Y(new_n5401_));
  NAND2X1  g05209(.A(new_n5345_), .B(new_n1469_), .Y(new_n5402_));
  OAI21X1  g05210(.A0(new_n5402_), .A1(new_n5400_), .B0(new_n5401_), .Y(new_n5403_));
  AOI21X1  g05211(.A0(new_n5403_), .A1(new_n5399_), .B0(new_n1277_), .Y(new_n5404_));
  AOI21X1  g05212(.A0(new_n5352_), .A1(\asqrt[50] ), .B0(\asqrt[51] ), .Y(new_n5405_));
  AOI21X1  g05213(.A0(new_n5405_), .A1(new_n5403_), .B0(new_n5376_), .Y(new_n5406_));
  OAI21X1  g05214(.A0(new_n5406_), .A1(new_n5404_), .B0(\asqrt[52] ), .Y(new_n5407_));
  NAND2X1  g05215(.A(new_n5407_), .B(new_n968_), .Y(new_n5408_));
  OAI21X1  g05216(.A0(new_n5408_), .A1(new_n5392_), .B0(new_n5398_), .Y(new_n5409_));
  AOI21X1  g05217(.A0(new_n5409_), .A1(new_n5391_), .B0(new_n902_), .Y(new_n5410_));
  NAND4X1  g05218(.A(\asqrt[36] ), .B(new_n5044_), .C(new_n5042_), .D(new_n5069_), .Y(new_n5411_));
  OR2X1    g05219(.A(new_n5070_), .B(new_n5037_), .Y(new_n5412_));
  OAI21X1  g05220(.A0(new_n5412_), .A1(new_n5176_), .B0(new_n5043_), .Y(new_n5413_));
  AND2X1   g05221(.A(new_n5413_), .B(new_n5411_), .Y(new_n5414_));
  NOR3X1   g05222(.A(new_n5406_), .B(new_n5404_), .C(\asqrt[52] ), .Y(new_n5415_));
  OAI21X1  g05223(.A0(new_n5415_), .A1(new_n5387_), .B0(new_n5407_), .Y(new_n5416_));
  AOI21X1  g05224(.A0(new_n5416_), .A1(\asqrt[53] ), .B0(\asqrt[54] ), .Y(new_n5417_));
  AOI21X1  g05225(.A0(new_n5417_), .A1(new_n5409_), .B0(new_n5414_), .Y(new_n5418_));
  OAI21X1  g05226(.A0(new_n5418_), .A1(new_n5410_), .B0(\asqrt[55] ), .Y(new_n5419_));
  AND2X1   g05227(.A(new_n5099_), .B(new_n5098_), .Y(new_n5420_));
  NOR3X1   g05228(.A(new_n5420_), .B(new_n5052_), .C(new_n5097_), .Y(new_n5421_));
  AOI22X1  g05229(.A0(new_n5099_), .A1(new_n5098_), .B0(new_n5071_), .B1(\asqrt[54] ), .Y(new_n5422_));
  AOI21X1  g05230(.A0(new_n5422_), .A1(\asqrt[36] ), .B0(new_n5051_), .Y(new_n5423_));
  AOI21X1  g05231(.A0(new_n5421_), .A1(\asqrt[36] ), .B0(new_n5423_), .Y(new_n5424_));
  NOR3X1   g05232(.A(new_n5418_), .B(new_n5410_), .C(\asqrt[55] ), .Y(new_n5425_));
  OAI21X1  g05233(.A0(new_n5425_), .A1(new_n5424_), .B0(new_n5419_), .Y(new_n5426_));
  AND2X1   g05234(.A(new_n5426_), .B(\asqrt[56] ), .Y(new_n5427_));
  INVX1    g05235(.A(new_n5424_), .Y(new_n5428_));
  AND2X1   g05236(.A(new_n5416_), .B(\asqrt[53] ), .Y(new_n5429_));
  NAND2X1  g05237(.A(new_n5389_), .B(new_n5388_), .Y(new_n5430_));
  AND2X1   g05238(.A(new_n5407_), .B(new_n968_), .Y(new_n5431_));
  AOI21X1  g05239(.A0(new_n5431_), .A1(new_n5430_), .B0(new_n5397_), .Y(new_n5432_));
  OAI21X1  g05240(.A0(new_n5432_), .A1(new_n5429_), .B0(\asqrt[54] ), .Y(new_n5433_));
  INVX1    g05241(.A(new_n5414_), .Y(new_n5434_));
  OAI21X1  g05242(.A0(new_n5390_), .A1(new_n968_), .B0(new_n902_), .Y(new_n5435_));
  OAI21X1  g05243(.A0(new_n5435_), .A1(new_n5432_), .B0(new_n5434_), .Y(new_n5436_));
  NAND3X1  g05244(.A(new_n5436_), .B(new_n5433_), .C(new_n697_), .Y(new_n5437_));
  NAND2X1  g05245(.A(new_n5437_), .B(new_n5428_), .Y(new_n5438_));
  AND2X1   g05246(.A(new_n5072_), .B(new_n5054_), .Y(new_n5439_));
  NOR3X1   g05247(.A(new_n5439_), .B(new_n5102_), .C(new_n5055_), .Y(new_n5440_));
  NOR2X1   g05248(.A(new_n5439_), .B(new_n5055_), .Y(new_n5441_));
  AOI21X1  g05249(.A0(new_n5441_), .A1(\asqrt[36] ), .B0(new_n5060_), .Y(new_n5442_));
  AOI21X1  g05250(.A0(new_n5440_), .A1(\asqrt[36] ), .B0(new_n5442_), .Y(new_n5443_));
  AND2X1   g05251(.A(new_n5419_), .B(new_n582_), .Y(new_n5444_));
  AOI21X1  g05252(.A0(new_n5444_), .A1(new_n5438_), .B0(new_n5443_), .Y(new_n5445_));
  OAI21X1  g05253(.A0(new_n5445_), .A1(new_n5427_), .B0(\asqrt[57] ), .Y(new_n5446_));
  OR4X1    g05254(.A(new_n5176_), .B(new_n5080_), .C(new_n5106_), .D(new_n5105_), .Y(new_n5447_));
  OR2X1    g05255(.A(new_n5080_), .B(new_n5105_), .Y(new_n5448_));
  OAI21X1  g05256(.A0(new_n5448_), .A1(new_n5176_), .B0(new_n5106_), .Y(new_n5449_));
  AND2X1   g05257(.A(new_n5449_), .B(new_n5447_), .Y(new_n5450_));
  INVX1    g05258(.A(new_n5450_), .Y(new_n5451_));
  AOI21X1  g05259(.A0(new_n5436_), .A1(new_n5433_), .B0(new_n697_), .Y(new_n5452_));
  AOI21X1  g05260(.A0(new_n5437_), .A1(new_n5428_), .B0(new_n5452_), .Y(new_n5453_));
  OAI21X1  g05261(.A0(new_n5453_), .A1(new_n582_), .B0(new_n481_), .Y(new_n5454_));
  OAI21X1  g05262(.A0(new_n5454_), .A1(new_n5445_), .B0(new_n5451_), .Y(new_n5455_));
  AOI21X1  g05263(.A0(new_n5455_), .A1(new_n5446_), .B0(new_n399_), .Y(new_n5456_));
  AOI21X1  g05264(.A0(new_n5088_), .A1(new_n5083_), .B0(new_n5123_), .Y(new_n5457_));
  AND2X1   g05265(.A(new_n5457_), .B(new_n5121_), .Y(new_n5458_));
  AOI22X1  g05266(.A0(new_n5088_), .A1(new_n5083_), .B0(new_n5081_), .B1(\asqrt[57] ), .Y(new_n5459_));
  AOI21X1  g05267(.A0(new_n5459_), .A1(\asqrt[36] ), .B0(new_n5087_), .Y(new_n5460_));
  AOI21X1  g05268(.A0(new_n5458_), .A1(\asqrt[36] ), .B0(new_n5460_), .Y(new_n5461_));
  INVX1    g05269(.A(new_n5461_), .Y(new_n5462_));
  NAND3X1  g05270(.A(new_n5455_), .B(new_n5446_), .C(new_n399_), .Y(new_n5463_));
  AOI21X1  g05271(.A0(new_n5463_), .A1(new_n5462_), .B0(new_n5456_), .Y(new_n5464_));
  OR2X1    g05272(.A(new_n5464_), .B(new_n328_), .Y(new_n5465_));
  AND2X1   g05273(.A(new_n5463_), .B(new_n5462_), .Y(new_n5466_));
  AND2X1   g05274(.A(new_n5127_), .B(new_n5125_), .Y(new_n5467_));
  NOR3X1   g05275(.A(new_n5467_), .B(new_n5096_), .C(new_n5126_), .Y(new_n5468_));
  NOR2X1   g05276(.A(new_n5467_), .B(new_n5126_), .Y(new_n5469_));
  AOI21X1  g05277(.A0(new_n5469_), .A1(\asqrt[36] ), .B0(new_n5095_), .Y(new_n5470_));
  AOI21X1  g05278(.A0(new_n5468_), .A1(\asqrt[36] ), .B0(new_n5470_), .Y(new_n5471_));
  INVX1    g05279(.A(new_n5471_), .Y(new_n5472_));
  OR2X1    g05280(.A(new_n5453_), .B(new_n582_), .Y(new_n5473_));
  AND2X1   g05281(.A(new_n5437_), .B(new_n5428_), .Y(new_n5474_));
  INVX1    g05282(.A(new_n5443_), .Y(new_n5475_));
  NAND2X1  g05283(.A(new_n5419_), .B(new_n582_), .Y(new_n5476_));
  OAI21X1  g05284(.A0(new_n5476_), .A1(new_n5474_), .B0(new_n5475_), .Y(new_n5477_));
  AOI21X1  g05285(.A0(new_n5477_), .A1(new_n5473_), .B0(new_n481_), .Y(new_n5478_));
  AOI21X1  g05286(.A0(new_n5426_), .A1(\asqrt[56] ), .B0(\asqrt[57] ), .Y(new_n5479_));
  AOI21X1  g05287(.A0(new_n5479_), .A1(new_n5477_), .B0(new_n5450_), .Y(new_n5480_));
  OAI21X1  g05288(.A0(new_n5480_), .A1(new_n5478_), .B0(\asqrt[58] ), .Y(new_n5481_));
  NAND2X1  g05289(.A(new_n5481_), .B(new_n328_), .Y(new_n5482_));
  OAI21X1  g05290(.A0(new_n5482_), .A1(new_n5466_), .B0(new_n5472_), .Y(new_n5483_));
  AOI21X1  g05291(.A0(new_n5483_), .A1(new_n5465_), .B0(new_n292_), .Y(new_n5484_));
  OR4X1    g05292(.A(new_n5176_), .B(new_n5129_), .C(new_n5117_), .D(new_n5111_), .Y(new_n5485_));
  OR2X1    g05293(.A(new_n5129_), .B(new_n5111_), .Y(new_n5486_));
  OAI21X1  g05294(.A0(new_n5486_), .A1(new_n5176_), .B0(new_n5117_), .Y(new_n5487_));
  AND2X1   g05295(.A(new_n5487_), .B(new_n5485_), .Y(new_n5488_));
  NOR3X1   g05296(.A(new_n5480_), .B(new_n5478_), .C(\asqrt[58] ), .Y(new_n5489_));
  OAI21X1  g05297(.A0(new_n5489_), .A1(new_n5461_), .B0(new_n5481_), .Y(new_n5490_));
  AOI21X1  g05298(.A0(new_n5490_), .A1(\asqrt[59] ), .B0(\asqrt[60] ), .Y(new_n5491_));
  AOI21X1  g05299(.A0(new_n5491_), .A1(new_n5483_), .B0(new_n5488_), .Y(new_n5492_));
  OAI21X1  g05300(.A0(new_n5492_), .A1(new_n5484_), .B0(\asqrt[61] ), .Y(new_n5493_));
  NOR3X1   g05301(.A(new_n5492_), .B(new_n5484_), .C(\asqrt[61] ), .Y(new_n5494_));
  AND2X1   g05302(.A(new_n5187_), .B(new_n5186_), .Y(new_n5495_));
  NOR3X1   g05303(.A(new_n5137_), .B(new_n5495_), .C(new_n5185_), .Y(new_n5496_));
  AOI22X1  g05304(.A0(new_n5187_), .A1(new_n5186_), .B0(new_n5145_), .B1(\asqrt[60] ), .Y(new_n5497_));
  AOI21X1  g05305(.A0(new_n5497_), .A1(\asqrt[36] ), .B0(new_n5136_), .Y(new_n5498_));
  AOI21X1  g05306(.A0(new_n5496_), .A1(\asqrt[36] ), .B0(new_n5498_), .Y(new_n5499_));
  OAI21X1  g05307(.A0(new_n5499_), .A1(new_n5494_), .B0(new_n5493_), .Y(new_n5500_));
  AND2X1   g05308(.A(new_n5500_), .B(\asqrt[62] ), .Y(new_n5501_));
  OR2X1    g05309(.A(new_n5499_), .B(new_n5494_), .Y(new_n5502_));
  AND2X1   g05310(.A(new_n5146_), .B(new_n5138_), .Y(new_n5503_));
  NOR3X1   g05311(.A(new_n5503_), .B(new_n5190_), .C(new_n5139_), .Y(new_n5504_));
  NOR2X1   g05312(.A(new_n5503_), .B(new_n5139_), .Y(new_n5505_));
  AOI21X1  g05313(.A0(new_n5505_), .A1(\asqrt[36] ), .B0(new_n5144_), .Y(new_n5506_));
  AOI21X1  g05314(.A0(new_n5504_), .A1(\asqrt[36] ), .B0(new_n5506_), .Y(new_n5507_));
  AND2X1   g05315(.A(new_n5493_), .B(new_n199_), .Y(new_n5508_));
  AOI21X1  g05316(.A0(new_n5508_), .A1(new_n5502_), .B0(new_n5507_), .Y(new_n5509_));
  NOR3X1   g05317(.A(new_n5154_), .B(new_n5194_), .C(new_n5193_), .Y(new_n5510_));
  AND2X1   g05318(.A(new_n5510_), .B(\asqrt[36] ), .Y(new_n5511_));
  NAND3X1  g05319(.A(\asqrt[36] ), .B(new_n5195_), .C(new_n5148_), .Y(new_n5512_));
  AOI21X1  g05320(.A0(new_n5512_), .A1(new_n5194_), .B0(new_n5511_), .Y(new_n5513_));
  INVX1    g05321(.A(new_n5513_), .Y(new_n5514_));
  AND2X1   g05322(.A(new_n5159_), .B(new_n5155_), .Y(new_n5515_));
  AOI22X1  g05323(.A0(new_n5515_), .A1(\asqrt[36] ), .B0(new_n5200_), .B1(new_n5199_), .Y(new_n5516_));
  AND2X1   g05324(.A(new_n5516_), .B(new_n5514_), .Y(new_n5517_));
  OAI21X1  g05325(.A0(new_n5509_), .A1(new_n5501_), .B0(new_n5517_), .Y(new_n5518_));
  AND2X1   g05326(.A(new_n5490_), .B(\asqrt[59] ), .Y(new_n5519_));
  OR2X1    g05327(.A(new_n5489_), .B(new_n5461_), .Y(new_n5520_));
  AND2X1   g05328(.A(new_n5481_), .B(new_n328_), .Y(new_n5521_));
  AOI21X1  g05329(.A0(new_n5521_), .A1(new_n5520_), .B0(new_n5471_), .Y(new_n5522_));
  OAI21X1  g05330(.A0(new_n5522_), .A1(new_n5519_), .B0(\asqrt[60] ), .Y(new_n5523_));
  INVX1    g05331(.A(new_n5488_), .Y(new_n5524_));
  OAI21X1  g05332(.A0(new_n5464_), .A1(new_n328_), .B0(new_n292_), .Y(new_n5525_));
  OAI21X1  g05333(.A0(new_n5525_), .A1(new_n5522_), .B0(new_n5524_), .Y(new_n5526_));
  AOI21X1  g05334(.A0(new_n5526_), .A1(new_n5523_), .B0(new_n217_), .Y(new_n5527_));
  NAND3X1  g05335(.A(new_n5526_), .B(new_n5523_), .C(new_n217_), .Y(new_n5528_));
  INVX1    g05336(.A(new_n5499_), .Y(new_n5529_));
  AOI21X1  g05337(.A0(new_n5529_), .A1(new_n5528_), .B0(new_n5527_), .Y(new_n5530_));
  OAI21X1  g05338(.A0(new_n5530_), .A1(new_n199_), .B0(new_n5513_), .Y(new_n5531_));
  AOI21X1  g05339(.A0(new_n5202_), .A1(new_n5198_), .B0(new_n5158_), .Y(new_n5532_));
  AOI21X1  g05340(.A0(new_n5159_), .A1(new_n5155_), .B0(new_n193_), .Y(new_n5533_));
  OAI21X1  g05341(.A0(new_n5532_), .A1(new_n5155_), .B0(new_n5533_), .Y(new_n5534_));
  OR2X1    g05342(.A(new_n5165_), .B(new_n5164_), .Y(new_n5535_));
  AND2X1   g05343(.A(new_n5157_), .B(new_n4841_), .Y(new_n5536_));
  NOR4X1   g05344(.A(new_n5172_), .B(new_n5212_), .C(new_n5536_), .D(new_n5156_), .Y(new_n5537_));
  NAND3X1  g05345(.A(new_n5537_), .B(new_n5535_), .C(new_n5198_), .Y(new_n5538_));
  AND2X1   g05346(.A(new_n5538_), .B(new_n5534_), .Y(new_n5539_));
  OAI21X1  g05347(.A0(new_n5531_), .A1(new_n5509_), .B0(new_n5539_), .Y(new_n5540_));
  AOI21X1  g05348(.A0(new_n5518_), .A1(new_n193_), .B0(new_n5540_), .Y(new_n5541_));
  NOR2X1   g05349(.A(\a[69] ), .B(\a[68] ), .Y(new_n5542_));
  INVX1    g05350(.A(new_n5542_), .Y(new_n5543_));
  MX2X1    g05351(.A(new_n5543_), .B(new_n5541_), .S0(\a[70] ), .Y(new_n5544_));
  OR2X1    g05352(.A(new_n5544_), .B(new_n5176_), .Y(new_n5545_));
  INVX1    g05353(.A(\a[70] ), .Y(new_n5546_));
  NOR3X1   g05354(.A(\a[70] ), .B(\a[69] ), .C(\a[68] ), .Y(new_n5547_));
  NOR3X1   g05355(.A(new_n5547_), .B(new_n5172_), .C(new_n5212_), .Y(new_n5548_));
  NAND3X1  g05356(.A(new_n5548_), .B(new_n5535_), .C(new_n5198_), .Y(new_n5549_));
  INVX1    g05357(.A(new_n5549_), .Y(new_n5550_));
  OAI21X1  g05358(.A0(new_n5541_), .A1(new_n5546_), .B0(new_n5550_), .Y(new_n5551_));
  OAI21X1  g05359(.A0(new_n5541_), .A1(\a[70] ), .B0(\a[71] ), .Y(new_n5552_));
  OR2X1    g05360(.A(new_n5541_), .B(new_n5178_), .Y(new_n5553_));
  NAND3X1  g05361(.A(new_n5553_), .B(new_n5552_), .C(new_n5551_), .Y(new_n5554_));
  AOI21X1  g05362(.A0(new_n5554_), .A1(new_n5545_), .B0(new_n4826_), .Y(new_n5555_));
  OR2X1    g05363(.A(new_n5530_), .B(new_n199_), .Y(new_n5556_));
  NOR2X1   g05364(.A(new_n5499_), .B(new_n5494_), .Y(new_n5557_));
  INVX1    g05365(.A(new_n5507_), .Y(new_n5558_));
  NAND2X1  g05366(.A(new_n5493_), .B(new_n199_), .Y(new_n5559_));
  OAI21X1  g05367(.A0(new_n5559_), .A1(new_n5557_), .B0(new_n5558_), .Y(new_n5560_));
  INVX1    g05368(.A(new_n5517_), .Y(new_n5561_));
  AOI21X1  g05369(.A0(new_n5560_), .A1(new_n5556_), .B0(new_n5561_), .Y(new_n5562_));
  AOI21X1  g05370(.A0(new_n5500_), .A1(\asqrt[62] ), .B0(new_n5514_), .Y(new_n5563_));
  INVX1    g05371(.A(new_n5539_), .Y(new_n5564_));
  AOI21X1  g05372(.A0(new_n5563_), .A1(new_n5560_), .B0(new_n5564_), .Y(new_n5565_));
  OAI21X1  g05373(.A0(new_n5562_), .A1(\asqrt[63] ), .B0(new_n5565_), .Y(\asqrt[35] ));
  MX2X1    g05374(.A(new_n5542_), .B(\asqrt[35] ), .S0(\a[70] ), .Y(new_n5567_));
  AOI21X1  g05375(.A0(new_n5567_), .A1(\asqrt[36] ), .B0(\asqrt[37] ), .Y(new_n5568_));
  NAND3X1  g05376(.A(new_n5538_), .B(new_n5534_), .C(\asqrt[36] ), .Y(new_n5569_));
  INVX1    g05377(.A(new_n5569_), .Y(new_n5570_));
  OAI21X1  g05378(.A0(new_n5531_), .A1(new_n5509_), .B0(new_n5570_), .Y(new_n5571_));
  AOI21X1  g05379(.A0(new_n5518_), .A1(new_n193_), .B0(new_n5571_), .Y(new_n5572_));
  AOI21X1  g05380(.A0(\asqrt[35] ), .A1(new_n5177_), .B0(new_n5572_), .Y(new_n5573_));
  OR2X1    g05381(.A(new_n5573_), .B(new_n5229_), .Y(new_n5574_));
  AND2X1   g05382(.A(\asqrt[35] ), .B(new_n5177_), .Y(new_n5575_));
  OR2X1    g05383(.A(new_n5572_), .B(\a[72] ), .Y(new_n5576_));
  OR2X1    g05384(.A(new_n5576_), .B(new_n5575_), .Y(new_n5577_));
  AOI22X1  g05385(.A0(new_n5577_), .A1(new_n5574_), .B0(new_n5568_), .B1(new_n5554_), .Y(new_n5578_));
  OAI21X1  g05386(.A0(new_n5578_), .A1(new_n5555_), .B0(\asqrt[38] ), .Y(new_n5579_));
  AOI21X1  g05387(.A0(new_n5210_), .A1(\asqrt[37] ), .B0(new_n5183_), .Y(new_n5580_));
  NAND3X1  g05388(.A(new_n5580_), .B(\asqrt[35] ), .C(new_n5205_), .Y(new_n5581_));
  INVX1    g05389(.A(new_n5580_), .Y(new_n5582_));
  OAI21X1  g05390(.A0(new_n5582_), .A1(new_n5541_), .B0(new_n5231_), .Y(new_n5583_));
  AND2X1   g05391(.A(new_n5583_), .B(new_n5581_), .Y(new_n5584_));
  NOR3X1   g05392(.A(new_n5578_), .B(new_n5555_), .C(\asqrt[38] ), .Y(new_n5585_));
  OAI21X1  g05393(.A0(new_n5585_), .A1(new_n5584_), .B0(new_n5579_), .Y(new_n5586_));
  AND2X1   g05394(.A(new_n5586_), .B(\asqrt[39] ), .Y(new_n5587_));
  INVX1    g05395(.A(new_n5584_), .Y(new_n5588_));
  AND2X1   g05396(.A(new_n5567_), .B(\asqrt[36] ), .Y(new_n5589_));
  AOI21X1  g05397(.A0(\asqrt[35] ), .A1(\a[70] ), .B0(new_n5549_), .Y(new_n5590_));
  INVX1    g05398(.A(\a[71] ), .Y(new_n5591_));
  AOI21X1  g05399(.A0(\asqrt[35] ), .A1(new_n5546_), .B0(new_n5591_), .Y(new_n5592_));
  NOR3X1   g05400(.A(new_n5575_), .B(new_n5592_), .C(new_n5590_), .Y(new_n5593_));
  OAI21X1  g05401(.A0(new_n5593_), .A1(new_n5589_), .B0(\asqrt[37] ), .Y(new_n5594_));
  OAI21X1  g05402(.A0(new_n5544_), .A1(new_n5176_), .B0(new_n4826_), .Y(new_n5595_));
  OAI22X1  g05403(.A0(new_n5576_), .A1(new_n5575_), .B0(new_n5573_), .B1(new_n5229_), .Y(new_n5596_));
  OAI21X1  g05404(.A0(new_n5595_), .A1(new_n5593_), .B0(new_n5596_), .Y(new_n5597_));
  NAND3X1  g05405(.A(new_n5597_), .B(new_n5594_), .C(new_n4493_), .Y(new_n5598_));
  NAND2X1  g05406(.A(new_n5598_), .B(new_n5588_), .Y(new_n5599_));
  OAI21X1  g05407(.A0(new_n5247_), .A1(new_n5246_), .B0(new_n5220_), .Y(new_n5600_));
  OR2X1    g05408(.A(new_n5600_), .B(new_n5207_), .Y(new_n5601_));
  OR2X1    g05409(.A(new_n5601_), .B(new_n5541_), .Y(new_n5602_));
  OAI22X1  g05410(.A0(new_n5247_), .A1(new_n5246_), .B0(new_n5232_), .B1(new_n4493_), .Y(new_n5603_));
  OAI21X1  g05411(.A0(new_n5603_), .A1(new_n5541_), .B0(new_n5248_), .Y(new_n5604_));
  AND2X1   g05412(.A(new_n5604_), .B(new_n5602_), .Y(new_n5605_));
  AOI21X1  g05413(.A0(new_n5597_), .A1(new_n5594_), .B0(new_n4493_), .Y(new_n5606_));
  NOR2X1   g05414(.A(new_n5606_), .B(\asqrt[39] ), .Y(new_n5607_));
  AOI21X1  g05415(.A0(new_n5607_), .A1(new_n5599_), .B0(new_n5605_), .Y(new_n5608_));
  OAI21X1  g05416(.A0(new_n5608_), .A1(new_n5587_), .B0(\asqrt[40] ), .Y(new_n5609_));
  AND2X1   g05417(.A(new_n5251_), .B(new_n5249_), .Y(new_n5610_));
  OR4X1    g05418(.A(new_n5541_), .B(new_n5610_), .C(new_n5227_), .D(new_n5250_), .Y(new_n5611_));
  OR2X1    g05419(.A(new_n5610_), .B(new_n5250_), .Y(new_n5612_));
  OAI21X1  g05420(.A0(new_n5612_), .A1(new_n5541_), .B0(new_n5227_), .Y(new_n5613_));
  AND2X1   g05421(.A(new_n5613_), .B(new_n5611_), .Y(new_n5614_));
  INVX1    g05422(.A(new_n5614_), .Y(new_n5615_));
  AOI21X1  g05423(.A0(new_n5598_), .A1(new_n5588_), .B0(new_n5606_), .Y(new_n5616_));
  OAI21X1  g05424(.A0(new_n5616_), .A1(new_n4165_), .B0(new_n3863_), .Y(new_n5617_));
  OAI21X1  g05425(.A0(new_n5617_), .A1(new_n5608_), .B0(new_n5615_), .Y(new_n5618_));
  AOI21X1  g05426(.A0(new_n5618_), .A1(new_n5609_), .B0(new_n3564_), .Y(new_n5619_));
  NAND3X1  g05427(.A(new_n5242_), .B(new_n5240_), .C(new_n5261_), .Y(new_n5620_));
  NOR3X1   g05428(.A(new_n5541_), .B(new_n5253_), .C(new_n5235_), .Y(new_n5621_));
  OAI22X1  g05429(.A0(new_n5621_), .A1(new_n5240_), .B0(new_n5620_), .B1(new_n5541_), .Y(new_n5622_));
  NAND3X1  g05430(.A(new_n5618_), .B(new_n5609_), .C(new_n3564_), .Y(new_n5623_));
  AOI21X1  g05431(.A0(new_n5623_), .A1(new_n5622_), .B0(new_n5619_), .Y(new_n5624_));
  OR2X1    g05432(.A(new_n5624_), .B(new_n3276_), .Y(new_n5625_));
  AND2X1   g05433(.A(new_n5623_), .B(new_n5622_), .Y(new_n5626_));
  AND2X1   g05434(.A(new_n5284_), .B(new_n5283_), .Y(new_n5627_));
  NOR4X1   g05435(.A(new_n5541_), .B(new_n5627_), .C(new_n5260_), .D(new_n5282_), .Y(new_n5628_));
  AOI22X1  g05436(.A0(new_n5284_), .A1(new_n5283_), .B0(new_n5269_), .B1(\asqrt[41] ), .Y(new_n5629_));
  AOI21X1  g05437(.A0(new_n5629_), .A1(\asqrt[35] ), .B0(new_n5259_), .Y(new_n5630_));
  NOR2X1   g05438(.A(new_n5630_), .B(new_n5628_), .Y(new_n5631_));
  INVX1    g05439(.A(new_n5631_), .Y(new_n5632_));
  OR2X1    g05440(.A(new_n5619_), .B(\asqrt[42] ), .Y(new_n5633_));
  OAI21X1  g05441(.A0(new_n5633_), .A1(new_n5626_), .B0(new_n5632_), .Y(new_n5634_));
  AOI21X1  g05442(.A0(new_n5634_), .A1(new_n5625_), .B0(new_n3008_), .Y(new_n5635_));
  AND2X1   g05443(.A(new_n5270_), .B(new_n5263_), .Y(new_n5636_));
  OR4X1    g05444(.A(new_n5541_), .B(new_n5636_), .C(new_n5267_), .D(new_n5264_), .Y(new_n5637_));
  OR2X1    g05445(.A(new_n5636_), .B(new_n5264_), .Y(new_n5638_));
  OAI21X1  g05446(.A0(new_n5638_), .A1(new_n5541_), .B0(new_n5267_), .Y(new_n5639_));
  AND2X1   g05447(.A(new_n5639_), .B(new_n5637_), .Y(new_n5640_));
  OR2X1    g05448(.A(new_n5616_), .B(new_n4165_), .Y(new_n5641_));
  AND2X1   g05449(.A(new_n5598_), .B(new_n5588_), .Y(new_n5642_));
  INVX1    g05450(.A(new_n5605_), .Y(new_n5643_));
  OR2X1    g05451(.A(new_n5606_), .B(\asqrt[39] ), .Y(new_n5644_));
  OAI21X1  g05452(.A0(new_n5644_), .A1(new_n5642_), .B0(new_n5643_), .Y(new_n5645_));
  AOI21X1  g05453(.A0(new_n5645_), .A1(new_n5641_), .B0(new_n3863_), .Y(new_n5646_));
  AOI21X1  g05454(.A0(new_n5586_), .A1(\asqrt[39] ), .B0(\asqrt[40] ), .Y(new_n5647_));
  AOI21X1  g05455(.A0(new_n5647_), .A1(new_n5645_), .B0(new_n5614_), .Y(new_n5648_));
  OAI21X1  g05456(.A0(new_n5648_), .A1(new_n5646_), .B0(\asqrt[41] ), .Y(new_n5649_));
  INVX1    g05457(.A(new_n5622_), .Y(new_n5650_));
  NOR3X1   g05458(.A(new_n5648_), .B(new_n5646_), .C(\asqrt[41] ), .Y(new_n5651_));
  OAI21X1  g05459(.A0(new_n5651_), .A1(new_n5650_), .B0(new_n5649_), .Y(new_n5652_));
  AOI21X1  g05460(.A0(new_n5652_), .A1(\asqrt[42] ), .B0(\asqrt[43] ), .Y(new_n5653_));
  AOI21X1  g05461(.A0(new_n5653_), .A1(new_n5634_), .B0(new_n5640_), .Y(new_n5654_));
  OAI21X1  g05462(.A0(new_n5654_), .A1(new_n5635_), .B0(\asqrt[44] ), .Y(new_n5655_));
  OR4X1    g05463(.A(new_n5541_), .B(new_n5278_), .C(new_n5281_), .D(new_n5304_), .Y(new_n5656_));
  NAND2X1  g05464(.A(new_n5289_), .B(new_n5272_), .Y(new_n5657_));
  OAI21X1  g05465(.A0(new_n5657_), .A1(new_n5541_), .B0(new_n5281_), .Y(new_n5658_));
  AND2X1   g05466(.A(new_n5658_), .B(new_n5656_), .Y(new_n5659_));
  NOR3X1   g05467(.A(new_n5654_), .B(new_n5635_), .C(\asqrt[44] ), .Y(new_n5660_));
  OAI21X1  g05468(.A0(new_n5660_), .A1(new_n5659_), .B0(new_n5655_), .Y(new_n5661_));
  AND2X1   g05469(.A(new_n5661_), .B(\asqrt[45] ), .Y(new_n5662_));
  INVX1    g05470(.A(new_n5659_), .Y(new_n5663_));
  AND2X1   g05471(.A(new_n5652_), .B(\asqrt[42] ), .Y(new_n5664_));
  NAND2X1  g05472(.A(new_n5623_), .B(new_n5622_), .Y(new_n5665_));
  NOR2X1   g05473(.A(new_n5619_), .B(\asqrt[42] ), .Y(new_n5666_));
  AOI21X1  g05474(.A0(new_n5666_), .A1(new_n5665_), .B0(new_n5631_), .Y(new_n5667_));
  OAI21X1  g05475(.A0(new_n5667_), .A1(new_n5664_), .B0(\asqrt[43] ), .Y(new_n5668_));
  INVX1    g05476(.A(new_n5640_), .Y(new_n5669_));
  OAI21X1  g05477(.A0(new_n5624_), .A1(new_n3276_), .B0(new_n3008_), .Y(new_n5670_));
  OAI21X1  g05478(.A0(new_n5670_), .A1(new_n5667_), .B0(new_n5669_), .Y(new_n5671_));
  NAND3X1  g05479(.A(new_n5671_), .B(new_n5668_), .C(new_n2769_), .Y(new_n5672_));
  NAND2X1  g05480(.A(new_n5672_), .B(new_n5663_), .Y(new_n5673_));
  OAI21X1  g05481(.A0(new_n5328_), .A1(new_n5326_), .B0(new_n5295_), .Y(new_n5674_));
  NOR3X1   g05482(.A(new_n5674_), .B(new_n5541_), .C(new_n5280_), .Y(new_n5675_));
  AOI22X1  g05483(.A0(new_n5296_), .A1(new_n5290_), .B0(new_n5279_), .B1(\asqrt[44] ), .Y(new_n5676_));
  AOI21X1  g05484(.A0(new_n5676_), .A1(\asqrt[35] ), .B0(new_n5295_), .Y(new_n5677_));
  NOR2X1   g05485(.A(new_n5677_), .B(new_n5675_), .Y(new_n5678_));
  AOI21X1  g05486(.A0(new_n5671_), .A1(new_n5668_), .B0(new_n2769_), .Y(new_n5679_));
  NOR2X1   g05487(.A(new_n5679_), .B(\asqrt[45] ), .Y(new_n5680_));
  AOI21X1  g05488(.A0(new_n5680_), .A1(new_n5673_), .B0(new_n5678_), .Y(new_n5681_));
  OAI21X1  g05489(.A0(new_n5681_), .A1(new_n5662_), .B0(\asqrt[46] ), .Y(new_n5682_));
  AND2X1   g05490(.A(new_n5331_), .B(new_n5329_), .Y(new_n5683_));
  NOR4X1   g05491(.A(new_n5541_), .B(new_n5683_), .C(new_n5303_), .D(new_n5330_), .Y(new_n5684_));
  NOR2X1   g05492(.A(new_n5683_), .B(new_n5330_), .Y(new_n5685_));
  AOI21X1  g05493(.A0(new_n5685_), .A1(\asqrt[35] ), .B0(new_n5302_), .Y(new_n5686_));
  NOR2X1   g05494(.A(new_n5686_), .B(new_n5684_), .Y(new_n5687_));
  INVX1    g05495(.A(new_n5687_), .Y(new_n5688_));
  AOI21X1  g05496(.A0(new_n5672_), .A1(new_n5663_), .B0(new_n5679_), .Y(new_n5689_));
  OAI21X1  g05497(.A0(new_n5689_), .A1(new_n2570_), .B0(new_n2263_), .Y(new_n5690_));
  OAI21X1  g05498(.A0(new_n5690_), .A1(new_n5681_), .B0(new_n5688_), .Y(new_n5691_));
  AOI21X1  g05499(.A0(new_n5691_), .A1(new_n5682_), .B0(new_n2040_), .Y(new_n5692_));
  OR4X1    g05500(.A(new_n5541_), .B(new_n5341_), .C(new_n5314_), .D(new_n5308_), .Y(new_n5693_));
  NAND2X1  g05501(.A(new_n5315_), .B(new_n5333_), .Y(new_n5694_));
  OAI21X1  g05502(.A0(new_n5694_), .A1(new_n5541_), .B0(new_n5314_), .Y(new_n5695_));
  AND2X1   g05503(.A(new_n5695_), .B(new_n5693_), .Y(new_n5696_));
  INVX1    g05504(.A(new_n5696_), .Y(new_n5697_));
  NAND3X1  g05505(.A(new_n5691_), .B(new_n5682_), .C(new_n2040_), .Y(new_n5698_));
  AOI21X1  g05506(.A0(new_n5698_), .A1(new_n5697_), .B0(new_n5692_), .Y(new_n5699_));
  OR2X1    g05507(.A(new_n5699_), .B(new_n1834_), .Y(new_n5700_));
  AND2X1   g05508(.A(new_n5698_), .B(new_n5697_), .Y(new_n5701_));
  AND2X1   g05509(.A(new_n5357_), .B(new_n5356_), .Y(new_n5702_));
  NOR4X1   g05510(.A(new_n5541_), .B(new_n5702_), .C(new_n5324_), .D(new_n5355_), .Y(new_n5703_));
  AOI22X1  g05511(.A0(new_n5357_), .A1(new_n5356_), .B0(new_n5342_), .B1(\asqrt[47] ), .Y(new_n5704_));
  AOI21X1  g05512(.A0(new_n5704_), .A1(\asqrt[35] ), .B0(new_n5323_), .Y(new_n5705_));
  NOR2X1   g05513(.A(new_n5705_), .B(new_n5703_), .Y(new_n5706_));
  INVX1    g05514(.A(new_n5706_), .Y(new_n5707_));
  OR2X1    g05515(.A(new_n5692_), .B(\asqrt[48] ), .Y(new_n5708_));
  OAI21X1  g05516(.A0(new_n5708_), .A1(new_n5701_), .B0(new_n5707_), .Y(new_n5709_));
  AOI21X1  g05517(.A0(new_n5709_), .A1(new_n5700_), .B0(new_n1632_), .Y(new_n5710_));
  OAI21X1  g05518(.A0(new_n5361_), .A1(new_n5358_), .B0(new_n5340_), .Y(new_n5711_));
  OR2X1    g05519(.A(new_n5711_), .B(new_n5336_), .Y(new_n5712_));
  OAI21X1  g05520(.A0(new_n5361_), .A1(new_n5358_), .B0(new_n5359_), .Y(new_n5713_));
  NOR2X1   g05521(.A(new_n5713_), .B(new_n5541_), .Y(new_n5714_));
  OAI22X1  g05522(.A0(new_n5714_), .A1(new_n5340_), .B0(new_n5712_), .B1(new_n5541_), .Y(new_n5715_));
  INVX1    g05523(.A(new_n5715_), .Y(new_n5716_));
  OR2X1    g05524(.A(new_n5689_), .B(new_n2570_), .Y(new_n5717_));
  AND2X1   g05525(.A(new_n5672_), .B(new_n5663_), .Y(new_n5718_));
  INVX1    g05526(.A(new_n5678_), .Y(new_n5719_));
  OR2X1    g05527(.A(new_n5679_), .B(\asqrt[45] ), .Y(new_n5720_));
  OAI21X1  g05528(.A0(new_n5720_), .A1(new_n5718_), .B0(new_n5719_), .Y(new_n5721_));
  AOI21X1  g05529(.A0(new_n5721_), .A1(new_n5717_), .B0(new_n2263_), .Y(new_n5722_));
  AOI21X1  g05530(.A0(new_n5661_), .A1(\asqrt[45] ), .B0(\asqrt[46] ), .Y(new_n5723_));
  AOI21X1  g05531(.A0(new_n5723_), .A1(new_n5721_), .B0(new_n5687_), .Y(new_n5724_));
  OAI21X1  g05532(.A0(new_n5724_), .A1(new_n5722_), .B0(\asqrt[47] ), .Y(new_n5725_));
  NOR3X1   g05533(.A(new_n5724_), .B(new_n5722_), .C(\asqrt[47] ), .Y(new_n5726_));
  OAI21X1  g05534(.A0(new_n5726_), .A1(new_n5696_), .B0(new_n5725_), .Y(new_n5727_));
  AOI21X1  g05535(.A0(new_n5727_), .A1(\asqrt[48] ), .B0(\asqrt[49] ), .Y(new_n5728_));
  AOI21X1  g05536(.A0(new_n5728_), .A1(new_n5709_), .B0(new_n5716_), .Y(new_n5729_));
  OAI21X1  g05537(.A0(new_n5729_), .A1(new_n5710_), .B0(\asqrt[50] ), .Y(new_n5730_));
  OR4X1    g05538(.A(new_n5541_), .B(new_n5351_), .C(new_n5354_), .D(new_n5378_), .Y(new_n5731_));
  NAND2X1  g05539(.A(new_n5363_), .B(new_n5345_), .Y(new_n5732_));
  OAI21X1  g05540(.A0(new_n5732_), .A1(new_n5541_), .B0(new_n5354_), .Y(new_n5733_));
  AND2X1   g05541(.A(new_n5733_), .B(new_n5731_), .Y(new_n5734_));
  NOR3X1   g05542(.A(new_n5729_), .B(new_n5710_), .C(\asqrt[50] ), .Y(new_n5735_));
  OAI21X1  g05543(.A0(new_n5735_), .A1(new_n5734_), .B0(new_n5730_), .Y(new_n5736_));
  AND2X1   g05544(.A(new_n5736_), .B(\asqrt[51] ), .Y(new_n5737_));
  INVX1    g05545(.A(new_n5734_), .Y(new_n5738_));
  AND2X1   g05546(.A(new_n5727_), .B(\asqrt[48] ), .Y(new_n5739_));
  NAND2X1  g05547(.A(new_n5698_), .B(new_n5697_), .Y(new_n5740_));
  NOR2X1   g05548(.A(new_n5692_), .B(\asqrt[48] ), .Y(new_n5741_));
  AOI21X1  g05549(.A0(new_n5741_), .A1(new_n5740_), .B0(new_n5706_), .Y(new_n5742_));
  OAI21X1  g05550(.A0(new_n5742_), .A1(new_n5739_), .B0(\asqrt[49] ), .Y(new_n5743_));
  OAI21X1  g05551(.A0(new_n5699_), .A1(new_n1834_), .B0(new_n1632_), .Y(new_n5744_));
  OAI21X1  g05552(.A0(new_n5744_), .A1(new_n5742_), .B0(new_n5715_), .Y(new_n5745_));
  NAND3X1  g05553(.A(new_n5745_), .B(new_n5743_), .C(new_n1469_), .Y(new_n5746_));
  NAND2X1  g05554(.A(new_n5746_), .B(new_n5738_), .Y(new_n5747_));
  OAI21X1  g05555(.A0(new_n5402_), .A1(new_n5400_), .B0(new_n5369_), .Y(new_n5748_));
  NOR3X1   g05556(.A(new_n5748_), .B(new_n5541_), .C(new_n5353_), .Y(new_n5749_));
  AOI22X1  g05557(.A0(new_n5370_), .A1(new_n5364_), .B0(new_n5352_), .B1(\asqrt[50] ), .Y(new_n5750_));
  AOI21X1  g05558(.A0(new_n5750_), .A1(\asqrt[35] ), .B0(new_n5369_), .Y(new_n5751_));
  NOR2X1   g05559(.A(new_n5751_), .B(new_n5749_), .Y(new_n5752_));
  AOI21X1  g05560(.A0(new_n5745_), .A1(new_n5743_), .B0(new_n1469_), .Y(new_n5753_));
  NOR2X1   g05561(.A(new_n5753_), .B(\asqrt[51] ), .Y(new_n5754_));
  AOI21X1  g05562(.A0(new_n5754_), .A1(new_n5747_), .B0(new_n5752_), .Y(new_n5755_));
  OAI21X1  g05563(.A0(new_n5755_), .A1(new_n5737_), .B0(\asqrt[52] ), .Y(new_n5756_));
  AND2X1   g05564(.A(new_n5405_), .B(new_n5403_), .Y(new_n5757_));
  OR4X1    g05565(.A(new_n5541_), .B(new_n5757_), .C(new_n5377_), .D(new_n5404_), .Y(new_n5758_));
  OR2X1    g05566(.A(new_n5757_), .B(new_n5404_), .Y(new_n5759_));
  OAI21X1  g05567(.A0(new_n5759_), .A1(new_n5541_), .B0(new_n5377_), .Y(new_n5760_));
  AND2X1   g05568(.A(new_n5760_), .B(new_n5758_), .Y(new_n5761_));
  INVX1    g05569(.A(new_n5761_), .Y(new_n5762_));
  AOI21X1  g05570(.A0(new_n5746_), .A1(new_n5738_), .B0(new_n5753_), .Y(new_n5763_));
  OAI21X1  g05571(.A0(new_n5763_), .A1(new_n1277_), .B0(new_n1111_), .Y(new_n5764_));
  OAI21X1  g05572(.A0(new_n5764_), .A1(new_n5755_), .B0(new_n5762_), .Y(new_n5765_));
  AOI21X1  g05573(.A0(new_n5765_), .A1(new_n5756_), .B0(new_n968_), .Y(new_n5766_));
  OR4X1    g05574(.A(new_n5541_), .B(new_n5415_), .C(new_n5388_), .D(new_n5382_), .Y(new_n5767_));
  NAND2X1  g05575(.A(new_n5389_), .B(new_n5407_), .Y(new_n5768_));
  OAI21X1  g05576(.A0(new_n5768_), .A1(new_n5541_), .B0(new_n5388_), .Y(new_n5769_));
  AND2X1   g05577(.A(new_n5769_), .B(new_n5767_), .Y(new_n5770_));
  INVX1    g05578(.A(new_n5770_), .Y(new_n5771_));
  NAND3X1  g05579(.A(new_n5765_), .B(new_n5756_), .C(new_n968_), .Y(new_n5772_));
  AOI21X1  g05580(.A0(new_n5772_), .A1(new_n5771_), .B0(new_n5766_), .Y(new_n5773_));
  OR2X1    g05581(.A(new_n5773_), .B(new_n902_), .Y(new_n5774_));
  AND2X1   g05582(.A(new_n5772_), .B(new_n5771_), .Y(new_n5775_));
  AND2X1   g05583(.A(new_n5431_), .B(new_n5430_), .Y(new_n5776_));
  NOR4X1   g05584(.A(new_n5541_), .B(new_n5776_), .C(new_n5398_), .D(new_n5429_), .Y(new_n5777_));
  AOI22X1  g05585(.A0(new_n5431_), .A1(new_n5430_), .B0(new_n5416_), .B1(\asqrt[53] ), .Y(new_n5778_));
  AOI21X1  g05586(.A0(new_n5778_), .A1(\asqrt[35] ), .B0(new_n5397_), .Y(new_n5779_));
  NOR2X1   g05587(.A(new_n5779_), .B(new_n5777_), .Y(new_n5780_));
  INVX1    g05588(.A(new_n5780_), .Y(new_n5781_));
  OR2X1    g05589(.A(new_n5766_), .B(\asqrt[54] ), .Y(new_n5782_));
  OAI21X1  g05590(.A0(new_n5782_), .A1(new_n5775_), .B0(new_n5781_), .Y(new_n5783_));
  AOI21X1  g05591(.A0(new_n5783_), .A1(new_n5774_), .B0(new_n697_), .Y(new_n5784_));
  AND2X1   g05592(.A(new_n5417_), .B(new_n5409_), .Y(new_n5785_));
  OR4X1    g05593(.A(new_n5541_), .B(new_n5785_), .C(new_n5434_), .D(new_n5410_), .Y(new_n5786_));
  OR2X1    g05594(.A(new_n5785_), .B(new_n5410_), .Y(new_n5787_));
  OAI21X1  g05595(.A0(new_n5787_), .A1(new_n5541_), .B0(new_n5434_), .Y(new_n5788_));
  AND2X1   g05596(.A(new_n5788_), .B(new_n5786_), .Y(new_n5789_));
  OR2X1    g05597(.A(new_n5763_), .B(new_n1277_), .Y(new_n5790_));
  AND2X1   g05598(.A(new_n5746_), .B(new_n5738_), .Y(new_n5791_));
  INVX1    g05599(.A(new_n5752_), .Y(new_n5792_));
  OR2X1    g05600(.A(new_n5753_), .B(\asqrt[51] ), .Y(new_n5793_));
  OAI21X1  g05601(.A0(new_n5793_), .A1(new_n5791_), .B0(new_n5792_), .Y(new_n5794_));
  AOI21X1  g05602(.A0(new_n5794_), .A1(new_n5790_), .B0(new_n1111_), .Y(new_n5795_));
  AOI21X1  g05603(.A0(new_n5736_), .A1(\asqrt[51] ), .B0(\asqrt[52] ), .Y(new_n5796_));
  AOI21X1  g05604(.A0(new_n5796_), .A1(new_n5794_), .B0(new_n5761_), .Y(new_n5797_));
  OAI21X1  g05605(.A0(new_n5797_), .A1(new_n5795_), .B0(\asqrt[53] ), .Y(new_n5798_));
  NOR3X1   g05606(.A(new_n5797_), .B(new_n5795_), .C(\asqrt[53] ), .Y(new_n5799_));
  OAI21X1  g05607(.A0(new_n5799_), .A1(new_n5770_), .B0(new_n5798_), .Y(new_n5800_));
  AOI21X1  g05608(.A0(new_n5800_), .A1(\asqrt[54] ), .B0(\asqrt[55] ), .Y(new_n5801_));
  AOI21X1  g05609(.A0(new_n5801_), .A1(new_n5783_), .B0(new_n5789_), .Y(new_n5802_));
  OAI21X1  g05610(.A0(new_n5802_), .A1(new_n5784_), .B0(\asqrt[56] ), .Y(new_n5803_));
  OR4X1    g05611(.A(new_n5541_), .B(new_n5425_), .C(new_n5428_), .D(new_n5452_), .Y(new_n5804_));
  NAND2X1  g05612(.A(new_n5437_), .B(new_n5419_), .Y(new_n5805_));
  OAI21X1  g05613(.A0(new_n5805_), .A1(new_n5541_), .B0(new_n5428_), .Y(new_n5806_));
  AND2X1   g05614(.A(new_n5806_), .B(new_n5804_), .Y(new_n5807_));
  NOR3X1   g05615(.A(new_n5802_), .B(new_n5784_), .C(\asqrt[56] ), .Y(new_n5808_));
  OAI21X1  g05616(.A0(new_n5808_), .A1(new_n5807_), .B0(new_n5803_), .Y(new_n5809_));
  AND2X1   g05617(.A(new_n5809_), .B(\asqrt[57] ), .Y(new_n5810_));
  OR2X1    g05618(.A(new_n5808_), .B(new_n5807_), .Y(new_n5811_));
  OAI21X1  g05619(.A0(new_n5476_), .A1(new_n5474_), .B0(new_n5443_), .Y(new_n5812_));
  NOR3X1   g05620(.A(new_n5812_), .B(new_n5541_), .C(new_n5427_), .Y(new_n5813_));
  AOI22X1  g05621(.A0(new_n5444_), .A1(new_n5438_), .B0(new_n5426_), .B1(\asqrt[56] ), .Y(new_n5814_));
  AOI21X1  g05622(.A0(new_n5814_), .A1(\asqrt[35] ), .B0(new_n5443_), .Y(new_n5815_));
  NOR2X1   g05623(.A(new_n5815_), .B(new_n5813_), .Y(new_n5816_));
  AND2X1   g05624(.A(new_n5803_), .B(new_n481_), .Y(new_n5817_));
  AOI21X1  g05625(.A0(new_n5817_), .A1(new_n5811_), .B0(new_n5816_), .Y(new_n5818_));
  OAI21X1  g05626(.A0(new_n5818_), .A1(new_n5810_), .B0(\asqrt[58] ), .Y(new_n5819_));
  AND2X1   g05627(.A(new_n5479_), .B(new_n5477_), .Y(new_n5820_));
  OR2X1    g05628(.A(new_n5451_), .B(new_n5478_), .Y(new_n5821_));
  OR2X1    g05629(.A(new_n5821_), .B(new_n5820_), .Y(new_n5822_));
  NOR3X1   g05630(.A(new_n5541_), .B(new_n5820_), .C(new_n5478_), .Y(new_n5823_));
  OAI22X1  g05631(.A0(new_n5823_), .A1(new_n5450_), .B0(new_n5822_), .B1(new_n5541_), .Y(new_n5824_));
  AND2X1   g05632(.A(new_n5800_), .B(\asqrt[54] ), .Y(new_n5825_));
  NAND2X1  g05633(.A(new_n5772_), .B(new_n5771_), .Y(new_n5826_));
  NOR2X1   g05634(.A(new_n5766_), .B(\asqrt[54] ), .Y(new_n5827_));
  AOI21X1  g05635(.A0(new_n5827_), .A1(new_n5826_), .B0(new_n5780_), .Y(new_n5828_));
  OAI21X1  g05636(.A0(new_n5828_), .A1(new_n5825_), .B0(\asqrt[55] ), .Y(new_n5829_));
  INVX1    g05637(.A(new_n5789_), .Y(new_n5830_));
  OAI21X1  g05638(.A0(new_n5773_), .A1(new_n902_), .B0(new_n697_), .Y(new_n5831_));
  OAI21X1  g05639(.A0(new_n5831_), .A1(new_n5828_), .B0(new_n5830_), .Y(new_n5832_));
  AOI21X1  g05640(.A0(new_n5832_), .A1(new_n5829_), .B0(new_n582_), .Y(new_n5833_));
  INVX1    g05641(.A(new_n5807_), .Y(new_n5834_));
  NAND3X1  g05642(.A(new_n5832_), .B(new_n5829_), .C(new_n582_), .Y(new_n5835_));
  AOI21X1  g05643(.A0(new_n5835_), .A1(new_n5834_), .B0(new_n5833_), .Y(new_n5836_));
  OAI21X1  g05644(.A0(new_n5836_), .A1(new_n481_), .B0(new_n399_), .Y(new_n5837_));
  OAI21X1  g05645(.A0(new_n5837_), .A1(new_n5818_), .B0(new_n5824_), .Y(new_n5838_));
  AOI21X1  g05646(.A0(new_n5838_), .A1(new_n5819_), .B0(new_n328_), .Y(new_n5839_));
  OR4X1    g05647(.A(new_n5541_), .B(new_n5489_), .C(new_n5462_), .D(new_n5456_), .Y(new_n5840_));
  OR2X1    g05648(.A(new_n5489_), .B(new_n5456_), .Y(new_n5841_));
  OAI21X1  g05649(.A0(new_n5841_), .A1(new_n5541_), .B0(new_n5462_), .Y(new_n5842_));
  AND2X1   g05650(.A(new_n5842_), .B(new_n5840_), .Y(new_n5843_));
  INVX1    g05651(.A(new_n5843_), .Y(new_n5844_));
  NAND3X1  g05652(.A(new_n5838_), .B(new_n5819_), .C(new_n328_), .Y(new_n5845_));
  AOI21X1  g05653(.A0(new_n5845_), .A1(new_n5844_), .B0(new_n5839_), .Y(new_n5846_));
  OR2X1    g05654(.A(new_n5846_), .B(new_n292_), .Y(new_n5847_));
  AND2X1   g05655(.A(new_n5845_), .B(new_n5844_), .Y(new_n5848_));
  AND2X1   g05656(.A(new_n5521_), .B(new_n5520_), .Y(new_n5849_));
  NOR4X1   g05657(.A(new_n5541_), .B(new_n5849_), .C(new_n5472_), .D(new_n5519_), .Y(new_n5850_));
  AOI22X1  g05658(.A0(new_n5521_), .A1(new_n5520_), .B0(new_n5490_), .B1(\asqrt[59] ), .Y(new_n5851_));
  AOI21X1  g05659(.A0(new_n5851_), .A1(\asqrt[35] ), .B0(new_n5471_), .Y(new_n5852_));
  NOR2X1   g05660(.A(new_n5852_), .B(new_n5850_), .Y(new_n5853_));
  INVX1    g05661(.A(new_n5853_), .Y(new_n5854_));
  OR2X1    g05662(.A(new_n5839_), .B(\asqrt[60] ), .Y(new_n5855_));
  OAI21X1  g05663(.A0(new_n5855_), .A1(new_n5848_), .B0(new_n5854_), .Y(new_n5856_));
  AOI21X1  g05664(.A0(new_n5856_), .A1(new_n5847_), .B0(new_n217_), .Y(new_n5857_));
  AND2X1   g05665(.A(new_n5491_), .B(new_n5483_), .Y(new_n5858_));
  OR4X1    g05666(.A(new_n5541_), .B(new_n5858_), .C(new_n5524_), .D(new_n5484_), .Y(new_n5859_));
  OR2X1    g05667(.A(new_n5858_), .B(new_n5484_), .Y(new_n5860_));
  OAI21X1  g05668(.A0(new_n5860_), .A1(new_n5541_), .B0(new_n5524_), .Y(new_n5861_));
  AND2X1   g05669(.A(new_n5861_), .B(new_n5859_), .Y(new_n5862_));
  OR2X1    g05670(.A(new_n5836_), .B(new_n481_), .Y(new_n5863_));
  AND2X1   g05671(.A(new_n5835_), .B(new_n5834_), .Y(new_n5864_));
  INVX1    g05672(.A(new_n5816_), .Y(new_n5865_));
  OR2X1    g05673(.A(new_n5833_), .B(\asqrt[57] ), .Y(new_n5866_));
  OAI21X1  g05674(.A0(new_n5866_), .A1(new_n5864_), .B0(new_n5865_), .Y(new_n5867_));
  AOI21X1  g05675(.A0(new_n5867_), .A1(new_n5863_), .B0(new_n399_), .Y(new_n5868_));
  INVX1    g05676(.A(new_n5824_), .Y(new_n5869_));
  AOI21X1  g05677(.A0(new_n5809_), .A1(\asqrt[57] ), .B0(\asqrt[58] ), .Y(new_n5870_));
  AOI21X1  g05678(.A0(new_n5870_), .A1(new_n5867_), .B0(new_n5869_), .Y(new_n5871_));
  OAI21X1  g05679(.A0(new_n5871_), .A1(new_n5868_), .B0(\asqrt[59] ), .Y(new_n5872_));
  NOR3X1   g05680(.A(new_n5871_), .B(new_n5868_), .C(\asqrt[59] ), .Y(new_n5873_));
  OAI21X1  g05681(.A0(new_n5873_), .A1(new_n5843_), .B0(new_n5872_), .Y(new_n5874_));
  AOI21X1  g05682(.A0(new_n5874_), .A1(\asqrt[60] ), .B0(\asqrt[61] ), .Y(new_n5875_));
  AOI21X1  g05683(.A0(new_n5875_), .A1(new_n5856_), .B0(new_n5862_), .Y(new_n5876_));
  OAI21X1  g05684(.A0(new_n5876_), .A1(new_n5857_), .B0(\asqrt[62] ), .Y(new_n5877_));
  NOR3X1   g05685(.A(new_n5876_), .B(new_n5857_), .C(\asqrt[62] ), .Y(new_n5878_));
  OR4X1    g05686(.A(new_n5541_), .B(new_n5529_), .C(new_n5494_), .D(new_n5527_), .Y(new_n5879_));
  OR2X1    g05687(.A(new_n5494_), .B(new_n5527_), .Y(new_n5880_));
  OAI21X1  g05688(.A0(new_n5880_), .A1(new_n5541_), .B0(new_n5529_), .Y(new_n5881_));
  AND2X1   g05689(.A(new_n5881_), .B(new_n5879_), .Y(new_n5882_));
  OAI21X1  g05690(.A0(new_n5882_), .A1(new_n5878_), .B0(new_n5877_), .Y(new_n5883_));
  AND2X1   g05691(.A(new_n5508_), .B(new_n5502_), .Y(new_n5884_));
  NOR4X1   g05692(.A(new_n5541_), .B(new_n5884_), .C(new_n5558_), .D(new_n5501_), .Y(new_n5885_));
  INVX1    g05693(.A(new_n5885_), .Y(new_n5886_));
  OAI22X1  g05694(.A0(new_n5559_), .A1(new_n5557_), .B0(new_n5530_), .B1(new_n199_), .Y(new_n5887_));
  OAI21X1  g05695(.A0(new_n5887_), .A1(new_n5541_), .B0(new_n5558_), .Y(new_n5888_));
  AND2X1   g05696(.A(new_n5888_), .B(new_n5886_), .Y(new_n5889_));
  INVX1    g05697(.A(new_n5889_), .Y(new_n5890_));
  AND2X1   g05698(.A(new_n5563_), .B(new_n5560_), .Y(new_n5891_));
  AOI21X1  g05699(.A0(new_n5560_), .A1(new_n5556_), .B0(new_n5513_), .Y(new_n5892_));
  AOI21X1  g05700(.A0(new_n5892_), .A1(\asqrt[35] ), .B0(new_n5891_), .Y(new_n5893_));
  AND2X1   g05701(.A(new_n5893_), .B(new_n5890_), .Y(new_n5894_));
  AOI21X1  g05702(.A0(new_n5894_), .A1(new_n5883_), .B0(\asqrt[63] ), .Y(new_n5895_));
  NOR2X1   g05703(.A(new_n5882_), .B(new_n5878_), .Y(new_n5896_));
  NAND2X1  g05704(.A(new_n5889_), .B(new_n5877_), .Y(new_n5897_));
  NAND2X1  g05705(.A(new_n5560_), .B(new_n5556_), .Y(new_n5898_));
  AOI21X1  g05706(.A0(\asqrt[35] ), .A1(new_n5514_), .B0(new_n5898_), .Y(new_n5899_));
  NOR3X1   g05707(.A(new_n5899_), .B(new_n5892_), .C(new_n193_), .Y(new_n5900_));
  AND2X1   g05708(.A(new_n5518_), .B(new_n193_), .Y(new_n5901_));
  AND2X1   g05709(.A(new_n5512_), .B(new_n5194_), .Y(new_n5902_));
  INVX1    g05710(.A(new_n5534_), .Y(new_n5903_));
  INVX1    g05711(.A(new_n5538_), .Y(new_n5904_));
  OR4X1    g05712(.A(new_n5904_), .B(new_n5903_), .C(new_n5902_), .D(new_n5511_), .Y(new_n5905_));
  NOR3X1   g05713(.A(new_n5905_), .B(new_n5891_), .C(new_n5901_), .Y(new_n5906_));
  NOR2X1   g05714(.A(new_n5906_), .B(new_n5900_), .Y(new_n5907_));
  OAI21X1  g05715(.A0(new_n5897_), .A1(new_n5896_), .B0(new_n5907_), .Y(new_n5908_));
  OR2X1    g05716(.A(new_n5908_), .B(new_n5895_), .Y(\asqrt[34] ));
  NOR2X1   g05717(.A(\a[67] ), .B(\a[66] ), .Y(new_n5910_));
  MX2X1    g05718(.A(new_n5910_), .B(\asqrt[34] ), .S0(\a[68] ), .Y(new_n5911_));
  INVX1    g05719(.A(\a[68] ), .Y(new_n5912_));
  AND2X1   g05720(.A(new_n5874_), .B(\asqrt[60] ), .Y(new_n5913_));
  NAND2X1  g05721(.A(new_n5845_), .B(new_n5844_), .Y(new_n5914_));
  NOR2X1   g05722(.A(new_n5839_), .B(\asqrt[60] ), .Y(new_n5915_));
  AOI21X1  g05723(.A0(new_n5915_), .A1(new_n5914_), .B0(new_n5853_), .Y(new_n5916_));
  OAI21X1  g05724(.A0(new_n5916_), .A1(new_n5913_), .B0(\asqrt[61] ), .Y(new_n5917_));
  INVX1    g05725(.A(new_n5862_), .Y(new_n5918_));
  OAI21X1  g05726(.A0(new_n5846_), .A1(new_n292_), .B0(new_n217_), .Y(new_n5919_));
  OAI21X1  g05727(.A0(new_n5919_), .A1(new_n5916_), .B0(new_n5918_), .Y(new_n5920_));
  AOI21X1  g05728(.A0(new_n5920_), .A1(new_n5917_), .B0(new_n199_), .Y(new_n5921_));
  NAND3X1  g05729(.A(new_n5920_), .B(new_n5917_), .C(new_n199_), .Y(new_n5922_));
  INVX1    g05730(.A(new_n5882_), .Y(new_n5923_));
  AOI21X1  g05731(.A0(new_n5923_), .A1(new_n5922_), .B0(new_n5921_), .Y(new_n5924_));
  INVX1    g05732(.A(new_n5894_), .Y(new_n5925_));
  OAI21X1  g05733(.A0(new_n5925_), .A1(new_n5924_), .B0(new_n193_), .Y(new_n5926_));
  OR2X1    g05734(.A(new_n5882_), .B(new_n5878_), .Y(new_n5927_));
  AND2X1   g05735(.A(new_n5889_), .B(new_n5877_), .Y(new_n5928_));
  INVX1    g05736(.A(new_n5907_), .Y(new_n5929_));
  AOI21X1  g05737(.A0(new_n5928_), .A1(new_n5927_), .B0(new_n5929_), .Y(new_n5930_));
  AOI21X1  g05738(.A0(new_n5930_), .A1(new_n5926_), .B0(new_n5912_), .Y(new_n5931_));
  NAND2X1  g05739(.A(new_n5910_), .B(new_n5912_), .Y(new_n5932_));
  NAND3X1  g05740(.A(new_n5932_), .B(new_n5538_), .C(new_n5534_), .Y(new_n5933_));
  OR4X1    g05741(.A(new_n5933_), .B(new_n5931_), .C(new_n5891_), .D(new_n5901_), .Y(new_n5934_));
  OAI21X1  g05742(.A0(new_n5908_), .A1(new_n5895_), .B0(new_n5912_), .Y(new_n5935_));
  AOI21X1  g05743(.A0(new_n5930_), .A1(new_n5926_), .B0(new_n5543_), .Y(new_n5936_));
  AOI21X1  g05744(.A0(new_n5935_), .A1(\a[69] ), .B0(new_n5936_), .Y(new_n5937_));
  AOI22X1  g05745(.A0(new_n5937_), .A1(new_n5934_), .B0(new_n5911_), .B1(\asqrt[35] ), .Y(new_n5938_));
  OR2X1    g05746(.A(new_n5938_), .B(new_n5176_), .Y(new_n5939_));
  AND2X1   g05747(.A(new_n5937_), .B(new_n5934_), .Y(new_n5940_));
  NOR2X1   g05748(.A(new_n5908_), .B(new_n5895_), .Y(new_n5941_));
  INVX1    g05749(.A(new_n5910_), .Y(new_n5942_));
  MX2X1    g05750(.A(new_n5942_), .B(new_n5941_), .S0(\a[68] ), .Y(new_n5943_));
  OAI21X1  g05751(.A0(new_n5943_), .A1(new_n5541_), .B0(new_n5176_), .Y(new_n5944_));
  OAI21X1  g05752(.A0(new_n5908_), .A1(new_n5895_), .B0(new_n5542_), .Y(new_n5945_));
  AND2X1   g05753(.A(new_n5928_), .B(new_n5927_), .Y(new_n5946_));
  OR2X1    g05754(.A(new_n5906_), .B(new_n5541_), .Y(new_n5947_));
  OR4X1    g05755(.A(new_n5947_), .B(new_n5900_), .C(new_n5946_), .D(new_n5895_), .Y(new_n5948_));
  AOI21X1  g05756(.A0(new_n5948_), .A1(new_n5945_), .B0(new_n5546_), .Y(new_n5949_));
  NOR4X1   g05757(.A(new_n5947_), .B(new_n5900_), .C(new_n5946_), .D(new_n5895_), .Y(new_n5950_));
  NOR3X1   g05758(.A(new_n5950_), .B(new_n5936_), .C(\a[70] ), .Y(new_n5951_));
  OR2X1    g05759(.A(new_n5951_), .B(new_n5949_), .Y(new_n5952_));
  OAI21X1  g05760(.A0(new_n5944_), .A1(new_n5940_), .B0(new_n5952_), .Y(new_n5953_));
  AOI21X1  g05761(.A0(new_n5953_), .A1(new_n5939_), .B0(new_n4826_), .Y(new_n5954_));
  AND2X1   g05762(.A(new_n5553_), .B(new_n5552_), .Y(new_n5955_));
  NOR3X1   g05763(.A(new_n5955_), .B(new_n5590_), .C(new_n5589_), .Y(new_n5956_));
  OAI21X1  g05764(.A0(new_n5908_), .A1(new_n5895_), .B0(new_n5956_), .Y(new_n5957_));
  NAND3X1  g05765(.A(\asqrt[34] ), .B(new_n5551_), .C(new_n5545_), .Y(new_n5958_));
  NAND2X1  g05766(.A(new_n5958_), .B(new_n5955_), .Y(new_n5959_));
  NOR4X1   g05767(.A(new_n5933_), .B(new_n5931_), .C(new_n5891_), .D(new_n5901_), .Y(new_n5960_));
  INVX1    g05768(.A(\a[69] ), .Y(new_n5961_));
  AOI21X1  g05769(.A0(new_n5930_), .A1(new_n5926_), .B0(\a[68] ), .Y(new_n5962_));
  OAI21X1  g05770(.A0(new_n5962_), .A1(new_n5961_), .B0(new_n5945_), .Y(new_n5963_));
  OAI22X1  g05771(.A0(new_n5963_), .A1(new_n5960_), .B0(new_n5943_), .B1(new_n5541_), .Y(new_n5964_));
  AOI21X1  g05772(.A0(new_n5964_), .A1(\asqrt[36] ), .B0(\asqrt[37] ), .Y(new_n5965_));
  AOI22X1  g05773(.A0(new_n5965_), .A1(new_n5953_), .B0(new_n5959_), .B1(new_n5957_), .Y(new_n5966_));
  OAI21X1  g05774(.A0(new_n5966_), .A1(new_n5954_), .B0(\asqrt[38] ), .Y(new_n5967_));
  AND2X1   g05775(.A(new_n5568_), .B(new_n5554_), .Y(new_n5968_));
  NOR3X1   g05776(.A(new_n5596_), .B(new_n5968_), .C(new_n5555_), .Y(new_n5969_));
  NOR2X1   g05777(.A(new_n5968_), .B(new_n5555_), .Y(new_n5970_));
  OAI21X1  g05778(.A0(new_n5908_), .A1(new_n5895_), .B0(new_n5970_), .Y(new_n5971_));
  AOI22X1  g05779(.A0(new_n5971_), .A1(new_n5596_), .B0(new_n5969_), .B1(\asqrt[34] ), .Y(new_n5972_));
  NOR3X1   g05780(.A(new_n5966_), .B(new_n5954_), .C(\asqrt[38] ), .Y(new_n5973_));
  OAI21X1  g05781(.A0(new_n5973_), .A1(new_n5972_), .B0(new_n5967_), .Y(new_n5974_));
  AND2X1   g05782(.A(new_n5974_), .B(\asqrt[39] ), .Y(new_n5975_));
  OR2X1    g05783(.A(new_n5973_), .B(new_n5972_), .Y(new_n5976_));
  NOR3X1   g05784(.A(new_n5585_), .B(new_n5588_), .C(new_n5606_), .Y(new_n5977_));
  OAI21X1  g05785(.A0(new_n5908_), .A1(new_n5895_), .B0(new_n5977_), .Y(new_n5978_));
  NOR3X1   g05786(.A(new_n5941_), .B(new_n5585_), .C(new_n5606_), .Y(new_n5979_));
  OR2X1    g05787(.A(new_n5979_), .B(new_n5584_), .Y(new_n5980_));
  AND2X1   g05788(.A(new_n5980_), .B(new_n5978_), .Y(new_n5981_));
  AND2X1   g05789(.A(new_n5964_), .B(\asqrt[36] ), .Y(new_n5982_));
  NAND2X1  g05790(.A(new_n5937_), .B(new_n5934_), .Y(new_n5983_));
  AOI21X1  g05791(.A0(new_n5911_), .A1(\asqrt[35] ), .B0(\asqrt[36] ), .Y(new_n5984_));
  NOR2X1   g05792(.A(new_n5951_), .B(new_n5949_), .Y(new_n5985_));
  AOI21X1  g05793(.A0(new_n5984_), .A1(new_n5983_), .B0(new_n5985_), .Y(new_n5986_));
  OAI21X1  g05794(.A0(new_n5986_), .A1(new_n5982_), .B0(\asqrt[37] ), .Y(new_n5987_));
  NAND2X1  g05795(.A(new_n5959_), .B(new_n5957_), .Y(new_n5988_));
  OAI21X1  g05796(.A0(new_n5938_), .A1(new_n5176_), .B0(new_n4826_), .Y(new_n5989_));
  OAI21X1  g05797(.A0(new_n5989_), .A1(new_n5986_), .B0(new_n5988_), .Y(new_n5990_));
  AOI21X1  g05798(.A0(new_n5990_), .A1(new_n5987_), .B0(new_n4493_), .Y(new_n5991_));
  NOR2X1   g05799(.A(new_n5991_), .B(\asqrt[39] ), .Y(new_n5992_));
  AOI21X1  g05800(.A0(new_n5992_), .A1(new_n5976_), .B0(new_n5981_), .Y(new_n5993_));
  OAI21X1  g05801(.A0(new_n5993_), .A1(new_n5975_), .B0(\asqrt[40] ), .Y(new_n5994_));
  AOI21X1  g05802(.A0(new_n5607_), .A1(new_n5599_), .B0(new_n5643_), .Y(new_n5995_));
  AND2X1   g05803(.A(new_n5995_), .B(new_n5641_), .Y(new_n5996_));
  AOI22X1  g05804(.A0(new_n5607_), .A1(new_n5599_), .B0(new_n5586_), .B1(\asqrt[39] ), .Y(new_n5997_));
  AOI21X1  g05805(.A0(new_n5997_), .A1(\asqrt[34] ), .B0(new_n5605_), .Y(new_n5998_));
  AOI21X1  g05806(.A0(new_n5996_), .A1(\asqrt[34] ), .B0(new_n5998_), .Y(new_n5999_));
  INVX1    g05807(.A(new_n5999_), .Y(new_n6000_));
  INVX1    g05808(.A(new_n5972_), .Y(new_n6001_));
  NAND3X1  g05809(.A(new_n5990_), .B(new_n5987_), .C(new_n4493_), .Y(new_n6002_));
  AOI21X1  g05810(.A0(new_n6002_), .A1(new_n6001_), .B0(new_n5991_), .Y(new_n6003_));
  OAI21X1  g05811(.A0(new_n6003_), .A1(new_n4165_), .B0(new_n3863_), .Y(new_n6004_));
  OAI21X1  g05812(.A0(new_n6004_), .A1(new_n5993_), .B0(new_n6000_), .Y(new_n6005_));
  AOI21X1  g05813(.A0(new_n6005_), .A1(new_n5994_), .B0(new_n3564_), .Y(new_n6006_));
  AND2X1   g05814(.A(new_n5647_), .B(new_n5645_), .Y(new_n6007_));
  NOR3X1   g05815(.A(new_n6007_), .B(new_n5615_), .C(new_n5646_), .Y(new_n6008_));
  NOR2X1   g05816(.A(new_n6007_), .B(new_n5646_), .Y(new_n6009_));
  AOI21X1  g05817(.A0(new_n6009_), .A1(\asqrt[34] ), .B0(new_n5614_), .Y(new_n6010_));
  AOI21X1  g05818(.A0(new_n6008_), .A1(\asqrt[34] ), .B0(new_n6010_), .Y(new_n6011_));
  INVX1    g05819(.A(new_n6011_), .Y(new_n6012_));
  NAND3X1  g05820(.A(new_n6005_), .B(new_n5994_), .C(new_n3564_), .Y(new_n6013_));
  AOI21X1  g05821(.A0(new_n6013_), .A1(new_n6012_), .B0(new_n6006_), .Y(new_n6014_));
  OR2X1    g05822(.A(new_n6014_), .B(new_n3276_), .Y(new_n6015_));
  OR2X1    g05823(.A(new_n6003_), .B(new_n4165_), .Y(new_n6016_));
  NOR2X1   g05824(.A(new_n5973_), .B(new_n5972_), .Y(new_n6017_));
  INVX1    g05825(.A(new_n5981_), .Y(new_n6018_));
  OR2X1    g05826(.A(new_n5991_), .B(\asqrt[39] ), .Y(new_n6019_));
  OAI21X1  g05827(.A0(new_n6019_), .A1(new_n6017_), .B0(new_n6018_), .Y(new_n6020_));
  AOI21X1  g05828(.A0(new_n6020_), .A1(new_n6016_), .B0(new_n3863_), .Y(new_n6021_));
  AOI21X1  g05829(.A0(new_n5974_), .A1(\asqrt[39] ), .B0(\asqrt[40] ), .Y(new_n6022_));
  AOI21X1  g05830(.A0(new_n6022_), .A1(new_n6020_), .B0(new_n5999_), .Y(new_n6023_));
  NOR3X1   g05831(.A(new_n6023_), .B(new_n6021_), .C(\asqrt[41] ), .Y(new_n6024_));
  NOR2X1   g05832(.A(new_n6024_), .B(new_n6011_), .Y(new_n6025_));
  OR4X1    g05833(.A(new_n5941_), .B(new_n5651_), .C(new_n5622_), .D(new_n5619_), .Y(new_n6026_));
  NAND2X1  g05834(.A(new_n5623_), .B(new_n5649_), .Y(new_n6027_));
  OAI21X1  g05835(.A0(new_n6027_), .A1(new_n5941_), .B0(new_n5622_), .Y(new_n6028_));
  AND2X1   g05836(.A(new_n6028_), .B(new_n6026_), .Y(new_n6029_));
  INVX1    g05837(.A(new_n6029_), .Y(new_n6030_));
  OAI21X1  g05838(.A0(new_n6023_), .A1(new_n6021_), .B0(\asqrt[41] ), .Y(new_n6031_));
  NAND2X1  g05839(.A(new_n6031_), .B(new_n3276_), .Y(new_n6032_));
  OAI21X1  g05840(.A0(new_n6032_), .A1(new_n6025_), .B0(new_n6030_), .Y(new_n6033_));
  AOI21X1  g05841(.A0(new_n6033_), .A1(new_n6015_), .B0(new_n3008_), .Y(new_n6034_));
  AND2X1   g05842(.A(new_n5666_), .B(new_n5665_), .Y(new_n6035_));
  NOR3X1   g05843(.A(new_n6035_), .B(new_n5632_), .C(new_n5664_), .Y(new_n6036_));
  AOI22X1  g05844(.A0(new_n5666_), .A1(new_n5665_), .B0(new_n5652_), .B1(\asqrt[42] ), .Y(new_n6037_));
  AOI21X1  g05845(.A0(new_n6037_), .A1(\asqrt[34] ), .B0(new_n5631_), .Y(new_n6038_));
  AOI21X1  g05846(.A0(new_n6036_), .A1(\asqrt[34] ), .B0(new_n6038_), .Y(new_n6039_));
  OAI21X1  g05847(.A0(new_n6024_), .A1(new_n6011_), .B0(new_n6031_), .Y(new_n6040_));
  AOI21X1  g05848(.A0(new_n6040_), .A1(\asqrt[42] ), .B0(\asqrt[43] ), .Y(new_n6041_));
  AOI21X1  g05849(.A0(new_n6041_), .A1(new_n6033_), .B0(new_n6039_), .Y(new_n6042_));
  OAI21X1  g05850(.A0(new_n6042_), .A1(new_n6034_), .B0(\asqrt[44] ), .Y(new_n6043_));
  AND2X1   g05851(.A(new_n5653_), .B(new_n5634_), .Y(new_n6044_));
  NOR3X1   g05852(.A(new_n6044_), .B(new_n5669_), .C(new_n5635_), .Y(new_n6045_));
  NOR2X1   g05853(.A(new_n6044_), .B(new_n5635_), .Y(new_n6046_));
  AOI21X1  g05854(.A0(new_n6046_), .A1(\asqrt[34] ), .B0(new_n5640_), .Y(new_n6047_));
  AOI21X1  g05855(.A0(new_n6045_), .A1(\asqrt[34] ), .B0(new_n6047_), .Y(new_n6048_));
  NOR3X1   g05856(.A(new_n6042_), .B(new_n6034_), .C(\asqrt[44] ), .Y(new_n6049_));
  OAI21X1  g05857(.A0(new_n6049_), .A1(new_n6048_), .B0(new_n6043_), .Y(new_n6050_));
  AND2X1   g05858(.A(new_n6050_), .B(\asqrt[45] ), .Y(new_n6051_));
  INVX1    g05859(.A(new_n6048_), .Y(new_n6052_));
  AND2X1   g05860(.A(new_n6040_), .B(\asqrt[42] ), .Y(new_n6053_));
  OR2X1    g05861(.A(new_n6024_), .B(new_n6011_), .Y(new_n6054_));
  AND2X1   g05862(.A(new_n6031_), .B(new_n3276_), .Y(new_n6055_));
  AOI21X1  g05863(.A0(new_n6055_), .A1(new_n6054_), .B0(new_n6029_), .Y(new_n6056_));
  OAI21X1  g05864(.A0(new_n6056_), .A1(new_n6053_), .B0(\asqrt[43] ), .Y(new_n6057_));
  INVX1    g05865(.A(new_n6039_), .Y(new_n6058_));
  OAI21X1  g05866(.A0(new_n6014_), .A1(new_n3276_), .B0(new_n3008_), .Y(new_n6059_));
  OAI21X1  g05867(.A0(new_n6059_), .A1(new_n6056_), .B0(new_n6058_), .Y(new_n6060_));
  NAND3X1  g05868(.A(new_n6060_), .B(new_n6057_), .C(new_n2769_), .Y(new_n6061_));
  NAND2X1  g05869(.A(new_n6061_), .B(new_n6052_), .Y(new_n6062_));
  NAND4X1  g05870(.A(\asqrt[34] ), .B(new_n5672_), .C(new_n5659_), .D(new_n5655_), .Y(new_n6063_));
  NAND2X1  g05871(.A(new_n5672_), .B(new_n5655_), .Y(new_n6064_));
  OAI21X1  g05872(.A0(new_n6064_), .A1(new_n5941_), .B0(new_n5663_), .Y(new_n6065_));
  AND2X1   g05873(.A(new_n6065_), .B(new_n6063_), .Y(new_n6066_));
  AOI21X1  g05874(.A0(new_n6060_), .A1(new_n6057_), .B0(new_n2769_), .Y(new_n6067_));
  NOR2X1   g05875(.A(new_n6067_), .B(\asqrt[45] ), .Y(new_n6068_));
  AOI21X1  g05876(.A0(new_n6068_), .A1(new_n6062_), .B0(new_n6066_), .Y(new_n6069_));
  OAI21X1  g05877(.A0(new_n6069_), .A1(new_n6051_), .B0(\asqrt[46] ), .Y(new_n6070_));
  AOI21X1  g05878(.A0(new_n5680_), .A1(new_n5673_), .B0(new_n5719_), .Y(new_n6071_));
  AND2X1   g05879(.A(new_n6071_), .B(new_n5717_), .Y(new_n6072_));
  AOI22X1  g05880(.A0(new_n5680_), .A1(new_n5673_), .B0(new_n5661_), .B1(\asqrt[45] ), .Y(new_n6073_));
  AOI21X1  g05881(.A0(new_n6073_), .A1(\asqrt[34] ), .B0(new_n5678_), .Y(new_n6074_));
  AOI21X1  g05882(.A0(new_n6072_), .A1(\asqrt[34] ), .B0(new_n6074_), .Y(new_n6075_));
  INVX1    g05883(.A(new_n6075_), .Y(new_n6076_));
  AOI21X1  g05884(.A0(new_n6061_), .A1(new_n6052_), .B0(new_n6067_), .Y(new_n6077_));
  OAI21X1  g05885(.A0(new_n6077_), .A1(new_n2570_), .B0(new_n2263_), .Y(new_n6078_));
  OAI21X1  g05886(.A0(new_n6078_), .A1(new_n6069_), .B0(new_n6076_), .Y(new_n6079_));
  AOI21X1  g05887(.A0(new_n6079_), .A1(new_n6070_), .B0(new_n2040_), .Y(new_n6080_));
  AND2X1   g05888(.A(new_n5723_), .B(new_n5721_), .Y(new_n6081_));
  NOR3X1   g05889(.A(new_n6081_), .B(new_n5688_), .C(new_n5722_), .Y(new_n6082_));
  NOR2X1   g05890(.A(new_n6081_), .B(new_n5722_), .Y(new_n6083_));
  AOI21X1  g05891(.A0(new_n6083_), .A1(\asqrt[34] ), .B0(new_n5687_), .Y(new_n6084_));
  AOI21X1  g05892(.A0(new_n6082_), .A1(\asqrt[34] ), .B0(new_n6084_), .Y(new_n6085_));
  INVX1    g05893(.A(new_n6085_), .Y(new_n6086_));
  NAND3X1  g05894(.A(new_n6079_), .B(new_n6070_), .C(new_n2040_), .Y(new_n6087_));
  AOI21X1  g05895(.A0(new_n6087_), .A1(new_n6086_), .B0(new_n6080_), .Y(new_n6088_));
  OR2X1    g05896(.A(new_n6088_), .B(new_n1834_), .Y(new_n6089_));
  OR2X1    g05897(.A(new_n6077_), .B(new_n2570_), .Y(new_n6090_));
  AND2X1   g05898(.A(new_n6061_), .B(new_n6052_), .Y(new_n6091_));
  INVX1    g05899(.A(new_n6066_), .Y(new_n6092_));
  OR2X1    g05900(.A(new_n6067_), .B(\asqrt[45] ), .Y(new_n6093_));
  OAI21X1  g05901(.A0(new_n6093_), .A1(new_n6091_), .B0(new_n6092_), .Y(new_n6094_));
  AOI21X1  g05902(.A0(new_n6094_), .A1(new_n6090_), .B0(new_n2263_), .Y(new_n6095_));
  AOI21X1  g05903(.A0(new_n6050_), .A1(\asqrt[45] ), .B0(\asqrt[46] ), .Y(new_n6096_));
  AOI21X1  g05904(.A0(new_n6096_), .A1(new_n6094_), .B0(new_n6075_), .Y(new_n6097_));
  NOR3X1   g05905(.A(new_n6097_), .B(new_n6095_), .C(\asqrt[47] ), .Y(new_n6098_));
  NOR2X1   g05906(.A(new_n6098_), .B(new_n6085_), .Y(new_n6099_));
  NAND4X1  g05907(.A(\asqrt[34] ), .B(new_n5698_), .C(new_n5696_), .D(new_n5725_), .Y(new_n6100_));
  NAND2X1  g05908(.A(new_n5698_), .B(new_n5725_), .Y(new_n6101_));
  OAI21X1  g05909(.A0(new_n6101_), .A1(new_n5941_), .B0(new_n5697_), .Y(new_n6102_));
  AND2X1   g05910(.A(new_n6102_), .B(new_n6100_), .Y(new_n6103_));
  INVX1    g05911(.A(new_n6103_), .Y(new_n6104_));
  OR2X1    g05912(.A(new_n6080_), .B(\asqrt[48] ), .Y(new_n6105_));
  OAI21X1  g05913(.A0(new_n6105_), .A1(new_n6099_), .B0(new_n6104_), .Y(new_n6106_));
  AOI21X1  g05914(.A0(new_n6106_), .A1(new_n6089_), .B0(new_n1632_), .Y(new_n6107_));
  AND2X1   g05915(.A(new_n5741_), .B(new_n5740_), .Y(new_n6108_));
  NOR3X1   g05916(.A(new_n6108_), .B(new_n5707_), .C(new_n5739_), .Y(new_n6109_));
  AOI22X1  g05917(.A0(new_n5741_), .A1(new_n5740_), .B0(new_n5727_), .B1(\asqrt[48] ), .Y(new_n6110_));
  AOI21X1  g05918(.A0(new_n6110_), .A1(\asqrt[34] ), .B0(new_n5706_), .Y(new_n6111_));
  AOI21X1  g05919(.A0(new_n6109_), .A1(\asqrt[34] ), .B0(new_n6111_), .Y(new_n6112_));
  OAI21X1  g05920(.A0(new_n6097_), .A1(new_n6095_), .B0(\asqrt[47] ), .Y(new_n6113_));
  OAI21X1  g05921(.A0(new_n6098_), .A1(new_n6085_), .B0(new_n6113_), .Y(new_n6114_));
  AOI21X1  g05922(.A0(new_n6114_), .A1(\asqrt[48] ), .B0(\asqrt[49] ), .Y(new_n6115_));
  AOI21X1  g05923(.A0(new_n6115_), .A1(new_n6106_), .B0(new_n6112_), .Y(new_n6116_));
  OAI21X1  g05924(.A0(new_n6116_), .A1(new_n6107_), .B0(\asqrt[50] ), .Y(new_n6117_));
  AND2X1   g05925(.A(new_n5728_), .B(new_n5709_), .Y(new_n6118_));
  NOR3X1   g05926(.A(new_n6118_), .B(new_n5715_), .C(new_n5710_), .Y(new_n6119_));
  NOR2X1   g05927(.A(new_n6118_), .B(new_n5710_), .Y(new_n6120_));
  AOI21X1  g05928(.A0(new_n6120_), .A1(\asqrt[34] ), .B0(new_n5716_), .Y(new_n6121_));
  AOI21X1  g05929(.A0(new_n6119_), .A1(\asqrt[34] ), .B0(new_n6121_), .Y(new_n6122_));
  NOR3X1   g05930(.A(new_n6116_), .B(new_n6107_), .C(\asqrt[50] ), .Y(new_n6123_));
  OAI21X1  g05931(.A0(new_n6123_), .A1(new_n6122_), .B0(new_n6117_), .Y(new_n6124_));
  AND2X1   g05932(.A(new_n6124_), .B(\asqrt[51] ), .Y(new_n6125_));
  OR2X1    g05933(.A(new_n6123_), .B(new_n6122_), .Y(new_n6126_));
  NAND4X1  g05934(.A(\asqrt[34] ), .B(new_n5746_), .C(new_n5734_), .D(new_n5730_), .Y(new_n6127_));
  NAND2X1  g05935(.A(new_n5746_), .B(new_n5730_), .Y(new_n6128_));
  OAI21X1  g05936(.A0(new_n6128_), .A1(new_n5941_), .B0(new_n5738_), .Y(new_n6129_));
  AND2X1   g05937(.A(new_n6129_), .B(new_n6127_), .Y(new_n6130_));
  AND2X1   g05938(.A(new_n6114_), .B(\asqrt[48] ), .Y(new_n6131_));
  OR2X1    g05939(.A(new_n6098_), .B(new_n6085_), .Y(new_n6132_));
  NOR2X1   g05940(.A(new_n6080_), .B(\asqrt[48] ), .Y(new_n6133_));
  AOI21X1  g05941(.A0(new_n6133_), .A1(new_n6132_), .B0(new_n6103_), .Y(new_n6134_));
  OAI21X1  g05942(.A0(new_n6134_), .A1(new_n6131_), .B0(\asqrt[49] ), .Y(new_n6135_));
  INVX1    g05943(.A(new_n6112_), .Y(new_n6136_));
  OAI21X1  g05944(.A0(new_n6088_), .A1(new_n1834_), .B0(new_n1632_), .Y(new_n6137_));
  OAI21X1  g05945(.A0(new_n6137_), .A1(new_n6134_), .B0(new_n6136_), .Y(new_n6138_));
  AOI21X1  g05946(.A0(new_n6138_), .A1(new_n6135_), .B0(new_n1469_), .Y(new_n6139_));
  NOR2X1   g05947(.A(new_n6139_), .B(\asqrt[51] ), .Y(new_n6140_));
  AOI21X1  g05948(.A0(new_n6140_), .A1(new_n6126_), .B0(new_n6130_), .Y(new_n6141_));
  OAI21X1  g05949(.A0(new_n6141_), .A1(new_n6125_), .B0(\asqrt[52] ), .Y(new_n6142_));
  AOI21X1  g05950(.A0(new_n5754_), .A1(new_n5747_), .B0(new_n5792_), .Y(new_n6143_));
  AND2X1   g05951(.A(new_n6143_), .B(new_n5790_), .Y(new_n6144_));
  AOI22X1  g05952(.A0(new_n5754_), .A1(new_n5747_), .B0(new_n5736_), .B1(\asqrt[51] ), .Y(new_n6145_));
  AOI21X1  g05953(.A0(new_n6145_), .A1(\asqrt[34] ), .B0(new_n5752_), .Y(new_n6146_));
  AOI21X1  g05954(.A0(new_n6144_), .A1(\asqrt[34] ), .B0(new_n6146_), .Y(new_n6147_));
  INVX1    g05955(.A(new_n6147_), .Y(new_n6148_));
  INVX1    g05956(.A(new_n6122_), .Y(new_n6149_));
  NAND3X1  g05957(.A(new_n6138_), .B(new_n6135_), .C(new_n1469_), .Y(new_n6150_));
  AOI21X1  g05958(.A0(new_n6150_), .A1(new_n6149_), .B0(new_n6139_), .Y(new_n6151_));
  OAI21X1  g05959(.A0(new_n6151_), .A1(new_n1277_), .B0(new_n1111_), .Y(new_n6152_));
  OAI21X1  g05960(.A0(new_n6152_), .A1(new_n6141_), .B0(new_n6148_), .Y(new_n6153_));
  AOI21X1  g05961(.A0(new_n6153_), .A1(new_n6142_), .B0(new_n968_), .Y(new_n6154_));
  AND2X1   g05962(.A(new_n5796_), .B(new_n5794_), .Y(new_n6155_));
  NOR3X1   g05963(.A(new_n6155_), .B(new_n5762_), .C(new_n5795_), .Y(new_n6156_));
  NOR2X1   g05964(.A(new_n6155_), .B(new_n5795_), .Y(new_n6157_));
  AOI21X1  g05965(.A0(new_n6157_), .A1(\asqrt[34] ), .B0(new_n5761_), .Y(new_n6158_));
  AOI21X1  g05966(.A0(new_n6156_), .A1(\asqrt[34] ), .B0(new_n6158_), .Y(new_n6159_));
  INVX1    g05967(.A(new_n6159_), .Y(new_n6160_));
  NAND3X1  g05968(.A(new_n6153_), .B(new_n6142_), .C(new_n968_), .Y(new_n6161_));
  AOI21X1  g05969(.A0(new_n6161_), .A1(new_n6160_), .B0(new_n6154_), .Y(new_n6162_));
  OR2X1    g05970(.A(new_n6162_), .B(new_n902_), .Y(new_n6163_));
  OR2X1    g05971(.A(new_n6151_), .B(new_n1277_), .Y(new_n6164_));
  NOR2X1   g05972(.A(new_n6123_), .B(new_n6122_), .Y(new_n6165_));
  INVX1    g05973(.A(new_n6130_), .Y(new_n6166_));
  OR2X1    g05974(.A(new_n6139_), .B(\asqrt[51] ), .Y(new_n6167_));
  OAI21X1  g05975(.A0(new_n6167_), .A1(new_n6165_), .B0(new_n6166_), .Y(new_n6168_));
  AOI21X1  g05976(.A0(new_n6168_), .A1(new_n6164_), .B0(new_n1111_), .Y(new_n6169_));
  AOI21X1  g05977(.A0(new_n6124_), .A1(\asqrt[51] ), .B0(\asqrt[52] ), .Y(new_n6170_));
  AOI21X1  g05978(.A0(new_n6170_), .A1(new_n6168_), .B0(new_n6147_), .Y(new_n6171_));
  NOR3X1   g05979(.A(new_n6171_), .B(new_n6169_), .C(\asqrt[53] ), .Y(new_n6172_));
  NOR2X1   g05980(.A(new_n6172_), .B(new_n6159_), .Y(new_n6173_));
  NAND4X1  g05981(.A(\asqrt[34] ), .B(new_n5772_), .C(new_n5770_), .D(new_n5798_), .Y(new_n6174_));
  NAND2X1  g05982(.A(new_n5772_), .B(new_n5798_), .Y(new_n6175_));
  OAI21X1  g05983(.A0(new_n6175_), .A1(new_n5941_), .B0(new_n5771_), .Y(new_n6176_));
  AND2X1   g05984(.A(new_n6176_), .B(new_n6174_), .Y(new_n6177_));
  INVX1    g05985(.A(new_n6177_), .Y(new_n6178_));
  OAI21X1  g05986(.A0(new_n6171_), .A1(new_n6169_), .B0(\asqrt[53] ), .Y(new_n6179_));
  NAND2X1  g05987(.A(new_n6179_), .B(new_n902_), .Y(new_n6180_));
  OAI21X1  g05988(.A0(new_n6180_), .A1(new_n6173_), .B0(new_n6178_), .Y(new_n6181_));
  AOI21X1  g05989(.A0(new_n6181_), .A1(new_n6163_), .B0(new_n697_), .Y(new_n6182_));
  AND2X1   g05990(.A(new_n5827_), .B(new_n5826_), .Y(new_n6183_));
  NOR3X1   g05991(.A(new_n6183_), .B(new_n5781_), .C(new_n5825_), .Y(new_n6184_));
  AOI22X1  g05992(.A0(new_n5827_), .A1(new_n5826_), .B0(new_n5800_), .B1(\asqrt[54] ), .Y(new_n6185_));
  AOI21X1  g05993(.A0(new_n6185_), .A1(\asqrt[34] ), .B0(new_n5780_), .Y(new_n6186_));
  AOI21X1  g05994(.A0(new_n6184_), .A1(\asqrt[34] ), .B0(new_n6186_), .Y(new_n6187_));
  OAI21X1  g05995(.A0(new_n6172_), .A1(new_n6159_), .B0(new_n6179_), .Y(new_n6188_));
  AOI21X1  g05996(.A0(new_n6188_), .A1(\asqrt[54] ), .B0(\asqrt[55] ), .Y(new_n6189_));
  AOI21X1  g05997(.A0(new_n6189_), .A1(new_n6181_), .B0(new_n6187_), .Y(new_n6190_));
  OAI21X1  g05998(.A0(new_n6190_), .A1(new_n6182_), .B0(\asqrt[56] ), .Y(new_n6191_));
  AND2X1   g05999(.A(new_n5801_), .B(new_n5783_), .Y(new_n6192_));
  NOR3X1   g06000(.A(new_n6192_), .B(new_n5830_), .C(new_n5784_), .Y(new_n6193_));
  NOR2X1   g06001(.A(new_n6192_), .B(new_n5784_), .Y(new_n6194_));
  AOI21X1  g06002(.A0(new_n6194_), .A1(\asqrt[34] ), .B0(new_n5789_), .Y(new_n6195_));
  AOI21X1  g06003(.A0(new_n6193_), .A1(\asqrt[34] ), .B0(new_n6195_), .Y(new_n6196_));
  NOR3X1   g06004(.A(new_n6190_), .B(new_n6182_), .C(\asqrt[56] ), .Y(new_n6197_));
  OAI21X1  g06005(.A0(new_n6197_), .A1(new_n6196_), .B0(new_n6191_), .Y(new_n6198_));
  AND2X1   g06006(.A(new_n6198_), .B(\asqrt[57] ), .Y(new_n6199_));
  OR2X1    g06007(.A(new_n6197_), .B(new_n6196_), .Y(new_n6200_));
  OR4X1    g06008(.A(new_n5941_), .B(new_n5808_), .C(new_n5834_), .D(new_n5833_), .Y(new_n6201_));
  OR2X1    g06009(.A(new_n5808_), .B(new_n5833_), .Y(new_n6202_));
  OAI21X1  g06010(.A0(new_n6202_), .A1(new_n5941_), .B0(new_n5834_), .Y(new_n6203_));
  AND2X1   g06011(.A(new_n6203_), .B(new_n6201_), .Y(new_n6204_));
  AND2X1   g06012(.A(new_n6191_), .B(new_n481_), .Y(new_n6205_));
  AOI21X1  g06013(.A0(new_n6205_), .A1(new_n6200_), .B0(new_n6204_), .Y(new_n6206_));
  OAI21X1  g06014(.A0(new_n6206_), .A1(new_n6199_), .B0(\asqrt[58] ), .Y(new_n6207_));
  AOI21X1  g06015(.A0(new_n5817_), .A1(new_n5811_), .B0(new_n5865_), .Y(new_n6208_));
  AND2X1   g06016(.A(new_n6208_), .B(new_n5863_), .Y(new_n6209_));
  AOI22X1  g06017(.A0(new_n5817_), .A1(new_n5811_), .B0(new_n5809_), .B1(\asqrt[57] ), .Y(new_n6210_));
  AOI21X1  g06018(.A0(new_n6210_), .A1(\asqrt[34] ), .B0(new_n5816_), .Y(new_n6211_));
  AOI21X1  g06019(.A0(new_n6209_), .A1(\asqrt[34] ), .B0(new_n6211_), .Y(new_n6212_));
  INVX1    g06020(.A(new_n6212_), .Y(new_n6213_));
  AND2X1   g06021(.A(new_n6188_), .B(\asqrt[54] ), .Y(new_n6214_));
  OR2X1    g06022(.A(new_n6172_), .B(new_n6159_), .Y(new_n6215_));
  AND2X1   g06023(.A(new_n6179_), .B(new_n902_), .Y(new_n6216_));
  AOI21X1  g06024(.A0(new_n6216_), .A1(new_n6215_), .B0(new_n6177_), .Y(new_n6217_));
  OAI21X1  g06025(.A0(new_n6217_), .A1(new_n6214_), .B0(\asqrt[55] ), .Y(new_n6218_));
  INVX1    g06026(.A(new_n6187_), .Y(new_n6219_));
  OAI21X1  g06027(.A0(new_n6162_), .A1(new_n902_), .B0(new_n697_), .Y(new_n6220_));
  OAI21X1  g06028(.A0(new_n6220_), .A1(new_n6217_), .B0(new_n6219_), .Y(new_n6221_));
  AOI21X1  g06029(.A0(new_n6221_), .A1(new_n6218_), .B0(new_n582_), .Y(new_n6222_));
  INVX1    g06030(.A(new_n6196_), .Y(new_n6223_));
  NAND3X1  g06031(.A(new_n6221_), .B(new_n6218_), .C(new_n582_), .Y(new_n6224_));
  AOI21X1  g06032(.A0(new_n6224_), .A1(new_n6223_), .B0(new_n6222_), .Y(new_n6225_));
  OAI21X1  g06033(.A0(new_n6225_), .A1(new_n481_), .B0(new_n399_), .Y(new_n6226_));
  OAI21X1  g06034(.A0(new_n6226_), .A1(new_n6206_), .B0(new_n6213_), .Y(new_n6227_));
  AOI21X1  g06035(.A0(new_n6227_), .A1(new_n6207_), .B0(new_n328_), .Y(new_n6228_));
  AND2X1   g06036(.A(new_n5870_), .B(new_n5867_), .Y(new_n6229_));
  NOR3X1   g06037(.A(new_n6229_), .B(new_n5824_), .C(new_n5868_), .Y(new_n6230_));
  NOR2X1   g06038(.A(new_n6229_), .B(new_n5868_), .Y(new_n6231_));
  AOI21X1  g06039(.A0(new_n6231_), .A1(\asqrt[34] ), .B0(new_n5869_), .Y(new_n6232_));
  AOI21X1  g06040(.A0(new_n6230_), .A1(\asqrt[34] ), .B0(new_n6232_), .Y(new_n6233_));
  INVX1    g06041(.A(new_n6233_), .Y(new_n6234_));
  NAND3X1  g06042(.A(new_n6227_), .B(new_n6207_), .C(new_n328_), .Y(new_n6235_));
  AOI21X1  g06043(.A0(new_n6235_), .A1(new_n6234_), .B0(new_n6228_), .Y(new_n6236_));
  OR2X1    g06044(.A(new_n6236_), .B(new_n292_), .Y(new_n6237_));
  OR2X1    g06045(.A(new_n6225_), .B(new_n481_), .Y(new_n6238_));
  NOR2X1   g06046(.A(new_n6197_), .B(new_n6196_), .Y(new_n6239_));
  INVX1    g06047(.A(new_n6204_), .Y(new_n6240_));
  NAND2X1  g06048(.A(new_n6191_), .B(new_n481_), .Y(new_n6241_));
  OAI21X1  g06049(.A0(new_n6241_), .A1(new_n6239_), .B0(new_n6240_), .Y(new_n6242_));
  AOI21X1  g06050(.A0(new_n6242_), .A1(new_n6238_), .B0(new_n399_), .Y(new_n6243_));
  AOI21X1  g06051(.A0(new_n6198_), .A1(\asqrt[57] ), .B0(\asqrt[58] ), .Y(new_n6244_));
  AOI21X1  g06052(.A0(new_n6244_), .A1(new_n6242_), .B0(new_n6212_), .Y(new_n6245_));
  NOR3X1   g06053(.A(new_n6245_), .B(new_n6243_), .C(\asqrt[59] ), .Y(new_n6246_));
  NOR2X1   g06054(.A(new_n6246_), .B(new_n6233_), .Y(new_n6247_));
  NAND4X1  g06055(.A(\asqrt[34] ), .B(new_n5845_), .C(new_n5843_), .D(new_n5872_), .Y(new_n6248_));
  NAND2X1  g06056(.A(new_n5845_), .B(new_n5872_), .Y(new_n6249_));
  OAI21X1  g06057(.A0(new_n6249_), .A1(new_n5941_), .B0(new_n5844_), .Y(new_n6250_));
  AND2X1   g06058(.A(new_n6250_), .B(new_n6248_), .Y(new_n6251_));
  INVX1    g06059(.A(new_n6251_), .Y(new_n6252_));
  OAI21X1  g06060(.A0(new_n6245_), .A1(new_n6243_), .B0(\asqrt[59] ), .Y(new_n6253_));
  NAND2X1  g06061(.A(new_n6253_), .B(new_n292_), .Y(new_n6254_));
  OAI21X1  g06062(.A0(new_n6254_), .A1(new_n6247_), .B0(new_n6252_), .Y(new_n6255_));
  AOI21X1  g06063(.A0(new_n6255_), .A1(new_n6237_), .B0(new_n217_), .Y(new_n6256_));
  AND2X1   g06064(.A(new_n5915_), .B(new_n5914_), .Y(new_n6257_));
  NOR3X1   g06065(.A(new_n6257_), .B(new_n5854_), .C(new_n5913_), .Y(new_n6258_));
  AOI22X1  g06066(.A0(new_n5915_), .A1(new_n5914_), .B0(new_n5874_), .B1(\asqrt[60] ), .Y(new_n6259_));
  AOI21X1  g06067(.A0(new_n6259_), .A1(\asqrt[34] ), .B0(new_n5853_), .Y(new_n6260_));
  AOI21X1  g06068(.A0(new_n6258_), .A1(\asqrt[34] ), .B0(new_n6260_), .Y(new_n6261_));
  OAI21X1  g06069(.A0(new_n6246_), .A1(new_n6233_), .B0(new_n6253_), .Y(new_n6262_));
  AOI21X1  g06070(.A0(new_n6262_), .A1(\asqrt[60] ), .B0(\asqrt[61] ), .Y(new_n6263_));
  AOI21X1  g06071(.A0(new_n6263_), .A1(new_n6255_), .B0(new_n6261_), .Y(new_n6264_));
  OAI21X1  g06072(.A0(new_n6264_), .A1(new_n6256_), .B0(\asqrt[62] ), .Y(new_n6265_));
  AND2X1   g06073(.A(new_n5875_), .B(new_n5856_), .Y(new_n6266_));
  NOR3X1   g06074(.A(new_n6266_), .B(new_n5918_), .C(new_n5857_), .Y(new_n6267_));
  NOR2X1   g06075(.A(new_n6266_), .B(new_n5857_), .Y(new_n6268_));
  AOI21X1  g06076(.A0(new_n6268_), .A1(\asqrt[34] ), .B0(new_n5862_), .Y(new_n6269_));
  AOI21X1  g06077(.A0(new_n6267_), .A1(\asqrt[34] ), .B0(new_n6269_), .Y(new_n6270_));
  NOR3X1   g06078(.A(new_n6264_), .B(new_n6256_), .C(\asqrt[62] ), .Y(new_n6271_));
  OAI21X1  g06079(.A0(new_n6271_), .A1(new_n6270_), .B0(new_n6265_), .Y(new_n6272_));
  NOR3X1   g06080(.A(new_n5923_), .B(new_n5878_), .C(new_n5921_), .Y(new_n6273_));
  AND2X1   g06081(.A(new_n6273_), .B(\asqrt[34] ), .Y(new_n6274_));
  NAND3X1  g06082(.A(\asqrt[34] ), .B(new_n5922_), .C(new_n5877_), .Y(new_n6275_));
  AOI21X1  g06083(.A0(new_n6275_), .A1(new_n5923_), .B0(new_n6274_), .Y(new_n6276_));
  INVX1    g06084(.A(new_n6276_), .Y(new_n6277_));
  AND2X1   g06085(.A(new_n5890_), .B(new_n5883_), .Y(new_n6278_));
  AOI21X1  g06086(.A0(new_n6278_), .A1(\asqrt[34] ), .B0(new_n5946_), .Y(new_n6279_));
  AND2X1   g06087(.A(new_n6279_), .B(new_n6277_), .Y(new_n6280_));
  AOI21X1  g06088(.A0(new_n6280_), .A1(new_n6272_), .B0(\asqrt[63] ), .Y(new_n6281_));
  NOR2X1   g06089(.A(new_n6271_), .B(new_n6270_), .Y(new_n6282_));
  NAND2X1  g06090(.A(new_n6276_), .B(new_n6265_), .Y(new_n6283_));
  AOI21X1  g06091(.A0(new_n5930_), .A1(new_n5926_), .B0(new_n5889_), .Y(new_n6284_));
  AOI21X1  g06092(.A0(new_n5890_), .A1(new_n5883_), .B0(new_n193_), .Y(new_n6285_));
  OAI21X1  g06093(.A0(new_n6284_), .A1(new_n5883_), .B0(new_n6285_), .Y(new_n6286_));
  INVX1    g06094(.A(new_n5888_), .Y(new_n6287_));
  NOR4X1   g06095(.A(new_n5906_), .B(new_n5900_), .C(new_n6287_), .D(new_n5885_), .Y(new_n6288_));
  OAI21X1  g06096(.A0(new_n5897_), .A1(new_n5896_), .B0(new_n6288_), .Y(new_n6289_));
  NOR2X1   g06097(.A(new_n6289_), .B(new_n5895_), .Y(new_n6290_));
  INVX1    g06098(.A(new_n6290_), .Y(new_n6291_));
  AND2X1   g06099(.A(new_n6291_), .B(new_n6286_), .Y(new_n6292_));
  OAI21X1  g06100(.A0(new_n6283_), .A1(new_n6282_), .B0(new_n6292_), .Y(new_n6293_));
  NOR2X1   g06101(.A(new_n6293_), .B(new_n6281_), .Y(new_n6294_));
  INVX1    g06102(.A(\a[66] ), .Y(new_n6295_));
  AND2X1   g06103(.A(new_n6262_), .B(\asqrt[60] ), .Y(new_n6296_));
  OR2X1    g06104(.A(new_n6246_), .B(new_n6233_), .Y(new_n6297_));
  AND2X1   g06105(.A(new_n6253_), .B(new_n292_), .Y(new_n6298_));
  AOI21X1  g06106(.A0(new_n6298_), .A1(new_n6297_), .B0(new_n6251_), .Y(new_n6299_));
  OAI21X1  g06107(.A0(new_n6299_), .A1(new_n6296_), .B0(\asqrt[61] ), .Y(new_n6300_));
  INVX1    g06108(.A(new_n6261_), .Y(new_n6301_));
  OAI21X1  g06109(.A0(new_n6236_), .A1(new_n292_), .B0(new_n217_), .Y(new_n6302_));
  OAI21X1  g06110(.A0(new_n6302_), .A1(new_n6299_), .B0(new_n6301_), .Y(new_n6303_));
  AOI21X1  g06111(.A0(new_n6303_), .A1(new_n6300_), .B0(new_n199_), .Y(new_n6304_));
  INVX1    g06112(.A(new_n6270_), .Y(new_n6305_));
  NAND3X1  g06113(.A(new_n6303_), .B(new_n6300_), .C(new_n199_), .Y(new_n6306_));
  AOI21X1  g06114(.A0(new_n6306_), .A1(new_n6305_), .B0(new_n6304_), .Y(new_n6307_));
  INVX1    g06115(.A(new_n6280_), .Y(new_n6308_));
  OAI21X1  g06116(.A0(new_n6308_), .A1(new_n6307_), .B0(new_n193_), .Y(new_n6309_));
  OR2X1    g06117(.A(new_n6271_), .B(new_n6270_), .Y(new_n6310_));
  AND2X1   g06118(.A(new_n6276_), .B(new_n6265_), .Y(new_n6311_));
  INVX1    g06119(.A(new_n6292_), .Y(new_n6312_));
  AOI21X1  g06120(.A0(new_n6311_), .A1(new_n6310_), .B0(new_n6312_), .Y(new_n6313_));
  AOI21X1  g06121(.A0(new_n6313_), .A1(new_n6309_), .B0(new_n6295_), .Y(new_n6314_));
  NOR3X1   g06122(.A(\a[66] ), .B(\a[65] ), .C(\a[64] ), .Y(new_n6315_));
  OR2X1    g06123(.A(new_n6315_), .B(new_n6314_), .Y(new_n6316_));
  OR2X1    g06124(.A(new_n6315_), .B(new_n5906_), .Y(new_n6317_));
  NOR4X1   g06125(.A(new_n6317_), .B(new_n5900_), .C(new_n5946_), .D(new_n5895_), .Y(new_n6318_));
  INVX1    g06126(.A(new_n6318_), .Y(new_n6319_));
  OR2X1    g06127(.A(new_n6319_), .B(new_n6314_), .Y(new_n6320_));
  OAI21X1  g06128(.A0(new_n6293_), .A1(new_n6281_), .B0(new_n6295_), .Y(new_n6321_));
  AOI21X1  g06129(.A0(new_n6313_), .A1(new_n6309_), .B0(new_n5942_), .Y(new_n6322_));
  AOI21X1  g06130(.A0(new_n6321_), .A1(\a[67] ), .B0(new_n6322_), .Y(new_n6323_));
  AOI22X1  g06131(.A0(new_n6323_), .A1(new_n6320_), .B0(new_n6316_), .B1(\asqrt[34] ), .Y(new_n6324_));
  OR2X1    g06132(.A(new_n6324_), .B(new_n5541_), .Y(new_n6325_));
  AND2X1   g06133(.A(new_n6323_), .B(new_n6320_), .Y(new_n6326_));
  OAI21X1  g06134(.A0(new_n6315_), .A1(new_n6314_), .B0(\asqrt[34] ), .Y(new_n6327_));
  NAND2X1  g06135(.A(new_n6327_), .B(new_n5541_), .Y(new_n6328_));
  OAI21X1  g06136(.A0(new_n6293_), .A1(new_n6281_), .B0(new_n5910_), .Y(new_n6329_));
  INVX1    g06137(.A(new_n6286_), .Y(new_n6330_));
  NOR3X1   g06138(.A(new_n6290_), .B(new_n6330_), .C(new_n5941_), .Y(new_n6331_));
  OAI21X1  g06139(.A0(new_n6283_), .A1(new_n6282_), .B0(new_n6331_), .Y(new_n6332_));
  OR2X1    g06140(.A(new_n6332_), .B(new_n6281_), .Y(new_n6333_));
  AOI21X1  g06141(.A0(new_n6333_), .A1(new_n6329_), .B0(new_n5912_), .Y(new_n6334_));
  OAI21X1  g06142(.A0(new_n6332_), .A1(new_n6281_), .B0(new_n5912_), .Y(new_n6335_));
  NOR2X1   g06143(.A(new_n6335_), .B(new_n6322_), .Y(new_n6336_));
  OR2X1    g06144(.A(new_n6336_), .B(new_n6334_), .Y(new_n6337_));
  OAI21X1  g06145(.A0(new_n6328_), .A1(new_n6326_), .B0(new_n6337_), .Y(new_n6338_));
  AOI21X1  g06146(.A0(new_n6338_), .A1(new_n6325_), .B0(new_n5176_), .Y(new_n6339_));
  AOI21X1  g06147(.A0(new_n5911_), .A1(\asqrt[35] ), .B0(new_n5960_), .Y(new_n6340_));
  AND2X1   g06148(.A(new_n6340_), .B(new_n5963_), .Y(new_n6341_));
  OAI21X1  g06149(.A0(new_n6293_), .A1(new_n6281_), .B0(new_n6341_), .Y(new_n6342_));
  OAI21X1  g06150(.A0(new_n6293_), .A1(new_n6281_), .B0(new_n6340_), .Y(new_n6343_));
  NAND2X1  g06151(.A(new_n6343_), .B(new_n5937_), .Y(new_n6344_));
  AND2X1   g06152(.A(new_n6344_), .B(new_n6342_), .Y(new_n6345_));
  NOR2X1   g06153(.A(new_n6319_), .B(new_n6314_), .Y(new_n6346_));
  INVX1    g06154(.A(\a[67] ), .Y(new_n6347_));
  AOI21X1  g06155(.A0(new_n6313_), .A1(new_n6309_), .B0(\a[66] ), .Y(new_n6348_));
  OAI21X1  g06156(.A0(new_n6348_), .A1(new_n6347_), .B0(new_n6329_), .Y(new_n6349_));
  OAI21X1  g06157(.A0(new_n6349_), .A1(new_n6346_), .B0(new_n6327_), .Y(new_n6350_));
  AOI21X1  g06158(.A0(new_n6350_), .A1(\asqrt[35] ), .B0(\asqrt[36] ), .Y(new_n6351_));
  AOI21X1  g06159(.A0(new_n6351_), .A1(new_n6338_), .B0(new_n6345_), .Y(new_n6352_));
  OAI21X1  g06160(.A0(new_n6352_), .A1(new_n6339_), .B0(\asqrt[37] ), .Y(new_n6353_));
  AOI21X1  g06161(.A0(new_n5984_), .A1(new_n5983_), .B0(new_n5952_), .Y(new_n6354_));
  AND2X1   g06162(.A(new_n6354_), .B(new_n5939_), .Y(new_n6355_));
  OAI21X1  g06163(.A0(new_n6293_), .A1(new_n6281_), .B0(new_n6355_), .Y(new_n6356_));
  AOI22X1  g06164(.A0(new_n5984_), .A1(new_n5983_), .B0(new_n5964_), .B1(\asqrt[36] ), .Y(new_n6357_));
  OAI21X1  g06165(.A0(new_n6293_), .A1(new_n6281_), .B0(new_n6357_), .Y(new_n6358_));
  NAND2X1  g06166(.A(new_n6358_), .B(new_n5952_), .Y(new_n6359_));
  AND2X1   g06167(.A(new_n6359_), .B(new_n6356_), .Y(new_n6360_));
  NOR3X1   g06168(.A(new_n6352_), .B(new_n6339_), .C(\asqrt[37] ), .Y(new_n6361_));
  OAI21X1  g06169(.A0(new_n6361_), .A1(new_n6360_), .B0(new_n6353_), .Y(new_n6362_));
  AND2X1   g06170(.A(new_n6362_), .B(\asqrt[38] ), .Y(new_n6363_));
  OR2X1    g06171(.A(new_n6361_), .B(new_n6360_), .Y(new_n6364_));
  INVX1    g06172(.A(new_n6294_), .Y(\asqrt[33] ));
  AND2X1   g06173(.A(new_n5965_), .B(new_n5953_), .Y(new_n6366_));
  NOR3X1   g06174(.A(new_n6366_), .B(new_n5988_), .C(new_n5954_), .Y(new_n6367_));
  NOR2X1   g06175(.A(new_n6366_), .B(new_n5954_), .Y(new_n6368_));
  OAI21X1  g06176(.A0(new_n6293_), .A1(new_n6281_), .B0(new_n6368_), .Y(new_n6369_));
  AOI22X1  g06177(.A0(new_n6369_), .A1(new_n5988_), .B0(new_n6367_), .B1(\asqrt[33] ), .Y(new_n6370_));
  AND2X1   g06178(.A(new_n6353_), .B(new_n4493_), .Y(new_n6371_));
  AOI21X1  g06179(.A0(new_n6371_), .A1(new_n6364_), .B0(new_n6370_), .Y(new_n6372_));
  OAI21X1  g06180(.A0(new_n6372_), .A1(new_n6363_), .B0(\asqrt[39] ), .Y(new_n6373_));
  NAND4X1  g06181(.A(\asqrt[33] ), .B(new_n6002_), .C(new_n5972_), .D(new_n5967_), .Y(new_n6374_));
  NOR3X1   g06182(.A(new_n6294_), .B(new_n5973_), .C(new_n5991_), .Y(new_n6375_));
  OAI21X1  g06183(.A0(new_n6375_), .A1(new_n5972_), .B0(new_n6374_), .Y(new_n6376_));
  AND2X1   g06184(.A(new_n6350_), .B(\asqrt[35] ), .Y(new_n6377_));
  OR2X1    g06185(.A(new_n6349_), .B(new_n6346_), .Y(new_n6378_));
  AND2X1   g06186(.A(new_n6327_), .B(new_n5541_), .Y(new_n6379_));
  NOR2X1   g06187(.A(new_n6336_), .B(new_n6334_), .Y(new_n6380_));
  AOI21X1  g06188(.A0(new_n6379_), .A1(new_n6378_), .B0(new_n6380_), .Y(new_n6381_));
  OAI21X1  g06189(.A0(new_n6381_), .A1(new_n6377_), .B0(\asqrt[36] ), .Y(new_n6382_));
  NAND2X1  g06190(.A(new_n6344_), .B(new_n6342_), .Y(new_n6383_));
  OAI21X1  g06191(.A0(new_n6324_), .A1(new_n5541_), .B0(new_n5176_), .Y(new_n6384_));
  OAI21X1  g06192(.A0(new_n6384_), .A1(new_n6381_), .B0(new_n6383_), .Y(new_n6385_));
  AOI21X1  g06193(.A0(new_n6385_), .A1(new_n6382_), .B0(new_n4826_), .Y(new_n6386_));
  INVX1    g06194(.A(new_n6360_), .Y(new_n6387_));
  NAND3X1  g06195(.A(new_n6385_), .B(new_n6382_), .C(new_n4826_), .Y(new_n6388_));
  AOI21X1  g06196(.A0(new_n6388_), .A1(new_n6387_), .B0(new_n6386_), .Y(new_n6389_));
  OAI21X1  g06197(.A0(new_n6389_), .A1(new_n4493_), .B0(new_n4165_), .Y(new_n6390_));
  OAI21X1  g06198(.A0(new_n6390_), .A1(new_n6372_), .B0(new_n6376_), .Y(new_n6391_));
  AOI21X1  g06199(.A0(new_n6391_), .A1(new_n6373_), .B0(new_n3863_), .Y(new_n6392_));
  AND2X1   g06200(.A(new_n5992_), .B(new_n5976_), .Y(new_n6393_));
  NOR3X1   g06201(.A(new_n6393_), .B(new_n6018_), .C(new_n5975_), .Y(new_n6394_));
  NOR3X1   g06202(.A(new_n6294_), .B(new_n6393_), .C(new_n5975_), .Y(new_n6395_));
  NOR2X1   g06203(.A(new_n6395_), .B(new_n5981_), .Y(new_n6396_));
  AOI21X1  g06204(.A0(new_n6394_), .A1(\asqrt[33] ), .B0(new_n6396_), .Y(new_n6397_));
  INVX1    g06205(.A(new_n6397_), .Y(new_n6398_));
  NAND3X1  g06206(.A(new_n6391_), .B(new_n6373_), .C(new_n3863_), .Y(new_n6399_));
  AOI21X1  g06207(.A0(new_n6399_), .A1(new_n6398_), .B0(new_n6392_), .Y(new_n6400_));
  OR2X1    g06208(.A(new_n6400_), .B(new_n3564_), .Y(new_n6401_));
  AND2X1   g06209(.A(new_n6399_), .B(new_n6398_), .Y(new_n6402_));
  AND2X1   g06210(.A(new_n6022_), .B(new_n6020_), .Y(new_n6403_));
  NOR3X1   g06211(.A(new_n6403_), .B(new_n6000_), .C(new_n6021_), .Y(new_n6404_));
  NOR3X1   g06212(.A(new_n6294_), .B(new_n6403_), .C(new_n6021_), .Y(new_n6405_));
  NOR2X1   g06213(.A(new_n6405_), .B(new_n5999_), .Y(new_n6406_));
  AOI21X1  g06214(.A0(new_n6404_), .A1(\asqrt[33] ), .B0(new_n6406_), .Y(new_n6407_));
  INVX1    g06215(.A(new_n6407_), .Y(new_n6408_));
  OR2X1    g06216(.A(new_n6389_), .B(new_n4493_), .Y(new_n6409_));
  NOR2X1   g06217(.A(new_n6361_), .B(new_n6360_), .Y(new_n6410_));
  INVX1    g06218(.A(new_n6370_), .Y(new_n6411_));
  NAND2X1  g06219(.A(new_n6353_), .B(new_n4493_), .Y(new_n6412_));
  OAI21X1  g06220(.A0(new_n6412_), .A1(new_n6410_), .B0(new_n6411_), .Y(new_n6413_));
  AOI21X1  g06221(.A0(new_n6413_), .A1(new_n6409_), .B0(new_n4165_), .Y(new_n6414_));
  INVX1    g06222(.A(new_n6376_), .Y(new_n6415_));
  AOI21X1  g06223(.A0(new_n6362_), .A1(\asqrt[38] ), .B0(\asqrt[39] ), .Y(new_n6416_));
  AOI21X1  g06224(.A0(new_n6416_), .A1(new_n6413_), .B0(new_n6415_), .Y(new_n6417_));
  OAI21X1  g06225(.A0(new_n6417_), .A1(new_n6414_), .B0(\asqrt[40] ), .Y(new_n6418_));
  NAND2X1  g06226(.A(new_n6418_), .B(new_n3564_), .Y(new_n6419_));
  OAI21X1  g06227(.A0(new_n6419_), .A1(new_n6402_), .B0(new_n6408_), .Y(new_n6420_));
  AOI21X1  g06228(.A0(new_n6420_), .A1(new_n6401_), .B0(new_n3276_), .Y(new_n6421_));
  OR4X1    g06229(.A(new_n6294_), .B(new_n6024_), .C(new_n6012_), .D(new_n6006_), .Y(new_n6422_));
  OR2X1    g06230(.A(new_n6024_), .B(new_n6006_), .Y(new_n6423_));
  OAI21X1  g06231(.A0(new_n6423_), .A1(new_n6294_), .B0(new_n6012_), .Y(new_n6424_));
  AND2X1   g06232(.A(new_n6424_), .B(new_n6422_), .Y(new_n6425_));
  NOR3X1   g06233(.A(new_n6417_), .B(new_n6414_), .C(\asqrt[40] ), .Y(new_n6426_));
  OAI21X1  g06234(.A0(new_n6426_), .A1(new_n6397_), .B0(new_n6418_), .Y(new_n6427_));
  AOI21X1  g06235(.A0(new_n6427_), .A1(\asqrt[41] ), .B0(\asqrt[42] ), .Y(new_n6428_));
  AOI21X1  g06236(.A0(new_n6428_), .A1(new_n6420_), .B0(new_n6425_), .Y(new_n6429_));
  OAI21X1  g06237(.A0(new_n6429_), .A1(new_n6421_), .B0(\asqrt[43] ), .Y(new_n6430_));
  AOI21X1  g06238(.A0(new_n6055_), .A1(new_n6054_), .B0(new_n6030_), .Y(new_n6431_));
  AND2X1   g06239(.A(new_n6431_), .B(new_n6015_), .Y(new_n6432_));
  AOI22X1  g06240(.A0(new_n6055_), .A1(new_n6054_), .B0(new_n6040_), .B1(\asqrt[42] ), .Y(new_n6433_));
  AOI21X1  g06241(.A0(new_n6433_), .A1(\asqrt[33] ), .B0(new_n6029_), .Y(new_n6434_));
  AOI21X1  g06242(.A0(new_n6432_), .A1(\asqrt[33] ), .B0(new_n6434_), .Y(new_n6435_));
  NOR3X1   g06243(.A(new_n6429_), .B(new_n6421_), .C(\asqrt[43] ), .Y(new_n6436_));
  OAI21X1  g06244(.A0(new_n6436_), .A1(new_n6435_), .B0(new_n6430_), .Y(new_n6437_));
  AND2X1   g06245(.A(new_n6437_), .B(\asqrt[44] ), .Y(new_n6438_));
  INVX1    g06246(.A(new_n6435_), .Y(new_n6439_));
  AND2X1   g06247(.A(new_n6427_), .B(\asqrt[41] ), .Y(new_n6440_));
  NAND2X1  g06248(.A(new_n6399_), .B(new_n6398_), .Y(new_n6441_));
  AND2X1   g06249(.A(new_n6418_), .B(new_n3564_), .Y(new_n6442_));
  AOI21X1  g06250(.A0(new_n6442_), .A1(new_n6441_), .B0(new_n6407_), .Y(new_n6443_));
  OAI21X1  g06251(.A0(new_n6443_), .A1(new_n6440_), .B0(\asqrt[42] ), .Y(new_n6444_));
  INVX1    g06252(.A(new_n6425_), .Y(new_n6445_));
  OAI21X1  g06253(.A0(new_n6400_), .A1(new_n3564_), .B0(new_n3276_), .Y(new_n6446_));
  OAI21X1  g06254(.A0(new_n6446_), .A1(new_n6443_), .B0(new_n6445_), .Y(new_n6447_));
  NAND3X1  g06255(.A(new_n6447_), .B(new_n6444_), .C(new_n3008_), .Y(new_n6448_));
  NAND2X1  g06256(.A(new_n6448_), .B(new_n6439_), .Y(new_n6449_));
  AND2X1   g06257(.A(new_n6041_), .B(new_n6033_), .Y(new_n6450_));
  NOR3X1   g06258(.A(new_n6450_), .B(new_n6058_), .C(new_n6034_), .Y(new_n6451_));
  NOR3X1   g06259(.A(new_n6294_), .B(new_n6450_), .C(new_n6034_), .Y(new_n6452_));
  NOR2X1   g06260(.A(new_n6452_), .B(new_n6039_), .Y(new_n6453_));
  AOI21X1  g06261(.A0(new_n6451_), .A1(\asqrt[33] ), .B0(new_n6453_), .Y(new_n6454_));
  AND2X1   g06262(.A(new_n6430_), .B(new_n2769_), .Y(new_n6455_));
  AOI21X1  g06263(.A0(new_n6455_), .A1(new_n6449_), .B0(new_n6454_), .Y(new_n6456_));
  OAI21X1  g06264(.A0(new_n6456_), .A1(new_n6438_), .B0(\asqrt[45] ), .Y(new_n6457_));
  NAND4X1  g06265(.A(\asqrt[33] ), .B(new_n6061_), .C(new_n6048_), .D(new_n6043_), .Y(new_n6458_));
  NAND2X1  g06266(.A(new_n6061_), .B(new_n6043_), .Y(new_n6459_));
  OAI21X1  g06267(.A0(new_n6459_), .A1(new_n6294_), .B0(new_n6052_), .Y(new_n6460_));
  AND2X1   g06268(.A(new_n6460_), .B(new_n6458_), .Y(new_n6461_));
  INVX1    g06269(.A(new_n6461_), .Y(new_n6462_));
  AOI21X1  g06270(.A0(new_n6447_), .A1(new_n6444_), .B0(new_n3008_), .Y(new_n6463_));
  AOI21X1  g06271(.A0(new_n6448_), .A1(new_n6439_), .B0(new_n6463_), .Y(new_n6464_));
  OAI21X1  g06272(.A0(new_n6464_), .A1(new_n2769_), .B0(new_n2570_), .Y(new_n6465_));
  OAI21X1  g06273(.A0(new_n6465_), .A1(new_n6456_), .B0(new_n6462_), .Y(new_n6466_));
  AOI21X1  g06274(.A0(new_n6466_), .A1(new_n6457_), .B0(new_n2263_), .Y(new_n6467_));
  AND2X1   g06275(.A(new_n6068_), .B(new_n6062_), .Y(new_n6468_));
  NOR3X1   g06276(.A(new_n6468_), .B(new_n6092_), .C(new_n6051_), .Y(new_n6469_));
  NOR3X1   g06277(.A(new_n6294_), .B(new_n6468_), .C(new_n6051_), .Y(new_n6470_));
  NOR2X1   g06278(.A(new_n6470_), .B(new_n6066_), .Y(new_n6471_));
  AOI21X1  g06279(.A0(new_n6469_), .A1(\asqrt[33] ), .B0(new_n6471_), .Y(new_n6472_));
  INVX1    g06280(.A(new_n6472_), .Y(new_n6473_));
  NAND3X1  g06281(.A(new_n6466_), .B(new_n6457_), .C(new_n2263_), .Y(new_n6474_));
  AOI21X1  g06282(.A0(new_n6474_), .A1(new_n6473_), .B0(new_n6467_), .Y(new_n6475_));
  OR2X1    g06283(.A(new_n6475_), .B(new_n2040_), .Y(new_n6476_));
  AND2X1   g06284(.A(new_n6474_), .B(new_n6473_), .Y(new_n6477_));
  AND2X1   g06285(.A(new_n6096_), .B(new_n6094_), .Y(new_n6478_));
  NOR3X1   g06286(.A(new_n6478_), .B(new_n6076_), .C(new_n6095_), .Y(new_n6479_));
  NOR3X1   g06287(.A(new_n6294_), .B(new_n6478_), .C(new_n6095_), .Y(new_n6480_));
  NOR2X1   g06288(.A(new_n6480_), .B(new_n6075_), .Y(new_n6481_));
  AOI21X1  g06289(.A0(new_n6479_), .A1(\asqrt[33] ), .B0(new_n6481_), .Y(new_n6482_));
  INVX1    g06290(.A(new_n6482_), .Y(new_n6483_));
  OR2X1    g06291(.A(new_n6464_), .B(new_n2769_), .Y(new_n6484_));
  AND2X1   g06292(.A(new_n6448_), .B(new_n6439_), .Y(new_n6485_));
  INVX1    g06293(.A(new_n6454_), .Y(new_n6486_));
  NAND2X1  g06294(.A(new_n6430_), .B(new_n2769_), .Y(new_n6487_));
  OAI21X1  g06295(.A0(new_n6487_), .A1(new_n6485_), .B0(new_n6486_), .Y(new_n6488_));
  AOI21X1  g06296(.A0(new_n6488_), .A1(new_n6484_), .B0(new_n2570_), .Y(new_n6489_));
  AOI21X1  g06297(.A0(new_n6437_), .A1(\asqrt[44] ), .B0(\asqrt[45] ), .Y(new_n6490_));
  AOI21X1  g06298(.A0(new_n6490_), .A1(new_n6488_), .B0(new_n6461_), .Y(new_n6491_));
  OAI21X1  g06299(.A0(new_n6491_), .A1(new_n6489_), .B0(\asqrt[46] ), .Y(new_n6492_));
  NAND2X1  g06300(.A(new_n6492_), .B(new_n2040_), .Y(new_n6493_));
  OAI21X1  g06301(.A0(new_n6493_), .A1(new_n6477_), .B0(new_n6483_), .Y(new_n6494_));
  AOI21X1  g06302(.A0(new_n6494_), .A1(new_n6476_), .B0(new_n1834_), .Y(new_n6495_));
  NAND4X1  g06303(.A(\asqrt[33] ), .B(new_n6087_), .C(new_n6085_), .D(new_n6113_), .Y(new_n6496_));
  NAND2X1  g06304(.A(new_n6087_), .B(new_n6113_), .Y(new_n6497_));
  OAI21X1  g06305(.A0(new_n6497_), .A1(new_n6294_), .B0(new_n6086_), .Y(new_n6498_));
  AND2X1   g06306(.A(new_n6498_), .B(new_n6496_), .Y(new_n6499_));
  NOR3X1   g06307(.A(new_n6491_), .B(new_n6489_), .C(\asqrt[46] ), .Y(new_n6500_));
  OAI21X1  g06308(.A0(new_n6500_), .A1(new_n6472_), .B0(new_n6492_), .Y(new_n6501_));
  AOI21X1  g06309(.A0(new_n6501_), .A1(\asqrt[47] ), .B0(\asqrt[48] ), .Y(new_n6502_));
  AOI21X1  g06310(.A0(new_n6502_), .A1(new_n6494_), .B0(new_n6499_), .Y(new_n6503_));
  OAI21X1  g06311(.A0(new_n6503_), .A1(new_n6495_), .B0(\asqrt[49] ), .Y(new_n6504_));
  AOI21X1  g06312(.A0(new_n6133_), .A1(new_n6132_), .B0(new_n6104_), .Y(new_n6505_));
  AND2X1   g06313(.A(new_n6505_), .B(new_n6089_), .Y(new_n6506_));
  AOI22X1  g06314(.A0(new_n6133_), .A1(new_n6132_), .B0(new_n6114_), .B1(\asqrt[48] ), .Y(new_n6507_));
  AOI21X1  g06315(.A0(new_n6507_), .A1(\asqrt[33] ), .B0(new_n6103_), .Y(new_n6508_));
  AOI21X1  g06316(.A0(new_n6506_), .A1(\asqrt[33] ), .B0(new_n6508_), .Y(new_n6509_));
  NOR3X1   g06317(.A(new_n6503_), .B(new_n6495_), .C(\asqrt[49] ), .Y(new_n6510_));
  OAI21X1  g06318(.A0(new_n6510_), .A1(new_n6509_), .B0(new_n6504_), .Y(new_n6511_));
  AND2X1   g06319(.A(new_n6511_), .B(\asqrt[50] ), .Y(new_n6512_));
  INVX1    g06320(.A(new_n6509_), .Y(new_n6513_));
  AND2X1   g06321(.A(new_n6501_), .B(\asqrt[47] ), .Y(new_n6514_));
  NAND2X1  g06322(.A(new_n6474_), .B(new_n6473_), .Y(new_n6515_));
  AND2X1   g06323(.A(new_n6492_), .B(new_n2040_), .Y(new_n6516_));
  AOI21X1  g06324(.A0(new_n6516_), .A1(new_n6515_), .B0(new_n6482_), .Y(new_n6517_));
  OAI21X1  g06325(.A0(new_n6517_), .A1(new_n6514_), .B0(\asqrt[48] ), .Y(new_n6518_));
  INVX1    g06326(.A(new_n6499_), .Y(new_n6519_));
  OAI21X1  g06327(.A0(new_n6475_), .A1(new_n2040_), .B0(new_n1834_), .Y(new_n6520_));
  OAI21X1  g06328(.A0(new_n6520_), .A1(new_n6517_), .B0(new_n6519_), .Y(new_n6521_));
  NAND3X1  g06329(.A(new_n6521_), .B(new_n6518_), .C(new_n1632_), .Y(new_n6522_));
  NAND2X1  g06330(.A(new_n6522_), .B(new_n6513_), .Y(new_n6523_));
  AND2X1   g06331(.A(new_n6115_), .B(new_n6106_), .Y(new_n6524_));
  NOR3X1   g06332(.A(new_n6524_), .B(new_n6136_), .C(new_n6107_), .Y(new_n6525_));
  NOR3X1   g06333(.A(new_n6294_), .B(new_n6524_), .C(new_n6107_), .Y(new_n6526_));
  NOR2X1   g06334(.A(new_n6526_), .B(new_n6112_), .Y(new_n6527_));
  AOI21X1  g06335(.A0(new_n6525_), .A1(\asqrt[33] ), .B0(new_n6527_), .Y(new_n6528_));
  AND2X1   g06336(.A(new_n6504_), .B(new_n1469_), .Y(new_n6529_));
  AOI21X1  g06337(.A0(new_n6529_), .A1(new_n6523_), .B0(new_n6528_), .Y(new_n6530_));
  OAI21X1  g06338(.A0(new_n6530_), .A1(new_n6512_), .B0(\asqrt[51] ), .Y(new_n6531_));
  NAND4X1  g06339(.A(\asqrt[33] ), .B(new_n6150_), .C(new_n6122_), .D(new_n6117_), .Y(new_n6532_));
  NAND2X1  g06340(.A(new_n6150_), .B(new_n6117_), .Y(new_n6533_));
  OAI21X1  g06341(.A0(new_n6533_), .A1(new_n6294_), .B0(new_n6149_), .Y(new_n6534_));
  AND2X1   g06342(.A(new_n6534_), .B(new_n6532_), .Y(new_n6535_));
  INVX1    g06343(.A(new_n6535_), .Y(new_n6536_));
  AOI21X1  g06344(.A0(new_n6521_), .A1(new_n6518_), .B0(new_n1632_), .Y(new_n6537_));
  AOI21X1  g06345(.A0(new_n6522_), .A1(new_n6513_), .B0(new_n6537_), .Y(new_n6538_));
  OAI21X1  g06346(.A0(new_n6538_), .A1(new_n1469_), .B0(new_n1277_), .Y(new_n6539_));
  OAI21X1  g06347(.A0(new_n6539_), .A1(new_n6530_), .B0(new_n6536_), .Y(new_n6540_));
  AOI21X1  g06348(.A0(new_n6540_), .A1(new_n6531_), .B0(new_n1111_), .Y(new_n6541_));
  AND2X1   g06349(.A(new_n6140_), .B(new_n6126_), .Y(new_n6542_));
  NOR3X1   g06350(.A(new_n6542_), .B(new_n6166_), .C(new_n6125_), .Y(new_n6543_));
  NOR3X1   g06351(.A(new_n6294_), .B(new_n6542_), .C(new_n6125_), .Y(new_n6544_));
  NOR2X1   g06352(.A(new_n6544_), .B(new_n6130_), .Y(new_n6545_));
  AOI21X1  g06353(.A0(new_n6543_), .A1(\asqrt[33] ), .B0(new_n6545_), .Y(new_n6546_));
  INVX1    g06354(.A(new_n6546_), .Y(new_n6547_));
  NAND3X1  g06355(.A(new_n6540_), .B(new_n6531_), .C(new_n1111_), .Y(new_n6548_));
  AOI21X1  g06356(.A0(new_n6548_), .A1(new_n6547_), .B0(new_n6541_), .Y(new_n6549_));
  OR2X1    g06357(.A(new_n6549_), .B(new_n968_), .Y(new_n6550_));
  AND2X1   g06358(.A(new_n6548_), .B(new_n6547_), .Y(new_n6551_));
  AND2X1   g06359(.A(new_n6170_), .B(new_n6168_), .Y(new_n6552_));
  NOR3X1   g06360(.A(new_n6552_), .B(new_n6148_), .C(new_n6169_), .Y(new_n6553_));
  NOR3X1   g06361(.A(new_n6294_), .B(new_n6552_), .C(new_n6169_), .Y(new_n6554_));
  NOR2X1   g06362(.A(new_n6554_), .B(new_n6147_), .Y(new_n6555_));
  AOI21X1  g06363(.A0(new_n6553_), .A1(\asqrt[33] ), .B0(new_n6555_), .Y(new_n6556_));
  INVX1    g06364(.A(new_n6556_), .Y(new_n6557_));
  OR2X1    g06365(.A(new_n6538_), .B(new_n1469_), .Y(new_n6558_));
  AND2X1   g06366(.A(new_n6522_), .B(new_n6513_), .Y(new_n6559_));
  INVX1    g06367(.A(new_n6528_), .Y(new_n6560_));
  NAND2X1  g06368(.A(new_n6504_), .B(new_n1469_), .Y(new_n6561_));
  OAI21X1  g06369(.A0(new_n6561_), .A1(new_n6559_), .B0(new_n6560_), .Y(new_n6562_));
  AOI21X1  g06370(.A0(new_n6562_), .A1(new_n6558_), .B0(new_n1277_), .Y(new_n6563_));
  AOI21X1  g06371(.A0(new_n6511_), .A1(\asqrt[50] ), .B0(\asqrt[51] ), .Y(new_n6564_));
  AOI21X1  g06372(.A0(new_n6564_), .A1(new_n6562_), .B0(new_n6535_), .Y(new_n6565_));
  OAI21X1  g06373(.A0(new_n6565_), .A1(new_n6563_), .B0(\asqrt[52] ), .Y(new_n6566_));
  NAND2X1  g06374(.A(new_n6566_), .B(new_n968_), .Y(new_n6567_));
  OAI21X1  g06375(.A0(new_n6567_), .A1(new_n6551_), .B0(new_n6557_), .Y(new_n6568_));
  AOI21X1  g06376(.A0(new_n6568_), .A1(new_n6550_), .B0(new_n902_), .Y(new_n6569_));
  OR4X1    g06377(.A(new_n6294_), .B(new_n6172_), .C(new_n6160_), .D(new_n6154_), .Y(new_n6570_));
  OR2X1    g06378(.A(new_n6172_), .B(new_n6154_), .Y(new_n6571_));
  OAI21X1  g06379(.A0(new_n6571_), .A1(new_n6294_), .B0(new_n6160_), .Y(new_n6572_));
  AND2X1   g06380(.A(new_n6572_), .B(new_n6570_), .Y(new_n6573_));
  NOR3X1   g06381(.A(new_n6565_), .B(new_n6563_), .C(\asqrt[52] ), .Y(new_n6574_));
  OAI21X1  g06382(.A0(new_n6574_), .A1(new_n6546_), .B0(new_n6566_), .Y(new_n6575_));
  AOI21X1  g06383(.A0(new_n6575_), .A1(\asqrt[53] ), .B0(\asqrt[54] ), .Y(new_n6576_));
  AOI21X1  g06384(.A0(new_n6576_), .A1(new_n6568_), .B0(new_n6573_), .Y(new_n6577_));
  OAI21X1  g06385(.A0(new_n6577_), .A1(new_n6569_), .B0(\asqrt[55] ), .Y(new_n6578_));
  AOI21X1  g06386(.A0(new_n6216_), .A1(new_n6215_), .B0(new_n6178_), .Y(new_n6579_));
  AND2X1   g06387(.A(new_n6579_), .B(new_n6163_), .Y(new_n6580_));
  AOI22X1  g06388(.A0(new_n6216_), .A1(new_n6215_), .B0(new_n6188_), .B1(\asqrt[54] ), .Y(new_n6581_));
  AOI21X1  g06389(.A0(new_n6581_), .A1(\asqrt[33] ), .B0(new_n6177_), .Y(new_n6582_));
  AOI21X1  g06390(.A0(new_n6580_), .A1(\asqrt[33] ), .B0(new_n6582_), .Y(new_n6583_));
  NOR3X1   g06391(.A(new_n6577_), .B(new_n6569_), .C(\asqrt[55] ), .Y(new_n6584_));
  OAI21X1  g06392(.A0(new_n6584_), .A1(new_n6583_), .B0(new_n6578_), .Y(new_n6585_));
  AND2X1   g06393(.A(new_n6585_), .B(\asqrt[56] ), .Y(new_n6586_));
  INVX1    g06394(.A(new_n6583_), .Y(new_n6587_));
  AND2X1   g06395(.A(new_n6575_), .B(\asqrt[53] ), .Y(new_n6588_));
  NAND2X1  g06396(.A(new_n6548_), .B(new_n6547_), .Y(new_n6589_));
  AND2X1   g06397(.A(new_n6566_), .B(new_n968_), .Y(new_n6590_));
  AOI21X1  g06398(.A0(new_n6590_), .A1(new_n6589_), .B0(new_n6556_), .Y(new_n6591_));
  OAI21X1  g06399(.A0(new_n6591_), .A1(new_n6588_), .B0(\asqrt[54] ), .Y(new_n6592_));
  INVX1    g06400(.A(new_n6573_), .Y(new_n6593_));
  OAI21X1  g06401(.A0(new_n6549_), .A1(new_n968_), .B0(new_n902_), .Y(new_n6594_));
  OAI21X1  g06402(.A0(new_n6594_), .A1(new_n6591_), .B0(new_n6593_), .Y(new_n6595_));
  NAND3X1  g06403(.A(new_n6595_), .B(new_n6592_), .C(new_n697_), .Y(new_n6596_));
  NAND2X1  g06404(.A(new_n6596_), .B(new_n6587_), .Y(new_n6597_));
  AND2X1   g06405(.A(new_n6189_), .B(new_n6181_), .Y(new_n6598_));
  NOR3X1   g06406(.A(new_n6598_), .B(new_n6219_), .C(new_n6182_), .Y(new_n6599_));
  NOR3X1   g06407(.A(new_n6294_), .B(new_n6598_), .C(new_n6182_), .Y(new_n6600_));
  NOR2X1   g06408(.A(new_n6600_), .B(new_n6187_), .Y(new_n6601_));
  AOI21X1  g06409(.A0(new_n6599_), .A1(\asqrt[33] ), .B0(new_n6601_), .Y(new_n6602_));
  AND2X1   g06410(.A(new_n6578_), .B(new_n582_), .Y(new_n6603_));
  AOI21X1  g06411(.A0(new_n6603_), .A1(new_n6597_), .B0(new_n6602_), .Y(new_n6604_));
  OAI21X1  g06412(.A0(new_n6604_), .A1(new_n6586_), .B0(\asqrt[57] ), .Y(new_n6605_));
  OR4X1    g06413(.A(new_n6294_), .B(new_n6197_), .C(new_n6223_), .D(new_n6222_), .Y(new_n6606_));
  OR2X1    g06414(.A(new_n6197_), .B(new_n6222_), .Y(new_n6607_));
  OAI21X1  g06415(.A0(new_n6607_), .A1(new_n6294_), .B0(new_n6223_), .Y(new_n6608_));
  AND2X1   g06416(.A(new_n6608_), .B(new_n6606_), .Y(new_n6609_));
  INVX1    g06417(.A(new_n6609_), .Y(new_n6610_));
  AOI21X1  g06418(.A0(new_n6595_), .A1(new_n6592_), .B0(new_n697_), .Y(new_n6611_));
  AOI21X1  g06419(.A0(new_n6596_), .A1(new_n6587_), .B0(new_n6611_), .Y(new_n6612_));
  OAI21X1  g06420(.A0(new_n6612_), .A1(new_n582_), .B0(new_n481_), .Y(new_n6613_));
  OAI21X1  g06421(.A0(new_n6613_), .A1(new_n6604_), .B0(new_n6610_), .Y(new_n6614_));
  AOI21X1  g06422(.A0(new_n6614_), .A1(new_n6605_), .B0(new_n399_), .Y(new_n6615_));
  AND2X1   g06423(.A(new_n6205_), .B(new_n6200_), .Y(new_n6616_));
  NOR3X1   g06424(.A(new_n6616_), .B(new_n6240_), .C(new_n6199_), .Y(new_n6617_));
  NOR3X1   g06425(.A(new_n6294_), .B(new_n6616_), .C(new_n6199_), .Y(new_n6618_));
  NOR2X1   g06426(.A(new_n6618_), .B(new_n6204_), .Y(new_n6619_));
  AOI21X1  g06427(.A0(new_n6617_), .A1(\asqrt[33] ), .B0(new_n6619_), .Y(new_n6620_));
  INVX1    g06428(.A(new_n6620_), .Y(new_n6621_));
  NAND3X1  g06429(.A(new_n6614_), .B(new_n6605_), .C(new_n399_), .Y(new_n6622_));
  AOI21X1  g06430(.A0(new_n6622_), .A1(new_n6621_), .B0(new_n6615_), .Y(new_n6623_));
  OR2X1    g06431(.A(new_n6623_), .B(new_n328_), .Y(new_n6624_));
  AND2X1   g06432(.A(new_n6622_), .B(new_n6621_), .Y(new_n6625_));
  AND2X1   g06433(.A(new_n6244_), .B(new_n6242_), .Y(new_n6626_));
  NOR3X1   g06434(.A(new_n6626_), .B(new_n6213_), .C(new_n6243_), .Y(new_n6627_));
  NOR3X1   g06435(.A(new_n6294_), .B(new_n6626_), .C(new_n6243_), .Y(new_n6628_));
  NOR2X1   g06436(.A(new_n6628_), .B(new_n6212_), .Y(new_n6629_));
  AOI21X1  g06437(.A0(new_n6627_), .A1(\asqrt[33] ), .B0(new_n6629_), .Y(new_n6630_));
  INVX1    g06438(.A(new_n6630_), .Y(new_n6631_));
  OR2X1    g06439(.A(new_n6612_), .B(new_n582_), .Y(new_n6632_));
  AND2X1   g06440(.A(new_n6596_), .B(new_n6587_), .Y(new_n6633_));
  INVX1    g06441(.A(new_n6602_), .Y(new_n6634_));
  NAND2X1  g06442(.A(new_n6578_), .B(new_n582_), .Y(new_n6635_));
  OAI21X1  g06443(.A0(new_n6635_), .A1(new_n6633_), .B0(new_n6634_), .Y(new_n6636_));
  AOI21X1  g06444(.A0(new_n6636_), .A1(new_n6632_), .B0(new_n481_), .Y(new_n6637_));
  AOI21X1  g06445(.A0(new_n6585_), .A1(\asqrt[56] ), .B0(\asqrt[57] ), .Y(new_n6638_));
  AOI21X1  g06446(.A0(new_n6638_), .A1(new_n6636_), .B0(new_n6609_), .Y(new_n6639_));
  OAI21X1  g06447(.A0(new_n6639_), .A1(new_n6637_), .B0(\asqrt[58] ), .Y(new_n6640_));
  NAND2X1  g06448(.A(new_n6640_), .B(new_n328_), .Y(new_n6641_));
  OAI21X1  g06449(.A0(new_n6641_), .A1(new_n6625_), .B0(new_n6631_), .Y(new_n6642_));
  AOI21X1  g06450(.A0(new_n6642_), .A1(new_n6624_), .B0(new_n292_), .Y(new_n6643_));
  NAND4X1  g06451(.A(\asqrt[33] ), .B(new_n6235_), .C(new_n6233_), .D(new_n6253_), .Y(new_n6644_));
  OR2X1    g06452(.A(new_n6246_), .B(new_n6228_), .Y(new_n6645_));
  OAI21X1  g06453(.A0(new_n6645_), .A1(new_n6294_), .B0(new_n6234_), .Y(new_n6646_));
  AND2X1   g06454(.A(new_n6646_), .B(new_n6644_), .Y(new_n6647_));
  NOR3X1   g06455(.A(new_n6639_), .B(new_n6637_), .C(\asqrt[58] ), .Y(new_n6648_));
  OAI21X1  g06456(.A0(new_n6648_), .A1(new_n6620_), .B0(new_n6640_), .Y(new_n6649_));
  AOI21X1  g06457(.A0(new_n6649_), .A1(\asqrt[59] ), .B0(\asqrt[60] ), .Y(new_n6650_));
  AOI21X1  g06458(.A0(new_n6650_), .A1(new_n6642_), .B0(new_n6647_), .Y(new_n6651_));
  OAI21X1  g06459(.A0(new_n6651_), .A1(new_n6643_), .B0(\asqrt[61] ), .Y(new_n6652_));
  AOI21X1  g06460(.A0(new_n6298_), .A1(new_n6297_), .B0(new_n6252_), .Y(new_n6653_));
  AND2X1   g06461(.A(new_n6653_), .B(new_n6237_), .Y(new_n6654_));
  AOI22X1  g06462(.A0(new_n6298_), .A1(new_n6297_), .B0(new_n6262_), .B1(\asqrt[60] ), .Y(new_n6655_));
  AOI21X1  g06463(.A0(new_n6655_), .A1(\asqrt[33] ), .B0(new_n6251_), .Y(new_n6656_));
  AOI21X1  g06464(.A0(new_n6654_), .A1(\asqrt[33] ), .B0(new_n6656_), .Y(new_n6657_));
  NOR3X1   g06465(.A(new_n6651_), .B(new_n6643_), .C(\asqrt[61] ), .Y(new_n6658_));
  OAI21X1  g06466(.A0(new_n6658_), .A1(new_n6657_), .B0(new_n6652_), .Y(new_n6659_));
  AND2X1   g06467(.A(new_n6659_), .B(\asqrt[62] ), .Y(new_n6660_));
  INVX1    g06468(.A(new_n6657_), .Y(new_n6661_));
  AND2X1   g06469(.A(new_n6649_), .B(\asqrt[59] ), .Y(new_n6662_));
  NAND2X1  g06470(.A(new_n6622_), .B(new_n6621_), .Y(new_n6663_));
  AND2X1   g06471(.A(new_n6640_), .B(new_n328_), .Y(new_n6664_));
  AOI21X1  g06472(.A0(new_n6664_), .A1(new_n6663_), .B0(new_n6630_), .Y(new_n6665_));
  OAI21X1  g06473(.A0(new_n6665_), .A1(new_n6662_), .B0(\asqrt[60] ), .Y(new_n6666_));
  INVX1    g06474(.A(new_n6647_), .Y(new_n6667_));
  OAI21X1  g06475(.A0(new_n6623_), .A1(new_n328_), .B0(new_n292_), .Y(new_n6668_));
  OAI21X1  g06476(.A0(new_n6668_), .A1(new_n6665_), .B0(new_n6667_), .Y(new_n6669_));
  NAND3X1  g06477(.A(new_n6669_), .B(new_n6666_), .C(new_n217_), .Y(new_n6670_));
  NAND2X1  g06478(.A(new_n6670_), .B(new_n6661_), .Y(new_n6671_));
  AND2X1   g06479(.A(new_n6263_), .B(new_n6255_), .Y(new_n6672_));
  NOR3X1   g06480(.A(new_n6672_), .B(new_n6301_), .C(new_n6256_), .Y(new_n6673_));
  NOR3X1   g06481(.A(new_n6294_), .B(new_n6672_), .C(new_n6256_), .Y(new_n6674_));
  NOR2X1   g06482(.A(new_n6674_), .B(new_n6261_), .Y(new_n6675_));
  AOI21X1  g06483(.A0(new_n6673_), .A1(\asqrt[33] ), .B0(new_n6675_), .Y(new_n6676_));
  AOI21X1  g06484(.A0(new_n6669_), .A1(new_n6666_), .B0(new_n217_), .Y(new_n6677_));
  NOR2X1   g06485(.A(new_n6677_), .B(\asqrt[62] ), .Y(new_n6678_));
  AOI21X1  g06486(.A0(new_n6678_), .A1(new_n6671_), .B0(new_n6676_), .Y(new_n6679_));
  NOR4X1   g06487(.A(new_n6294_), .B(new_n6271_), .C(new_n6305_), .D(new_n6304_), .Y(new_n6680_));
  NAND3X1  g06488(.A(\asqrt[33] ), .B(new_n6306_), .C(new_n6265_), .Y(new_n6681_));
  AOI21X1  g06489(.A0(new_n6681_), .A1(new_n6305_), .B0(new_n6680_), .Y(new_n6682_));
  INVX1    g06490(.A(new_n6682_), .Y(new_n6683_));
  NOR3X1   g06491(.A(new_n6294_), .B(new_n6276_), .C(new_n6307_), .Y(new_n6684_));
  AOI21X1  g06492(.A0(new_n6311_), .A1(new_n6310_), .B0(new_n6684_), .Y(new_n6685_));
  AND2X1   g06493(.A(new_n6685_), .B(new_n6683_), .Y(new_n6686_));
  OAI21X1  g06494(.A0(new_n6679_), .A1(new_n6660_), .B0(new_n6686_), .Y(new_n6687_));
  AOI21X1  g06495(.A0(new_n6670_), .A1(new_n6661_), .B0(new_n6677_), .Y(new_n6688_));
  OAI21X1  g06496(.A0(new_n6688_), .A1(new_n199_), .B0(new_n6682_), .Y(new_n6689_));
  AOI21X1  g06497(.A0(new_n6313_), .A1(new_n6309_), .B0(new_n6276_), .Y(new_n6690_));
  AOI21X1  g06498(.A0(new_n6277_), .A1(new_n6272_), .B0(new_n193_), .Y(new_n6691_));
  OAI21X1  g06499(.A0(new_n6690_), .A1(new_n6272_), .B0(new_n6691_), .Y(new_n6692_));
  OR2X1    g06500(.A(new_n6283_), .B(new_n6282_), .Y(new_n6693_));
  AND2X1   g06501(.A(new_n6275_), .B(new_n5923_), .Y(new_n6694_));
  NOR4X1   g06502(.A(new_n6290_), .B(new_n6330_), .C(new_n6694_), .D(new_n6274_), .Y(new_n6695_));
  NAND3X1  g06503(.A(new_n6695_), .B(new_n6693_), .C(new_n6309_), .Y(new_n6696_));
  AND2X1   g06504(.A(new_n6696_), .B(new_n6692_), .Y(new_n6697_));
  OAI21X1  g06505(.A0(new_n6689_), .A1(new_n6679_), .B0(new_n6697_), .Y(new_n6698_));
  AOI21X1  g06506(.A0(new_n6687_), .A1(new_n193_), .B0(new_n6698_), .Y(new_n6699_));
  OR2X1    g06507(.A(new_n6688_), .B(new_n199_), .Y(new_n6700_));
  AND2X1   g06508(.A(new_n6670_), .B(new_n6661_), .Y(new_n6701_));
  INVX1    g06509(.A(new_n6676_), .Y(new_n6702_));
  OR2X1    g06510(.A(new_n6677_), .B(\asqrt[62] ), .Y(new_n6703_));
  OAI21X1  g06511(.A0(new_n6703_), .A1(new_n6701_), .B0(new_n6702_), .Y(new_n6704_));
  INVX1    g06512(.A(new_n6686_), .Y(new_n6705_));
  AOI21X1  g06513(.A0(new_n6704_), .A1(new_n6700_), .B0(new_n6705_), .Y(new_n6706_));
  AOI21X1  g06514(.A0(new_n6659_), .A1(\asqrt[62] ), .B0(new_n6683_), .Y(new_n6707_));
  INVX1    g06515(.A(new_n6697_), .Y(new_n6708_));
  AOI21X1  g06516(.A0(new_n6707_), .A1(new_n6704_), .B0(new_n6708_), .Y(new_n6709_));
  OAI21X1  g06517(.A0(new_n6706_), .A1(\asqrt[63] ), .B0(new_n6709_), .Y(\asqrt[32] ));
  NOR2X1   g06518(.A(\a[63] ), .B(\a[62] ), .Y(new_n6711_));
  MX2X1    g06519(.A(new_n6711_), .B(\asqrt[32] ), .S0(\a[64] ), .Y(new_n6712_));
  AND2X1   g06520(.A(new_n6712_), .B(\asqrt[33] ), .Y(new_n6713_));
  INVX1    g06521(.A(\a[64] ), .Y(new_n6714_));
  INVX1    g06522(.A(\a[65] ), .Y(new_n6715_));
  AOI21X1  g06523(.A0(\asqrt[32] ), .A1(new_n6714_), .B0(new_n6715_), .Y(new_n6716_));
  NOR2X1   g06524(.A(\a[65] ), .B(\a[64] ), .Y(new_n6717_));
  AND2X1   g06525(.A(\asqrt[32] ), .B(new_n6717_), .Y(new_n6718_));
  NOR3X1   g06526(.A(\a[64] ), .B(\a[63] ), .C(\a[62] ), .Y(new_n6719_));
  NOR3X1   g06527(.A(new_n6719_), .B(new_n6290_), .C(new_n6330_), .Y(new_n6720_));
  NAND3X1  g06528(.A(new_n6720_), .B(new_n6693_), .C(new_n6309_), .Y(new_n6721_));
  AOI21X1  g06529(.A0(\asqrt[32] ), .A1(\a[64] ), .B0(new_n6721_), .Y(new_n6722_));
  NOR3X1   g06530(.A(new_n6722_), .B(new_n6718_), .C(new_n6716_), .Y(new_n6723_));
  OAI21X1  g06531(.A0(new_n6723_), .A1(new_n6713_), .B0(\asqrt[34] ), .Y(new_n6724_));
  INVX1    g06532(.A(new_n6711_), .Y(new_n6725_));
  MX2X1    g06533(.A(new_n6725_), .B(new_n6699_), .S0(\a[64] ), .Y(new_n6726_));
  OAI21X1  g06534(.A0(new_n6726_), .A1(new_n6294_), .B0(new_n5941_), .Y(new_n6727_));
  NAND3X1  g06535(.A(new_n6696_), .B(new_n6692_), .C(\asqrt[33] ), .Y(new_n6728_));
  INVX1    g06536(.A(new_n6728_), .Y(new_n6729_));
  OAI21X1  g06537(.A0(new_n6689_), .A1(new_n6679_), .B0(new_n6729_), .Y(new_n6730_));
  AOI21X1  g06538(.A0(new_n6687_), .A1(new_n193_), .B0(new_n6730_), .Y(new_n6731_));
  AOI21X1  g06539(.A0(\asqrt[32] ), .A1(new_n6717_), .B0(new_n6731_), .Y(new_n6732_));
  OR2X1    g06540(.A(new_n6731_), .B(\a[66] ), .Y(new_n6733_));
  OAI22X1  g06541(.A0(new_n6733_), .A1(new_n6718_), .B0(new_n6732_), .B1(new_n6295_), .Y(new_n6734_));
  OAI21X1  g06542(.A0(new_n6727_), .A1(new_n6723_), .B0(new_n6734_), .Y(new_n6735_));
  AOI21X1  g06543(.A0(new_n6735_), .A1(new_n6724_), .B0(new_n5541_), .Y(new_n6736_));
  AND2X1   g06544(.A(new_n6320_), .B(new_n6327_), .Y(new_n6737_));
  NAND3X1  g06545(.A(new_n6737_), .B(\asqrt[32] ), .C(new_n6349_), .Y(new_n6738_));
  INVX1    g06546(.A(new_n6737_), .Y(new_n6739_));
  OAI21X1  g06547(.A0(new_n6739_), .A1(new_n6699_), .B0(new_n6323_), .Y(new_n6740_));
  AND2X1   g06548(.A(new_n6740_), .B(new_n6738_), .Y(new_n6741_));
  INVX1    g06549(.A(new_n6741_), .Y(new_n6742_));
  NAND3X1  g06550(.A(new_n6735_), .B(new_n6724_), .C(new_n5541_), .Y(new_n6743_));
  AOI21X1  g06551(.A0(new_n6743_), .A1(new_n6742_), .B0(new_n6736_), .Y(new_n6744_));
  OR2X1    g06552(.A(new_n6744_), .B(new_n5176_), .Y(new_n6745_));
  AND2X1   g06553(.A(new_n6743_), .B(new_n6742_), .Y(new_n6746_));
  AOI21X1  g06554(.A0(new_n6379_), .A1(new_n6378_), .B0(new_n6337_), .Y(new_n6747_));
  NAND3X1  g06555(.A(new_n6747_), .B(\asqrt[32] ), .C(new_n6325_), .Y(new_n6748_));
  OAI22X1  g06556(.A0(new_n6328_), .A1(new_n6326_), .B0(new_n6324_), .B1(new_n5541_), .Y(new_n6749_));
  OAI21X1  g06557(.A0(new_n6749_), .A1(new_n6699_), .B0(new_n6337_), .Y(new_n6750_));
  AND2X1   g06558(.A(new_n6750_), .B(new_n6748_), .Y(new_n6751_));
  INVX1    g06559(.A(new_n6751_), .Y(new_n6752_));
  OR2X1    g06560(.A(new_n6736_), .B(\asqrt[36] ), .Y(new_n6753_));
  OAI21X1  g06561(.A0(new_n6753_), .A1(new_n6746_), .B0(new_n6752_), .Y(new_n6754_));
  AOI21X1  g06562(.A0(new_n6754_), .A1(new_n6745_), .B0(new_n4826_), .Y(new_n6755_));
  AND2X1   g06563(.A(new_n6351_), .B(new_n6338_), .Y(new_n6756_));
  OR4X1    g06564(.A(new_n6699_), .B(new_n6756_), .C(new_n6383_), .D(new_n6339_), .Y(new_n6757_));
  OR2X1    g06565(.A(new_n6756_), .B(new_n6339_), .Y(new_n6758_));
  OAI21X1  g06566(.A0(new_n6758_), .A1(new_n6699_), .B0(new_n6383_), .Y(new_n6759_));
  AND2X1   g06567(.A(new_n6759_), .B(new_n6757_), .Y(new_n6760_));
  OR2X1    g06568(.A(new_n6726_), .B(new_n6294_), .Y(new_n6761_));
  OAI21X1  g06569(.A0(new_n6699_), .A1(\a[64] ), .B0(\a[65] ), .Y(new_n6762_));
  INVX1    g06570(.A(new_n6717_), .Y(new_n6763_));
  OR2X1    g06571(.A(new_n6699_), .B(new_n6763_), .Y(new_n6764_));
  INVX1    g06572(.A(new_n6721_), .Y(new_n6765_));
  OAI21X1  g06573(.A0(new_n6699_), .A1(new_n6714_), .B0(new_n6765_), .Y(new_n6766_));
  NAND3X1  g06574(.A(new_n6766_), .B(new_n6764_), .C(new_n6762_), .Y(new_n6767_));
  AOI21X1  g06575(.A0(new_n6767_), .A1(new_n6761_), .B0(new_n5941_), .Y(new_n6768_));
  AOI21X1  g06576(.A0(new_n6712_), .A1(\asqrt[33] ), .B0(\asqrt[34] ), .Y(new_n6769_));
  OR2X1    g06577(.A(new_n6732_), .B(new_n6295_), .Y(new_n6770_));
  OR2X1    g06578(.A(new_n6733_), .B(new_n6718_), .Y(new_n6771_));
  AOI22X1  g06579(.A0(new_n6771_), .A1(new_n6770_), .B0(new_n6769_), .B1(new_n6767_), .Y(new_n6772_));
  OAI21X1  g06580(.A0(new_n6772_), .A1(new_n6768_), .B0(\asqrt[35] ), .Y(new_n6773_));
  NOR3X1   g06581(.A(new_n6772_), .B(new_n6768_), .C(\asqrt[35] ), .Y(new_n6774_));
  OAI21X1  g06582(.A0(new_n6774_), .A1(new_n6741_), .B0(new_n6773_), .Y(new_n6775_));
  AOI21X1  g06583(.A0(new_n6775_), .A1(\asqrt[36] ), .B0(\asqrt[37] ), .Y(new_n6776_));
  AOI21X1  g06584(.A0(new_n6776_), .A1(new_n6754_), .B0(new_n6760_), .Y(new_n6777_));
  OAI21X1  g06585(.A0(new_n6777_), .A1(new_n6755_), .B0(\asqrt[38] ), .Y(new_n6778_));
  NAND3X1  g06586(.A(new_n6388_), .B(new_n6360_), .C(new_n6353_), .Y(new_n6779_));
  NOR3X1   g06587(.A(new_n6699_), .B(new_n6361_), .C(new_n6386_), .Y(new_n6780_));
  OAI22X1  g06588(.A0(new_n6780_), .A1(new_n6360_), .B0(new_n6779_), .B1(new_n6699_), .Y(new_n6781_));
  INVX1    g06589(.A(new_n6781_), .Y(new_n6782_));
  NOR3X1   g06590(.A(new_n6777_), .B(new_n6755_), .C(\asqrt[38] ), .Y(new_n6783_));
  OAI21X1  g06591(.A0(new_n6783_), .A1(new_n6782_), .B0(new_n6778_), .Y(new_n6784_));
  AND2X1   g06592(.A(new_n6784_), .B(\asqrt[39] ), .Y(new_n6785_));
  AND2X1   g06593(.A(new_n6775_), .B(\asqrt[36] ), .Y(new_n6786_));
  NAND2X1  g06594(.A(new_n6743_), .B(new_n6742_), .Y(new_n6787_));
  NOR2X1   g06595(.A(new_n6736_), .B(\asqrt[36] ), .Y(new_n6788_));
  AOI21X1  g06596(.A0(new_n6788_), .A1(new_n6787_), .B0(new_n6751_), .Y(new_n6789_));
  OAI21X1  g06597(.A0(new_n6789_), .A1(new_n6786_), .B0(\asqrt[37] ), .Y(new_n6790_));
  INVX1    g06598(.A(new_n6760_), .Y(new_n6791_));
  OAI21X1  g06599(.A0(new_n6744_), .A1(new_n5176_), .B0(new_n4826_), .Y(new_n6792_));
  OAI21X1  g06600(.A0(new_n6792_), .A1(new_n6789_), .B0(new_n6791_), .Y(new_n6793_));
  NAND3X1  g06601(.A(new_n6793_), .B(new_n6790_), .C(new_n4493_), .Y(new_n6794_));
  NAND2X1  g06602(.A(new_n6794_), .B(new_n6781_), .Y(new_n6795_));
  AND2X1   g06603(.A(new_n6371_), .B(new_n6364_), .Y(new_n6796_));
  NOR4X1   g06604(.A(new_n6699_), .B(new_n6796_), .C(new_n6411_), .D(new_n6363_), .Y(new_n6797_));
  AOI22X1  g06605(.A0(new_n6371_), .A1(new_n6364_), .B0(new_n6362_), .B1(\asqrt[38] ), .Y(new_n6798_));
  AOI21X1  g06606(.A0(new_n6798_), .A1(\asqrt[32] ), .B0(new_n6370_), .Y(new_n6799_));
  NOR2X1   g06607(.A(new_n6799_), .B(new_n6797_), .Y(new_n6800_));
  AOI21X1  g06608(.A0(new_n6793_), .A1(new_n6790_), .B0(new_n4493_), .Y(new_n6801_));
  NOR2X1   g06609(.A(new_n6801_), .B(\asqrt[39] ), .Y(new_n6802_));
  AOI21X1  g06610(.A0(new_n6802_), .A1(new_n6795_), .B0(new_n6800_), .Y(new_n6803_));
  OAI21X1  g06611(.A0(new_n6803_), .A1(new_n6785_), .B0(\asqrt[40] ), .Y(new_n6804_));
  AND2X1   g06612(.A(new_n6416_), .B(new_n6413_), .Y(new_n6805_));
  OR4X1    g06613(.A(new_n6699_), .B(new_n6805_), .C(new_n6376_), .D(new_n6414_), .Y(new_n6806_));
  OR2X1    g06614(.A(new_n6805_), .B(new_n6414_), .Y(new_n6807_));
  OAI21X1  g06615(.A0(new_n6807_), .A1(new_n6699_), .B0(new_n6376_), .Y(new_n6808_));
  AND2X1   g06616(.A(new_n6808_), .B(new_n6806_), .Y(new_n6809_));
  INVX1    g06617(.A(new_n6809_), .Y(new_n6810_));
  AOI21X1  g06618(.A0(new_n6794_), .A1(new_n6781_), .B0(new_n6801_), .Y(new_n6811_));
  OAI21X1  g06619(.A0(new_n6811_), .A1(new_n4165_), .B0(new_n3863_), .Y(new_n6812_));
  OAI21X1  g06620(.A0(new_n6812_), .A1(new_n6803_), .B0(new_n6810_), .Y(new_n6813_));
  AOI21X1  g06621(.A0(new_n6813_), .A1(new_n6804_), .B0(new_n3564_), .Y(new_n6814_));
  OR4X1    g06622(.A(new_n6699_), .B(new_n6426_), .C(new_n6398_), .D(new_n6392_), .Y(new_n6815_));
  NAND2X1  g06623(.A(new_n6399_), .B(new_n6418_), .Y(new_n6816_));
  OAI21X1  g06624(.A0(new_n6816_), .A1(new_n6699_), .B0(new_n6398_), .Y(new_n6817_));
  AND2X1   g06625(.A(new_n6817_), .B(new_n6815_), .Y(new_n6818_));
  INVX1    g06626(.A(new_n6818_), .Y(new_n6819_));
  NAND3X1  g06627(.A(new_n6813_), .B(new_n6804_), .C(new_n3564_), .Y(new_n6820_));
  AOI21X1  g06628(.A0(new_n6820_), .A1(new_n6819_), .B0(new_n6814_), .Y(new_n6821_));
  OR2X1    g06629(.A(new_n6821_), .B(new_n3276_), .Y(new_n6822_));
  AND2X1   g06630(.A(new_n6820_), .B(new_n6819_), .Y(new_n6823_));
  OAI21X1  g06631(.A0(new_n6419_), .A1(new_n6402_), .B0(new_n6407_), .Y(new_n6824_));
  NOR3X1   g06632(.A(new_n6824_), .B(new_n6699_), .C(new_n6440_), .Y(new_n6825_));
  AOI22X1  g06633(.A0(new_n6442_), .A1(new_n6441_), .B0(new_n6427_), .B1(\asqrt[41] ), .Y(new_n6826_));
  AOI21X1  g06634(.A0(new_n6826_), .A1(\asqrt[32] ), .B0(new_n6407_), .Y(new_n6827_));
  NOR2X1   g06635(.A(new_n6827_), .B(new_n6825_), .Y(new_n6828_));
  INVX1    g06636(.A(new_n6828_), .Y(new_n6829_));
  OR2X1    g06637(.A(new_n6814_), .B(\asqrt[42] ), .Y(new_n6830_));
  OAI21X1  g06638(.A0(new_n6830_), .A1(new_n6823_), .B0(new_n6829_), .Y(new_n6831_));
  AOI21X1  g06639(.A0(new_n6831_), .A1(new_n6822_), .B0(new_n3008_), .Y(new_n6832_));
  AND2X1   g06640(.A(new_n6428_), .B(new_n6420_), .Y(new_n6833_));
  OR4X1    g06641(.A(new_n6699_), .B(new_n6833_), .C(new_n6445_), .D(new_n6421_), .Y(new_n6834_));
  OR2X1    g06642(.A(new_n6833_), .B(new_n6421_), .Y(new_n6835_));
  OAI21X1  g06643(.A0(new_n6835_), .A1(new_n6699_), .B0(new_n6445_), .Y(new_n6836_));
  AND2X1   g06644(.A(new_n6836_), .B(new_n6834_), .Y(new_n6837_));
  OR2X1    g06645(.A(new_n6811_), .B(new_n4165_), .Y(new_n6838_));
  AND2X1   g06646(.A(new_n6794_), .B(new_n6781_), .Y(new_n6839_));
  INVX1    g06647(.A(new_n6800_), .Y(new_n6840_));
  OR2X1    g06648(.A(new_n6801_), .B(\asqrt[39] ), .Y(new_n6841_));
  OAI21X1  g06649(.A0(new_n6841_), .A1(new_n6839_), .B0(new_n6840_), .Y(new_n6842_));
  AOI21X1  g06650(.A0(new_n6842_), .A1(new_n6838_), .B0(new_n3863_), .Y(new_n6843_));
  AOI21X1  g06651(.A0(new_n6784_), .A1(\asqrt[39] ), .B0(\asqrt[40] ), .Y(new_n6844_));
  AOI21X1  g06652(.A0(new_n6844_), .A1(new_n6842_), .B0(new_n6809_), .Y(new_n6845_));
  OAI21X1  g06653(.A0(new_n6845_), .A1(new_n6843_), .B0(\asqrt[41] ), .Y(new_n6846_));
  NOR3X1   g06654(.A(new_n6845_), .B(new_n6843_), .C(\asqrt[41] ), .Y(new_n6847_));
  OAI21X1  g06655(.A0(new_n6847_), .A1(new_n6818_), .B0(new_n6846_), .Y(new_n6848_));
  AOI21X1  g06656(.A0(new_n6848_), .A1(\asqrt[42] ), .B0(\asqrt[43] ), .Y(new_n6849_));
  AOI21X1  g06657(.A0(new_n6849_), .A1(new_n6831_), .B0(new_n6837_), .Y(new_n6850_));
  OAI21X1  g06658(.A0(new_n6850_), .A1(new_n6832_), .B0(\asqrt[44] ), .Y(new_n6851_));
  OR4X1    g06659(.A(new_n6699_), .B(new_n6436_), .C(new_n6439_), .D(new_n6463_), .Y(new_n6852_));
  NAND2X1  g06660(.A(new_n6448_), .B(new_n6430_), .Y(new_n6853_));
  OAI21X1  g06661(.A0(new_n6853_), .A1(new_n6699_), .B0(new_n6439_), .Y(new_n6854_));
  AND2X1   g06662(.A(new_n6854_), .B(new_n6852_), .Y(new_n6855_));
  NOR3X1   g06663(.A(new_n6850_), .B(new_n6832_), .C(\asqrt[44] ), .Y(new_n6856_));
  OAI21X1  g06664(.A0(new_n6856_), .A1(new_n6855_), .B0(new_n6851_), .Y(new_n6857_));
  AND2X1   g06665(.A(new_n6857_), .B(\asqrt[45] ), .Y(new_n6858_));
  INVX1    g06666(.A(new_n6855_), .Y(new_n6859_));
  AND2X1   g06667(.A(new_n6848_), .B(\asqrt[42] ), .Y(new_n6860_));
  NAND2X1  g06668(.A(new_n6820_), .B(new_n6819_), .Y(new_n6861_));
  NOR2X1   g06669(.A(new_n6814_), .B(\asqrt[42] ), .Y(new_n6862_));
  AOI21X1  g06670(.A0(new_n6862_), .A1(new_n6861_), .B0(new_n6828_), .Y(new_n6863_));
  OAI21X1  g06671(.A0(new_n6863_), .A1(new_n6860_), .B0(\asqrt[43] ), .Y(new_n6864_));
  INVX1    g06672(.A(new_n6837_), .Y(new_n6865_));
  OAI21X1  g06673(.A0(new_n6821_), .A1(new_n3276_), .B0(new_n3008_), .Y(new_n6866_));
  OAI21X1  g06674(.A0(new_n6866_), .A1(new_n6863_), .B0(new_n6865_), .Y(new_n6867_));
  NAND3X1  g06675(.A(new_n6867_), .B(new_n6864_), .C(new_n2769_), .Y(new_n6868_));
  NAND2X1  g06676(.A(new_n6868_), .B(new_n6859_), .Y(new_n6869_));
  AND2X1   g06677(.A(new_n6455_), .B(new_n6449_), .Y(new_n6870_));
  NOR4X1   g06678(.A(new_n6699_), .B(new_n6870_), .C(new_n6486_), .D(new_n6438_), .Y(new_n6871_));
  AOI22X1  g06679(.A0(new_n6455_), .A1(new_n6449_), .B0(new_n6437_), .B1(\asqrt[44] ), .Y(new_n6872_));
  AOI21X1  g06680(.A0(new_n6872_), .A1(\asqrt[32] ), .B0(new_n6454_), .Y(new_n6873_));
  NOR2X1   g06681(.A(new_n6873_), .B(new_n6871_), .Y(new_n6874_));
  AOI21X1  g06682(.A0(new_n6867_), .A1(new_n6864_), .B0(new_n2769_), .Y(new_n6875_));
  NOR2X1   g06683(.A(new_n6875_), .B(\asqrt[45] ), .Y(new_n6876_));
  AOI21X1  g06684(.A0(new_n6876_), .A1(new_n6869_), .B0(new_n6874_), .Y(new_n6877_));
  OAI21X1  g06685(.A0(new_n6877_), .A1(new_n6858_), .B0(\asqrt[46] ), .Y(new_n6878_));
  AND2X1   g06686(.A(new_n6490_), .B(new_n6488_), .Y(new_n6879_));
  OR4X1    g06687(.A(new_n6699_), .B(new_n6879_), .C(new_n6462_), .D(new_n6489_), .Y(new_n6880_));
  OR2X1    g06688(.A(new_n6879_), .B(new_n6489_), .Y(new_n6881_));
  OAI21X1  g06689(.A0(new_n6881_), .A1(new_n6699_), .B0(new_n6462_), .Y(new_n6882_));
  AND2X1   g06690(.A(new_n6882_), .B(new_n6880_), .Y(new_n6883_));
  INVX1    g06691(.A(new_n6883_), .Y(new_n6884_));
  AOI21X1  g06692(.A0(new_n6868_), .A1(new_n6859_), .B0(new_n6875_), .Y(new_n6885_));
  OAI21X1  g06693(.A0(new_n6885_), .A1(new_n2570_), .B0(new_n2263_), .Y(new_n6886_));
  OAI21X1  g06694(.A0(new_n6886_), .A1(new_n6877_), .B0(new_n6884_), .Y(new_n6887_));
  AOI21X1  g06695(.A0(new_n6887_), .A1(new_n6878_), .B0(new_n2040_), .Y(new_n6888_));
  OR4X1    g06696(.A(new_n6699_), .B(new_n6500_), .C(new_n6473_), .D(new_n6467_), .Y(new_n6889_));
  NAND2X1  g06697(.A(new_n6474_), .B(new_n6492_), .Y(new_n6890_));
  OAI21X1  g06698(.A0(new_n6890_), .A1(new_n6699_), .B0(new_n6473_), .Y(new_n6891_));
  AND2X1   g06699(.A(new_n6891_), .B(new_n6889_), .Y(new_n6892_));
  INVX1    g06700(.A(new_n6892_), .Y(new_n6893_));
  NAND3X1  g06701(.A(new_n6887_), .B(new_n6878_), .C(new_n2040_), .Y(new_n6894_));
  AOI21X1  g06702(.A0(new_n6894_), .A1(new_n6893_), .B0(new_n6888_), .Y(new_n6895_));
  OR2X1    g06703(.A(new_n6895_), .B(new_n1834_), .Y(new_n6896_));
  AND2X1   g06704(.A(new_n6894_), .B(new_n6893_), .Y(new_n6897_));
  OAI21X1  g06705(.A0(new_n6493_), .A1(new_n6477_), .B0(new_n6482_), .Y(new_n6898_));
  NOR3X1   g06706(.A(new_n6898_), .B(new_n6699_), .C(new_n6514_), .Y(new_n6899_));
  AOI22X1  g06707(.A0(new_n6516_), .A1(new_n6515_), .B0(new_n6501_), .B1(\asqrt[47] ), .Y(new_n6900_));
  AOI21X1  g06708(.A0(new_n6900_), .A1(\asqrt[32] ), .B0(new_n6482_), .Y(new_n6901_));
  NOR2X1   g06709(.A(new_n6901_), .B(new_n6899_), .Y(new_n6902_));
  INVX1    g06710(.A(new_n6902_), .Y(new_n6903_));
  OR2X1    g06711(.A(new_n6888_), .B(\asqrt[48] ), .Y(new_n6904_));
  OAI21X1  g06712(.A0(new_n6904_), .A1(new_n6897_), .B0(new_n6903_), .Y(new_n6905_));
  AOI21X1  g06713(.A0(new_n6905_), .A1(new_n6896_), .B0(new_n1632_), .Y(new_n6906_));
  AND2X1   g06714(.A(new_n6502_), .B(new_n6494_), .Y(new_n6907_));
  OR4X1    g06715(.A(new_n6699_), .B(new_n6907_), .C(new_n6519_), .D(new_n6495_), .Y(new_n6908_));
  OR2X1    g06716(.A(new_n6907_), .B(new_n6495_), .Y(new_n6909_));
  OAI21X1  g06717(.A0(new_n6909_), .A1(new_n6699_), .B0(new_n6519_), .Y(new_n6910_));
  AND2X1   g06718(.A(new_n6910_), .B(new_n6908_), .Y(new_n6911_));
  OR2X1    g06719(.A(new_n6885_), .B(new_n2570_), .Y(new_n6912_));
  AND2X1   g06720(.A(new_n6868_), .B(new_n6859_), .Y(new_n6913_));
  INVX1    g06721(.A(new_n6874_), .Y(new_n6914_));
  OR2X1    g06722(.A(new_n6875_), .B(\asqrt[45] ), .Y(new_n6915_));
  OAI21X1  g06723(.A0(new_n6915_), .A1(new_n6913_), .B0(new_n6914_), .Y(new_n6916_));
  AOI21X1  g06724(.A0(new_n6916_), .A1(new_n6912_), .B0(new_n2263_), .Y(new_n6917_));
  AOI21X1  g06725(.A0(new_n6857_), .A1(\asqrt[45] ), .B0(\asqrt[46] ), .Y(new_n6918_));
  AOI21X1  g06726(.A0(new_n6918_), .A1(new_n6916_), .B0(new_n6883_), .Y(new_n6919_));
  OAI21X1  g06727(.A0(new_n6919_), .A1(new_n6917_), .B0(\asqrt[47] ), .Y(new_n6920_));
  NOR3X1   g06728(.A(new_n6919_), .B(new_n6917_), .C(\asqrt[47] ), .Y(new_n6921_));
  OAI21X1  g06729(.A0(new_n6921_), .A1(new_n6892_), .B0(new_n6920_), .Y(new_n6922_));
  AOI21X1  g06730(.A0(new_n6922_), .A1(\asqrt[48] ), .B0(\asqrt[49] ), .Y(new_n6923_));
  AOI21X1  g06731(.A0(new_n6923_), .A1(new_n6905_), .B0(new_n6911_), .Y(new_n6924_));
  OAI21X1  g06732(.A0(new_n6924_), .A1(new_n6906_), .B0(\asqrt[50] ), .Y(new_n6925_));
  OR4X1    g06733(.A(new_n6699_), .B(new_n6510_), .C(new_n6513_), .D(new_n6537_), .Y(new_n6926_));
  NAND2X1  g06734(.A(new_n6522_), .B(new_n6504_), .Y(new_n6927_));
  OAI21X1  g06735(.A0(new_n6927_), .A1(new_n6699_), .B0(new_n6513_), .Y(new_n6928_));
  AND2X1   g06736(.A(new_n6928_), .B(new_n6926_), .Y(new_n6929_));
  NOR3X1   g06737(.A(new_n6924_), .B(new_n6906_), .C(\asqrt[50] ), .Y(new_n6930_));
  OAI21X1  g06738(.A0(new_n6930_), .A1(new_n6929_), .B0(new_n6925_), .Y(new_n6931_));
  AND2X1   g06739(.A(new_n6931_), .B(\asqrt[51] ), .Y(new_n6932_));
  INVX1    g06740(.A(new_n6929_), .Y(new_n6933_));
  AND2X1   g06741(.A(new_n6922_), .B(\asqrt[48] ), .Y(new_n6934_));
  NAND2X1  g06742(.A(new_n6894_), .B(new_n6893_), .Y(new_n6935_));
  NOR2X1   g06743(.A(new_n6888_), .B(\asqrt[48] ), .Y(new_n6936_));
  AOI21X1  g06744(.A0(new_n6936_), .A1(new_n6935_), .B0(new_n6902_), .Y(new_n6937_));
  OAI21X1  g06745(.A0(new_n6937_), .A1(new_n6934_), .B0(\asqrt[49] ), .Y(new_n6938_));
  INVX1    g06746(.A(new_n6911_), .Y(new_n6939_));
  OAI21X1  g06747(.A0(new_n6895_), .A1(new_n1834_), .B0(new_n1632_), .Y(new_n6940_));
  OAI21X1  g06748(.A0(new_n6940_), .A1(new_n6937_), .B0(new_n6939_), .Y(new_n6941_));
  NAND3X1  g06749(.A(new_n6941_), .B(new_n6938_), .C(new_n1469_), .Y(new_n6942_));
  NAND2X1  g06750(.A(new_n6942_), .B(new_n6933_), .Y(new_n6943_));
  AND2X1   g06751(.A(new_n6529_), .B(new_n6523_), .Y(new_n6944_));
  NOR4X1   g06752(.A(new_n6699_), .B(new_n6944_), .C(new_n6560_), .D(new_n6512_), .Y(new_n6945_));
  AOI22X1  g06753(.A0(new_n6529_), .A1(new_n6523_), .B0(new_n6511_), .B1(\asqrt[50] ), .Y(new_n6946_));
  AOI21X1  g06754(.A0(new_n6946_), .A1(\asqrt[32] ), .B0(new_n6528_), .Y(new_n6947_));
  NOR2X1   g06755(.A(new_n6947_), .B(new_n6945_), .Y(new_n6948_));
  AOI21X1  g06756(.A0(new_n6941_), .A1(new_n6938_), .B0(new_n1469_), .Y(new_n6949_));
  NOR2X1   g06757(.A(new_n6949_), .B(\asqrt[51] ), .Y(new_n6950_));
  AOI21X1  g06758(.A0(new_n6950_), .A1(new_n6943_), .B0(new_n6948_), .Y(new_n6951_));
  OAI21X1  g06759(.A0(new_n6951_), .A1(new_n6932_), .B0(\asqrt[52] ), .Y(new_n6952_));
  AND2X1   g06760(.A(new_n6564_), .B(new_n6562_), .Y(new_n6953_));
  NOR4X1   g06761(.A(new_n6699_), .B(new_n6953_), .C(new_n6536_), .D(new_n6563_), .Y(new_n6954_));
  NOR2X1   g06762(.A(new_n6953_), .B(new_n6563_), .Y(new_n6955_));
  AOI21X1  g06763(.A0(new_n6955_), .A1(\asqrt[32] ), .B0(new_n6535_), .Y(new_n6956_));
  NOR2X1   g06764(.A(new_n6956_), .B(new_n6954_), .Y(new_n6957_));
  INVX1    g06765(.A(new_n6957_), .Y(new_n6958_));
  AOI21X1  g06766(.A0(new_n6942_), .A1(new_n6933_), .B0(new_n6949_), .Y(new_n6959_));
  OAI21X1  g06767(.A0(new_n6959_), .A1(new_n1277_), .B0(new_n1111_), .Y(new_n6960_));
  OAI21X1  g06768(.A0(new_n6960_), .A1(new_n6951_), .B0(new_n6958_), .Y(new_n6961_));
  AOI21X1  g06769(.A0(new_n6961_), .A1(new_n6952_), .B0(new_n968_), .Y(new_n6962_));
  OR4X1    g06770(.A(new_n6699_), .B(new_n6574_), .C(new_n6547_), .D(new_n6541_), .Y(new_n6963_));
  NAND2X1  g06771(.A(new_n6548_), .B(new_n6566_), .Y(new_n6964_));
  OAI21X1  g06772(.A0(new_n6964_), .A1(new_n6699_), .B0(new_n6547_), .Y(new_n6965_));
  AND2X1   g06773(.A(new_n6965_), .B(new_n6963_), .Y(new_n6966_));
  INVX1    g06774(.A(new_n6966_), .Y(new_n6967_));
  NAND3X1  g06775(.A(new_n6961_), .B(new_n6952_), .C(new_n968_), .Y(new_n6968_));
  AOI21X1  g06776(.A0(new_n6968_), .A1(new_n6967_), .B0(new_n6962_), .Y(new_n6969_));
  OR2X1    g06777(.A(new_n6969_), .B(new_n902_), .Y(new_n6970_));
  AND2X1   g06778(.A(new_n6968_), .B(new_n6967_), .Y(new_n6971_));
  OAI21X1  g06779(.A0(new_n6567_), .A1(new_n6551_), .B0(new_n6556_), .Y(new_n6972_));
  NOR3X1   g06780(.A(new_n6972_), .B(new_n6699_), .C(new_n6588_), .Y(new_n6973_));
  AOI22X1  g06781(.A0(new_n6590_), .A1(new_n6589_), .B0(new_n6575_), .B1(\asqrt[53] ), .Y(new_n6974_));
  AOI21X1  g06782(.A0(new_n6974_), .A1(\asqrt[32] ), .B0(new_n6556_), .Y(new_n6975_));
  NOR2X1   g06783(.A(new_n6975_), .B(new_n6973_), .Y(new_n6976_));
  INVX1    g06784(.A(new_n6976_), .Y(new_n6977_));
  OR2X1    g06785(.A(new_n6962_), .B(\asqrt[54] ), .Y(new_n6978_));
  OAI21X1  g06786(.A0(new_n6978_), .A1(new_n6971_), .B0(new_n6977_), .Y(new_n6979_));
  AOI21X1  g06787(.A0(new_n6979_), .A1(new_n6970_), .B0(new_n697_), .Y(new_n6980_));
  AND2X1   g06788(.A(new_n6576_), .B(new_n6568_), .Y(new_n6981_));
  OR4X1    g06789(.A(new_n6699_), .B(new_n6981_), .C(new_n6593_), .D(new_n6569_), .Y(new_n6982_));
  OR2X1    g06790(.A(new_n6981_), .B(new_n6569_), .Y(new_n6983_));
  OAI21X1  g06791(.A0(new_n6983_), .A1(new_n6699_), .B0(new_n6593_), .Y(new_n6984_));
  AND2X1   g06792(.A(new_n6984_), .B(new_n6982_), .Y(new_n6985_));
  OR2X1    g06793(.A(new_n6959_), .B(new_n1277_), .Y(new_n6986_));
  AND2X1   g06794(.A(new_n6942_), .B(new_n6933_), .Y(new_n6987_));
  INVX1    g06795(.A(new_n6948_), .Y(new_n6988_));
  OR2X1    g06796(.A(new_n6949_), .B(\asqrt[51] ), .Y(new_n6989_));
  OAI21X1  g06797(.A0(new_n6989_), .A1(new_n6987_), .B0(new_n6988_), .Y(new_n6990_));
  AOI21X1  g06798(.A0(new_n6990_), .A1(new_n6986_), .B0(new_n1111_), .Y(new_n6991_));
  AOI21X1  g06799(.A0(new_n6931_), .A1(\asqrt[51] ), .B0(\asqrt[52] ), .Y(new_n6992_));
  AOI21X1  g06800(.A0(new_n6992_), .A1(new_n6990_), .B0(new_n6957_), .Y(new_n6993_));
  OAI21X1  g06801(.A0(new_n6993_), .A1(new_n6991_), .B0(\asqrt[53] ), .Y(new_n6994_));
  NOR3X1   g06802(.A(new_n6993_), .B(new_n6991_), .C(\asqrt[53] ), .Y(new_n6995_));
  OAI21X1  g06803(.A0(new_n6995_), .A1(new_n6966_), .B0(new_n6994_), .Y(new_n6996_));
  AOI21X1  g06804(.A0(new_n6996_), .A1(\asqrt[54] ), .B0(\asqrt[55] ), .Y(new_n6997_));
  AOI21X1  g06805(.A0(new_n6997_), .A1(new_n6979_), .B0(new_n6985_), .Y(new_n6998_));
  OAI21X1  g06806(.A0(new_n6998_), .A1(new_n6980_), .B0(\asqrt[56] ), .Y(new_n6999_));
  NAND3X1  g06807(.A(new_n6596_), .B(new_n6583_), .C(new_n6578_), .Y(new_n7000_));
  NOR3X1   g06808(.A(new_n6699_), .B(new_n6584_), .C(new_n6611_), .Y(new_n7001_));
  OAI22X1  g06809(.A0(new_n7001_), .A1(new_n6583_), .B0(new_n7000_), .B1(new_n6699_), .Y(new_n7002_));
  INVX1    g06810(.A(new_n7002_), .Y(new_n7003_));
  NOR3X1   g06811(.A(new_n6998_), .B(new_n6980_), .C(\asqrt[56] ), .Y(new_n7004_));
  OAI21X1  g06812(.A0(new_n7004_), .A1(new_n7003_), .B0(new_n6999_), .Y(new_n7005_));
  AND2X1   g06813(.A(new_n7005_), .B(\asqrt[57] ), .Y(new_n7006_));
  AND2X1   g06814(.A(new_n6996_), .B(\asqrt[54] ), .Y(new_n7007_));
  NAND2X1  g06815(.A(new_n6968_), .B(new_n6967_), .Y(new_n7008_));
  NOR2X1   g06816(.A(new_n6962_), .B(\asqrt[54] ), .Y(new_n7009_));
  AOI21X1  g06817(.A0(new_n7009_), .A1(new_n7008_), .B0(new_n6976_), .Y(new_n7010_));
  OAI21X1  g06818(.A0(new_n7010_), .A1(new_n7007_), .B0(\asqrt[55] ), .Y(new_n7011_));
  INVX1    g06819(.A(new_n6985_), .Y(new_n7012_));
  OAI21X1  g06820(.A0(new_n6969_), .A1(new_n902_), .B0(new_n697_), .Y(new_n7013_));
  OAI21X1  g06821(.A0(new_n7013_), .A1(new_n7010_), .B0(new_n7012_), .Y(new_n7014_));
  NAND3X1  g06822(.A(new_n7014_), .B(new_n7011_), .C(new_n582_), .Y(new_n7015_));
  NAND2X1  g06823(.A(new_n7015_), .B(new_n7002_), .Y(new_n7016_));
  AND2X1   g06824(.A(new_n6603_), .B(new_n6597_), .Y(new_n7017_));
  NOR4X1   g06825(.A(new_n6699_), .B(new_n7017_), .C(new_n6634_), .D(new_n6586_), .Y(new_n7018_));
  AOI22X1  g06826(.A0(new_n6603_), .A1(new_n6597_), .B0(new_n6585_), .B1(\asqrt[56] ), .Y(new_n7019_));
  AOI21X1  g06827(.A0(new_n7019_), .A1(\asqrt[32] ), .B0(new_n6602_), .Y(new_n7020_));
  NOR2X1   g06828(.A(new_n7020_), .B(new_n7018_), .Y(new_n7021_));
  AND2X1   g06829(.A(new_n6999_), .B(new_n481_), .Y(new_n7022_));
  AOI21X1  g06830(.A0(new_n7022_), .A1(new_n7016_), .B0(new_n7021_), .Y(new_n7023_));
  OAI21X1  g06831(.A0(new_n7023_), .A1(new_n7006_), .B0(\asqrt[58] ), .Y(new_n7024_));
  AND2X1   g06832(.A(new_n6638_), .B(new_n6636_), .Y(new_n7025_));
  OR4X1    g06833(.A(new_n6699_), .B(new_n7025_), .C(new_n6610_), .D(new_n6637_), .Y(new_n7026_));
  OR2X1    g06834(.A(new_n7025_), .B(new_n6637_), .Y(new_n7027_));
  OAI21X1  g06835(.A0(new_n7027_), .A1(new_n6699_), .B0(new_n6610_), .Y(new_n7028_));
  AND2X1   g06836(.A(new_n7028_), .B(new_n7026_), .Y(new_n7029_));
  INVX1    g06837(.A(new_n7029_), .Y(new_n7030_));
  AOI21X1  g06838(.A0(new_n7014_), .A1(new_n7011_), .B0(new_n582_), .Y(new_n7031_));
  AOI21X1  g06839(.A0(new_n7015_), .A1(new_n7002_), .B0(new_n7031_), .Y(new_n7032_));
  OAI21X1  g06840(.A0(new_n7032_), .A1(new_n481_), .B0(new_n399_), .Y(new_n7033_));
  OAI21X1  g06841(.A0(new_n7033_), .A1(new_n7023_), .B0(new_n7030_), .Y(new_n7034_));
  AOI21X1  g06842(.A0(new_n7034_), .A1(new_n7024_), .B0(new_n328_), .Y(new_n7035_));
  OR4X1    g06843(.A(new_n6699_), .B(new_n6648_), .C(new_n6621_), .D(new_n6615_), .Y(new_n7036_));
  NAND2X1  g06844(.A(new_n6622_), .B(new_n6640_), .Y(new_n7037_));
  OAI21X1  g06845(.A0(new_n7037_), .A1(new_n6699_), .B0(new_n6621_), .Y(new_n7038_));
  AND2X1   g06846(.A(new_n7038_), .B(new_n7036_), .Y(new_n7039_));
  INVX1    g06847(.A(new_n7039_), .Y(new_n7040_));
  NAND3X1  g06848(.A(new_n7034_), .B(new_n7024_), .C(new_n328_), .Y(new_n7041_));
  AOI21X1  g06849(.A0(new_n7041_), .A1(new_n7040_), .B0(new_n7035_), .Y(new_n7042_));
  OR2X1    g06850(.A(new_n7042_), .B(new_n292_), .Y(new_n7043_));
  OR2X1    g06851(.A(new_n7032_), .B(new_n481_), .Y(new_n7044_));
  AND2X1   g06852(.A(new_n7015_), .B(new_n7002_), .Y(new_n7045_));
  INVX1    g06853(.A(new_n7021_), .Y(new_n7046_));
  NAND2X1  g06854(.A(new_n6999_), .B(new_n481_), .Y(new_n7047_));
  OAI21X1  g06855(.A0(new_n7047_), .A1(new_n7045_), .B0(new_n7046_), .Y(new_n7048_));
  AOI21X1  g06856(.A0(new_n7048_), .A1(new_n7044_), .B0(new_n399_), .Y(new_n7049_));
  AOI21X1  g06857(.A0(new_n7005_), .A1(\asqrt[57] ), .B0(\asqrt[58] ), .Y(new_n7050_));
  AOI21X1  g06858(.A0(new_n7050_), .A1(new_n7048_), .B0(new_n7029_), .Y(new_n7051_));
  NOR3X1   g06859(.A(new_n7051_), .B(new_n7049_), .C(\asqrt[59] ), .Y(new_n7052_));
  NOR2X1   g06860(.A(new_n7052_), .B(new_n7039_), .Y(new_n7053_));
  OAI21X1  g06861(.A0(new_n6641_), .A1(new_n6625_), .B0(new_n6630_), .Y(new_n7054_));
  NOR3X1   g06862(.A(new_n7054_), .B(new_n6699_), .C(new_n6662_), .Y(new_n7055_));
  AOI22X1  g06863(.A0(new_n6664_), .A1(new_n6663_), .B0(new_n6649_), .B1(\asqrt[59] ), .Y(new_n7056_));
  AOI21X1  g06864(.A0(new_n7056_), .A1(\asqrt[32] ), .B0(new_n6630_), .Y(new_n7057_));
  NOR2X1   g06865(.A(new_n7057_), .B(new_n7055_), .Y(new_n7058_));
  INVX1    g06866(.A(new_n7058_), .Y(new_n7059_));
  OAI21X1  g06867(.A0(new_n7051_), .A1(new_n7049_), .B0(\asqrt[59] ), .Y(new_n7060_));
  NAND2X1  g06868(.A(new_n7060_), .B(new_n292_), .Y(new_n7061_));
  OAI21X1  g06869(.A0(new_n7061_), .A1(new_n7053_), .B0(new_n7059_), .Y(new_n7062_));
  AOI21X1  g06870(.A0(new_n7062_), .A1(new_n7043_), .B0(new_n217_), .Y(new_n7063_));
  AND2X1   g06871(.A(new_n6650_), .B(new_n6642_), .Y(new_n7064_));
  OR4X1    g06872(.A(new_n6699_), .B(new_n7064_), .C(new_n6667_), .D(new_n6643_), .Y(new_n7065_));
  OR2X1    g06873(.A(new_n7064_), .B(new_n6643_), .Y(new_n7066_));
  OAI21X1  g06874(.A0(new_n7066_), .A1(new_n6699_), .B0(new_n6667_), .Y(new_n7067_));
  AND2X1   g06875(.A(new_n7067_), .B(new_n7065_), .Y(new_n7068_));
  OAI21X1  g06876(.A0(new_n7052_), .A1(new_n7039_), .B0(new_n7060_), .Y(new_n7069_));
  AOI21X1  g06877(.A0(new_n7069_), .A1(\asqrt[60] ), .B0(\asqrt[61] ), .Y(new_n7070_));
  AOI21X1  g06878(.A0(new_n7070_), .A1(new_n7062_), .B0(new_n7068_), .Y(new_n7071_));
  OAI21X1  g06879(.A0(new_n7071_), .A1(new_n7063_), .B0(\asqrt[62] ), .Y(new_n7072_));
  OR4X1    g06880(.A(new_n6699_), .B(new_n6658_), .C(new_n6661_), .D(new_n6677_), .Y(new_n7073_));
  NAND2X1  g06881(.A(new_n6670_), .B(new_n6652_), .Y(new_n7074_));
  OAI21X1  g06882(.A0(new_n7074_), .A1(new_n6699_), .B0(new_n6661_), .Y(new_n7075_));
  AND2X1   g06883(.A(new_n7075_), .B(new_n7073_), .Y(new_n7076_));
  NOR3X1   g06884(.A(new_n7071_), .B(new_n7063_), .C(\asqrt[62] ), .Y(new_n7077_));
  OAI21X1  g06885(.A0(new_n7077_), .A1(new_n7076_), .B0(new_n7072_), .Y(new_n7078_));
  AND2X1   g06886(.A(new_n6678_), .B(new_n6671_), .Y(new_n7079_));
  NOR4X1   g06887(.A(new_n6699_), .B(new_n7079_), .C(new_n6702_), .D(new_n6660_), .Y(new_n7080_));
  AOI22X1  g06888(.A0(new_n6678_), .A1(new_n6671_), .B0(new_n6659_), .B1(\asqrt[62] ), .Y(new_n7081_));
  AOI21X1  g06889(.A0(new_n7081_), .A1(\asqrt[32] ), .B0(new_n6676_), .Y(new_n7082_));
  NOR2X1   g06890(.A(new_n7082_), .B(new_n7080_), .Y(new_n7083_));
  INVX1    g06891(.A(new_n7083_), .Y(new_n7084_));
  AND2X1   g06892(.A(new_n6707_), .B(new_n6704_), .Y(new_n7085_));
  AOI21X1  g06893(.A0(new_n6704_), .A1(new_n6700_), .B0(new_n6682_), .Y(new_n7086_));
  AOI21X1  g06894(.A0(new_n7086_), .A1(\asqrt[32] ), .B0(new_n7085_), .Y(new_n7087_));
  AND2X1   g06895(.A(new_n7087_), .B(new_n7084_), .Y(new_n7088_));
  AOI21X1  g06896(.A0(new_n7088_), .A1(new_n7078_), .B0(\asqrt[63] ), .Y(new_n7089_));
  NOR2X1   g06897(.A(new_n7077_), .B(new_n7076_), .Y(new_n7090_));
  NAND2X1  g06898(.A(new_n7083_), .B(new_n7072_), .Y(new_n7091_));
  AND2X1   g06899(.A(new_n6704_), .B(new_n6700_), .Y(new_n7092_));
  OAI21X1  g06900(.A0(new_n6699_), .A1(new_n6682_), .B0(new_n7092_), .Y(new_n7093_));
  NOR2X1   g06901(.A(new_n7086_), .B(new_n193_), .Y(new_n7094_));
  AND2X1   g06902(.A(new_n6687_), .B(new_n193_), .Y(new_n7095_));
  INVX1    g06903(.A(new_n6696_), .Y(new_n7096_));
  OR2X1    g06904(.A(new_n7096_), .B(new_n6680_), .Y(new_n7097_));
  AOI21X1  g06905(.A0(new_n6681_), .A1(new_n6305_), .B0(new_n7097_), .Y(new_n7098_));
  NAND2X1  g06906(.A(new_n7098_), .B(new_n6692_), .Y(new_n7099_));
  NOR3X1   g06907(.A(new_n7099_), .B(new_n7085_), .C(new_n7095_), .Y(new_n7100_));
  AOI21X1  g06908(.A0(new_n7094_), .A1(new_n7093_), .B0(new_n7100_), .Y(new_n7101_));
  OAI21X1  g06909(.A0(new_n7091_), .A1(new_n7090_), .B0(new_n7101_), .Y(new_n7102_));
  NOR2X1   g06910(.A(new_n7102_), .B(new_n7089_), .Y(new_n7103_));
  INVX1    g06911(.A(new_n7103_), .Y(\asqrt[31] ));
  OAI21X1  g06912(.A0(new_n7102_), .A1(new_n7089_), .B0(\a[62] ), .Y(new_n7105_));
  INVX1    g06913(.A(\a[62] ), .Y(new_n7106_));
  NOR2X1   g06914(.A(\a[61] ), .B(\a[60] ), .Y(new_n7107_));
  NAND2X1  g06915(.A(new_n7107_), .B(new_n7106_), .Y(new_n7108_));
  AND2X1   g06916(.A(new_n7108_), .B(new_n7105_), .Y(new_n7109_));
  AND2X1   g06917(.A(new_n7069_), .B(\asqrt[60] ), .Y(new_n7110_));
  OR2X1    g06918(.A(new_n7052_), .B(new_n7039_), .Y(new_n7111_));
  AND2X1   g06919(.A(new_n7060_), .B(new_n292_), .Y(new_n7112_));
  AOI21X1  g06920(.A0(new_n7112_), .A1(new_n7111_), .B0(new_n7058_), .Y(new_n7113_));
  OAI21X1  g06921(.A0(new_n7113_), .A1(new_n7110_), .B0(\asqrt[61] ), .Y(new_n7114_));
  INVX1    g06922(.A(new_n7068_), .Y(new_n7115_));
  OAI21X1  g06923(.A0(new_n7042_), .A1(new_n292_), .B0(new_n217_), .Y(new_n7116_));
  OAI21X1  g06924(.A0(new_n7116_), .A1(new_n7113_), .B0(new_n7115_), .Y(new_n7117_));
  AOI21X1  g06925(.A0(new_n7117_), .A1(new_n7114_), .B0(new_n199_), .Y(new_n7118_));
  INVX1    g06926(.A(new_n7076_), .Y(new_n7119_));
  NAND3X1  g06927(.A(new_n7117_), .B(new_n7114_), .C(new_n199_), .Y(new_n7120_));
  AOI21X1  g06928(.A0(new_n7120_), .A1(new_n7119_), .B0(new_n7118_), .Y(new_n7121_));
  INVX1    g06929(.A(new_n7088_), .Y(new_n7122_));
  OAI21X1  g06930(.A0(new_n7122_), .A1(new_n7121_), .B0(new_n193_), .Y(new_n7123_));
  OR2X1    g06931(.A(new_n7077_), .B(new_n7076_), .Y(new_n7124_));
  AND2X1   g06932(.A(new_n7083_), .B(new_n7072_), .Y(new_n7125_));
  INVX1    g06933(.A(new_n7101_), .Y(new_n7126_));
  AOI21X1  g06934(.A0(new_n7125_), .A1(new_n7124_), .B0(new_n7126_), .Y(new_n7127_));
  AOI21X1  g06935(.A0(new_n7127_), .A1(new_n7123_), .B0(new_n7106_), .Y(new_n7128_));
  NAND3X1  g06936(.A(new_n7108_), .B(new_n6696_), .C(new_n6692_), .Y(new_n7129_));
  NOR4X1   g06937(.A(new_n7129_), .B(new_n7128_), .C(new_n7085_), .D(new_n7095_), .Y(new_n7130_));
  INVX1    g06938(.A(\a[63] ), .Y(new_n7131_));
  AOI21X1  g06939(.A0(new_n7127_), .A1(new_n7123_), .B0(\a[62] ), .Y(new_n7132_));
  OAI21X1  g06940(.A0(new_n7102_), .A1(new_n7089_), .B0(new_n6711_), .Y(new_n7133_));
  OAI21X1  g06941(.A0(new_n7132_), .A1(new_n7131_), .B0(new_n7133_), .Y(new_n7134_));
  OAI22X1  g06942(.A0(new_n7134_), .A1(new_n7130_), .B0(new_n7109_), .B1(new_n6699_), .Y(new_n7135_));
  AND2X1   g06943(.A(new_n7135_), .B(\asqrt[33] ), .Y(new_n7136_));
  OR4X1    g06944(.A(new_n7129_), .B(new_n7128_), .C(new_n7085_), .D(new_n7095_), .Y(new_n7137_));
  OAI21X1  g06945(.A0(new_n7102_), .A1(new_n7089_), .B0(new_n7106_), .Y(new_n7138_));
  AOI21X1  g06946(.A0(new_n7127_), .A1(new_n7123_), .B0(new_n6725_), .Y(new_n7139_));
  AOI21X1  g06947(.A0(new_n7138_), .A1(\a[63] ), .B0(new_n7139_), .Y(new_n7140_));
  NAND2X1  g06948(.A(new_n7140_), .B(new_n7137_), .Y(new_n7141_));
  AOI21X1  g06949(.A0(new_n7108_), .A1(new_n7105_), .B0(new_n6699_), .Y(new_n7142_));
  NOR2X1   g06950(.A(new_n7142_), .B(\asqrt[33] ), .Y(new_n7143_));
  AND2X1   g06951(.A(new_n7125_), .B(new_n7124_), .Y(new_n7144_));
  AND2X1   g06952(.A(new_n7094_), .B(new_n7093_), .Y(new_n7145_));
  OR2X1    g06953(.A(new_n7100_), .B(new_n6699_), .Y(new_n7146_));
  OR4X1    g06954(.A(new_n7146_), .B(new_n7145_), .C(new_n7144_), .D(new_n7089_), .Y(new_n7147_));
  AOI21X1  g06955(.A0(new_n7147_), .A1(new_n7133_), .B0(new_n6714_), .Y(new_n7148_));
  NOR4X1   g06956(.A(new_n7146_), .B(new_n7145_), .C(new_n7144_), .D(new_n7089_), .Y(new_n7149_));
  NOR3X1   g06957(.A(new_n7149_), .B(new_n7139_), .C(\a[64] ), .Y(new_n7150_));
  NOR2X1   g06958(.A(new_n7150_), .B(new_n7148_), .Y(new_n7151_));
  AOI21X1  g06959(.A0(new_n7143_), .A1(new_n7141_), .B0(new_n7151_), .Y(new_n7152_));
  OAI21X1  g06960(.A0(new_n7152_), .A1(new_n7136_), .B0(\asqrt[34] ), .Y(new_n7153_));
  AOI21X1  g06961(.A0(new_n7140_), .A1(new_n7137_), .B0(new_n7142_), .Y(new_n7154_));
  OAI21X1  g06962(.A0(new_n7154_), .A1(new_n6294_), .B0(new_n5941_), .Y(new_n7155_));
  AND2X1   g06963(.A(new_n6764_), .B(new_n6762_), .Y(new_n7156_));
  NOR3X1   g06964(.A(new_n6722_), .B(new_n7156_), .C(new_n6713_), .Y(new_n7157_));
  OAI21X1  g06965(.A0(new_n7102_), .A1(new_n7089_), .B0(new_n7157_), .Y(new_n7158_));
  AOI21X1  g06966(.A0(new_n6712_), .A1(\asqrt[33] ), .B0(new_n6722_), .Y(new_n7159_));
  OAI21X1  g06967(.A0(new_n7102_), .A1(new_n7089_), .B0(new_n7159_), .Y(new_n7160_));
  NAND2X1  g06968(.A(new_n7160_), .B(new_n7156_), .Y(new_n7161_));
  NAND2X1  g06969(.A(new_n7161_), .B(new_n7158_), .Y(new_n7162_));
  OAI21X1  g06970(.A0(new_n7155_), .A1(new_n7152_), .B0(new_n7162_), .Y(new_n7163_));
  AOI21X1  g06971(.A0(new_n7163_), .A1(new_n7153_), .B0(new_n5541_), .Y(new_n7164_));
  AND2X1   g06972(.A(new_n6769_), .B(new_n6767_), .Y(new_n7165_));
  NOR3X1   g06973(.A(new_n6734_), .B(new_n7165_), .C(new_n6768_), .Y(new_n7166_));
  OAI21X1  g06974(.A0(new_n7102_), .A1(new_n7089_), .B0(new_n7166_), .Y(new_n7167_));
  NOR2X1   g06975(.A(new_n7165_), .B(new_n6768_), .Y(new_n7168_));
  OAI21X1  g06976(.A0(new_n7102_), .A1(new_n7089_), .B0(new_n7168_), .Y(new_n7169_));
  NAND2X1  g06977(.A(new_n7169_), .B(new_n6734_), .Y(new_n7170_));
  AND2X1   g06978(.A(new_n7170_), .B(new_n7167_), .Y(new_n7171_));
  INVX1    g06979(.A(new_n7171_), .Y(new_n7172_));
  NAND3X1  g06980(.A(new_n7163_), .B(new_n7153_), .C(new_n5541_), .Y(new_n7173_));
  AOI21X1  g06981(.A0(new_n7173_), .A1(new_n7172_), .B0(new_n7164_), .Y(new_n7174_));
  OR2X1    g06982(.A(new_n7174_), .B(new_n5176_), .Y(new_n7175_));
  OR2X1    g06983(.A(new_n7154_), .B(new_n6294_), .Y(new_n7176_));
  AND2X1   g06984(.A(new_n7140_), .B(new_n7137_), .Y(new_n7177_));
  OR2X1    g06985(.A(new_n7142_), .B(\asqrt[33] ), .Y(new_n7178_));
  OR2X1    g06986(.A(new_n7150_), .B(new_n7148_), .Y(new_n7179_));
  OAI21X1  g06987(.A0(new_n7178_), .A1(new_n7177_), .B0(new_n7179_), .Y(new_n7180_));
  AOI21X1  g06988(.A0(new_n7180_), .A1(new_n7176_), .B0(new_n5941_), .Y(new_n7181_));
  AOI21X1  g06989(.A0(new_n7135_), .A1(\asqrt[33] ), .B0(\asqrt[34] ), .Y(new_n7182_));
  AOI22X1  g06990(.A0(new_n7161_), .A1(new_n7158_), .B0(new_n7182_), .B1(new_n7180_), .Y(new_n7183_));
  NOR3X1   g06991(.A(new_n7183_), .B(new_n7181_), .C(\asqrt[35] ), .Y(new_n7184_));
  NOR2X1   g06992(.A(new_n7184_), .B(new_n7171_), .Y(new_n7185_));
  NOR3X1   g06993(.A(new_n6774_), .B(new_n6742_), .C(new_n6736_), .Y(new_n7186_));
  OAI21X1  g06994(.A0(new_n7102_), .A1(new_n7089_), .B0(new_n7186_), .Y(new_n7187_));
  NOR3X1   g06995(.A(new_n7103_), .B(new_n6774_), .C(new_n6736_), .Y(new_n7188_));
  OR2X1    g06996(.A(new_n7188_), .B(new_n6741_), .Y(new_n7189_));
  AND2X1   g06997(.A(new_n7189_), .B(new_n7187_), .Y(new_n7190_));
  INVX1    g06998(.A(new_n7190_), .Y(new_n7191_));
  OR2X1    g06999(.A(new_n7164_), .B(\asqrt[36] ), .Y(new_n7192_));
  OAI21X1  g07000(.A0(new_n7192_), .A1(new_n7185_), .B0(new_n7191_), .Y(new_n7193_));
  AOI21X1  g07001(.A0(new_n7193_), .A1(new_n7175_), .B0(new_n4826_), .Y(new_n7194_));
  AOI21X1  g07002(.A0(new_n6788_), .A1(new_n6787_), .B0(new_n6752_), .Y(new_n7195_));
  AND2X1   g07003(.A(new_n7195_), .B(new_n6745_), .Y(new_n7196_));
  AOI22X1  g07004(.A0(new_n6788_), .A1(new_n6787_), .B0(new_n6775_), .B1(\asqrt[36] ), .Y(new_n7197_));
  AOI21X1  g07005(.A0(new_n7197_), .A1(\asqrt[31] ), .B0(new_n6751_), .Y(new_n7198_));
  AOI21X1  g07006(.A0(new_n7196_), .A1(\asqrt[31] ), .B0(new_n7198_), .Y(new_n7199_));
  OAI21X1  g07007(.A0(new_n7183_), .A1(new_n7181_), .B0(\asqrt[35] ), .Y(new_n7200_));
  OAI21X1  g07008(.A0(new_n7184_), .A1(new_n7171_), .B0(new_n7200_), .Y(new_n7201_));
  AOI21X1  g07009(.A0(new_n7201_), .A1(\asqrt[36] ), .B0(\asqrt[37] ), .Y(new_n7202_));
  AOI21X1  g07010(.A0(new_n7202_), .A1(new_n7193_), .B0(new_n7199_), .Y(new_n7203_));
  OAI21X1  g07011(.A0(new_n7203_), .A1(new_n7194_), .B0(\asqrt[38] ), .Y(new_n7204_));
  AND2X1   g07012(.A(new_n6776_), .B(new_n6754_), .Y(new_n7205_));
  NOR3X1   g07013(.A(new_n7205_), .B(new_n6791_), .C(new_n6755_), .Y(new_n7206_));
  NOR3X1   g07014(.A(new_n7103_), .B(new_n7205_), .C(new_n6755_), .Y(new_n7207_));
  NOR2X1   g07015(.A(new_n7207_), .B(new_n6760_), .Y(new_n7208_));
  AOI21X1  g07016(.A0(new_n7206_), .A1(\asqrt[31] ), .B0(new_n7208_), .Y(new_n7209_));
  NOR3X1   g07017(.A(new_n7203_), .B(new_n7194_), .C(\asqrt[38] ), .Y(new_n7210_));
  OAI21X1  g07018(.A0(new_n7210_), .A1(new_n7209_), .B0(new_n7204_), .Y(new_n7211_));
  AND2X1   g07019(.A(new_n7211_), .B(\asqrt[39] ), .Y(new_n7212_));
  OR2X1    g07020(.A(new_n7210_), .B(new_n7209_), .Y(new_n7213_));
  OR4X1    g07021(.A(new_n7103_), .B(new_n6783_), .C(new_n6781_), .D(new_n6801_), .Y(new_n7214_));
  NAND2X1  g07022(.A(new_n6794_), .B(new_n6778_), .Y(new_n7215_));
  OAI21X1  g07023(.A0(new_n7215_), .A1(new_n7103_), .B0(new_n6781_), .Y(new_n7216_));
  AND2X1   g07024(.A(new_n7216_), .B(new_n7214_), .Y(new_n7217_));
  AND2X1   g07025(.A(new_n7204_), .B(new_n4165_), .Y(new_n7218_));
  AOI21X1  g07026(.A0(new_n7218_), .A1(new_n7213_), .B0(new_n7217_), .Y(new_n7219_));
  OAI21X1  g07027(.A0(new_n7219_), .A1(new_n7212_), .B0(\asqrt[40] ), .Y(new_n7220_));
  AND2X1   g07028(.A(new_n6802_), .B(new_n6795_), .Y(new_n7221_));
  NOR3X1   g07029(.A(new_n7221_), .B(new_n6840_), .C(new_n6785_), .Y(new_n7222_));
  NOR3X1   g07030(.A(new_n7103_), .B(new_n7221_), .C(new_n6785_), .Y(new_n7223_));
  NOR2X1   g07031(.A(new_n7223_), .B(new_n6800_), .Y(new_n7224_));
  AOI21X1  g07032(.A0(new_n7222_), .A1(\asqrt[31] ), .B0(new_n7224_), .Y(new_n7225_));
  INVX1    g07033(.A(new_n7225_), .Y(new_n7226_));
  AND2X1   g07034(.A(new_n7201_), .B(\asqrt[36] ), .Y(new_n7227_));
  OR2X1    g07035(.A(new_n7184_), .B(new_n7171_), .Y(new_n7228_));
  NOR2X1   g07036(.A(new_n7164_), .B(\asqrt[36] ), .Y(new_n7229_));
  AOI21X1  g07037(.A0(new_n7229_), .A1(new_n7228_), .B0(new_n7190_), .Y(new_n7230_));
  OAI21X1  g07038(.A0(new_n7230_), .A1(new_n7227_), .B0(\asqrt[37] ), .Y(new_n7231_));
  INVX1    g07039(.A(new_n7199_), .Y(new_n7232_));
  OAI21X1  g07040(.A0(new_n7174_), .A1(new_n5176_), .B0(new_n4826_), .Y(new_n7233_));
  OAI21X1  g07041(.A0(new_n7233_), .A1(new_n7230_), .B0(new_n7232_), .Y(new_n7234_));
  AOI21X1  g07042(.A0(new_n7234_), .A1(new_n7231_), .B0(new_n4493_), .Y(new_n7235_));
  INVX1    g07043(.A(new_n7209_), .Y(new_n7236_));
  NAND3X1  g07044(.A(new_n7234_), .B(new_n7231_), .C(new_n4493_), .Y(new_n7237_));
  AOI21X1  g07045(.A0(new_n7237_), .A1(new_n7236_), .B0(new_n7235_), .Y(new_n7238_));
  OAI21X1  g07046(.A0(new_n7238_), .A1(new_n4165_), .B0(new_n3863_), .Y(new_n7239_));
  OAI21X1  g07047(.A0(new_n7239_), .A1(new_n7219_), .B0(new_n7226_), .Y(new_n7240_));
  AOI21X1  g07048(.A0(new_n7240_), .A1(new_n7220_), .B0(new_n3564_), .Y(new_n7241_));
  AND2X1   g07049(.A(new_n6844_), .B(new_n6842_), .Y(new_n7242_));
  NOR3X1   g07050(.A(new_n7242_), .B(new_n6810_), .C(new_n6843_), .Y(new_n7243_));
  NOR3X1   g07051(.A(new_n7103_), .B(new_n7242_), .C(new_n6843_), .Y(new_n7244_));
  NOR2X1   g07052(.A(new_n7244_), .B(new_n6809_), .Y(new_n7245_));
  AOI21X1  g07053(.A0(new_n7243_), .A1(\asqrt[31] ), .B0(new_n7245_), .Y(new_n7246_));
  INVX1    g07054(.A(new_n7246_), .Y(new_n7247_));
  NAND3X1  g07055(.A(new_n7240_), .B(new_n7220_), .C(new_n3564_), .Y(new_n7248_));
  AOI21X1  g07056(.A0(new_n7248_), .A1(new_n7247_), .B0(new_n7241_), .Y(new_n7249_));
  OR2X1    g07057(.A(new_n7249_), .B(new_n3276_), .Y(new_n7250_));
  AND2X1   g07058(.A(new_n7248_), .B(new_n7247_), .Y(new_n7251_));
  NAND4X1  g07059(.A(\asqrt[31] ), .B(new_n6820_), .C(new_n6818_), .D(new_n6846_), .Y(new_n7252_));
  NAND2X1  g07060(.A(new_n6820_), .B(new_n6846_), .Y(new_n7253_));
  OAI21X1  g07061(.A0(new_n7253_), .A1(new_n7103_), .B0(new_n6819_), .Y(new_n7254_));
  AND2X1   g07062(.A(new_n7254_), .B(new_n7252_), .Y(new_n7255_));
  INVX1    g07063(.A(new_n7255_), .Y(new_n7256_));
  OR2X1    g07064(.A(new_n7241_), .B(\asqrt[42] ), .Y(new_n7257_));
  OAI21X1  g07065(.A0(new_n7257_), .A1(new_n7251_), .B0(new_n7256_), .Y(new_n7258_));
  AOI21X1  g07066(.A0(new_n7258_), .A1(new_n7250_), .B0(new_n3008_), .Y(new_n7259_));
  AOI21X1  g07067(.A0(new_n6862_), .A1(new_n6861_), .B0(new_n6829_), .Y(new_n7260_));
  AND2X1   g07068(.A(new_n7260_), .B(new_n6822_), .Y(new_n7261_));
  AOI22X1  g07069(.A0(new_n6862_), .A1(new_n6861_), .B0(new_n6848_), .B1(\asqrt[42] ), .Y(new_n7262_));
  AOI21X1  g07070(.A0(new_n7262_), .A1(\asqrt[31] ), .B0(new_n6828_), .Y(new_n7263_));
  AOI21X1  g07071(.A0(new_n7261_), .A1(\asqrt[31] ), .B0(new_n7263_), .Y(new_n7264_));
  OR2X1    g07072(.A(new_n7238_), .B(new_n4165_), .Y(new_n7265_));
  NOR2X1   g07073(.A(new_n7210_), .B(new_n7209_), .Y(new_n7266_));
  INVX1    g07074(.A(new_n7217_), .Y(new_n7267_));
  NAND2X1  g07075(.A(new_n7204_), .B(new_n4165_), .Y(new_n7268_));
  OAI21X1  g07076(.A0(new_n7268_), .A1(new_n7266_), .B0(new_n7267_), .Y(new_n7269_));
  AOI21X1  g07077(.A0(new_n7269_), .A1(new_n7265_), .B0(new_n3863_), .Y(new_n7270_));
  AOI21X1  g07078(.A0(new_n7211_), .A1(\asqrt[39] ), .B0(\asqrt[40] ), .Y(new_n7271_));
  AOI21X1  g07079(.A0(new_n7271_), .A1(new_n7269_), .B0(new_n7225_), .Y(new_n7272_));
  OAI21X1  g07080(.A0(new_n7272_), .A1(new_n7270_), .B0(\asqrt[41] ), .Y(new_n7273_));
  NOR3X1   g07081(.A(new_n7272_), .B(new_n7270_), .C(\asqrt[41] ), .Y(new_n7274_));
  OAI21X1  g07082(.A0(new_n7274_), .A1(new_n7246_), .B0(new_n7273_), .Y(new_n7275_));
  AOI21X1  g07083(.A0(new_n7275_), .A1(\asqrt[42] ), .B0(\asqrt[43] ), .Y(new_n7276_));
  AOI21X1  g07084(.A0(new_n7276_), .A1(new_n7258_), .B0(new_n7264_), .Y(new_n7277_));
  OAI21X1  g07085(.A0(new_n7277_), .A1(new_n7259_), .B0(\asqrt[44] ), .Y(new_n7278_));
  AND2X1   g07086(.A(new_n6849_), .B(new_n6831_), .Y(new_n7279_));
  NOR3X1   g07087(.A(new_n7279_), .B(new_n6865_), .C(new_n6832_), .Y(new_n7280_));
  NOR3X1   g07088(.A(new_n7103_), .B(new_n7279_), .C(new_n6832_), .Y(new_n7281_));
  NOR2X1   g07089(.A(new_n7281_), .B(new_n6837_), .Y(new_n7282_));
  AOI21X1  g07090(.A0(new_n7280_), .A1(\asqrt[31] ), .B0(new_n7282_), .Y(new_n7283_));
  NOR3X1   g07091(.A(new_n7277_), .B(new_n7259_), .C(\asqrt[44] ), .Y(new_n7284_));
  OAI21X1  g07092(.A0(new_n7284_), .A1(new_n7283_), .B0(new_n7278_), .Y(new_n7285_));
  AND2X1   g07093(.A(new_n7285_), .B(\asqrt[45] ), .Y(new_n7286_));
  INVX1    g07094(.A(new_n7283_), .Y(new_n7287_));
  AND2X1   g07095(.A(new_n7275_), .B(\asqrt[42] ), .Y(new_n7288_));
  NAND2X1  g07096(.A(new_n7248_), .B(new_n7247_), .Y(new_n7289_));
  NOR2X1   g07097(.A(new_n7241_), .B(\asqrt[42] ), .Y(new_n7290_));
  AOI21X1  g07098(.A0(new_n7290_), .A1(new_n7289_), .B0(new_n7255_), .Y(new_n7291_));
  OAI21X1  g07099(.A0(new_n7291_), .A1(new_n7288_), .B0(\asqrt[43] ), .Y(new_n7292_));
  INVX1    g07100(.A(new_n7264_), .Y(new_n7293_));
  OAI21X1  g07101(.A0(new_n7249_), .A1(new_n3276_), .B0(new_n3008_), .Y(new_n7294_));
  OAI21X1  g07102(.A0(new_n7294_), .A1(new_n7291_), .B0(new_n7293_), .Y(new_n7295_));
  NAND3X1  g07103(.A(new_n7295_), .B(new_n7292_), .C(new_n2769_), .Y(new_n7296_));
  NAND2X1  g07104(.A(new_n7296_), .B(new_n7287_), .Y(new_n7297_));
  NAND4X1  g07105(.A(\asqrt[31] ), .B(new_n6868_), .C(new_n6855_), .D(new_n6851_), .Y(new_n7298_));
  NAND2X1  g07106(.A(new_n6868_), .B(new_n6851_), .Y(new_n7299_));
  OAI21X1  g07107(.A0(new_n7299_), .A1(new_n7103_), .B0(new_n6859_), .Y(new_n7300_));
  AND2X1   g07108(.A(new_n7300_), .B(new_n7298_), .Y(new_n7301_));
  AOI21X1  g07109(.A0(new_n7295_), .A1(new_n7292_), .B0(new_n2769_), .Y(new_n7302_));
  NOR2X1   g07110(.A(new_n7302_), .B(\asqrt[45] ), .Y(new_n7303_));
  AOI21X1  g07111(.A0(new_n7303_), .A1(new_n7297_), .B0(new_n7301_), .Y(new_n7304_));
  OAI21X1  g07112(.A0(new_n7304_), .A1(new_n7286_), .B0(\asqrt[46] ), .Y(new_n7305_));
  AND2X1   g07113(.A(new_n6876_), .B(new_n6869_), .Y(new_n7306_));
  NOR3X1   g07114(.A(new_n7306_), .B(new_n6914_), .C(new_n6858_), .Y(new_n7307_));
  NOR3X1   g07115(.A(new_n7103_), .B(new_n7306_), .C(new_n6858_), .Y(new_n7308_));
  NOR2X1   g07116(.A(new_n7308_), .B(new_n6874_), .Y(new_n7309_));
  AOI21X1  g07117(.A0(new_n7307_), .A1(\asqrt[31] ), .B0(new_n7309_), .Y(new_n7310_));
  INVX1    g07118(.A(new_n7310_), .Y(new_n7311_));
  AOI21X1  g07119(.A0(new_n7296_), .A1(new_n7287_), .B0(new_n7302_), .Y(new_n7312_));
  OAI21X1  g07120(.A0(new_n7312_), .A1(new_n2570_), .B0(new_n2263_), .Y(new_n7313_));
  OAI21X1  g07121(.A0(new_n7313_), .A1(new_n7304_), .B0(new_n7311_), .Y(new_n7314_));
  AOI21X1  g07122(.A0(new_n7314_), .A1(new_n7305_), .B0(new_n2040_), .Y(new_n7315_));
  AND2X1   g07123(.A(new_n6918_), .B(new_n6916_), .Y(new_n7316_));
  NOR3X1   g07124(.A(new_n7316_), .B(new_n6884_), .C(new_n6917_), .Y(new_n7317_));
  NOR3X1   g07125(.A(new_n7103_), .B(new_n7316_), .C(new_n6917_), .Y(new_n7318_));
  NOR2X1   g07126(.A(new_n7318_), .B(new_n6883_), .Y(new_n7319_));
  AOI21X1  g07127(.A0(new_n7317_), .A1(\asqrt[31] ), .B0(new_n7319_), .Y(new_n7320_));
  INVX1    g07128(.A(new_n7320_), .Y(new_n7321_));
  NAND3X1  g07129(.A(new_n7314_), .B(new_n7305_), .C(new_n2040_), .Y(new_n7322_));
  AOI21X1  g07130(.A0(new_n7322_), .A1(new_n7321_), .B0(new_n7315_), .Y(new_n7323_));
  OR2X1    g07131(.A(new_n7323_), .B(new_n1834_), .Y(new_n7324_));
  AND2X1   g07132(.A(new_n7322_), .B(new_n7321_), .Y(new_n7325_));
  NAND4X1  g07133(.A(\asqrt[31] ), .B(new_n6894_), .C(new_n6892_), .D(new_n6920_), .Y(new_n7326_));
  NAND2X1  g07134(.A(new_n6894_), .B(new_n6920_), .Y(new_n7327_));
  OAI21X1  g07135(.A0(new_n7327_), .A1(new_n7103_), .B0(new_n6893_), .Y(new_n7328_));
  AND2X1   g07136(.A(new_n7328_), .B(new_n7326_), .Y(new_n7329_));
  INVX1    g07137(.A(new_n7329_), .Y(new_n7330_));
  OR2X1    g07138(.A(new_n7315_), .B(\asqrt[48] ), .Y(new_n7331_));
  OAI21X1  g07139(.A0(new_n7331_), .A1(new_n7325_), .B0(new_n7330_), .Y(new_n7332_));
  AOI21X1  g07140(.A0(new_n7332_), .A1(new_n7324_), .B0(new_n1632_), .Y(new_n7333_));
  AOI21X1  g07141(.A0(new_n6936_), .A1(new_n6935_), .B0(new_n6903_), .Y(new_n7334_));
  AND2X1   g07142(.A(new_n7334_), .B(new_n6896_), .Y(new_n7335_));
  AOI22X1  g07143(.A0(new_n6936_), .A1(new_n6935_), .B0(new_n6922_), .B1(\asqrt[48] ), .Y(new_n7336_));
  AOI21X1  g07144(.A0(new_n7336_), .A1(\asqrt[31] ), .B0(new_n6902_), .Y(new_n7337_));
  AOI21X1  g07145(.A0(new_n7335_), .A1(\asqrt[31] ), .B0(new_n7337_), .Y(new_n7338_));
  OR2X1    g07146(.A(new_n7312_), .B(new_n2570_), .Y(new_n7339_));
  AND2X1   g07147(.A(new_n7296_), .B(new_n7287_), .Y(new_n7340_));
  INVX1    g07148(.A(new_n7301_), .Y(new_n7341_));
  OR2X1    g07149(.A(new_n7302_), .B(\asqrt[45] ), .Y(new_n7342_));
  OAI21X1  g07150(.A0(new_n7342_), .A1(new_n7340_), .B0(new_n7341_), .Y(new_n7343_));
  AOI21X1  g07151(.A0(new_n7343_), .A1(new_n7339_), .B0(new_n2263_), .Y(new_n7344_));
  AOI21X1  g07152(.A0(new_n7285_), .A1(\asqrt[45] ), .B0(\asqrt[46] ), .Y(new_n7345_));
  AOI21X1  g07153(.A0(new_n7345_), .A1(new_n7343_), .B0(new_n7310_), .Y(new_n7346_));
  OAI21X1  g07154(.A0(new_n7346_), .A1(new_n7344_), .B0(\asqrt[47] ), .Y(new_n7347_));
  NOR3X1   g07155(.A(new_n7346_), .B(new_n7344_), .C(\asqrt[47] ), .Y(new_n7348_));
  OAI21X1  g07156(.A0(new_n7348_), .A1(new_n7320_), .B0(new_n7347_), .Y(new_n7349_));
  AOI21X1  g07157(.A0(new_n7349_), .A1(\asqrt[48] ), .B0(\asqrt[49] ), .Y(new_n7350_));
  AOI21X1  g07158(.A0(new_n7350_), .A1(new_n7332_), .B0(new_n7338_), .Y(new_n7351_));
  OAI21X1  g07159(.A0(new_n7351_), .A1(new_n7333_), .B0(\asqrt[50] ), .Y(new_n7352_));
  AND2X1   g07160(.A(new_n6923_), .B(new_n6905_), .Y(new_n7353_));
  NOR3X1   g07161(.A(new_n7353_), .B(new_n6939_), .C(new_n6906_), .Y(new_n7354_));
  NOR3X1   g07162(.A(new_n7103_), .B(new_n7353_), .C(new_n6906_), .Y(new_n7355_));
  NOR2X1   g07163(.A(new_n7355_), .B(new_n6911_), .Y(new_n7356_));
  AOI21X1  g07164(.A0(new_n7354_), .A1(\asqrt[31] ), .B0(new_n7356_), .Y(new_n7357_));
  NOR3X1   g07165(.A(new_n7351_), .B(new_n7333_), .C(\asqrt[50] ), .Y(new_n7358_));
  OAI21X1  g07166(.A0(new_n7358_), .A1(new_n7357_), .B0(new_n7352_), .Y(new_n7359_));
  AND2X1   g07167(.A(new_n7359_), .B(\asqrt[51] ), .Y(new_n7360_));
  INVX1    g07168(.A(new_n7357_), .Y(new_n7361_));
  AND2X1   g07169(.A(new_n7349_), .B(\asqrt[48] ), .Y(new_n7362_));
  NAND2X1  g07170(.A(new_n7322_), .B(new_n7321_), .Y(new_n7363_));
  NOR2X1   g07171(.A(new_n7315_), .B(\asqrt[48] ), .Y(new_n7364_));
  AOI21X1  g07172(.A0(new_n7364_), .A1(new_n7363_), .B0(new_n7329_), .Y(new_n7365_));
  OAI21X1  g07173(.A0(new_n7365_), .A1(new_n7362_), .B0(\asqrt[49] ), .Y(new_n7366_));
  INVX1    g07174(.A(new_n7338_), .Y(new_n7367_));
  OAI21X1  g07175(.A0(new_n7323_), .A1(new_n1834_), .B0(new_n1632_), .Y(new_n7368_));
  OAI21X1  g07176(.A0(new_n7368_), .A1(new_n7365_), .B0(new_n7367_), .Y(new_n7369_));
  NAND3X1  g07177(.A(new_n7369_), .B(new_n7366_), .C(new_n1469_), .Y(new_n7370_));
  NAND2X1  g07178(.A(new_n7370_), .B(new_n7361_), .Y(new_n7371_));
  NAND4X1  g07179(.A(\asqrt[31] ), .B(new_n6942_), .C(new_n6929_), .D(new_n6925_), .Y(new_n7372_));
  NAND2X1  g07180(.A(new_n6942_), .B(new_n6925_), .Y(new_n7373_));
  OAI21X1  g07181(.A0(new_n7373_), .A1(new_n7103_), .B0(new_n6933_), .Y(new_n7374_));
  AND2X1   g07182(.A(new_n7374_), .B(new_n7372_), .Y(new_n7375_));
  AOI21X1  g07183(.A0(new_n7369_), .A1(new_n7366_), .B0(new_n1469_), .Y(new_n7376_));
  NOR2X1   g07184(.A(new_n7376_), .B(\asqrt[51] ), .Y(new_n7377_));
  AOI21X1  g07185(.A0(new_n7377_), .A1(new_n7371_), .B0(new_n7375_), .Y(new_n7378_));
  OAI21X1  g07186(.A0(new_n7378_), .A1(new_n7360_), .B0(\asqrt[52] ), .Y(new_n7379_));
  AND2X1   g07187(.A(new_n6950_), .B(new_n6943_), .Y(new_n7380_));
  NOR3X1   g07188(.A(new_n7380_), .B(new_n6988_), .C(new_n6932_), .Y(new_n7381_));
  NOR3X1   g07189(.A(new_n7103_), .B(new_n7380_), .C(new_n6932_), .Y(new_n7382_));
  NOR2X1   g07190(.A(new_n7382_), .B(new_n6948_), .Y(new_n7383_));
  AOI21X1  g07191(.A0(new_n7381_), .A1(\asqrt[31] ), .B0(new_n7383_), .Y(new_n7384_));
  INVX1    g07192(.A(new_n7384_), .Y(new_n7385_));
  AOI21X1  g07193(.A0(new_n7370_), .A1(new_n7361_), .B0(new_n7376_), .Y(new_n7386_));
  OAI21X1  g07194(.A0(new_n7386_), .A1(new_n1277_), .B0(new_n1111_), .Y(new_n7387_));
  OAI21X1  g07195(.A0(new_n7387_), .A1(new_n7378_), .B0(new_n7385_), .Y(new_n7388_));
  AOI21X1  g07196(.A0(new_n7388_), .A1(new_n7379_), .B0(new_n968_), .Y(new_n7389_));
  AND2X1   g07197(.A(new_n6992_), .B(new_n6990_), .Y(new_n7390_));
  NOR3X1   g07198(.A(new_n7390_), .B(new_n6958_), .C(new_n6991_), .Y(new_n7391_));
  NOR3X1   g07199(.A(new_n7103_), .B(new_n7390_), .C(new_n6991_), .Y(new_n7392_));
  NOR2X1   g07200(.A(new_n7392_), .B(new_n6957_), .Y(new_n7393_));
  AOI21X1  g07201(.A0(new_n7391_), .A1(\asqrt[31] ), .B0(new_n7393_), .Y(new_n7394_));
  INVX1    g07202(.A(new_n7394_), .Y(new_n7395_));
  NAND3X1  g07203(.A(new_n7388_), .B(new_n7379_), .C(new_n968_), .Y(new_n7396_));
  AOI21X1  g07204(.A0(new_n7396_), .A1(new_n7395_), .B0(new_n7389_), .Y(new_n7397_));
  OR2X1    g07205(.A(new_n7397_), .B(new_n902_), .Y(new_n7398_));
  OR2X1    g07206(.A(new_n7386_), .B(new_n1277_), .Y(new_n7399_));
  AND2X1   g07207(.A(new_n7370_), .B(new_n7361_), .Y(new_n7400_));
  INVX1    g07208(.A(new_n7375_), .Y(new_n7401_));
  OR2X1    g07209(.A(new_n7376_), .B(\asqrt[51] ), .Y(new_n7402_));
  OAI21X1  g07210(.A0(new_n7402_), .A1(new_n7400_), .B0(new_n7401_), .Y(new_n7403_));
  AOI21X1  g07211(.A0(new_n7403_), .A1(new_n7399_), .B0(new_n1111_), .Y(new_n7404_));
  AOI21X1  g07212(.A0(new_n7359_), .A1(\asqrt[51] ), .B0(\asqrt[52] ), .Y(new_n7405_));
  AOI21X1  g07213(.A0(new_n7405_), .A1(new_n7403_), .B0(new_n7384_), .Y(new_n7406_));
  NOR3X1   g07214(.A(new_n7406_), .B(new_n7404_), .C(\asqrt[53] ), .Y(new_n7407_));
  NOR2X1   g07215(.A(new_n7407_), .B(new_n7394_), .Y(new_n7408_));
  NAND4X1  g07216(.A(\asqrt[31] ), .B(new_n6968_), .C(new_n6966_), .D(new_n6994_), .Y(new_n7409_));
  NAND2X1  g07217(.A(new_n6968_), .B(new_n6994_), .Y(new_n7410_));
  OAI21X1  g07218(.A0(new_n7410_), .A1(new_n7103_), .B0(new_n6967_), .Y(new_n7411_));
  AND2X1   g07219(.A(new_n7411_), .B(new_n7409_), .Y(new_n7412_));
  INVX1    g07220(.A(new_n7412_), .Y(new_n7413_));
  OAI21X1  g07221(.A0(new_n7406_), .A1(new_n7404_), .B0(\asqrt[53] ), .Y(new_n7414_));
  NAND2X1  g07222(.A(new_n7414_), .B(new_n902_), .Y(new_n7415_));
  OAI21X1  g07223(.A0(new_n7415_), .A1(new_n7408_), .B0(new_n7413_), .Y(new_n7416_));
  AOI21X1  g07224(.A0(new_n7416_), .A1(new_n7398_), .B0(new_n697_), .Y(new_n7417_));
  AOI21X1  g07225(.A0(new_n7009_), .A1(new_n7008_), .B0(new_n6977_), .Y(new_n7418_));
  AND2X1   g07226(.A(new_n7418_), .B(new_n6970_), .Y(new_n7419_));
  AOI22X1  g07227(.A0(new_n7009_), .A1(new_n7008_), .B0(new_n6996_), .B1(\asqrt[54] ), .Y(new_n7420_));
  AOI21X1  g07228(.A0(new_n7420_), .A1(\asqrt[31] ), .B0(new_n6976_), .Y(new_n7421_));
  AOI21X1  g07229(.A0(new_n7419_), .A1(\asqrt[31] ), .B0(new_n7421_), .Y(new_n7422_));
  OAI21X1  g07230(.A0(new_n7407_), .A1(new_n7394_), .B0(new_n7414_), .Y(new_n7423_));
  AOI21X1  g07231(.A0(new_n7423_), .A1(\asqrt[54] ), .B0(\asqrt[55] ), .Y(new_n7424_));
  AOI21X1  g07232(.A0(new_n7424_), .A1(new_n7416_), .B0(new_n7422_), .Y(new_n7425_));
  OAI21X1  g07233(.A0(new_n7425_), .A1(new_n7417_), .B0(\asqrt[56] ), .Y(new_n7426_));
  AND2X1   g07234(.A(new_n6997_), .B(new_n6979_), .Y(new_n7427_));
  NOR3X1   g07235(.A(new_n7427_), .B(new_n7012_), .C(new_n6980_), .Y(new_n7428_));
  NOR3X1   g07236(.A(new_n7103_), .B(new_n7427_), .C(new_n6980_), .Y(new_n7429_));
  NOR2X1   g07237(.A(new_n7429_), .B(new_n6985_), .Y(new_n7430_));
  AOI21X1  g07238(.A0(new_n7428_), .A1(\asqrt[31] ), .B0(new_n7430_), .Y(new_n7431_));
  NOR3X1   g07239(.A(new_n7425_), .B(new_n7417_), .C(\asqrt[56] ), .Y(new_n7432_));
  OAI21X1  g07240(.A0(new_n7432_), .A1(new_n7431_), .B0(new_n7426_), .Y(new_n7433_));
  AND2X1   g07241(.A(new_n7433_), .B(\asqrt[57] ), .Y(new_n7434_));
  OR2X1    g07242(.A(new_n7432_), .B(new_n7431_), .Y(new_n7435_));
  OR4X1    g07243(.A(new_n7103_), .B(new_n7004_), .C(new_n7002_), .D(new_n7031_), .Y(new_n7436_));
  OR2X1    g07244(.A(new_n7004_), .B(new_n7031_), .Y(new_n7437_));
  OAI21X1  g07245(.A0(new_n7437_), .A1(new_n7103_), .B0(new_n7002_), .Y(new_n7438_));
  AND2X1   g07246(.A(new_n7438_), .B(new_n7436_), .Y(new_n7439_));
  AND2X1   g07247(.A(new_n7426_), .B(new_n481_), .Y(new_n7440_));
  AOI21X1  g07248(.A0(new_n7440_), .A1(new_n7435_), .B0(new_n7439_), .Y(new_n7441_));
  OAI21X1  g07249(.A0(new_n7441_), .A1(new_n7434_), .B0(\asqrt[58] ), .Y(new_n7442_));
  AND2X1   g07250(.A(new_n7022_), .B(new_n7016_), .Y(new_n7443_));
  NOR3X1   g07251(.A(new_n7443_), .B(new_n7046_), .C(new_n7006_), .Y(new_n7444_));
  NOR3X1   g07252(.A(new_n7103_), .B(new_n7443_), .C(new_n7006_), .Y(new_n7445_));
  NOR2X1   g07253(.A(new_n7445_), .B(new_n7021_), .Y(new_n7446_));
  AOI21X1  g07254(.A0(new_n7444_), .A1(\asqrt[31] ), .B0(new_n7446_), .Y(new_n7447_));
  INVX1    g07255(.A(new_n7447_), .Y(new_n7448_));
  AND2X1   g07256(.A(new_n7423_), .B(\asqrt[54] ), .Y(new_n7449_));
  OR2X1    g07257(.A(new_n7407_), .B(new_n7394_), .Y(new_n7450_));
  AND2X1   g07258(.A(new_n7414_), .B(new_n902_), .Y(new_n7451_));
  AOI21X1  g07259(.A0(new_n7451_), .A1(new_n7450_), .B0(new_n7412_), .Y(new_n7452_));
  OAI21X1  g07260(.A0(new_n7452_), .A1(new_n7449_), .B0(\asqrt[55] ), .Y(new_n7453_));
  INVX1    g07261(.A(new_n7422_), .Y(new_n7454_));
  OAI21X1  g07262(.A0(new_n7397_), .A1(new_n902_), .B0(new_n697_), .Y(new_n7455_));
  OAI21X1  g07263(.A0(new_n7455_), .A1(new_n7452_), .B0(new_n7454_), .Y(new_n7456_));
  AOI21X1  g07264(.A0(new_n7456_), .A1(new_n7453_), .B0(new_n582_), .Y(new_n7457_));
  INVX1    g07265(.A(new_n7431_), .Y(new_n7458_));
  NAND3X1  g07266(.A(new_n7456_), .B(new_n7453_), .C(new_n582_), .Y(new_n7459_));
  AOI21X1  g07267(.A0(new_n7459_), .A1(new_n7458_), .B0(new_n7457_), .Y(new_n7460_));
  OAI21X1  g07268(.A0(new_n7460_), .A1(new_n481_), .B0(new_n399_), .Y(new_n7461_));
  OAI21X1  g07269(.A0(new_n7461_), .A1(new_n7441_), .B0(new_n7448_), .Y(new_n7462_));
  AOI21X1  g07270(.A0(new_n7462_), .A1(new_n7442_), .B0(new_n328_), .Y(new_n7463_));
  AND2X1   g07271(.A(new_n7050_), .B(new_n7048_), .Y(new_n7464_));
  NOR3X1   g07272(.A(new_n7464_), .B(new_n7030_), .C(new_n7049_), .Y(new_n7465_));
  NOR3X1   g07273(.A(new_n7103_), .B(new_n7464_), .C(new_n7049_), .Y(new_n7466_));
  NOR2X1   g07274(.A(new_n7466_), .B(new_n7029_), .Y(new_n7467_));
  AOI21X1  g07275(.A0(new_n7465_), .A1(\asqrt[31] ), .B0(new_n7467_), .Y(new_n7468_));
  INVX1    g07276(.A(new_n7468_), .Y(new_n7469_));
  NAND3X1  g07277(.A(new_n7462_), .B(new_n7442_), .C(new_n328_), .Y(new_n7470_));
  AOI21X1  g07278(.A0(new_n7470_), .A1(new_n7469_), .B0(new_n7463_), .Y(new_n7471_));
  OR2X1    g07279(.A(new_n7471_), .B(new_n292_), .Y(new_n7472_));
  OR2X1    g07280(.A(new_n7460_), .B(new_n481_), .Y(new_n7473_));
  NOR2X1   g07281(.A(new_n7432_), .B(new_n7431_), .Y(new_n7474_));
  INVX1    g07282(.A(new_n7439_), .Y(new_n7475_));
  NAND2X1  g07283(.A(new_n7426_), .B(new_n481_), .Y(new_n7476_));
  OAI21X1  g07284(.A0(new_n7476_), .A1(new_n7474_), .B0(new_n7475_), .Y(new_n7477_));
  AOI21X1  g07285(.A0(new_n7477_), .A1(new_n7473_), .B0(new_n399_), .Y(new_n7478_));
  AOI21X1  g07286(.A0(new_n7433_), .A1(\asqrt[57] ), .B0(\asqrt[58] ), .Y(new_n7479_));
  AOI21X1  g07287(.A0(new_n7479_), .A1(new_n7477_), .B0(new_n7447_), .Y(new_n7480_));
  NOR3X1   g07288(.A(new_n7480_), .B(new_n7478_), .C(\asqrt[59] ), .Y(new_n7481_));
  NOR2X1   g07289(.A(new_n7481_), .B(new_n7468_), .Y(new_n7482_));
  OR4X1    g07290(.A(new_n7103_), .B(new_n7052_), .C(new_n7040_), .D(new_n7035_), .Y(new_n7483_));
  OR2X1    g07291(.A(new_n7052_), .B(new_n7035_), .Y(new_n7484_));
  OAI21X1  g07292(.A0(new_n7484_), .A1(new_n7103_), .B0(new_n7040_), .Y(new_n7485_));
  AND2X1   g07293(.A(new_n7485_), .B(new_n7483_), .Y(new_n7486_));
  INVX1    g07294(.A(new_n7486_), .Y(new_n7487_));
  OAI21X1  g07295(.A0(new_n7480_), .A1(new_n7478_), .B0(\asqrt[59] ), .Y(new_n7488_));
  NAND2X1  g07296(.A(new_n7488_), .B(new_n292_), .Y(new_n7489_));
  OAI21X1  g07297(.A0(new_n7489_), .A1(new_n7482_), .B0(new_n7487_), .Y(new_n7490_));
  AOI21X1  g07298(.A0(new_n7490_), .A1(new_n7472_), .B0(new_n217_), .Y(new_n7491_));
  AOI21X1  g07299(.A0(new_n7112_), .A1(new_n7111_), .B0(new_n7059_), .Y(new_n7492_));
  AND2X1   g07300(.A(new_n7492_), .B(new_n7043_), .Y(new_n7493_));
  AOI22X1  g07301(.A0(new_n7112_), .A1(new_n7111_), .B0(new_n7069_), .B1(\asqrt[60] ), .Y(new_n7494_));
  AOI21X1  g07302(.A0(new_n7494_), .A1(\asqrt[31] ), .B0(new_n7058_), .Y(new_n7495_));
  AOI21X1  g07303(.A0(new_n7493_), .A1(\asqrt[31] ), .B0(new_n7495_), .Y(new_n7496_));
  OAI21X1  g07304(.A0(new_n7481_), .A1(new_n7468_), .B0(new_n7488_), .Y(new_n7497_));
  AOI21X1  g07305(.A0(new_n7497_), .A1(\asqrt[60] ), .B0(\asqrt[61] ), .Y(new_n7498_));
  AOI21X1  g07306(.A0(new_n7498_), .A1(new_n7490_), .B0(new_n7496_), .Y(new_n7499_));
  OAI21X1  g07307(.A0(new_n7499_), .A1(new_n7491_), .B0(\asqrt[62] ), .Y(new_n7500_));
  AND2X1   g07308(.A(new_n7070_), .B(new_n7062_), .Y(new_n7501_));
  NOR3X1   g07309(.A(new_n7501_), .B(new_n7115_), .C(new_n7063_), .Y(new_n7502_));
  NOR3X1   g07310(.A(new_n7103_), .B(new_n7501_), .C(new_n7063_), .Y(new_n7503_));
  NOR2X1   g07311(.A(new_n7503_), .B(new_n7068_), .Y(new_n7504_));
  AOI21X1  g07312(.A0(new_n7502_), .A1(\asqrt[31] ), .B0(new_n7504_), .Y(new_n7505_));
  NOR3X1   g07313(.A(new_n7499_), .B(new_n7491_), .C(\asqrt[62] ), .Y(new_n7506_));
  OAI21X1  g07314(.A0(new_n7506_), .A1(new_n7505_), .B0(new_n7500_), .Y(new_n7507_));
  NOR4X1   g07315(.A(new_n7103_), .B(new_n7077_), .C(new_n7119_), .D(new_n7118_), .Y(new_n7508_));
  NAND3X1  g07316(.A(\asqrt[31] ), .B(new_n7120_), .C(new_n7072_), .Y(new_n7509_));
  AOI21X1  g07317(.A0(new_n7509_), .A1(new_n7119_), .B0(new_n7508_), .Y(new_n7510_));
  INVX1    g07318(.A(new_n7510_), .Y(new_n7511_));
  AND2X1   g07319(.A(new_n7084_), .B(new_n7078_), .Y(new_n7512_));
  AOI21X1  g07320(.A0(new_n7512_), .A1(\asqrt[31] ), .B0(new_n7144_), .Y(new_n7513_));
  AND2X1   g07321(.A(new_n7513_), .B(new_n7511_), .Y(new_n7514_));
  AOI21X1  g07322(.A0(new_n7514_), .A1(new_n7507_), .B0(\asqrt[63] ), .Y(new_n7515_));
  NOR2X1   g07323(.A(new_n7506_), .B(new_n7505_), .Y(new_n7516_));
  NAND2X1  g07324(.A(new_n7510_), .B(new_n7500_), .Y(new_n7517_));
  AOI21X1  g07325(.A0(new_n7127_), .A1(new_n7123_), .B0(new_n7083_), .Y(new_n7518_));
  AOI21X1  g07326(.A0(new_n7084_), .A1(new_n7078_), .B0(new_n193_), .Y(new_n7519_));
  OAI21X1  g07327(.A0(new_n7518_), .A1(new_n7078_), .B0(new_n7519_), .Y(new_n7520_));
  NOR4X1   g07328(.A(new_n7100_), .B(new_n7145_), .C(new_n7082_), .D(new_n7080_), .Y(new_n7521_));
  OAI21X1  g07329(.A0(new_n7091_), .A1(new_n7090_), .B0(new_n7521_), .Y(new_n7522_));
  NOR2X1   g07330(.A(new_n7522_), .B(new_n7089_), .Y(new_n7523_));
  INVX1    g07331(.A(new_n7523_), .Y(new_n7524_));
  AND2X1   g07332(.A(new_n7524_), .B(new_n7520_), .Y(new_n7525_));
  OAI21X1  g07333(.A0(new_n7517_), .A1(new_n7516_), .B0(new_n7525_), .Y(new_n7526_));
  NOR2X1   g07334(.A(new_n7526_), .B(new_n7515_), .Y(new_n7527_));
  INVX1    g07335(.A(\a[60] ), .Y(new_n7528_));
  AND2X1   g07336(.A(new_n7497_), .B(\asqrt[60] ), .Y(new_n7529_));
  OR2X1    g07337(.A(new_n7481_), .B(new_n7468_), .Y(new_n7530_));
  AND2X1   g07338(.A(new_n7488_), .B(new_n292_), .Y(new_n7531_));
  AOI21X1  g07339(.A0(new_n7531_), .A1(new_n7530_), .B0(new_n7486_), .Y(new_n7532_));
  OAI21X1  g07340(.A0(new_n7532_), .A1(new_n7529_), .B0(\asqrt[61] ), .Y(new_n7533_));
  INVX1    g07341(.A(new_n7496_), .Y(new_n7534_));
  OAI21X1  g07342(.A0(new_n7471_), .A1(new_n292_), .B0(new_n217_), .Y(new_n7535_));
  OAI21X1  g07343(.A0(new_n7535_), .A1(new_n7532_), .B0(new_n7534_), .Y(new_n7536_));
  AOI21X1  g07344(.A0(new_n7536_), .A1(new_n7533_), .B0(new_n199_), .Y(new_n7537_));
  INVX1    g07345(.A(new_n7505_), .Y(new_n7538_));
  NAND3X1  g07346(.A(new_n7536_), .B(new_n7533_), .C(new_n199_), .Y(new_n7539_));
  AOI21X1  g07347(.A0(new_n7539_), .A1(new_n7538_), .B0(new_n7537_), .Y(new_n7540_));
  INVX1    g07348(.A(new_n7514_), .Y(new_n7541_));
  OAI21X1  g07349(.A0(new_n7541_), .A1(new_n7540_), .B0(new_n193_), .Y(new_n7542_));
  OR2X1    g07350(.A(new_n7506_), .B(new_n7505_), .Y(new_n7543_));
  AND2X1   g07351(.A(new_n7510_), .B(new_n7500_), .Y(new_n7544_));
  INVX1    g07352(.A(new_n7525_), .Y(new_n7545_));
  AOI21X1  g07353(.A0(new_n7544_), .A1(new_n7543_), .B0(new_n7545_), .Y(new_n7546_));
  AOI21X1  g07354(.A0(new_n7546_), .A1(new_n7542_), .B0(new_n7528_), .Y(new_n7547_));
  NOR3X1   g07355(.A(\a[60] ), .B(\a[59] ), .C(\a[58] ), .Y(new_n7548_));
  OAI21X1  g07356(.A0(new_n7548_), .A1(new_n7547_), .B0(\asqrt[31] ), .Y(new_n7549_));
  OR2X1    g07357(.A(new_n7548_), .B(new_n7100_), .Y(new_n7550_));
  NOR4X1   g07358(.A(new_n7550_), .B(new_n7145_), .C(new_n7144_), .D(new_n7089_), .Y(new_n7551_));
  INVX1    g07359(.A(new_n7551_), .Y(new_n7552_));
  NOR2X1   g07360(.A(new_n7552_), .B(new_n7547_), .Y(new_n7553_));
  INVX1    g07361(.A(\a[61] ), .Y(new_n7554_));
  AOI21X1  g07362(.A0(new_n7546_), .A1(new_n7542_), .B0(\a[60] ), .Y(new_n7555_));
  OAI21X1  g07363(.A0(new_n7526_), .A1(new_n7515_), .B0(new_n7107_), .Y(new_n7556_));
  OAI21X1  g07364(.A0(new_n7555_), .A1(new_n7554_), .B0(new_n7556_), .Y(new_n7557_));
  OAI21X1  g07365(.A0(new_n7557_), .A1(new_n7553_), .B0(new_n7549_), .Y(new_n7558_));
  AND2X1   g07366(.A(new_n7558_), .B(\asqrt[32] ), .Y(new_n7559_));
  OR2X1    g07367(.A(new_n7557_), .B(new_n7553_), .Y(new_n7560_));
  AND2X1   g07368(.A(new_n7549_), .B(new_n6699_), .Y(new_n7561_));
  INVX1    g07369(.A(new_n7520_), .Y(new_n7562_));
  NOR3X1   g07370(.A(new_n7523_), .B(new_n7562_), .C(new_n7103_), .Y(new_n7563_));
  OAI21X1  g07371(.A0(new_n7517_), .A1(new_n7516_), .B0(new_n7563_), .Y(new_n7564_));
  OR2X1    g07372(.A(new_n7564_), .B(new_n7515_), .Y(new_n7565_));
  AOI21X1  g07373(.A0(new_n7565_), .A1(new_n7556_), .B0(new_n7106_), .Y(new_n7566_));
  INVX1    g07374(.A(new_n7107_), .Y(new_n7567_));
  AOI21X1  g07375(.A0(new_n7546_), .A1(new_n7542_), .B0(new_n7567_), .Y(new_n7568_));
  OAI21X1  g07376(.A0(new_n7564_), .A1(new_n7515_), .B0(new_n7106_), .Y(new_n7569_));
  NOR2X1   g07377(.A(new_n7569_), .B(new_n7568_), .Y(new_n7570_));
  NOR2X1   g07378(.A(new_n7570_), .B(new_n7566_), .Y(new_n7571_));
  AOI21X1  g07379(.A0(new_n7561_), .A1(new_n7560_), .B0(new_n7571_), .Y(new_n7572_));
  OAI21X1  g07380(.A0(new_n7572_), .A1(new_n7559_), .B0(\asqrt[33] ), .Y(new_n7573_));
  NOR3X1   g07381(.A(new_n7140_), .B(new_n7130_), .C(new_n7142_), .Y(new_n7574_));
  OAI21X1  g07382(.A0(new_n7526_), .A1(new_n7515_), .B0(new_n7574_), .Y(new_n7575_));
  NOR2X1   g07383(.A(new_n7130_), .B(new_n7142_), .Y(new_n7576_));
  OAI21X1  g07384(.A0(new_n7526_), .A1(new_n7515_), .B0(new_n7576_), .Y(new_n7577_));
  NAND2X1  g07385(.A(new_n7577_), .B(new_n7140_), .Y(new_n7578_));
  NAND2X1  g07386(.A(new_n7578_), .B(new_n7575_), .Y(new_n7579_));
  OR2X1    g07387(.A(new_n7548_), .B(new_n7547_), .Y(new_n7580_));
  OR2X1    g07388(.A(new_n7552_), .B(new_n7547_), .Y(new_n7581_));
  OAI21X1  g07389(.A0(new_n7526_), .A1(new_n7515_), .B0(new_n7528_), .Y(new_n7582_));
  AOI21X1  g07390(.A0(new_n7582_), .A1(\a[61] ), .B0(new_n7568_), .Y(new_n7583_));
  AOI22X1  g07391(.A0(new_n7583_), .A1(new_n7581_), .B0(new_n7580_), .B1(\asqrt[31] ), .Y(new_n7584_));
  OAI21X1  g07392(.A0(new_n7584_), .A1(new_n6699_), .B0(new_n6294_), .Y(new_n7585_));
  OAI21X1  g07393(.A0(new_n7585_), .A1(new_n7572_), .B0(new_n7579_), .Y(new_n7586_));
  AOI21X1  g07394(.A0(new_n7586_), .A1(new_n7573_), .B0(new_n5941_), .Y(new_n7587_));
  AOI21X1  g07395(.A0(new_n7143_), .A1(new_n7141_), .B0(new_n7179_), .Y(new_n7588_));
  AND2X1   g07396(.A(new_n7588_), .B(new_n7176_), .Y(new_n7589_));
  OAI21X1  g07397(.A0(new_n7526_), .A1(new_n7515_), .B0(new_n7589_), .Y(new_n7590_));
  AOI22X1  g07398(.A0(new_n7143_), .A1(new_n7141_), .B0(new_n7135_), .B1(\asqrt[33] ), .Y(new_n7591_));
  OAI21X1  g07399(.A0(new_n7526_), .A1(new_n7515_), .B0(new_n7591_), .Y(new_n7592_));
  NAND2X1  g07400(.A(new_n7592_), .B(new_n7179_), .Y(new_n7593_));
  AND2X1   g07401(.A(new_n7593_), .B(new_n7590_), .Y(new_n7594_));
  INVX1    g07402(.A(new_n7594_), .Y(new_n7595_));
  NAND3X1  g07403(.A(new_n7586_), .B(new_n7573_), .C(new_n5941_), .Y(new_n7596_));
  AOI21X1  g07404(.A0(new_n7596_), .A1(new_n7595_), .B0(new_n7587_), .Y(new_n7597_));
  OR2X1    g07405(.A(new_n7597_), .B(new_n5541_), .Y(new_n7598_));
  OR2X1    g07406(.A(new_n7584_), .B(new_n6699_), .Y(new_n7599_));
  AND2X1   g07407(.A(new_n7583_), .B(new_n7581_), .Y(new_n7600_));
  NAND2X1  g07408(.A(new_n7549_), .B(new_n6699_), .Y(new_n7601_));
  OR2X1    g07409(.A(new_n7570_), .B(new_n7566_), .Y(new_n7602_));
  OAI21X1  g07410(.A0(new_n7601_), .A1(new_n7600_), .B0(new_n7602_), .Y(new_n7603_));
  AOI21X1  g07411(.A0(new_n7603_), .A1(new_n7599_), .B0(new_n6294_), .Y(new_n7604_));
  AND2X1   g07412(.A(new_n7578_), .B(new_n7575_), .Y(new_n7605_));
  AOI21X1  g07413(.A0(new_n7558_), .A1(\asqrt[32] ), .B0(\asqrt[33] ), .Y(new_n7606_));
  AOI21X1  g07414(.A0(new_n7606_), .A1(new_n7603_), .B0(new_n7605_), .Y(new_n7607_));
  NOR3X1   g07415(.A(new_n7607_), .B(new_n7604_), .C(\asqrt[34] ), .Y(new_n7608_));
  NOR2X1   g07416(.A(new_n7608_), .B(new_n7594_), .Y(new_n7609_));
  OAI21X1  g07417(.A0(new_n7607_), .A1(new_n7604_), .B0(\asqrt[34] ), .Y(new_n7610_));
  NAND2X1  g07418(.A(new_n7610_), .B(new_n5541_), .Y(new_n7611_));
  INVX1    g07419(.A(new_n7527_), .Y(\asqrt[30] ));
  AND2X1   g07420(.A(new_n7182_), .B(new_n7180_), .Y(new_n7613_));
  NOR3X1   g07421(.A(new_n7162_), .B(new_n7613_), .C(new_n7181_), .Y(new_n7614_));
  NOR2X1   g07422(.A(new_n7613_), .B(new_n7181_), .Y(new_n7615_));
  OAI21X1  g07423(.A0(new_n7526_), .A1(new_n7515_), .B0(new_n7615_), .Y(new_n7616_));
  AOI22X1  g07424(.A0(new_n7616_), .A1(new_n7162_), .B0(new_n7614_), .B1(\asqrt[30] ), .Y(new_n7617_));
  INVX1    g07425(.A(new_n7617_), .Y(new_n7618_));
  OAI21X1  g07426(.A0(new_n7611_), .A1(new_n7609_), .B0(new_n7618_), .Y(new_n7619_));
  AOI21X1  g07427(.A0(new_n7619_), .A1(new_n7598_), .B0(new_n5176_), .Y(new_n7620_));
  NAND4X1  g07428(.A(\asqrt[30] ), .B(new_n7173_), .C(new_n7171_), .D(new_n7200_), .Y(new_n7621_));
  NOR3X1   g07429(.A(new_n7527_), .B(new_n7184_), .C(new_n7164_), .Y(new_n7622_));
  OAI21X1  g07430(.A0(new_n7622_), .A1(new_n7171_), .B0(new_n7621_), .Y(new_n7623_));
  INVX1    g07431(.A(new_n7623_), .Y(new_n7624_));
  OAI21X1  g07432(.A0(new_n7608_), .A1(new_n7594_), .B0(new_n7610_), .Y(new_n7625_));
  AOI21X1  g07433(.A0(new_n7625_), .A1(\asqrt[35] ), .B0(\asqrt[36] ), .Y(new_n7626_));
  AOI21X1  g07434(.A0(new_n7626_), .A1(new_n7619_), .B0(new_n7624_), .Y(new_n7627_));
  OAI21X1  g07435(.A0(new_n7627_), .A1(new_n7620_), .B0(\asqrt[37] ), .Y(new_n7628_));
  AND2X1   g07436(.A(new_n7229_), .B(new_n7228_), .Y(new_n7629_));
  NOR3X1   g07437(.A(new_n7629_), .B(new_n7191_), .C(new_n7227_), .Y(new_n7630_));
  NOR3X1   g07438(.A(new_n7527_), .B(new_n7629_), .C(new_n7227_), .Y(new_n7631_));
  NOR2X1   g07439(.A(new_n7631_), .B(new_n7190_), .Y(new_n7632_));
  AOI21X1  g07440(.A0(new_n7630_), .A1(\asqrt[30] ), .B0(new_n7632_), .Y(new_n7633_));
  NOR3X1   g07441(.A(new_n7627_), .B(new_n7620_), .C(\asqrt[37] ), .Y(new_n7634_));
  OAI21X1  g07442(.A0(new_n7634_), .A1(new_n7633_), .B0(new_n7628_), .Y(new_n7635_));
  AND2X1   g07443(.A(new_n7635_), .B(\asqrt[38] ), .Y(new_n7636_));
  INVX1    g07444(.A(new_n7633_), .Y(new_n7637_));
  AND2X1   g07445(.A(new_n7625_), .B(\asqrt[35] ), .Y(new_n7638_));
  OR2X1    g07446(.A(new_n7608_), .B(new_n7594_), .Y(new_n7639_));
  AND2X1   g07447(.A(new_n7610_), .B(new_n5541_), .Y(new_n7640_));
  AOI21X1  g07448(.A0(new_n7640_), .A1(new_n7639_), .B0(new_n7617_), .Y(new_n7641_));
  OAI21X1  g07449(.A0(new_n7641_), .A1(new_n7638_), .B0(\asqrt[36] ), .Y(new_n7642_));
  OAI21X1  g07450(.A0(new_n7597_), .A1(new_n5541_), .B0(new_n5176_), .Y(new_n7643_));
  OAI21X1  g07451(.A0(new_n7643_), .A1(new_n7641_), .B0(new_n7623_), .Y(new_n7644_));
  NAND3X1  g07452(.A(new_n7644_), .B(new_n7642_), .C(new_n4826_), .Y(new_n7645_));
  NAND2X1  g07453(.A(new_n7645_), .B(new_n7637_), .Y(new_n7646_));
  AND2X1   g07454(.A(new_n7202_), .B(new_n7193_), .Y(new_n7647_));
  NOR3X1   g07455(.A(new_n7647_), .B(new_n7232_), .C(new_n7194_), .Y(new_n7648_));
  NOR3X1   g07456(.A(new_n7527_), .B(new_n7647_), .C(new_n7194_), .Y(new_n7649_));
  NOR2X1   g07457(.A(new_n7649_), .B(new_n7199_), .Y(new_n7650_));
  AOI21X1  g07458(.A0(new_n7648_), .A1(\asqrt[30] ), .B0(new_n7650_), .Y(new_n7651_));
  AND2X1   g07459(.A(new_n7628_), .B(new_n4493_), .Y(new_n7652_));
  AOI21X1  g07460(.A0(new_n7652_), .A1(new_n7646_), .B0(new_n7651_), .Y(new_n7653_));
  OAI21X1  g07461(.A0(new_n7653_), .A1(new_n7636_), .B0(\asqrt[39] ), .Y(new_n7654_));
  OR4X1    g07462(.A(new_n7527_), .B(new_n7210_), .C(new_n7236_), .D(new_n7235_), .Y(new_n7655_));
  OR2X1    g07463(.A(new_n7210_), .B(new_n7235_), .Y(new_n7656_));
  OAI21X1  g07464(.A0(new_n7656_), .A1(new_n7527_), .B0(new_n7236_), .Y(new_n7657_));
  AND2X1   g07465(.A(new_n7657_), .B(new_n7655_), .Y(new_n7658_));
  INVX1    g07466(.A(new_n7658_), .Y(new_n7659_));
  AOI21X1  g07467(.A0(new_n7644_), .A1(new_n7642_), .B0(new_n4826_), .Y(new_n7660_));
  AOI21X1  g07468(.A0(new_n7645_), .A1(new_n7637_), .B0(new_n7660_), .Y(new_n7661_));
  OAI21X1  g07469(.A0(new_n7661_), .A1(new_n4493_), .B0(new_n4165_), .Y(new_n7662_));
  OAI21X1  g07470(.A0(new_n7662_), .A1(new_n7653_), .B0(new_n7659_), .Y(new_n7663_));
  AOI21X1  g07471(.A0(new_n7663_), .A1(new_n7654_), .B0(new_n3863_), .Y(new_n7664_));
  AOI21X1  g07472(.A0(new_n7218_), .A1(new_n7213_), .B0(new_n7267_), .Y(new_n7665_));
  AND2X1   g07473(.A(new_n7665_), .B(new_n7265_), .Y(new_n7666_));
  AOI22X1  g07474(.A0(new_n7218_), .A1(new_n7213_), .B0(new_n7211_), .B1(\asqrt[39] ), .Y(new_n7667_));
  AOI21X1  g07475(.A0(new_n7667_), .A1(\asqrt[30] ), .B0(new_n7217_), .Y(new_n7668_));
  AOI21X1  g07476(.A0(new_n7666_), .A1(\asqrt[30] ), .B0(new_n7668_), .Y(new_n7669_));
  INVX1    g07477(.A(new_n7669_), .Y(new_n7670_));
  NAND3X1  g07478(.A(new_n7663_), .B(new_n7654_), .C(new_n3863_), .Y(new_n7671_));
  AOI21X1  g07479(.A0(new_n7671_), .A1(new_n7670_), .B0(new_n7664_), .Y(new_n7672_));
  OR2X1    g07480(.A(new_n7672_), .B(new_n3564_), .Y(new_n7673_));
  AND2X1   g07481(.A(new_n7671_), .B(new_n7670_), .Y(new_n7674_));
  AND2X1   g07482(.A(new_n7271_), .B(new_n7269_), .Y(new_n7675_));
  NOR3X1   g07483(.A(new_n7675_), .B(new_n7226_), .C(new_n7270_), .Y(new_n7676_));
  NOR3X1   g07484(.A(new_n7527_), .B(new_n7675_), .C(new_n7270_), .Y(new_n7677_));
  NOR2X1   g07485(.A(new_n7677_), .B(new_n7225_), .Y(new_n7678_));
  AOI21X1  g07486(.A0(new_n7676_), .A1(\asqrt[30] ), .B0(new_n7678_), .Y(new_n7679_));
  INVX1    g07487(.A(new_n7679_), .Y(new_n7680_));
  OR2X1    g07488(.A(new_n7661_), .B(new_n4493_), .Y(new_n7681_));
  AND2X1   g07489(.A(new_n7645_), .B(new_n7637_), .Y(new_n7682_));
  INVX1    g07490(.A(new_n7651_), .Y(new_n7683_));
  NAND2X1  g07491(.A(new_n7628_), .B(new_n4493_), .Y(new_n7684_));
  OAI21X1  g07492(.A0(new_n7684_), .A1(new_n7682_), .B0(new_n7683_), .Y(new_n7685_));
  AOI21X1  g07493(.A0(new_n7685_), .A1(new_n7681_), .B0(new_n4165_), .Y(new_n7686_));
  AOI21X1  g07494(.A0(new_n7635_), .A1(\asqrt[38] ), .B0(\asqrt[39] ), .Y(new_n7687_));
  AOI21X1  g07495(.A0(new_n7687_), .A1(new_n7685_), .B0(new_n7658_), .Y(new_n7688_));
  OAI21X1  g07496(.A0(new_n7688_), .A1(new_n7686_), .B0(\asqrt[40] ), .Y(new_n7689_));
  NAND2X1  g07497(.A(new_n7689_), .B(new_n3564_), .Y(new_n7690_));
  OAI21X1  g07498(.A0(new_n7690_), .A1(new_n7674_), .B0(new_n7680_), .Y(new_n7691_));
  AOI21X1  g07499(.A0(new_n7691_), .A1(new_n7673_), .B0(new_n3276_), .Y(new_n7692_));
  NAND4X1  g07500(.A(\asqrt[30] ), .B(new_n7248_), .C(new_n7246_), .D(new_n7273_), .Y(new_n7693_));
  NAND2X1  g07501(.A(new_n7248_), .B(new_n7273_), .Y(new_n7694_));
  OAI21X1  g07502(.A0(new_n7694_), .A1(new_n7527_), .B0(new_n7247_), .Y(new_n7695_));
  AND2X1   g07503(.A(new_n7695_), .B(new_n7693_), .Y(new_n7696_));
  NOR3X1   g07504(.A(new_n7688_), .B(new_n7686_), .C(\asqrt[40] ), .Y(new_n7697_));
  OAI21X1  g07505(.A0(new_n7697_), .A1(new_n7669_), .B0(new_n7689_), .Y(new_n7698_));
  AOI21X1  g07506(.A0(new_n7698_), .A1(\asqrt[41] ), .B0(\asqrt[42] ), .Y(new_n7699_));
  AOI21X1  g07507(.A0(new_n7699_), .A1(new_n7691_), .B0(new_n7696_), .Y(new_n7700_));
  OAI21X1  g07508(.A0(new_n7700_), .A1(new_n7692_), .B0(\asqrt[43] ), .Y(new_n7701_));
  AND2X1   g07509(.A(new_n7290_), .B(new_n7289_), .Y(new_n7702_));
  NOR3X1   g07510(.A(new_n7702_), .B(new_n7256_), .C(new_n7288_), .Y(new_n7703_));
  NOR3X1   g07511(.A(new_n7527_), .B(new_n7702_), .C(new_n7288_), .Y(new_n7704_));
  NOR2X1   g07512(.A(new_n7704_), .B(new_n7255_), .Y(new_n7705_));
  AOI21X1  g07513(.A0(new_n7703_), .A1(\asqrt[30] ), .B0(new_n7705_), .Y(new_n7706_));
  NOR3X1   g07514(.A(new_n7700_), .B(new_n7692_), .C(\asqrt[43] ), .Y(new_n7707_));
  OAI21X1  g07515(.A0(new_n7707_), .A1(new_n7706_), .B0(new_n7701_), .Y(new_n7708_));
  AND2X1   g07516(.A(new_n7708_), .B(\asqrt[44] ), .Y(new_n7709_));
  INVX1    g07517(.A(new_n7706_), .Y(new_n7710_));
  AND2X1   g07518(.A(new_n7698_), .B(\asqrt[41] ), .Y(new_n7711_));
  NAND2X1  g07519(.A(new_n7671_), .B(new_n7670_), .Y(new_n7712_));
  AND2X1   g07520(.A(new_n7689_), .B(new_n3564_), .Y(new_n7713_));
  AOI21X1  g07521(.A0(new_n7713_), .A1(new_n7712_), .B0(new_n7679_), .Y(new_n7714_));
  OAI21X1  g07522(.A0(new_n7714_), .A1(new_n7711_), .B0(\asqrt[42] ), .Y(new_n7715_));
  INVX1    g07523(.A(new_n7696_), .Y(new_n7716_));
  OAI21X1  g07524(.A0(new_n7672_), .A1(new_n3564_), .B0(new_n3276_), .Y(new_n7717_));
  OAI21X1  g07525(.A0(new_n7717_), .A1(new_n7714_), .B0(new_n7716_), .Y(new_n7718_));
  NAND3X1  g07526(.A(new_n7718_), .B(new_n7715_), .C(new_n3008_), .Y(new_n7719_));
  NAND2X1  g07527(.A(new_n7719_), .B(new_n7710_), .Y(new_n7720_));
  AND2X1   g07528(.A(new_n7276_), .B(new_n7258_), .Y(new_n7721_));
  NOR3X1   g07529(.A(new_n7721_), .B(new_n7293_), .C(new_n7259_), .Y(new_n7722_));
  NOR3X1   g07530(.A(new_n7527_), .B(new_n7721_), .C(new_n7259_), .Y(new_n7723_));
  NOR2X1   g07531(.A(new_n7723_), .B(new_n7264_), .Y(new_n7724_));
  AOI21X1  g07532(.A0(new_n7722_), .A1(\asqrt[30] ), .B0(new_n7724_), .Y(new_n7725_));
  AND2X1   g07533(.A(new_n7701_), .B(new_n2769_), .Y(new_n7726_));
  AOI21X1  g07534(.A0(new_n7726_), .A1(new_n7720_), .B0(new_n7725_), .Y(new_n7727_));
  OAI21X1  g07535(.A0(new_n7727_), .A1(new_n7709_), .B0(\asqrt[45] ), .Y(new_n7728_));
  NAND4X1  g07536(.A(\asqrt[30] ), .B(new_n7296_), .C(new_n7283_), .D(new_n7278_), .Y(new_n7729_));
  NAND2X1  g07537(.A(new_n7296_), .B(new_n7278_), .Y(new_n7730_));
  OAI21X1  g07538(.A0(new_n7730_), .A1(new_n7527_), .B0(new_n7287_), .Y(new_n7731_));
  AND2X1   g07539(.A(new_n7731_), .B(new_n7729_), .Y(new_n7732_));
  INVX1    g07540(.A(new_n7732_), .Y(new_n7733_));
  AOI21X1  g07541(.A0(new_n7718_), .A1(new_n7715_), .B0(new_n3008_), .Y(new_n7734_));
  AOI21X1  g07542(.A0(new_n7719_), .A1(new_n7710_), .B0(new_n7734_), .Y(new_n7735_));
  OAI21X1  g07543(.A0(new_n7735_), .A1(new_n2769_), .B0(new_n2570_), .Y(new_n7736_));
  OAI21X1  g07544(.A0(new_n7736_), .A1(new_n7727_), .B0(new_n7733_), .Y(new_n7737_));
  AOI21X1  g07545(.A0(new_n7737_), .A1(new_n7728_), .B0(new_n2263_), .Y(new_n7738_));
  AOI21X1  g07546(.A0(new_n7303_), .A1(new_n7297_), .B0(new_n7341_), .Y(new_n7739_));
  AND2X1   g07547(.A(new_n7739_), .B(new_n7339_), .Y(new_n7740_));
  AOI22X1  g07548(.A0(new_n7303_), .A1(new_n7297_), .B0(new_n7285_), .B1(\asqrt[45] ), .Y(new_n7741_));
  AOI21X1  g07549(.A0(new_n7741_), .A1(\asqrt[30] ), .B0(new_n7301_), .Y(new_n7742_));
  AOI21X1  g07550(.A0(new_n7740_), .A1(\asqrt[30] ), .B0(new_n7742_), .Y(new_n7743_));
  INVX1    g07551(.A(new_n7743_), .Y(new_n7744_));
  NAND3X1  g07552(.A(new_n7737_), .B(new_n7728_), .C(new_n2263_), .Y(new_n7745_));
  AOI21X1  g07553(.A0(new_n7745_), .A1(new_n7744_), .B0(new_n7738_), .Y(new_n7746_));
  OR2X1    g07554(.A(new_n7746_), .B(new_n2040_), .Y(new_n7747_));
  AND2X1   g07555(.A(new_n7745_), .B(new_n7744_), .Y(new_n7748_));
  AND2X1   g07556(.A(new_n7345_), .B(new_n7343_), .Y(new_n7749_));
  NOR3X1   g07557(.A(new_n7749_), .B(new_n7311_), .C(new_n7344_), .Y(new_n7750_));
  NOR3X1   g07558(.A(new_n7527_), .B(new_n7749_), .C(new_n7344_), .Y(new_n7751_));
  NOR2X1   g07559(.A(new_n7751_), .B(new_n7310_), .Y(new_n7752_));
  AOI21X1  g07560(.A0(new_n7750_), .A1(\asqrt[30] ), .B0(new_n7752_), .Y(new_n7753_));
  INVX1    g07561(.A(new_n7753_), .Y(new_n7754_));
  OR2X1    g07562(.A(new_n7735_), .B(new_n2769_), .Y(new_n7755_));
  AND2X1   g07563(.A(new_n7719_), .B(new_n7710_), .Y(new_n7756_));
  INVX1    g07564(.A(new_n7725_), .Y(new_n7757_));
  NAND2X1  g07565(.A(new_n7701_), .B(new_n2769_), .Y(new_n7758_));
  OAI21X1  g07566(.A0(new_n7758_), .A1(new_n7756_), .B0(new_n7757_), .Y(new_n7759_));
  AOI21X1  g07567(.A0(new_n7759_), .A1(new_n7755_), .B0(new_n2570_), .Y(new_n7760_));
  AOI21X1  g07568(.A0(new_n7708_), .A1(\asqrt[44] ), .B0(\asqrt[45] ), .Y(new_n7761_));
  AOI21X1  g07569(.A0(new_n7761_), .A1(new_n7759_), .B0(new_n7732_), .Y(new_n7762_));
  OAI21X1  g07570(.A0(new_n7762_), .A1(new_n7760_), .B0(\asqrt[46] ), .Y(new_n7763_));
  NAND2X1  g07571(.A(new_n7763_), .B(new_n2040_), .Y(new_n7764_));
  OAI21X1  g07572(.A0(new_n7764_), .A1(new_n7748_), .B0(new_n7754_), .Y(new_n7765_));
  AOI21X1  g07573(.A0(new_n7765_), .A1(new_n7747_), .B0(new_n1834_), .Y(new_n7766_));
  NAND4X1  g07574(.A(\asqrt[30] ), .B(new_n7322_), .C(new_n7320_), .D(new_n7347_), .Y(new_n7767_));
  NAND2X1  g07575(.A(new_n7322_), .B(new_n7347_), .Y(new_n7768_));
  OAI21X1  g07576(.A0(new_n7768_), .A1(new_n7527_), .B0(new_n7321_), .Y(new_n7769_));
  AND2X1   g07577(.A(new_n7769_), .B(new_n7767_), .Y(new_n7770_));
  NOR3X1   g07578(.A(new_n7762_), .B(new_n7760_), .C(\asqrt[46] ), .Y(new_n7771_));
  OAI21X1  g07579(.A0(new_n7771_), .A1(new_n7743_), .B0(new_n7763_), .Y(new_n7772_));
  AOI21X1  g07580(.A0(new_n7772_), .A1(\asqrt[47] ), .B0(\asqrt[48] ), .Y(new_n7773_));
  AOI21X1  g07581(.A0(new_n7773_), .A1(new_n7765_), .B0(new_n7770_), .Y(new_n7774_));
  OAI21X1  g07582(.A0(new_n7774_), .A1(new_n7766_), .B0(\asqrt[49] ), .Y(new_n7775_));
  AND2X1   g07583(.A(new_n7364_), .B(new_n7363_), .Y(new_n7776_));
  NOR3X1   g07584(.A(new_n7776_), .B(new_n7330_), .C(new_n7362_), .Y(new_n7777_));
  NOR3X1   g07585(.A(new_n7527_), .B(new_n7776_), .C(new_n7362_), .Y(new_n7778_));
  NOR2X1   g07586(.A(new_n7778_), .B(new_n7329_), .Y(new_n7779_));
  AOI21X1  g07587(.A0(new_n7777_), .A1(\asqrt[30] ), .B0(new_n7779_), .Y(new_n7780_));
  NOR3X1   g07588(.A(new_n7774_), .B(new_n7766_), .C(\asqrt[49] ), .Y(new_n7781_));
  OAI21X1  g07589(.A0(new_n7781_), .A1(new_n7780_), .B0(new_n7775_), .Y(new_n7782_));
  AND2X1   g07590(.A(new_n7782_), .B(\asqrt[50] ), .Y(new_n7783_));
  INVX1    g07591(.A(new_n7780_), .Y(new_n7784_));
  AND2X1   g07592(.A(new_n7772_), .B(\asqrt[47] ), .Y(new_n7785_));
  NAND2X1  g07593(.A(new_n7745_), .B(new_n7744_), .Y(new_n7786_));
  AND2X1   g07594(.A(new_n7763_), .B(new_n2040_), .Y(new_n7787_));
  AOI21X1  g07595(.A0(new_n7787_), .A1(new_n7786_), .B0(new_n7753_), .Y(new_n7788_));
  OAI21X1  g07596(.A0(new_n7788_), .A1(new_n7785_), .B0(\asqrt[48] ), .Y(new_n7789_));
  INVX1    g07597(.A(new_n7770_), .Y(new_n7790_));
  OAI21X1  g07598(.A0(new_n7746_), .A1(new_n2040_), .B0(new_n1834_), .Y(new_n7791_));
  OAI21X1  g07599(.A0(new_n7791_), .A1(new_n7788_), .B0(new_n7790_), .Y(new_n7792_));
  NAND3X1  g07600(.A(new_n7792_), .B(new_n7789_), .C(new_n1632_), .Y(new_n7793_));
  NAND2X1  g07601(.A(new_n7793_), .B(new_n7784_), .Y(new_n7794_));
  AND2X1   g07602(.A(new_n7350_), .B(new_n7332_), .Y(new_n7795_));
  NOR3X1   g07603(.A(new_n7795_), .B(new_n7367_), .C(new_n7333_), .Y(new_n7796_));
  NOR3X1   g07604(.A(new_n7527_), .B(new_n7795_), .C(new_n7333_), .Y(new_n7797_));
  NOR2X1   g07605(.A(new_n7797_), .B(new_n7338_), .Y(new_n7798_));
  AOI21X1  g07606(.A0(new_n7796_), .A1(\asqrt[30] ), .B0(new_n7798_), .Y(new_n7799_));
  AND2X1   g07607(.A(new_n7775_), .B(new_n1469_), .Y(new_n7800_));
  AOI21X1  g07608(.A0(new_n7800_), .A1(new_n7794_), .B0(new_n7799_), .Y(new_n7801_));
  OAI21X1  g07609(.A0(new_n7801_), .A1(new_n7783_), .B0(\asqrt[51] ), .Y(new_n7802_));
  NAND4X1  g07610(.A(\asqrt[30] ), .B(new_n7370_), .C(new_n7357_), .D(new_n7352_), .Y(new_n7803_));
  NAND2X1  g07611(.A(new_n7370_), .B(new_n7352_), .Y(new_n7804_));
  OAI21X1  g07612(.A0(new_n7804_), .A1(new_n7527_), .B0(new_n7361_), .Y(new_n7805_));
  AND2X1   g07613(.A(new_n7805_), .B(new_n7803_), .Y(new_n7806_));
  INVX1    g07614(.A(new_n7806_), .Y(new_n7807_));
  AOI21X1  g07615(.A0(new_n7792_), .A1(new_n7789_), .B0(new_n1632_), .Y(new_n7808_));
  AOI21X1  g07616(.A0(new_n7793_), .A1(new_n7784_), .B0(new_n7808_), .Y(new_n7809_));
  OAI21X1  g07617(.A0(new_n7809_), .A1(new_n1469_), .B0(new_n1277_), .Y(new_n7810_));
  OAI21X1  g07618(.A0(new_n7810_), .A1(new_n7801_), .B0(new_n7807_), .Y(new_n7811_));
  AOI21X1  g07619(.A0(new_n7811_), .A1(new_n7802_), .B0(new_n1111_), .Y(new_n7812_));
  AOI21X1  g07620(.A0(new_n7377_), .A1(new_n7371_), .B0(new_n7401_), .Y(new_n7813_));
  AND2X1   g07621(.A(new_n7813_), .B(new_n7399_), .Y(new_n7814_));
  AOI22X1  g07622(.A0(new_n7377_), .A1(new_n7371_), .B0(new_n7359_), .B1(\asqrt[51] ), .Y(new_n7815_));
  AOI21X1  g07623(.A0(new_n7815_), .A1(\asqrt[30] ), .B0(new_n7375_), .Y(new_n7816_));
  AOI21X1  g07624(.A0(new_n7814_), .A1(\asqrt[30] ), .B0(new_n7816_), .Y(new_n7817_));
  INVX1    g07625(.A(new_n7817_), .Y(new_n7818_));
  NAND3X1  g07626(.A(new_n7811_), .B(new_n7802_), .C(new_n1111_), .Y(new_n7819_));
  AOI21X1  g07627(.A0(new_n7819_), .A1(new_n7818_), .B0(new_n7812_), .Y(new_n7820_));
  OR2X1    g07628(.A(new_n7820_), .B(new_n968_), .Y(new_n7821_));
  AND2X1   g07629(.A(new_n7819_), .B(new_n7818_), .Y(new_n7822_));
  AND2X1   g07630(.A(new_n7405_), .B(new_n7403_), .Y(new_n7823_));
  NOR3X1   g07631(.A(new_n7823_), .B(new_n7385_), .C(new_n7404_), .Y(new_n7824_));
  NOR3X1   g07632(.A(new_n7527_), .B(new_n7823_), .C(new_n7404_), .Y(new_n7825_));
  NOR2X1   g07633(.A(new_n7825_), .B(new_n7384_), .Y(new_n7826_));
  AOI21X1  g07634(.A0(new_n7824_), .A1(\asqrt[30] ), .B0(new_n7826_), .Y(new_n7827_));
  INVX1    g07635(.A(new_n7827_), .Y(new_n7828_));
  OR2X1    g07636(.A(new_n7809_), .B(new_n1469_), .Y(new_n7829_));
  AND2X1   g07637(.A(new_n7793_), .B(new_n7784_), .Y(new_n7830_));
  INVX1    g07638(.A(new_n7799_), .Y(new_n7831_));
  NAND2X1  g07639(.A(new_n7775_), .B(new_n1469_), .Y(new_n7832_));
  OAI21X1  g07640(.A0(new_n7832_), .A1(new_n7830_), .B0(new_n7831_), .Y(new_n7833_));
  AOI21X1  g07641(.A0(new_n7833_), .A1(new_n7829_), .B0(new_n1277_), .Y(new_n7834_));
  AOI21X1  g07642(.A0(new_n7782_), .A1(\asqrt[50] ), .B0(\asqrt[51] ), .Y(new_n7835_));
  AOI21X1  g07643(.A0(new_n7835_), .A1(new_n7833_), .B0(new_n7806_), .Y(new_n7836_));
  OAI21X1  g07644(.A0(new_n7836_), .A1(new_n7834_), .B0(\asqrt[52] ), .Y(new_n7837_));
  NAND2X1  g07645(.A(new_n7837_), .B(new_n968_), .Y(new_n7838_));
  OAI21X1  g07646(.A0(new_n7838_), .A1(new_n7822_), .B0(new_n7828_), .Y(new_n7839_));
  AOI21X1  g07647(.A0(new_n7839_), .A1(new_n7821_), .B0(new_n902_), .Y(new_n7840_));
  NAND4X1  g07648(.A(\asqrt[30] ), .B(new_n7396_), .C(new_n7394_), .D(new_n7414_), .Y(new_n7841_));
  OR2X1    g07649(.A(new_n7407_), .B(new_n7389_), .Y(new_n7842_));
  OAI21X1  g07650(.A0(new_n7842_), .A1(new_n7527_), .B0(new_n7395_), .Y(new_n7843_));
  AND2X1   g07651(.A(new_n7843_), .B(new_n7841_), .Y(new_n7844_));
  NOR3X1   g07652(.A(new_n7836_), .B(new_n7834_), .C(\asqrt[52] ), .Y(new_n7845_));
  OAI21X1  g07653(.A0(new_n7845_), .A1(new_n7817_), .B0(new_n7837_), .Y(new_n7846_));
  AOI21X1  g07654(.A0(new_n7846_), .A1(\asqrt[53] ), .B0(\asqrt[54] ), .Y(new_n7847_));
  AOI21X1  g07655(.A0(new_n7847_), .A1(new_n7839_), .B0(new_n7844_), .Y(new_n7848_));
  OAI21X1  g07656(.A0(new_n7848_), .A1(new_n7840_), .B0(\asqrt[55] ), .Y(new_n7849_));
  AND2X1   g07657(.A(new_n7451_), .B(new_n7450_), .Y(new_n7850_));
  NOR3X1   g07658(.A(new_n7850_), .B(new_n7413_), .C(new_n7449_), .Y(new_n7851_));
  NOR3X1   g07659(.A(new_n7527_), .B(new_n7850_), .C(new_n7449_), .Y(new_n7852_));
  NOR2X1   g07660(.A(new_n7852_), .B(new_n7412_), .Y(new_n7853_));
  AOI21X1  g07661(.A0(new_n7851_), .A1(\asqrt[30] ), .B0(new_n7853_), .Y(new_n7854_));
  NOR3X1   g07662(.A(new_n7848_), .B(new_n7840_), .C(\asqrt[55] ), .Y(new_n7855_));
  OAI21X1  g07663(.A0(new_n7855_), .A1(new_n7854_), .B0(new_n7849_), .Y(new_n7856_));
  AND2X1   g07664(.A(new_n7856_), .B(\asqrt[56] ), .Y(new_n7857_));
  INVX1    g07665(.A(new_n7854_), .Y(new_n7858_));
  AND2X1   g07666(.A(new_n7846_), .B(\asqrt[53] ), .Y(new_n7859_));
  NAND2X1  g07667(.A(new_n7819_), .B(new_n7818_), .Y(new_n7860_));
  AND2X1   g07668(.A(new_n7837_), .B(new_n968_), .Y(new_n7861_));
  AOI21X1  g07669(.A0(new_n7861_), .A1(new_n7860_), .B0(new_n7827_), .Y(new_n7862_));
  OAI21X1  g07670(.A0(new_n7862_), .A1(new_n7859_), .B0(\asqrt[54] ), .Y(new_n7863_));
  INVX1    g07671(.A(new_n7844_), .Y(new_n7864_));
  OAI21X1  g07672(.A0(new_n7820_), .A1(new_n968_), .B0(new_n902_), .Y(new_n7865_));
  OAI21X1  g07673(.A0(new_n7865_), .A1(new_n7862_), .B0(new_n7864_), .Y(new_n7866_));
  NAND3X1  g07674(.A(new_n7866_), .B(new_n7863_), .C(new_n697_), .Y(new_n7867_));
  NAND2X1  g07675(.A(new_n7867_), .B(new_n7858_), .Y(new_n7868_));
  AND2X1   g07676(.A(new_n7424_), .B(new_n7416_), .Y(new_n7869_));
  NOR3X1   g07677(.A(new_n7869_), .B(new_n7454_), .C(new_n7417_), .Y(new_n7870_));
  NOR3X1   g07678(.A(new_n7527_), .B(new_n7869_), .C(new_n7417_), .Y(new_n7871_));
  NOR2X1   g07679(.A(new_n7871_), .B(new_n7422_), .Y(new_n7872_));
  AOI21X1  g07680(.A0(new_n7870_), .A1(\asqrt[30] ), .B0(new_n7872_), .Y(new_n7873_));
  AND2X1   g07681(.A(new_n7849_), .B(new_n582_), .Y(new_n7874_));
  AOI21X1  g07682(.A0(new_n7874_), .A1(new_n7868_), .B0(new_n7873_), .Y(new_n7875_));
  OAI21X1  g07683(.A0(new_n7875_), .A1(new_n7857_), .B0(\asqrt[57] ), .Y(new_n7876_));
  OR4X1    g07684(.A(new_n7527_), .B(new_n7432_), .C(new_n7458_), .D(new_n7457_), .Y(new_n7877_));
  OR2X1    g07685(.A(new_n7432_), .B(new_n7457_), .Y(new_n7878_));
  OAI21X1  g07686(.A0(new_n7878_), .A1(new_n7527_), .B0(new_n7458_), .Y(new_n7879_));
  AND2X1   g07687(.A(new_n7879_), .B(new_n7877_), .Y(new_n7880_));
  INVX1    g07688(.A(new_n7880_), .Y(new_n7881_));
  AOI21X1  g07689(.A0(new_n7866_), .A1(new_n7863_), .B0(new_n697_), .Y(new_n7882_));
  AOI21X1  g07690(.A0(new_n7867_), .A1(new_n7858_), .B0(new_n7882_), .Y(new_n7883_));
  OAI21X1  g07691(.A0(new_n7883_), .A1(new_n582_), .B0(new_n481_), .Y(new_n7884_));
  OAI21X1  g07692(.A0(new_n7884_), .A1(new_n7875_), .B0(new_n7881_), .Y(new_n7885_));
  AOI21X1  g07693(.A0(new_n7885_), .A1(new_n7876_), .B0(new_n399_), .Y(new_n7886_));
  AOI21X1  g07694(.A0(new_n7440_), .A1(new_n7435_), .B0(new_n7475_), .Y(new_n7887_));
  AND2X1   g07695(.A(new_n7887_), .B(new_n7473_), .Y(new_n7888_));
  AOI22X1  g07696(.A0(new_n7440_), .A1(new_n7435_), .B0(new_n7433_), .B1(\asqrt[57] ), .Y(new_n7889_));
  AOI21X1  g07697(.A0(new_n7889_), .A1(\asqrt[30] ), .B0(new_n7439_), .Y(new_n7890_));
  AOI21X1  g07698(.A0(new_n7888_), .A1(\asqrt[30] ), .B0(new_n7890_), .Y(new_n7891_));
  INVX1    g07699(.A(new_n7891_), .Y(new_n7892_));
  NAND3X1  g07700(.A(new_n7885_), .B(new_n7876_), .C(new_n399_), .Y(new_n7893_));
  AOI21X1  g07701(.A0(new_n7893_), .A1(new_n7892_), .B0(new_n7886_), .Y(new_n7894_));
  OR2X1    g07702(.A(new_n7894_), .B(new_n328_), .Y(new_n7895_));
  AND2X1   g07703(.A(new_n7893_), .B(new_n7892_), .Y(new_n7896_));
  AND2X1   g07704(.A(new_n7479_), .B(new_n7477_), .Y(new_n7897_));
  NOR3X1   g07705(.A(new_n7897_), .B(new_n7448_), .C(new_n7478_), .Y(new_n7898_));
  NOR3X1   g07706(.A(new_n7527_), .B(new_n7897_), .C(new_n7478_), .Y(new_n7899_));
  NOR2X1   g07707(.A(new_n7899_), .B(new_n7447_), .Y(new_n7900_));
  AOI21X1  g07708(.A0(new_n7898_), .A1(\asqrt[30] ), .B0(new_n7900_), .Y(new_n7901_));
  INVX1    g07709(.A(new_n7901_), .Y(new_n7902_));
  OR2X1    g07710(.A(new_n7883_), .B(new_n582_), .Y(new_n7903_));
  AND2X1   g07711(.A(new_n7867_), .B(new_n7858_), .Y(new_n7904_));
  INVX1    g07712(.A(new_n7873_), .Y(new_n7905_));
  NAND2X1  g07713(.A(new_n7849_), .B(new_n582_), .Y(new_n7906_));
  OAI21X1  g07714(.A0(new_n7906_), .A1(new_n7904_), .B0(new_n7905_), .Y(new_n7907_));
  AOI21X1  g07715(.A0(new_n7907_), .A1(new_n7903_), .B0(new_n481_), .Y(new_n7908_));
  AOI21X1  g07716(.A0(new_n7856_), .A1(\asqrt[56] ), .B0(\asqrt[57] ), .Y(new_n7909_));
  AOI21X1  g07717(.A0(new_n7909_), .A1(new_n7907_), .B0(new_n7880_), .Y(new_n7910_));
  OAI21X1  g07718(.A0(new_n7910_), .A1(new_n7908_), .B0(\asqrt[58] ), .Y(new_n7911_));
  NAND2X1  g07719(.A(new_n7911_), .B(new_n328_), .Y(new_n7912_));
  OAI21X1  g07720(.A0(new_n7912_), .A1(new_n7896_), .B0(new_n7902_), .Y(new_n7913_));
  AOI21X1  g07721(.A0(new_n7913_), .A1(new_n7895_), .B0(new_n292_), .Y(new_n7914_));
  OR4X1    g07722(.A(new_n7527_), .B(new_n7481_), .C(new_n7469_), .D(new_n7463_), .Y(new_n7915_));
  OR2X1    g07723(.A(new_n7481_), .B(new_n7463_), .Y(new_n7916_));
  OAI21X1  g07724(.A0(new_n7916_), .A1(new_n7527_), .B0(new_n7469_), .Y(new_n7917_));
  AND2X1   g07725(.A(new_n7917_), .B(new_n7915_), .Y(new_n7918_));
  NOR3X1   g07726(.A(new_n7910_), .B(new_n7908_), .C(\asqrt[58] ), .Y(new_n7919_));
  OAI21X1  g07727(.A0(new_n7919_), .A1(new_n7891_), .B0(new_n7911_), .Y(new_n7920_));
  AOI21X1  g07728(.A0(new_n7920_), .A1(\asqrt[59] ), .B0(\asqrt[60] ), .Y(new_n7921_));
  AOI21X1  g07729(.A0(new_n7921_), .A1(new_n7913_), .B0(new_n7918_), .Y(new_n7922_));
  OAI21X1  g07730(.A0(new_n7922_), .A1(new_n7914_), .B0(\asqrt[61] ), .Y(new_n7923_));
  AND2X1   g07731(.A(new_n7531_), .B(new_n7530_), .Y(new_n7924_));
  NOR3X1   g07732(.A(new_n7924_), .B(new_n7487_), .C(new_n7529_), .Y(new_n7925_));
  NOR3X1   g07733(.A(new_n7527_), .B(new_n7924_), .C(new_n7529_), .Y(new_n7926_));
  NOR2X1   g07734(.A(new_n7926_), .B(new_n7486_), .Y(new_n7927_));
  AOI21X1  g07735(.A0(new_n7925_), .A1(\asqrt[30] ), .B0(new_n7927_), .Y(new_n7928_));
  NOR3X1   g07736(.A(new_n7922_), .B(new_n7914_), .C(\asqrt[61] ), .Y(new_n7929_));
  OAI21X1  g07737(.A0(new_n7929_), .A1(new_n7928_), .B0(new_n7923_), .Y(new_n7930_));
  AND2X1   g07738(.A(new_n7930_), .B(\asqrt[62] ), .Y(new_n7931_));
  INVX1    g07739(.A(new_n7928_), .Y(new_n7932_));
  AND2X1   g07740(.A(new_n7920_), .B(\asqrt[59] ), .Y(new_n7933_));
  NAND2X1  g07741(.A(new_n7893_), .B(new_n7892_), .Y(new_n7934_));
  AND2X1   g07742(.A(new_n7911_), .B(new_n328_), .Y(new_n7935_));
  AOI21X1  g07743(.A0(new_n7935_), .A1(new_n7934_), .B0(new_n7901_), .Y(new_n7936_));
  OAI21X1  g07744(.A0(new_n7936_), .A1(new_n7933_), .B0(\asqrt[60] ), .Y(new_n7937_));
  INVX1    g07745(.A(new_n7918_), .Y(new_n7938_));
  OAI21X1  g07746(.A0(new_n7894_), .A1(new_n328_), .B0(new_n292_), .Y(new_n7939_));
  OAI21X1  g07747(.A0(new_n7939_), .A1(new_n7936_), .B0(new_n7938_), .Y(new_n7940_));
  NAND3X1  g07748(.A(new_n7940_), .B(new_n7937_), .C(new_n217_), .Y(new_n7941_));
  NAND2X1  g07749(.A(new_n7941_), .B(new_n7932_), .Y(new_n7942_));
  AND2X1   g07750(.A(new_n7498_), .B(new_n7490_), .Y(new_n7943_));
  NOR3X1   g07751(.A(new_n7943_), .B(new_n7534_), .C(new_n7491_), .Y(new_n7944_));
  NOR3X1   g07752(.A(new_n7527_), .B(new_n7943_), .C(new_n7491_), .Y(new_n7945_));
  NOR2X1   g07753(.A(new_n7945_), .B(new_n7496_), .Y(new_n7946_));
  AOI21X1  g07754(.A0(new_n7944_), .A1(\asqrt[30] ), .B0(new_n7946_), .Y(new_n7947_));
  AOI21X1  g07755(.A0(new_n7940_), .A1(new_n7937_), .B0(new_n217_), .Y(new_n7948_));
  NOR2X1   g07756(.A(new_n7948_), .B(\asqrt[62] ), .Y(new_n7949_));
  AOI21X1  g07757(.A0(new_n7949_), .A1(new_n7942_), .B0(new_n7947_), .Y(new_n7950_));
  NOR4X1   g07758(.A(new_n7527_), .B(new_n7506_), .C(new_n7538_), .D(new_n7537_), .Y(new_n7951_));
  NAND3X1  g07759(.A(\asqrt[30] ), .B(new_n7539_), .C(new_n7500_), .Y(new_n7952_));
  AOI21X1  g07760(.A0(new_n7952_), .A1(new_n7538_), .B0(new_n7951_), .Y(new_n7953_));
  INVX1    g07761(.A(new_n7953_), .Y(new_n7954_));
  NOR3X1   g07762(.A(new_n7527_), .B(new_n7510_), .C(new_n7540_), .Y(new_n7955_));
  AOI21X1  g07763(.A0(new_n7544_), .A1(new_n7543_), .B0(new_n7955_), .Y(new_n7956_));
  AND2X1   g07764(.A(new_n7956_), .B(new_n7954_), .Y(new_n7957_));
  OAI21X1  g07765(.A0(new_n7950_), .A1(new_n7931_), .B0(new_n7957_), .Y(new_n7958_));
  AOI21X1  g07766(.A0(new_n7941_), .A1(new_n7932_), .B0(new_n7948_), .Y(new_n7959_));
  OAI21X1  g07767(.A0(new_n7959_), .A1(new_n199_), .B0(new_n7953_), .Y(new_n7960_));
  AOI21X1  g07768(.A0(new_n7546_), .A1(new_n7542_), .B0(new_n7510_), .Y(new_n7961_));
  AOI21X1  g07769(.A0(new_n7511_), .A1(new_n7507_), .B0(new_n193_), .Y(new_n7962_));
  OAI21X1  g07770(.A0(new_n7961_), .A1(new_n7507_), .B0(new_n7962_), .Y(new_n7963_));
  OR2X1    g07771(.A(new_n7517_), .B(new_n7516_), .Y(new_n7964_));
  AND2X1   g07772(.A(new_n7509_), .B(new_n7119_), .Y(new_n7965_));
  NOR4X1   g07773(.A(new_n7523_), .B(new_n7562_), .C(new_n7965_), .D(new_n7508_), .Y(new_n7966_));
  NAND3X1  g07774(.A(new_n7966_), .B(new_n7964_), .C(new_n7542_), .Y(new_n7967_));
  AND2X1   g07775(.A(new_n7967_), .B(new_n7963_), .Y(new_n7968_));
  OAI21X1  g07776(.A0(new_n7960_), .A1(new_n7950_), .B0(new_n7968_), .Y(new_n7969_));
  AOI21X1  g07777(.A0(new_n7958_), .A1(new_n193_), .B0(new_n7969_), .Y(new_n7970_));
  NOR2X1   g07778(.A(\a[57] ), .B(\a[56] ), .Y(new_n7971_));
  INVX1    g07779(.A(new_n7971_), .Y(new_n7972_));
  MX2X1    g07780(.A(new_n7972_), .B(new_n7970_), .S0(\a[58] ), .Y(new_n7973_));
  OR2X1    g07781(.A(new_n7973_), .B(new_n7527_), .Y(new_n7974_));
  INVX1    g07782(.A(\a[58] ), .Y(new_n7975_));
  NOR3X1   g07783(.A(\a[58] ), .B(\a[57] ), .C(\a[56] ), .Y(new_n7976_));
  NOR3X1   g07784(.A(new_n7976_), .B(new_n7523_), .C(new_n7562_), .Y(new_n7977_));
  NAND3X1  g07785(.A(new_n7977_), .B(new_n7964_), .C(new_n7542_), .Y(new_n7978_));
  INVX1    g07786(.A(new_n7978_), .Y(new_n7979_));
  OAI21X1  g07787(.A0(new_n7970_), .A1(new_n7975_), .B0(new_n7979_), .Y(new_n7980_));
  OAI21X1  g07788(.A0(new_n7970_), .A1(\a[58] ), .B0(\a[59] ), .Y(new_n7981_));
  NOR2X1   g07789(.A(\a[59] ), .B(\a[58] ), .Y(new_n7982_));
  INVX1    g07790(.A(new_n7982_), .Y(new_n7983_));
  OR2X1    g07791(.A(new_n7970_), .B(new_n7983_), .Y(new_n7984_));
  NAND3X1  g07792(.A(new_n7984_), .B(new_n7981_), .C(new_n7980_), .Y(new_n7985_));
  AOI21X1  g07793(.A0(new_n7985_), .A1(new_n7974_), .B0(new_n7103_), .Y(new_n7986_));
  OR2X1    g07794(.A(new_n7959_), .B(new_n199_), .Y(new_n7987_));
  AND2X1   g07795(.A(new_n7941_), .B(new_n7932_), .Y(new_n7988_));
  INVX1    g07796(.A(new_n7947_), .Y(new_n7989_));
  OR2X1    g07797(.A(new_n7948_), .B(\asqrt[62] ), .Y(new_n7990_));
  OAI21X1  g07798(.A0(new_n7990_), .A1(new_n7988_), .B0(new_n7989_), .Y(new_n7991_));
  INVX1    g07799(.A(new_n7957_), .Y(new_n7992_));
  AOI21X1  g07800(.A0(new_n7991_), .A1(new_n7987_), .B0(new_n7992_), .Y(new_n7993_));
  AOI21X1  g07801(.A0(new_n7930_), .A1(\asqrt[62] ), .B0(new_n7954_), .Y(new_n7994_));
  INVX1    g07802(.A(new_n7968_), .Y(new_n7995_));
  AOI21X1  g07803(.A0(new_n7994_), .A1(new_n7991_), .B0(new_n7995_), .Y(new_n7996_));
  OAI21X1  g07804(.A0(new_n7993_), .A1(\asqrt[63] ), .B0(new_n7996_), .Y(\asqrt[29] ));
  MX2X1    g07805(.A(new_n7971_), .B(\asqrt[29] ), .S0(\a[58] ), .Y(new_n7998_));
  AOI21X1  g07806(.A0(new_n7998_), .A1(\asqrt[30] ), .B0(\asqrt[31] ), .Y(new_n7999_));
  NAND3X1  g07807(.A(new_n7967_), .B(new_n7963_), .C(\asqrt[30] ), .Y(new_n8000_));
  INVX1    g07808(.A(new_n8000_), .Y(new_n8001_));
  OAI21X1  g07809(.A0(new_n7960_), .A1(new_n7950_), .B0(new_n8001_), .Y(new_n8002_));
  AOI21X1  g07810(.A0(new_n7958_), .A1(new_n193_), .B0(new_n8002_), .Y(new_n8003_));
  AOI21X1  g07811(.A0(\asqrt[29] ), .A1(new_n7982_), .B0(new_n8003_), .Y(new_n8004_));
  OR2X1    g07812(.A(new_n8004_), .B(new_n7528_), .Y(new_n8005_));
  AND2X1   g07813(.A(\asqrt[29] ), .B(new_n7982_), .Y(new_n8006_));
  OR2X1    g07814(.A(new_n8003_), .B(\a[60] ), .Y(new_n8007_));
  OR2X1    g07815(.A(new_n8007_), .B(new_n8006_), .Y(new_n8008_));
  AOI22X1  g07816(.A0(new_n8008_), .A1(new_n8005_), .B0(new_n7999_), .B1(new_n7985_), .Y(new_n8009_));
  OAI21X1  g07817(.A0(new_n8009_), .A1(new_n7986_), .B0(\asqrt[32] ), .Y(new_n8010_));
  AND2X1   g07818(.A(new_n7581_), .B(new_n7549_), .Y(new_n8011_));
  NAND3X1  g07819(.A(new_n8011_), .B(\asqrt[29] ), .C(new_n7557_), .Y(new_n8012_));
  INVX1    g07820(.A(new_n8011_), .Y(new_n8013_));
  OAI21X1  g07821(.A0(new_n8013_), .A1(new_n7970_), .B0(new_n7583_), .Y(new_n8014_));
  AND2X1   g07822(.A(new_n8014_), .B(new_n8012_), .Y(new_n8015_));
  NOR3X1   g07823(.A(new_n8009_), .B(new_n7986_), .C(\asqrt[32] ), .Y(new_n8016_));
  OAI21X1  g07824(.A0(new_n8016_), .A1(new_n8015_), .B0(new_n8010_), .Y(new_n8017_));
  AND2X1   g07825(.A(new_n8017_), .B(\asqrt[33] ), .Y(new_n8018_));
  INVX1    g07826(.A(new_n8015_), .Y(new_n8019_));
  AND2X1   g07827(.A(new_n7998_), .B(\asqrt[30] ), .Y(new_n8020_));
  AOI21X1  g07828(.A0(\asqrt[29] ), .A1(\a[58] ), .B0(new_n7978_), .Y(new_n8021_));
  INVX1    g07829(.A(\a[59] ), .Y(new_n8022_));
  AOI21X1  g07830(.A0(\asqrt[29] ), .A1(new_n7975_), .B0(new_n8022_), .Y(new_n8023_));
  NOR3X1   g07831(.A(new_n8006_), .B(new_n8023_), .C(new_n8021_), .Y(new_n8024_));
  OAI21X1  g07832(.A0(new_n8024_), .A1(new_n8020_), .B0(\asqrt[31] ), .Y(new_n8025_));
  OAI21X1  g07833(.A0(new_n7973_), .A1(new_n7527_), .B0(new_n7103_), .Y(new_n8026_));
  OAI22X1  g07834(.A0(new_n8007_), .A1(new_n8006_), .B0(new_n8004_), .B1(new_n7528_), .Y(new_n8027_));
  OAI21X1  g07835(.A0(new_n8026_), .A1(new_n8024_), .B0(new_n8027_), .Y(new_n8028_));
  NAND3X1  g07836(.A(new_n8028_), .B(new_n8025_), .C(new_n6699_), .Y(new_n8029_));
  NAND2X1  g07837(.A(new_n8029_), .B(new_n8019_), .Y(new_n8030_));
  AOI21X1  g07838(.A0(new_n7561_), .A1(new_n7560_), .B0(new_n7602_), .Y(new_n8031_));
  NAND3X1  g07839(.A(new_n8031_), .B(\asqrt[29] ), .C(new_n7599_), .Y(new_n8032_));
  OAI22X1  g07840(.A0(new_n7601_), .A1(new_n7600_), .B0(new_n7584_), .B1(new_n6699_), .Y(new_n8033_));
  OAI21X1  g07841(.A0(new_n8033_), .A1(new_n7970_), .B0(new_n7602_), .Y(new_n8034_));
  AND2X1   g07842(.A(new_n8034_), .B(new_n8032_), .Y(new_n8035_));
  AOI21X1  g07843(.A0(new_n8028_), .A1(new_n8025_), .B0(new_n6699_), .Y(new_n8036_));
  NOR2X1   g07844(.A(new_n8036_), .B(\asqrt[33] ), .Y(new_n8037_));
  AOI21X1  g07845(.A0(new_n8037_), .A1(new_n8030_), .B0(new_n8035_), .Y(new_n8038_));
  OAI21X1  g07846(.A0(new_n8038_), .A1(new_n8018_), .B0(\asqrt[34] ), .Y(new_n8039_));
  AND2X1   g07847(.A(new_n7606_), .B(new_n7603_), .Y(new_n8040_));
  OR4X1    g07848(.A(new_n7970_), .B(new_n8040_), .C(new_n7579_), .D(new_n7604_), .Y(new_n8041_));
  OR2X1    g07849(.A(new_n8040_), .B(new_n7604_), .Y(new_n8042_));
  OAI21X1  g07850(.A0(new_n8042_), .A1(new_n7970_), .B0(new_n7579_), .Y(new_n8043_));
  AND2X1   g07851(.A(new_n8043_), .B(new_n8041_), .Y(new_n8044_));
  INVX1    g07852(.A(new_n8044_), .Y(new_n8045_));
  AOI21X1  g07853(.A0(new_n8029_), .A1(new_n8019_), .B0(new_n8036_), .Y(new_n8046_));
  OAI21X1  g07854(.A0(new_n8046_), .A1(new_n6294_), .B0(new_n5941_), .Y(new_n8047_));
  OAI21X1  g07855(.A0(new_n8047_), .A1(new_n8038_), .B0(new_n8045_), .Y(new_n8048_));
  AOI21X1  g07856(.A0(new_n8048_), .A1(new_n8039_), .B0(new_n5541_), .Y(new_n8049_));
  OR4X1    g07857(.A(new_n7970_), .B(new_n7608_), .C(new_n7595_), .D(new_n7587_), .Y(new_n8050_));
  NAND2X1  g07858(.A(new_n7596_), .B(new_n7610_), .Y(new_n8051_));
  OAI21X1  g07859(.A0(new_n8051_), .A1(new_n7970_), .B0(new_n7595_), .Y(new_n8052_));
  AND2X1   g07860(.A(new_n8052_), .B(new_n8050_), .Y(new_n8053_));
  INVX1    g07861(.A(new_n8053_), .Y(new_n8054_));
  NAND3X1  g07862(.A(new_n8048_), .B(new_n8039_), .C(new_n5541_), .Y(new_n8055_));
  AOI21X1  g07863(.A0(new_n8055_), .A1(new_n8054_), .B0(new_n8049_), .Y(new_n8056_));
  OR2X1    g07864(.A(new_n8056_), .B(new_n5176_), .Y(new_n8057_));
  AND2X1   g07865(.A(new_n8055_), .B(new_n8054_), .Y(new_n8058_));
  OR2X1    g07866(.A(new_n8049_), .B(\asqrt[36] ), .Y(new_n8059_));
  AND2X1   g07867(.A(new_n7640_), .B(new_n7639_), .Y(new_n8060_));
  NOR4X1   g07868(.A(new_n7970_), .B(new_n7618_), .C(new_n8060_), .D(new_n7638_), .Y(new_n8061_));
  AOI22X1  g07869(.A0(new_n7640_), .A1(new_n7639_), .B0(new_n7625_), .B1(\asqrt[35] ), .Y(new_n8062_));
  AOI21X1  g07870(.A0(new_n8062_), .A1(\asqrt[29] ), .B0(new_n7617_), .Y(new_n8063_));
  NOR2X1   g07871(.A(new_n8063_), .B(new_n8061_), .Y(new_n8064_));
  INVX1    g07872(.A(new_n8064_), .Y(new_n8065_));
  OAI21X1  g07873(.A0(new_n8059_), .A1(new_n8058_), .B0(new_n8065_), .Y(new_n8066_));
  AOI21X1  g07874(.A0(new_n8066_), .A1(new_n8057_), .B0(new_n4826_), .Y(new_n8067_));
  AND2X1   g07875(.A(new_n7626_), .B(new_n7619_), .Y(new_n8068_));
  OR4X1    g07876(.A(new_n7970_), .B(new_n8068_), .C(new_n7623_), .D(new_n7620_), .Y(new_n8069_));
  OR2X1    g07877(.A(new_n8068_), .B(new_n7620_), .Y(new_n8070_));
  OAI21X1  g07878(.A0(new_n8070_), .A1(new_n7970_), .B0(new_n7623_), .Y(new_n8071_));
  AND2X1   g07879(.A(new_n8071_), .B(new_n8069_), .Y(new_n8072_));
  OR2X1    g07880(.A(new_n8046_), .B(new_n6294_), .Y(new_n8073_));
  AND2X1   g07881(.A(new_n8029_), .B(new_n8019_), .Y(new_n8074_));
  INVX1    g07882(.A(new_n8035_), .Y(new_n8075_));
  OR2X1    g07883(.A(new_n8036_), .B(\asqrt[33] ), .Y(new_n8076_));
  OAI21X1  g07884(.A0(new_n8076_), .A1(new_n8074_), .B0(new_n8075_), .Y(new_n8077_));
  AOI21X1  g07885(.A0(new_n8077_), .A1(new_n8073_), .B0(new_n5941_), .Y(new_n8078_));
  AOI21X1  g07886(.A0(new_n8017_), .A1(\asqrt[33] ), .B0(\asqrt[34] ), .Y(new_n8079_));
  AOI21X1  g07887(.A0(new_n8079_), .A1(new_n8077_), .B0(new_n8044_), .Y(new_n8080_));
  OAI21X1  g07888(.A0(new_n8080_), .A1(new_n8078_), .B0(\asqrt[35] ), .Y(new_n8081_));
  NOR3X1   g07889(.A(new_n8080_), .B(new_n8078_), .C(\asqrt[35] ), .Y(new_n8082_));
  OAI21X1  g07890(.A0(new_n8082_), .A1(new_n8053_), .B0(new_n8081_), .Y(new_n8083_));
  AOI21X1  g07891(.A0(new_n8083_), .A1(\asqrt[36] ), .B0(\asqrt[37] ), .Y(new_n8084_));
  AOI21X1  g07892(.A0(new_n8084_), .A1(new_n8066_), .B0(new_n8072_), .Y(new_n8085_));
  OAI21X1  g07893(.A0(new_n8085_), .A1(new_n8067_), .B0(\asqrt[38] ), .Y(new_n8086_));
  OR4X1    g07894(.A(new_n7970_), .B(new_n7634_), .C(new_n7637_), .D(new_n7660_), .Y(new_n8087_));
  NAND2X1  g07895(.A(new_n7645_), .B(new_n7628_), .Y(new_n8088_));
  OAI21X1  g07896(.A0(new_n8088_), .A1(new_n7970_), .B0(new_n7637_), .Y(new_n8089_));
  AND2X1   g07897(.A(new_n8089_), .B(new_n8087_), .Y(new_n8090_));
  NOR3X1   g07898(.A(new_n8085_), .B(new_n8067_), .C(\asqrt[38] ), .Y(new_n8091_));
  OAI21X1  g07899(.A0(new_n8091_), .A1(new_n8090_), .B0(new_n8086_), .Y(new_n8092_));
  AND2X1   g07900(.A(new_n8092_), .B(\asqrt[39] ), .Y(new_n8093_));
  INVX1    g07901(.A(new_n8090_), .Y(new_n8094_));
  AND2X1   g07902(.A(new_n8083_), .B(\asqrt[36] ), .Y(new_n8095_));
  NAND2X1  g07903(.A(new_n8055_), .B(new_n8054_), .Y(new_n8096_));
  NOR2X1   g07904(.A(new_n8049_), .B(\asqrt[36] ), .Y(new_n8097_));
  AOI21X1  g07905(.A0(new_n8097_), .A1(new_n8096_), .B0(new_n8064_), .Y(new_n8098_));
  OAI21X1  g07906(.A0(new_n8098_), .A1(new_n8095_), .B0(\asqrt[37] ), .Y(new_n8099_));
  INVX1    g07907(.A(new_n8072_), .Y(new_n8100_));
  OAI21X1  g07908(.A0(new_n8056_), .A1(new_n5176_), .B0(new_n4826_), .Y(new_n8101_));
  OAI21X1  g07909(.A0(new_n8101_), .A1(new_n8098_), .B0(new_n8100_), .Y(new_n8102_));
  NAND3X1  g07910(.A(new_n8102_), .B(new_n8099_), .C(new_n4493_), .Y(new_n8103_));
  NAND2X1  g07911(.A(new_n8103_), .B(new_n8094_), .Y(new_n8104_));
  OAI21X1  g07912(.A0(new_n7684_), .A1(new_n7682_), .B0(new_n7651_), .Y(new_n8105_));
  NOR3X1   g07913(.A(new_n8105_), .B(new_n7970_), .C(new_n7636_), .Y(new_n8106_));
  AOI22X1  g07914(.A0(new_n7652_), .A1(new_n7646_), .B0(new_n7635_), .B1(\asqrt[38] ), .Y(new_n8107_));
  AOI21X1  g07915(.A0(new_n8107_), .A1(\asqrt[29] ), .B0(new_n7651_), .Y(new_n8108_));
  NOR2X1   g07916(.A(new_n8108_), .B(new_n8106_), .Y(new_n8109_));
  AOI21X1  g07917(.A0(new_n8102_), .A1(new_n8099_), .B0(new_n4493_), .Y(new_n8110_));
  NOR2X1   g07918(.A(new_n8110_), .B(\asqrt[39] ), .Y(new_n8111_));
  AOI21X1  g07919(.A0(new_n8111_), .A1(new_n8104_), .B0(new_n8109_), .Y(new_n8112_));
  OAI21X1  g07920(.A0(new_n8112_), .A1(new_n8093_), .B0(\asqrt[40] ), .Y(new_n8113_));
  AND2X1   g07921(.A(new_n7687_), .B(new_n7685_), .Y(new_n8114_));
  OR4X1    g07922(.A(new_n7970_), .B(new_n8114_), .C(new_n7659_), .D(new_n7686_), .Y(new_n8115_));
  OR2X1    g07923(.A(new_n8114_), .B(new_n7686_), .Y(new_n8116_));
  OAI21X1  g07924(.A0(new_n8116_), .A1(new_n7970_), .B0(new_n7659_), .Y(new_n8117_));
  AND2X1   g07925(.A(new_n8117_), .B(new_n8115_), .Y(new_n8118_));
  INVX1    g07926(.A(new_n8118_), .Y(new_n8119_));
  AOI21X1  g07927(.A0(new_n8103_), .A1(new_n8094_), .B0(new_n8110_), .Y(new_n8120_));
  OAI21X1  g07928(.A0(new_n8120_), .A1(new_n4165_), .B0(new_n3863_), .Y(new_n8121_));
  OAI21X1  g07929(.A0(new_n8121_), .A1(new_n8112_), .B0(new_n8119_), .Y(new_n8122_));
  AOI21X1  g07930(.A0(new_n8122_), .A1(new_n8113_), .B0(new_n3564_), .Y(new_n8123_));
  OR4X1    g07931(.A(new_n7970_), .B(new_n7697_), .C(new_n7670_), .D(new_n7664_), .Y(new_n8124_));
  NAND2X1  g07932(.A(new_n7671_), .B(new_n7689_), .Y(new_n8125_));
  OAI21X1  g07933(.A0(new_n8125_), .A1(new_n7970_), .B0(new_n7670_), .Y(new_n8126_));
  AND2X1   g07934(.A(new_n8126_), .B(new_n8124_), .Y(new_n8127_));
  INVX1    g07935(.A(new_n8127_), .Y(new_n8128_));
  NAND3X1  g07936(.A(new_n8122_), .B(new_n8113_), .C(new_n3564_), .Y(new_n8129_));
  AOI21X1  g07937(.A0(new_n8129_), .A1(new_n8128_), .B0(new_n8123_), .Y(new_n8130_));
  OR2X1    g07938(.A(new_n8130_), .B(new_n3276_), .Y(new_n8131_));
  AND2X1   g07939(.A(new_n8129_), .B(new_n8128_), .Y(new_n8132_));
  AND2X1   g07940(.A(new_n7713_), .B(new_n7712_), .Y(new_n8133_));
  NOR4X1   g07941(.A(new_n7970_), .B(new_n8133_), .C(new_n7680_), .D(new_n7711_), .Y(new_n8134_));
  AOI22X1  g07942(.A0(new_n7713_), .A1(new_n7712_), .B0(new_n7698_), .B1(\asqrt[41] ), .Y(new_n8135_));
  AOI21X1  g07943(.A0(new_n8135_), .A1(\asqrt[29] ), .B0(new_n7679_), .Y(new_n8136_));
  NOR2X1   g07944(.A(new_n8136_), .B(new_n8134_), .Y(new_n8137_));
  INVX1    g07945(.A(new_n8137_), .Y(new_n8138_));
  OR2X1    g07946(.A(new_n8123_), .B(\asqrt[42] ), .Y(new_n8139_));
  OAI21X1  g07947(.A0(new_n8139_), .A1(new_n8132_), .B0(new_n8138_), .Y(new_n8140_));
  AOI21X1  g07948(.A0(new_n8140_), .A1(new_n8131_), .B0(new_n3008_), .Y(new_n8141_));
  AND2X1   g07949(.A(new_n7699_), .B(new_n7691_), .Y(new_n8142_));
  OR4X1    g07950(.A(new_n7970_), .B(new_n8142_), .C(new_n7716_), .D(new_n7692_), .Y(new_n8143_));
  OR2X1    g07951(.A(new_n8142_), .B(new_n7692_), .Y(new_n8144_));
  OAI21X1  g07952(.A0(new_n8144_), .A1(new_n7970_), .B0(new_n7716_), .Y(new_n8145_));
  AND2X1   g07953(.A(new_n8145_), .B(new_n8143_), .Y(new_n8146_));
  OR2X1    g07954(.A(new_n8120_), .B(new_n4165_), .Y(new_n8147_));
  AND2X1   g07955(.A(new_n8103_), .B(new_n8094_), .Y(new_n8148_));
  INVX1    g07956(.A(new_n8109_), .Y(new_n8149_));
  OR2X1    g07957(.A(new_n8110_), .B(\asqrt[39] ), .Y(new_n8150_));
  OAI21X1  g07958(.A0(new_n8150_), .A1(new_n8148_), .B0(new_n8149_), .Y(new_n8151_));
  AOI21X1  g07959(.A0(new_n8151_), .A1(new_n8147_), .B0(new_n3863_), .Y(new_n8152_));
  AOI21X1  g07960(.A0(new_n8092_), .A1(\asqrt[39] ), .B0(\asqrt[40] ), .Y(new_n8153_));
  AOI21X1  g07961(.A0(new_n8153_), .A1(new_n8151_), .B0(new_n8118_), .Y(new_n8154_));
  OAI21X1  g07962(.A0(new_n8154_), .A1(new_n8152_), .B0(\asqrt[41] ), .Y(new_n8155_));
  NOR3X1   g07963(.A(new_n8154_), .B(new_n8152_), .C(\asqrt[41] ), .Y(new_n8156_));
  OAI21X1  g07964(.A0(new_n8156_), .A1(new_n8127_), .B0(new_n8155_), .Y(new_n8157_));
  AOI21X1  g07965(.A0(new_n8157_), .A1(\asqrt[42] ), .B0(\asqrt[43] ), .Y(new_n8158_));
  AOI21X1  g07966(.A0(new_n8158_), .A1(new_n8140_), .B0(new_n8146_), .Y(new_n8159_));
  OAI21X1  g07967(.A0(new_n8159_), .A1(new_n8141_), .B0(\asqrt[44] ), .Y(new_n8160_));
  OR4X1    g07968(.A(new_n7970_), .B(new_n7707_), .C(new_n7710_), .D(new_n7734_), .Y(new_n8161_));
  NAND2X1  g07969(.A(new_n7719_), .B(new_n7701_), .Y(new_n8162_));
  OAI21X1  g07970(.A0(new_n8162_), .A1(new_n7970_), .B0(new_n7710_), .Y(new_n8163_));
  AND2X1   g07971(.A(new_n8163_), .B(new_n8161_), .Y(new_n8164_));
  NOR3X1   g07972(.A(new_n8159_), .B(new_n8141_), .C(\asqrt[44] ), .Y(new_n8165_));
  OAI21X1  g07973(.A0(new_n8165_), .A1(new_n8164_), .B0(new_n8160_), .Y(new_n8166_));
  AND2X1   g07974(.A(new_n8166_), .B(\asqrt[45] ), .Y(new_n8167_));
  INVX1    g07975(.A(new_n8164_), .Y(new_n8168_));
  AND2X1   g07976(.A(new_n8157_), .B(\asqrt[42] ), .Y(new_n8169_));
  NAND2X1  g07977(.A(new_n8129_), .B(new_n8128_), .Y(new_n8170_));
  NOR2X1   g07978(.A(new_n8123_), .B(\asqrt[42] ), .Y(new_n8171_));
  AOI21X1  g07979(.A0(new_n8171_), .A1(new_n8170_), .B0(new_n8137_), .Y(new_n8172_));
  OAI21X1  g07980(.A0(new_n8172_), .A1(new_n8169_), .B0(\asqrt[43] ), .Y(new_n8173_));
  INVX1    g07981(.A(new_n8146_), .Y(new_n8174_));
  OAI21X1  g07982(.A0(new_n8130_), .A1(new_n3276_), .B0(new_n3008_), .Y(new_n8175_));
  OAI21X1  g07983(.A0(new_n8175_), .A1(new_n8172_), .B0(new_n8174_), .Y(new_n8176_));
  NAND3X1  g07984(.A(new_n8176_), .B(new_n8173_), .C(new_n2769_), .Y(new_n8177_));
  NAND2X1  g07985(.A(new_n8177_), .B(new_n8168_), .Y(new_n8178_));
  OAI21X1  g07986(.A0(new_n7758_), .A1(new_n7756_), .B0(new_n7725_), .Y(new_n8179_));
  NOR3X1   g07987(.A(new_n8179_), .B(new_n7970_), .C(new_n7709_), .Y(new_n8180_));
  AOI22X1  g07988(.A0(new_n7726_), .A1(new_n7720_), .B0(new_n7708_), .B1(\asqrt[44] ), .Y(new_n8181_));
  AOI21X1  g07989(.A0(new_n8181_), .A1(\asqrt[29] ), .B0(new_n7725_), .Y(new_n8182_));
  NOR2X1   g07990(.A(new_n8182_), .B(new_n8180_), .Y(new_n8183_));
  AOI21X1  g07991(.A0(new_n8176_), .A1(new_n8173_), .B0(new_n2769_), .Y(new_n8184_));
  NOR2X1   g07992(.A(new_n8184_), .B(\asqrt[45] ), .Y(new_n8185_));
  AOI21X1  g07993(.A0(new_n8185_), .A1(new_n8178_), .B0(new_n8183_), .Y(new_n8186_));
  OAI21X1  g07994(.A0(new_n8186_), .A1(new_n8167_), .B0(\asqrt[46] ), .Y(new_n8187_));
  AND2X1   g07995(.A(new_n7761_), .B(new_n7759_), .Y(new_n8188_));
  OR4X1    g07996(.A(new_n7970_), .B(new_n8188_), .C(new_n7733_), .D(new_n7760_), .Y(new_n8189_));
  OR2X1    g07997(.A(new_n8188_), .B(new_n7760_), .Y(new_n8190_));
  OAI21X1  g07998(.A0(new_n8190_), .A1(new_n7970_), .B0(new_n7733_), .Y(new_n8191_));
  AND2X1   g07999(.A(new_n8191_), .B(new_n8189_), .Y(new_n8192_));
  INVX1    g08000(.A(new_n8192_), .Y(new_n8193_));
  AOI21X1  g08001(.A0(new_n8177_), .A1(new_n8168_), .B0(new_n8184_), .Y(new_n8194_));
  OAI21X1  g08002(.A0(new_n8194_), .A1(new_n2570_), .B0(new_n2263_), .Y(new_n8195_));
  OAI21X1  g08003(.A0(new_n8195_), .A1(new_n8186_), .B0(new_n8193_), .Y(new_n8196_));
  AOI21X1  g08004(.A0(new_n8196_), .A1(new_n8187_), .B0(new_n2040_), .Y(new_n8197_));
  NAND3X1  g08005(.A(new_n7745_), .B(new_n7743_), .C(new_n7763_), .Y(new_n8198_));
  NOR3X1   g08006(.A(new_n7970_), .B(new_n7771_), .C(new_n7738_), .Y(new_n8199_));
  OAI22X1  g08007(.A0(new_n8199_), .A1(new_n7743_), .B0(new_n8198_), .B1(new_n7970_), .Y(new_n8200_));
  NAND3X1  g08008(.A(new_n8196_), .B(new_n8187_), .C(new_n2040_), .Y(new_n8201_));
  AOI21X1  g08009(.A0(new_n8201_), .A1(new_n8200_), .B0(new_n8197_), .Y(new_n8202_));
  OR2X1    g08010(.A(new_n8202_), .B(new_n1834_), .Y(new_n8203_));
  AND2X1   g08011(.A(new_n8201_), .B(new_n8200_), .Y(new_n8204_));
  AND2X1   g08012(.A(new_n7787_), .B(new_n7786_), .Y(new_n8205_));
  NOR4X1   g08013(.A(new_n7970_), .B(new_n8205_), .C(new_n7754_), .D(new_n7785_), .Y(new_n8206_));
  AOI22X1  g08014(.A0(new_n7787_), .A1(new_n7786_), .B0(new_n7772_), .B1(\asqrt[47] ), .Y(new_n8207_));
  AOI21X1  g08015(.A0(new_n8207_), .A1(\asqrt[29] ), .B0(new_n7753_), .Y(new_n8208_));
  NOR2X1   g08016(.A(new_n8208_), .B(new_n8206_), .Y(new_n8209_));
  INVX1    g08017(.A(new_n8209_), .Y(new_n8210_));
  OR2X1    g08018(.A(new_n8197_), .B(\asqrt[48] ), .Y(new_n8211_));
  OAI21X1  g08019(.A0(new_n8211_), .A1(new_n8204_), .B0(new_n8210_), .Y(new_n8212_));
  AOI21X1  g08020(.A0(new_n8212_), .A1(new_n8203_), .B0(new_n1632_), .Y(new_n8213_));
  AND2X1   g08021(.A(new_n7773_), .B(new_n7765_), .Y(new_n8214_));
  OR4X1    g08022(.A(new_n7970_), .B(new_n8214_), .C(new_n7790_), .D(new_n7766_), .Y(new_n8215_));
  OR2X1    g08023(.A(new_n8214_), .B(new_n7766_), .Y(new_n8216_));
  OAI21X1  g08024(.A0(new_n8216_), .A1(new_n7970_), .B0(new_n7790_), .Y(new_n8217_));
  AND2X1   g08025(.A(new_n8217_), .B(new_n8215_), .Y(new_n8218_));
  OR2X1    g08026(.A(new_n8194_), .B(new_n2570_), .Y(new_n8219_));
  AND2X1   g08027(.A(new_n8177_), .B(new_n8168_), .Y(new_n8220_));
  INVX1    g08028(.A(new_n8183_), .Y(new_n8221_));
  OR2X1    g08029(.A(new_n8184_), .B(\asqrt[45] ), .Y(new_n8222_));
  OAI21X1  g08030(.A0(new_n8222_), .A1(new_n8220_), .B0(new_n8221_), .Y(new_n8223_));
  AOI21X1  g08031(.A0(new_n8223_), .A1(new_n8219_), .B0(new_n2263_), .Y(new_n8224_));
  AOI21X1  g08032(.A0(new_n8166_), .A1(\asqrt[45] ), .B0(\asqrt[46] ), .Y(new_n8225_));
  AOI21X1  g08033(.A0(new_n8225_), .A1(new_n8223_), .B0(new_n8192_), .Y(new_n8226_));
  OAI21X1  g08034(.A0(new_n8226_), .A1(new_n8224_), .B0(\asqrt[47] ), .Y(new_n8227_));
  INVX1    g08035(.A(new_n8200_), .Y(new_n8228_));
  NOR3X1   g08036(.A(new_n8226_), .B(new_n8224_), .C(\asqrt[47] ), .Y(new_n8229_));
  OAI21X1  g08037(.A0(new_n8229_), .A1(new_n8228_), .B0(new_n8227_), .Y(new_n8230_));
  AOI21X1  g08038(.A0(new_n8230_), .A1(\asqrt[48] ), .B0(\asqrt[49] ), .Y(new_n8231_));
  AOI21X1  g08039(.A0(new_n8231_), .A1(new_n8212_), .B0(new_n8218_), .Y(new_n8232_));
  OAI21X1  g08040(.A0(new_n8232_), .A1(new_n8213_), .B0(\asqrt[50] ), .Y(new_n8233_));
  OR4X1    g08041(.A(new_n7970_), .B(new_n7781_), .C(new_n7784_), .D(new_n7808_), .Y(new_n8234_));
  NAND2X1  g08042(.A(new_n7793_), .B(new_n7775_), .Y(new_n8235_));
  OAI21X1  g08043(.A0(new_n8235_), .A1(new_n7970_), .B0(new_n7784_), .Y(new_n8236_));
  AND2X1   g08044(.A(new_n8236_), .B(new_n8234_), .Y(new_n8237_));
  NOR3X1   g08045(.A(new_n8232_), .B(new_n8213_), .C(\asqrt[50] ), .Y(new_n8238_));
  OAI21X1  g08046(.A0(new_n8238_), .A1(new_n8237_), .B0(new_n8233_), .Y(new_n8239_));
  AND2X1   g08047(.A(new_n8239_), .B(\asqrt[51] ), .Y(new_n8240_));
  INVX1    g08048(.A(new_n8237_), .Y(new_n8241_));
  AND2X1   g08049(.A(new_n8230_), .B(\asqrt[48] ), .Y(new_n8242_));
  NAND2X1  g08050(.A(new_n8201_), .B(new_n8200_), .Y(new_n8243_));
  NOR2X1   g08051(.A(new_n8197_), .B(\asqrt[48] ), .Y(new_n8244_));
  AOI21X1  g08052(.A0(new_n8244_), .A1(new_n8243_), .B0(new_n8209_), .Y(new_n8245_));
  OAI21X1  g08053(.A0(new_n8245_), .A1(new_n8242_), .B0(\asqrt[49] ), .Y(new_n8246_));
  INVX1    g08054(.A(new_n8218_), .Y(new_n8247_));
  OAI21X1  g08055(.A0(new_n8202_), .A1(new_n1834_), .B0(new_n1632_), .Y(new_n8248_));
  OAI21X1  g08056(.A0(new_n8248_), .A1(new_n8245_), .B0(new_n8247_), .Y(new_n8249_));
  NAND3X1  g08057(.A(new_n8249_), .B(new_n8246_), .C(new_n1469_), .Y(new_n8250_));
  NAND2X1  g08058(.A(new_n8250_), .B(new_n8241_), .Y(new_n8251_));
  OAI21X1  g08059(.A0(new_n7832_), .A1(new_n7830_), .B0(new_n7799_), .Y(new_n8252_));
  NOR3X1   g08060(.A(new_n8252_), .B(new_n7970_), .C(new_n7783_), .Y(new_n8253_));
  AOI22X1  g08061(.A0(new_n7800_), .A1(new_n7794_), .B0(new_n7782_), .B1(\asqrt[50] ), .Y(new_n8254_));
  AOI21X1  g08062(.A0(new_n8254_), .A1(\asqrt[29] ), .B0(new_n7799_), .Y(new_n8255_));
  NOR2X1   g08063(.A(new_n8255_), .B(new_n8253_), .Y(new_n8256_));
  AOI21X1  g08064(.A0(new_n8249_), .A1(new_n8246_), .B0(new_n1469_), .Y(new_n8257_));
  NOR2X1   g08065(.A(new_n8257_), .B(\asqrt[51] ), .Y(new_n8258_));
  AOI21X1  g08066(.A0(new_n8258_), .A1(new_n8251_), .B0(new_n8256_), .Y(new_n8259_));
  OAI21X1  g08067(.A0(new_n8259_), .A1(new_n8240_), .B0(\asqrt[52] ), .Y(new_n8260_));
  AND2X1   g08068(.A(new_n7835_), .B(new_n7833_), .Y(new_n8261_));
  OR4X1    g08069(.A(new_n7970_), .B(new_n8261_), .C(new_n7807_), .D(new_n7834_), .Y(new_n8262_));
  OR2X1    g08070(.A(new_n8261_), .B(new_n7834_), .Y(new_n8263_));
  OAI21X1  g08071(.A0(new_n8263_), .A1(new_n7970_), .B0(new_n7807_), .Y(new_n8264_));
  AND2X1   g08072(.A(new_n8264_), .B(new_n8262_), .Y(new_n8265_));
  INVX1    g08073(.A(new_n8265_), .Y(new_n8266_));
  AOI21X1  g08074(.A0(new_n8250_), .A1(new_n8241_), .B0(new_n8257_), .Y(new_n8267_));
  OAI21X1  g08075(.A0(new_n8267_), .A1(new_n1277_), .B0(new_n1111_), .Y(new_n8268_));
  OAI21X1  g08076(.A0(new_n8268_), .A1(new_n8259_), .B0(new_n8266_), .Y(new_n8269_));
  AOI21X1  g08077(.A0(new_n8269_), .A1(new_n8260_), .B0(new_n968_), .Y(new_n8270_));
  OR4X1    g08078(.A(new_n7970_), .B(new_n7845_), .C(new_n7818_), .D(new_n7812_), .Y(new_n8271_));
  NAND2X1  g08079(.A(new_n7819_), .B(new_n7837_), .Y(new_n8272_));
  OAI21X1  g08080(.A0(new_n8272_), .A1(new_n7970_), .B0(new_n7818_), .Y(new_n8273_));
  AND2X1   g08081(.A(new_n8273_), .B(new_n8271_), .Y(new_n8274_));
  INVX1    g08082(.A(new_n8274_), .Y(new_n8275_));
  NAND3X1  g08083(.A(new_n8269_), .B(new_n8260_), .C(new_n968_), .Y(new_n8276_));
  AOI21X1  g08084(.A0(new_n8276_), .A1(new_n8275_), .B0(new_n8270_), .Y(new_n8277_));
  OR2X1    g08085(.A(new_n8277_), .B(new_n902_), .Y(new_n8278_));
  OR2X1    g08086(.A(new_n8267_), .B(new_n1277_), .Y(new_n8279_));
  AND2X1   g08087(.A(new_n8250_), .B(new_n8241_), .Y(new_n8280_));
  INVX1    g08088(.A(new_n8256_), .Y(new_n8281_));
  OR2X1    g08089(.A(new_n8257_), .B(\asqrt[51] ), .Y(new_n8282_));
  OAI21X1  g08090(.A0(new_n8282_), .A1(new_n8280_), .B0(new_n8281_), .Y(new_n8283_));
  AOI21X1  g08091(.A0(new_n8283_), .A1(new_n8279_), .B0(new_n1111_), .Y(new_n8284_));
  AOI21X1  g08092(.A0(new_n8239_), .A1(\asqrt[51] ), .B0(\asqrt[52] ), .Y(new_n8285_));
  AOI21X1  g08093(.A0(new_n8285_), .A1(new_n8283_), .B0(new_n8265_), .Y(new_n8286_));
  NOR3X1   g08094(.A(new_n8286_), .B(new_n8284_), .C(\asqrt[53] ), .Y(new_n8287_));
  NOR2X1   g08095(.A(new_n8287_), .B(new_n8274_), .Y(new_n8288_));
  AND2X1   g08096(.A(new_n7861_), .B(new_n7860_), .Y(new_n8289_));
  NOR4X1   g08097(.A(new_n7970_), .B(new_n8289_), .C(new_n7828_), .D(new_n7859_), .Y(new_n8290_));
  AOI22X1  g08098(.A0(new_n7861_), .A1(new_n7860_), .B0(new_n7846_), .B1(\asqrt[53] ), .Y(new_n8291_));
  AOI21X1  g08099(.A0(new_n8291_), .A1(\asqrt[29] ), .B0(new_n7827_), .Y(new_n8292_));
  NOR2X1   g08100(.A(new_n8292_), .B(new_n8290_), .Y(new_n8293_));
  INVX1    g08101(.A(new_n8293_), .Y(new_n8294_));
  OAI21X1  g08102(.A0(new_n8286_), .A1(new_n8284_), .B0(\asqrt[53] ), .Y(new_n8295_));
  NAND2X1  g08103(.A(new_n8295_), .B(new_n902_), .Y(new_n8296_));
  OAI21X1  g08104(.A0(new_n8296_), .A1(new_n8288_), .B0(new_n8294_), .Y(new_n8297_));
  AOI21X1  g08105(.A0(new_n8297_), .A1(new_n8278_), .B0(new_n697_), .Y(new_n8298_));
  AND2X1   g08106(.A(new_n7847_), .B(new_n7839_), .Y(new_n8299_));
  OR4X1    g08107(.A(new_n7970_), .B(new_n8299_), .C(new_n7864_), .D(new_n7840_), .Y(new_n8300_));
  OR2X1    g08108(.A(new_n8299_), .B(new_n7840_), .Y(new_n8301_));
  OAI21X1  g08109(.A0(new_n8301_), .A1(new_n7970_), .B0(new_n7864_), .Y(new_n8302_));
  AND2X1   g08110(.A(new_n8302_), .B(new_n8300_), .Y(new_n8303_));
  OAI21X1  g08111(.A0(new_n8287_), .A1(new_n8274_), .B0(new_n8295_), .Y(new_n8304_));
  AOI21X1  g08112(.A0(new_n8304_), .A1(\asqrt[54] ), .B0(\asqrt[55] ), .Y(new_n8305_));
  AOI21X1  g08113(.A0(new_n8305_), .A1(new_n8297_), .B0(new_n8303_), .Y(new_n8306_));
  OAI21X1  g08114(.A0(new_n8306_), .A1(new_n8298_), .B0(\asqrt[56] ), .Y(new_n8307_));
  NAND3X1  g08115(.A(new_n7867_), .B(new_n7854_), .C(new_n7849_), .Y(new_n8308_));
  NOR3X1   g08116(.A(new_n7970_), .B(new_n7855_), .C(new_n7882_), .Y(new_n8309_));
  OAI22X1  g08117(.A0(new_n8309_), .A1(new_n7854_), .B0(new_n8308_), .B1(new_n7970_), .Y(new_n8310_));
  INVX1    g08118(.A(new_n8310_), .Y(new_n8311_));
  NOR3X1   g08119(.A(new_n8306_), .B(new_n8298_), .C(\asqrt[56] ), .Y(new_n8312_));
  OAI21X1  g08120(.A0(new_n8312_), .A1(new_n8311_), .B0(new_n8307_), .Y(new_n8313_));
  AND2X1   g08121(.A(new_n8313_), .B(\asqrt[57] ), .Y(new_n8314_));
  AND2X1   g08122(.A(new_n8304_), .B(\asqrt[54] ), .Y(new_n8315_));
  OR2X1    g08123(.A(new_n8287_), .B(new_n8274_), .Y(new_n8316_));
  AND2X1   g08124(.A(new_n8295_), .B(new_n902_), .Y(new_n8317_));
  AOI21X1  g08125(.A0(new_n8317_), .A1(new_n8316_), .B0(new_n8293_), .Y(new_n8318_));
  OAI21X1  g08126(.A0(new_n8318_), .A1(new_n8315_), .B0(\asqrt[55] ), .Y(new_n8319_));
  INVX1    g08127(.A(new_n8303_), .Y(new_n8320_));
  OAI21X1  g08128(.A0(new_n8277_), .A1(new_n902_), .B0(new_n697_), .Y(new_n8321_));
  OAI21X1  g08129(.A0(new_n8321_), .A1(new_n8318_), .B0(new_n8320_), .Y(new_n8322_));
  NAND3X1  g08130(.A(new_n8322_), .B(new_n8319_), .C(new_n582_), .Y(new_n8323_));
  NAND2X1  g08131(.A(new_n8323_), .B(new_n8310_), .Y(new_n8324_));
  OAI21X1  g08132(.A0(new_n7906_), .A1(new_n7904_), .B0(new_n7873_), .Y(new_n8325_));
  NOR3X1   g08133(.A(new_n8325_), .B(new_n7970_), .C(new_n7857_), .Y(new_n8326_));
  AOI22X1  g08134(.A0(new_n7874_), .A1(new_n7868_), .B0(new_n7856_), .B1(\asqrt[56] ), .Y(new_n8327_));
  AOI21X1  g08135(.A0(new_n8327_), .A1(\asqrt[29] ), .B0(new_n7873_), .Y(new_n8328_));
  NOR2X1   g08136(.A(new_n8328_), .B(new_n8326_), .Y(new_n8329_));
  AND2X1   g08137(.A(new_n8307_), .B(new_n481_), .Y(new_n8330_));
  AOI21X1  g08138(.A0(new_n8330_), .A1(new_n8324_), .B0(new_n8329_), .Y(new_n8331_));
  OAI21X1  g08139(.A0(new_n8331_), .A1(new_n8314_), .B0(\asqrt[58] ), .Y(new_n8332_));
  AND2X1   g08140(.A(new_n7909_), .B(new_n7907_), .Y(new_n8333_));
  OR4X1    g08141(.A(new_n7970_), .B(new_n8333_), .C(new_n7881_), .D(new_n7908_), .Y(new_n8334_));
  OR2X1    g08142(.A(new_n8333_), .B(new_n7908_), .Y(new_n8335_));
  OAI21X1  g08143(.A0(new_n8335_), .A1(new_n7970_), .B0(new_n7881_), .Y(new_n8336_));
  AND2X1   g08144(.A(new_n8336_), .B(new_n8334_), .Y(new_n8337_));
  INVX1    g08145(.A(new_n8337_), .Y(new_n8338_));
  AOI21X1  g08146(.A0(new_n8322_), .A1(new_n8319_), .B0(new_n582_), .Y(new_n8339_));
  AOI21X1  g08147(.A0(new_n8323_), .A1(new_n8310_), .B0(new_n8339_), .Y(new_n8340_));
  OAI21X1  g08148(.A0(new_n8340_), .A1(new_n481_), .B0(new_n399_), .Y(new_n8341_));
  OAI21X1  g08149(.A0(new_n8341_), .A1(new_n8331_), .B0(new_n8338_), .Y(new_n8342_));
  AOI21X1  g08150(.A0(new_n8342_), .A1(new_n8332_), .B0(new_n328_), .Y(new_n8343_));
  OR4X1    g08151(.A(new_n7970_), .B(new_n7919_), .C(new_n7892_), .D(new_n7886_), .Y(new_n8344_));
  OR2X1    g08152(.A(new_n7919_), .B(new_n7886_), .Y(new_n8345_));
  OAI21X1  g08153(.A0(new_n8345_), .A1(new_n7970_), .B0(new_n7892_), .Y(new_n8346_));
  AND2X1   g08154(.A(new_n8346_), .B(new_n8344_), .Y(new_n8347_));
  INVX1    g08155(.A(new_n8347_), .Y(new_n8348_));
  NAND3X1  g08156(.A(new_n8342_), .B(new_n8332_), .C(new_n328_), .Y(new_n8349_));
  AOI21X1  g08157(.A0(new_n8349_), .A1(new_n8348_), .B0(new_n8343_), .Y(new_n8350_));
  OR2X1    g08158(.A(new_n8350_), .B(new_n292_), .Y(new_n8351_));
  OR2X1    g08159(.A(new_n8340_), .B(new_n481_), .Y(new_n8352_));
  AND2X1   g08160(.A(new_n8323_), .B(new_n8310_), .Y(new_n8353_));
  INVX1    g08161(.A(new_n8329_), .Y(new_n8354_));
  NAND2X1  g08162(.A(new_n8307_), .B(new_n481_), .Y(new_n8355_));
  OAI21X1  g08163(.A0(new_n8355_), .A1(new_n8353_), .B0(new_n8354_), .Y(new_n8356_));
  AOI21X1  g08164(.A0(new_n8356_), .A1(new_n8352_), .B0(new_n399_), .Y(new_n8357_));
  AOI21X1  g08165(.A0(new_n8313_), .A1(\asqrt[57] ), .B0(\asqrt[58] ), .Y(new_n8358_));
  AOI21X1  g08166(.A0(new_n8358_), .A1(new_n8356_), .B0(new_n8337_), .Y(new_n8359_));
  NOR3X1   g08167(.A(new_n8359_), .B(new_n8357_), .C(\asqrt[59] ), .Y(new_n8360_));
  NOR2X1   g08168(.A(new_n8360_), .B(new_n8347_), .Y(new_n8361_));
  AND2X1   g08169(.A(new_n7935_), .B(new_n7934_), .Y(new_n8362_));
  NOR4X1   g08170(.A(new_n7970_), .B(new_n8362_), .C(new_n7902_), .D(new_n7933_), .Y(new_n8363_));
  AOI22X1  g08171(.A0(new_n7935_), .A1(new_n7934_), .B0(new_n7920_), .B1(\asqrt[59] ), .Y(new_n8364_));
  AOI21X1  g08172(.A0(new_n8364_), .A1(\asqrt[29] ), .B0(new_n7901_), .Y(new_n8365_));
  NOR2X1   g08173(.A(new_n8365_), .B(new_n8363_), .Y(new_n8366_));
  INVX1    g08174(.A(new_n8366_), .Y(new_n8367_));
  OAI21X1  g08175(.A0(new_n8359_), .A1(new_n8357_), .B0(\asqrt[59] ), .Y(new_n8368_));
  NAND2X1  g08176(.A(new_n8368_), .B(new_n292_), .Y(new_n8369_));
  OAI21X1  g08177(.A0(new_n8369_), .A1(new_n8361_), .B0(new_n8367_), .Y(new_n8370_));
  AOI21X1  g08178(.A0(new_n8370_), .A1(new_n8351_), .B0(new_n217_), .Y(new_n8371_));
  AND2X1   g08179(.A(new_n7921_), .B(new_n7913_), .Y(new_n8372_));
  OR4X1    g08180(.A(new_n7970_), .B(new_n8372_), .C(new_n7938_), .D(new_n7914_), .Y(new_n8373_));
  OR2X1    g08181(.A(new_n8372_), .B(new_n7914_), .Y(new_n8374_));
  OAI21X1  g08182(.A0(new_n8374_), .A1(new_n7970_), .B0(new_n7938_), .Y(new_n8375_));
  AND2X1   g08183(.A(new_n8375_), .B(new_n8373_), .Y(new_n8376_));
  OAI21X1  g08184(.A0(new_n8360_), .A1(new_n8347_), .B0(new_n8368_), .Y(new_n8377_));
  AOI21X1  g08185(.A0(new_n8377_), .A1(\asqrt[60] ), .B0(\asqrt[61] ), .Y(new_n8378_));
  AOI21X1  g08186(.A0(new_n8378_), .A1(new_n8370_), .B0(new_n8376_), .Y(new_n8379_));
  OAI21X1  g08187(.A0(new_n8379_), .A1(new_n8371_), .B0(\asqrt[62] ), .Y(new_n8380_));
  OR4X1    g08188(.A(new_n7970_), .B(new_n7929_), .C(new_n7932_), .D(new_n7948_), .Y(new_n8381_));
  OR2X1    g08189(.A(new_n7929_), .B(new_n7948_), .Y(new_n8382_));
  OAI21X1  g08190(.A0(new_n8382_), .A1(new_n7970_), .B0(new_n7932_), .Y(new_n8383_));
  AND2X1   g08191(.A(new_n8383_), .B(new_n8381_), .Y(new_n8384_));
  NOR3X1   g08192(.A(new_n8379_), .B(new_n8371_), .C(\asqrt[62] ), .Y(new_n8385_));
  OAI21X1  g08193(.A0(new_n8385_), .A1(new_n8384_), .B0(new_n8380_), .Y(new_n8386_));
  AND2X1   g08194(.A(new_n7949_), .B(new_n7942_), .Y(new_n8387_));
  NOR4X1   g08195(.A(new_n7970_), .B(new_n8387_), .C(new_n7989_), .D(new_n7931_), .Y(new_n8388_));
  INVX1    g08196(.A(new_n8388_), .Y(new_n8389_));
  OAI22X1  g08197(.A0(new_n7990_), .A1(new_n7988_), .B0(new_n7959_), .B1(new_n199_), .Y(new_n8390_));
  OAI21X1  g08198(.A0(new_n8390_), .A1(new_n7970_), .B0(new_n7989_), .Y(new_n8391_));
  AND2X1   g08199(.A(new_n8391_), .B(new_n8389_), .Y(new_n8392_));
  INVX1    g08200(.A(new_n8392_), .Y(new_n8393_));
  AND2X1   g08201(.A(new_n7994_), .B(new_n7991_), .Y(new_n8394_));
  AOI21X1  g08202(.A0(new_n7991_), .A1(new_n7987_), .B0(new_n7953_), .Y(new_n8395_));
  AOI21X1  g08203(.A0(new_n8395_), .A1(\asqrt[29] ), .B0(new_n8394_), .Y(new_n8396_));
  AND2X1   g08204(.A(new_n8396_), .B(new_n8393_), .Y(new_n8397_));
  AOI21X1  g08205(.A0(new_n8397_), .A1(new_n8386_), .B0(\asqrt[63] ), .Y(new_n8398_));
  NOR2X1   g08206(.A(new_n8385_), .B(new_n8384_), .Y(new_n8399_));
  NAND2X1  g08207(.A(new_n8392_), .B(new_n8380_), .Y(new_n8400_));
  NAND2X1  g08208(.A(new_n7991_), .B(new_n7987_), .Y(new_n8401_));
  AOI21X1  g08209(.A0(\asqrt[29] ), .A1(new_n7954_), .B0(new_n8401_), .Y(new_n8402_));
  NOR3X1   g08210(.A(new_n8402_), .B(new_n8395_), .C(new_n193_), .Y(new_n8403_));
  AND2X1   g08211(.A(new_n7958_), .B(new_n193_), .Y(new_n8404_));
  INVX1    g08212(.A(new_n7967_), .Y(new_n8405_));
  OR2X1    g08213(.A(new_n8405_), .B(new_n7951_), .Y(new_n8406_));
  AOI21X1  g08214(.A0(new_n7952_), .A1(new_n7538_), .B0(new_n8406_), .Y(new_n8407_));
  NAND2X1  g08215(.A(new_n8407_), .B(new_n7963_), .Y(new_n8408_));
  NOR3X1   g08216(.A(new_n8408_), .B(new_n8394_), .C(new_n8404_), .Y(new_n8409_));
  NOR2X1   g08217(.A(new_n8409_), .B(new_n8403_), .Y(new_n8410_));
  OAI21X1  g08218(.A0(new_n8400_), .A1(new_n8399_), .B0(new_n8410_), .Y(new_n8411_));
  NOR2X1   g08219(.A(new_n8411_), .B(new_n8398_), .Y(new_n8412_));
  INVX1    g08220(.A(new_n8412_), .Y(\asqrt[28] ));
  OAI21X1  g08221(.A0(new_n8411_), .A1(new_n8398_), .B0(\a[56] ), .Y(new_n8414_));
  INVX1    g08222(.A(\a[56] ), .Y(new_n8415_));
  NOR2X1   g08223(.A(\a[55] ), .B(\a[54] ), .Y(new_n8416_));
  NAND2X1  g08224(.A(new_n8416_), .B(new_n8415_), .Y(new_n8417_));
  AOI21X1  g08225(.A0(new_n8417_), .A1(new_n8414_), .B0(new_n7970_), .Y(new_n8418_));
  AND2X1   g08226(.A(new_n8377_), .B(\asqrt[60] ), .Y(new_n8419_));
  OR2X1    g08227(.A(new_n8360_), .B(new_n8347_), .Y(new_n8420_));
  AND2X1   g08228(.A(new_n8368_), .B(new_n292_), .Y(new_n8421_));
  AOI21X1  g08229(.A0(new_n8421_), .A1(new_n8420_), .B0(new_n8366_), .Y(new_n8422_));
  OAI21X1  g08230(.A0(new_n8422_), .A1(new_n8419_), .B0(\asqrt[61] ), .Y(new_n8423_));
  INVX1    g08231(.A(new_n8376_), .Y(new_n8424_));
  OAI21X1  g08232(.A0(new_n8350_), .A1(new_n292_), .B0(new_n217_), .Y(new_n8425_));
  OAI21X1  g08233(.A0(new_n8425_), .A1(new_n8422_), .B0(new_n8424_), .Y(new_n8426_));
  AOI21X1  g08234(.A0(new_n8426_), .A1(new_n8423_), .B0(new_n199_), .Y(new_n8427_));
  INVX1    g08235(.A(new_n8384_), .Y(new_n8428_));
  NAND3X1  g08236(.A(new_n8426_), .B(new_n8423_), .C(new_n199_), .Y(new_n8429_));
  AOI21X1  g08237(.A0(new_n8429_), .A1(new_n8428_), .B0(new_n8427_), .Y(new_n8430_));
  INVX1    g08238(.A(new_n8397_), .Y(new_n8431_));
  OAI21X1  g08239(.A0(new_n8431_), .A1(new_n8430_), .B0(new_n193_), .Y(new_n8432_));
  OR2X1    g08240(.A(new_n8385_), .B(new_n8384_), .Y(new_n8433_));
  AND2X1   g08241(.A(new_n8392_), .B(new_n8380_), .Y(new_n8434_));
  INVX1    g08242(.A(new_n8410_), .Y(new_n8435_));
  AOI21X1  g08243(.A0(new_n8434_), .A1(new_n8433_), .B0(new_n8435_), .Y(new_n8436_));
  AOI21X1  g08244(.A0(new_n8436_), .A1(new_n8432_), .B0(new_n8415_), .Y(new_n8437_));
  NAND3X1  g08245(.A(new_n8417_), .B(new_n7967_), .C(new_n7963_), .Y(new_n8438_));
  OR4X1    g08246(.A(new_n8438_), .B(new_n8437_), .C(new_n8394_), .D(new_n8404_), .Y(new_n8439_));
  OAI21X1  g08247(.A0(new_n8411_), .A1(new_n8398_), .B0(new_n8415_), .Y(new_n8440_));
  AOI21X1  g08248(.A0(new_n8436_), .A1(new_n8432_), .B0(new_n7972_), .Y(new_n8441_));
  AOI21X1  g08249(.A0(new_n8440_), .A1(\a[57] ), .B0(new_n8441_), .Y(new_n8442_));
  AOI21X1  g08250(.A0(new_n8442_), .A1(new_n8439_), .B0(new_n8418_), .Y(new_n8443_));
  OR2X1    g08251(.A(new_n8443_), .B(new_n7527_), .Y(new_n8444_));
  AND2X1   g08252(.A(new_n8442_), .B(new_n8439_), .Y(new_n8445_));
  OR2X1    g08253(.A(new_n8418_), .B(\asqrt[30] ), .Y(new_n8446_));
  OAI21X1  g08254(.A0(new_n8411_), .A1(new_n8398_), .B0(new_n7971_), .Y(new_n8447_));
  AND2X1   g08255(.A(new_n8434_), .B(new_n8433_), .Y(new_n8448_));
  OR2X1    g08256(.A(new_n8409_), .B(new_n7970_), .Y(new_n8449_));
  OR4X1    g08257(.A(new_n8449_), .B(new_n8403_), .C(new_n8448_), .D(new_n8398_), .Y(new_n8450_));
  AOI21X1  g08258(.A0(new_n8450_), .A1(new_n8447_), .B0(new_n7975_), .Y(new_n8451_));
  NOR4X1   g08259(.A(new_n8449_), .B(new_n8403_), .C(new_n8448_), .D(new_n8398_), .Y(new_n8452_));
  NOR3X1   g08260(.A(new_n8452_), .B(new_n8441_), .C(\a[58] ), .Y(new_n8453_));
  OR2X1    g08261(.A(new_n8453_), .B(new_n8451_), .Y(new_n8454_));
  OAI21X1  g08262(.A0(new_n8446_), .A1(new_n8445_), .B0(new_n8454_), .Y(new_n8455_));
  AOI21X1  g08263(.A0(new_n8455_), .A1(new_n8444_), .B0(new_n7103_), .Y(new_n8456_));
  AND2X1   g08264(.A(new_n7984_), .B(new_n7981_), .Y(new_n8457_));
  NOR3X1   g08265(.A(new_n8457_), .B(new_n8021_), .C(new_n8020_), .Y(new_n8458_));
  OAI21X1  g08266(.A0(new_n8411_), .A1(new_n8398_), .B0(new_n8458_), .Y(new_n8459_));
  AOI21X1  g08267(.A0(new_n7998_), .A1(\asqrt[30] ), .B0(new_n8021_), .Y(new_n8460_));
  OAI21X1  g08268(.A0(new_n8411_), .A1(new_n8398_), .B0(new_n8460_), .Y(new_n8461_));
  NAND2X1  g08269(.A(new_n8461_), .B(new_n8457_), .Y(new_n8462_));
  AND2X1   g08270(.A(new_n8417_), .B(new_n8414_), .Y(new_n8463_));
  NOR4X1   g08271(.A(new_n8438_), .B(new_n8437_), .C(new_n8394_), .D(new_n8404_), .Y(new_n8464_));
  INVX1    g08272(.A(\a[57] ), .Y(new_n8465_));
  AOI21X1  g08273(.A0(new_n8436_), .A1(new_n8432_), .B0(\a[56] ), .Y(new_n8466_));
  OAI21X1  g08274(.A0(new_n8466_), .A1(new_n8465_), .B0(new_n8447_), .Y(new_n8467_));
  OAI22X1  g08275(.A0(new_n8467_), .A1(new_n8464_), .B0(new_n8463_), .B1(new_n7970_), .Y(new_n8468_));
  AOI21X1  g08276(.A0(new_n8468_), .A1(\asqrt[30] ), .B0(\asqrt[31] ), .Y(new_n8469_));
  AOI22X1  g08277(.A0(new_n8469_), .A1(new_n8455_), .B0(new_n8462_), .B1(new_n8459_), .Y(new_n8470_));
  OAI21X1  g08278(.A0(new_n8470_), .A1(new_n8456_), .B0(\asqrt[32] ), .Y(new_n8471_));
  AND2X1   g08279(.A(new_n7999_), .B(new_n7985_), .Y(new_n8472_));
  NOR3X1   g08280(.A(new_n8027_), .B(new_n8472_), .C(new_n7986_), .Y(new_n8473_));
  OAI21X1  g08281(.A0(new_n8411_), .A1(new_n8398_), .B0(new_n8473_), .Y(new_n8474_));
  NOR2X1   g08282(.A(new_n8472_), .B(new_n7986_), .Y(new_n8475_));
  OAI21X1  g08283(.A0(new_n8411_), .A1(new_n8398_), .B0(new_n8475_), .Y(new_n8476_));
  NAND2X1  g08284(.A(new_n8476_), .B(new_n8027_), .Y(new_n8477_));
  AND2X1   g08285(.A(new_n8477_), .B(new_n8474_), .Y(new_n8478_));
  NOR3X1   g08286(.A(new_n8470_), .B(new_n8456_), .C(\asqrt[32] ), .Y(new_n8479_));
  OAI21X1  g08287(.A0(new_n8479_), .A1(new_n8478_), .B0(new_n8471_), .Y(new_n8480_));
  AND2X1   g08288(.A(new_n8480_), .B(\asqrt[33] ), .Y(new_n8481_));
  OR2X1    g08289(.A(new_n8479_), .B(new_n8478_), .Y(new_n8482_));
  NOR3X1   g08290(.A(new_n8016_), .B(new_n8019_), .C(new_n8036_), .Y(new_n8483_));
  OAI21X1  g08291(.A0(new_n8411_), .A1(new_n8398_), .B0(new_n8483_), .Y(new_n8484_));
  NOR3X1   g08292(.A(new_n8412_), .B(new_n8016_), .C(new_n8036_), .Y(new_n8485_));
  OR2X1    g08293(.A(new_n8485_), .B(new_n8015_), .Y(new_n8486_));
  AND2X1   g08294(.A(new_n8486_), .B(new_n8484_), .Y(new_n8487_));
  AND2X1   g08295(.A(new_n8468_), .B(\asqrt[30] ), .Y(new_n8488_));
  NAND2X1  g08296(.A(new_n8442_), .B(new_n8439_), .Y(new_n8489_));
  NOR2X1   g08297(.A(new_n8418_), .B(\asqrt[30] ), .Y(new_n8490_));
  NOR2X1   g08298(.A(new_n8453_), .B(new_n8451_), .Y(new_n8491_));
  AOI21X1  g08299(.A0(new_n8490_), .A1(new_n8489_), .B0(new_n8491_), .Y(new_n8492_));
  OAI21X1  g08300(.A0(new_n8492_), .A1(new_n8488_), .B0(\asqrt[31] ), .Y(new_n8493_));
  NAND2X1  g08301(.A(new_n8462_), .B(new_n8459_), .Y(new_n8494_));
  OAI21X1  g08302(.A0(new_n8443_), .A1(new_n7527_), .B0(new_n7103_), .Y(new_n8495_));
  OAI21X1  g08303(.A0(new_n8495_), .A1(new_n8492_), .B0(new_n8494_), .Y(new_n8496_));
  AOI21X1  g08304(.A0(new_n8496_), .A1(new_n8493_), .B0(new_n6699_), .Y(new_n8497_));
  NOR2X1   g08305(.A(new_n8497_), .B(\asqrt[33] ), .Y(new_n8498_));
  AOI21X1  g08306(.A0(new_n8498_), .A1(new_n8482_), .B0(new_n8487_), .Y(new_n8499_));
  OAI21X1  g08307(.A0(new_n8499_), .A1(new_n8481_), .B0(\asqrt[34] ), .Y(new_n8500_));
  AOI21X1  g08308(.A0(new_n8037_), .A1(new_n8030_), .B0(new_n8075_), .Y(new_n8501_));
  AND2X1   g08309(.A(new_n8501_), .B(new_n8073_), .Y(new_n8502_));
  AOI22X1  g08310(.A0(new_n8037_), .A1(new_n8030_), .B0(new_n8017_), .B1(\asqrt[33] ), .Y(new_n8503_));
  AOI21X1  g08311(.A0(new_n8503_), .A1(\asqrt[28] ), .B0(new_n8035_), .Y(new_n8504_));
  AOI21X1  g08312(.A0(new_n8502_), .A1(\asqrt[28] ), .B0(new_n8504_), .Y(new_n8505_));
  INVX1    g08313(.A(new_n8505_), .Y(new_n8506_));
  INVX1    g08314(.A(new_n8478_), .Y(new_n8507_));
  NAND3X1  g08315(.A(new_n8496_), .B(new_n8493_), .C(new_n6699_), .Y(new_n8508_));
  AOI21X1  g08316(.A0(new_n8508_), .A1(new_n8507_), .B0(new_n8497_), .Y(new_n8509_));
  OAI21X1  g08317(.A0(new_n8509_), .A1(new_n6294_), .B0(new_n5941_), .Y(new_n8510_));
  OAI21X1  g08318(.A0(new_n8510_), .A1(new_n8499_), .B0(new_n8506_), .Y(new_n8511_));
  AOI21X1  g08319(.A0(new_n8511_), .A1(new_n8500_), .B0(new_n5541_), .Y(new_n8512_));
  AND2X1   g08320(.A(new_n8079_), .B(new_n8077_), .Y(new_n8513_));
  NOR3X1   g08321(.A(new_n8513_), .B(new_n8045_), .C(new_n8078_), .Y(new_n8514_));
  NOR3X1   g08322(.A(new_n8412_), .B(new_n8513_), .C(new_n8078_), .Y(new_n8515_));
  NOR2X1   g08323(.A(new_n8515_), .B(new_n8044_), .Y(new_n8516_));
  AOI21X1  g08324(.A0(new_n8514_), .A1(\asqrt[28] ), .B0(new_n8516_), .Y(new_n8517_));
  INVX1    g08325(.A(new_n8517_), .Y(new_n8518_));
  NAND3X1  g08326(.A(new_n8511_), .B(new_n8500_), .C(new_n5541_), .Y(new_n8519_));
  AOI21X1  g08327(.A0(new_n8519_), .A1(new_n8518_), .B0(new_n8512_), .Y(new_n8520_));
  OR2X1    g08328(.A(new_n8520_), .B(new_n5176_), .Y(new_n8521_));
  OR2X1    g08329(.A(new_n8509_), .B(new_n6294_), .Y(new_n8522_));
  NOR2X1   g08330(.A(new_n8479_), .B(new_n8478_), .Y(new_n8523_));
  INVX1    g08331(.A(new_n8487_), .Y(new_n8524_));
  OR2X1    g08332(.A(new_n8497_), .B(\asqrt[33] ), .Y(new_n8525_));
  OAI21X1  g08333(.A0(new_n8525_), .A1(new_n8523_), .B0(new_n8524_), .Y(new_n8526_));
  AOI21X1  g08334(.A0(new_n8526_), .A1(new_n8522_), .B0(new_n5941_), .Y(new_n8527_));
  AOI21X1  g08335(.A0(new_n8480_), .A1(\asqrt[33] ), .B0(\asqrt[34] ), .Y(new_n8528_));
  AOI21X1  g08336(.A0(new_n8528_), .A1(new_n8526_), .B0(new_n8505_), .Y(new_n8529_));
  NOR3X1   g08337(.A(new_n8529_), .B(new_n8527_), .C(\asqrt[35] ), .Y(new_n8530_));
  NOR2X1   g08338(.A(new_n8530_), .B(new_n8517_), .Y(new_n8531_));
  NAND4X1  g08339(.A(\asqrt[28] ), .B(new_n8055_), .C(new_n8053_), .D(new_n8081_), .Y(new_n8532_));
  NAND2X1  g08340(.A(new_n8055_), .B(new_n8081_), .Y(new_n8533_));
  OAI21X1  g08341(.A0(new_n8533_), .A1(new_n8412_), .B0(new_n8054_), .Y(new_n8534_));
  AND2X1   g08342(.A(new_n8534_), .B(new_n8532_), .Y(new_n8535_));
  INVX1    g08343(.A(new_n8535_), .Y(new_n8536_));
  OAI21X1  g08344(.A0(new_n8529_), .A1(new_n8527_), .B0(\asqrt[35] ), .Y(new_n8537_));
  NAND2X1  g08345(.A(new_n8537_), .B(new_n5176_), .Y(new_n8538_));
  OAI21X1  g08346(.A0(new_n8538_), .A1(new_n8531_), .B0(new_n8536_), .Y(new_n8539_));
  AOI21X1  g08347(.A0(new_n8539_), .A1(new_n8521_), .B0(new_n4826_), .Y(new_n8540_));
  OAI21X1  g08348(.A0(new_n8530_), .A1(new_n8517_), .B0(new_n8537_), .Y(new_n8541_));
  AOI21X1  g08349(.A0(new_n8541_), .A1(\asqrt[36] ), .B0(\asqrt[37] ), .Y(new_n8542_));
  AND2X1   g08350(.A(new_n8097_), .B(new_n8096_), .Y(new_n8543_));
  NOR3X1   g08351(.A(new_n8065_), .B(new_n8543_), .C(new_n8095_), .Y(new_n8544_));
  NOR3X1   g08352(.A(new_n8412_), .B(new_n8543_), .C(new_n8095_), .Y(new_n8545_));
  NOR2X1   g08353(.A(new_n8545_), .B(new_n8064_), .Y(new_n8546_));
  AOI21X1  g08354(.A0(new_n8544_), .A1(\asqrt[28] ), .B0(new_n8546_), .Y(new_n8547_));
  AOI21X1  g08355(.A0(new_n8542_), .A1(new_n8539_), .B0(new_n8547_), .Y(new_n8548_));
  OAI21X1  g08356(.A0(new_n8548_), .A1(new_n8540_), .B0(\asqrt[38] ), .Y(new_n8549_));
  AND2X1   g08357(.A(new_n8084_), .B(new_n8066_), .Y(new_n8550_));
  NOR3X1   g08358(.A(new_n8550_), .B(new_n8100_), .C(new_n8067_), .Y(new_n8551_));
  NOR3X1   g08359(.A(new_n8412_), .B(new_n8550_), .C(new_n8067_), .Y(new_n8552_));
  NOR2X1   g08360(.A(new_n8552_), .B(new_n8072_), .Y(new_n8553_));
  AOI21X1  g08361(.A0(new_n8551_), .A1(\asqrt[28] ), .B0(new_n8553_), .Y(new_n8554_));
  NOR3X1   g08362(.A(new_n8548_), .B(new_n8540_), .C(\asqrt[38] ), .Y(new_n8555_));
  OAI21X1  g08363(.A0(new_n8555_), .A1(new_n8554_), .B0(new_n8549_), .Y(new_n8556_));
  AND2X1   g08364(.A(new_n8556_), .B(\asqrt[39] ), .Y(new_n8557_));
  OR2X1    g08365(.A(new_n8555_), .B(new_n8554_), .Y(new_n8558_));
  NAND4X1  g08366(.A(\asqrt[28] ), .B(new_n8103_), .C(new_n8090_), .D(new_n8086_), .Y(new_n8559_));
  NAND2X1  g08367(.A(new_n8103_), .B(new_n8086_), .Y(new_n8560_));
  OAI21X1  g08368(.A0(new_n8560_), .A1(new_n8412_), .B0(new_n8094_), .Y(new_n8561_));
  AND2X1   g08369(.A(new_n8561_), .B(new_n8559_), .Y(new_n8562_));
  AND2X1   g08370(.A(new_n8549_), .B(new_n4165_), .Y(new_n8563_));
  AOI21X1  g08371(.A0(new_n8563_), .A1(new_n8558_), .B0(new_n8562_), .Y(new_n8564_));
  OAI21X1  g08372(.A0(new_n8564_), .A1(new_n8557_), .B0(\asqrt[40] ), .Y(new_n8565_));
  AOI21X1  g08373(.A0(new_n8111_), .A1(new_n8104_), .B0(new_n8149_), .Y(new_n8566_));
  AND2X1   g08374(.A(new_n8566_), .B(new_n8147_), .Y(new_n8567_));
  AOI22X1  g08375(.A0(new_n8111_), .A1(new_n8104_), .B0(new_n8092_), .B1(\asqrt[39] ), .Y(new_n8568_));
  AOI21X1  g08376(.A0(new_n8568_), .A1(\asqrt[28] ), .B0(new_n8109_), .Y(new_n8569_));
  AOI21X1  g08377(.A0(new_n8567_), .A1(\asqrt[28] ), .B0(new_n8569_), .Y(new_n8570_));
  INVX1    g08378(.A(new_n8570_), .Y(new_n8571_));
  AND2X1   g08379(.A(new_n8541_), .B(\asqrt[36] ), .Y(new_n8572_));
  OR2X1    g08380(.A(new_n8530_), .B(new_n8517_), .Y(new_n8573_));
  AND2X1   g08381(.A(new_n8537_), .B(new_n5176_), .Y(new_n8574_));
  AOI21X1  g08382(.A0(new_n8574_), .A1(new_n8573_), .B0(new_n8535_), .Y(new_n8575_));
  OAI21X1  g08383(.A0(new_n8575_), .A1(new_n8572_), .B0(\asqrt[37] ), .Y(new_n8576_));
  OAI21X1  g08384(.A0(new_n8520_), .A1(new_n5176_), .B0(new_n4826_), .Y(new_n8577_));
  INVX1    g08385(.A(new_n8547_), .Y(new_n8578_));
  OAI21X1  g08386(.A0(new_n8577_), .A1(new_n8575_), .B0(new_n8578_), .Y(new_n8579_));
  AOI21X1  g08387(.A0(new_n8579_), .A1(new_n8576_), .B0(new_n4493_), .Y(new_n8580_));
  INVX1    g08388(.A(new_n8554_), .Y(new_n8581_));
  NAND3X1  g08389(.A(new_n8579_), .B(new_n8576_), .C(new_n4493_), .Y(new_n8582_));
  AOI21X1  g08390(.A0(new_n8582_), .A1(new_n8581_), .B0(new_n8580_), .Y(new_n8583_));
  OAI21X1  g08391(.A0(new_n8583_), .A1(new_n4165_), .B0(new_n3863_), .Y(new_n8584_));
  OAI21X1  g08392(.A0(new_n8584_), .A1(new_n8564_), .B0(new_n8571_), .Y(new_n8585_));
  AOI21X1  g08393(.A0(new_n8585_), .A1(new_n8565_), .B0(new_n3564_), .Y(new_n8586_));
  AND2X1   g08394(.A(new_n8153_), .B(new_n8151_), .Y(new_n8587_));
  NOR3X1   g08395(.A(new_n8587_), .B(new_n8119_), .C(new_n8152_), .Y(new_n8588_));
  NOR3X1   g08396(.A(new_n8412_), .B(new_n8587_), .C(new_n8152_), .Y(new_n8589_));
  NOR2X1   g08397(.A(new_n8589_), .B(new_n8118_), .Y(new_n8590_));
  AOI21X1  g08398(.A0(new_n8588_), .A1(\asqrt[28] ), .B0(new_n8590_), .Y(new_n8591_));
  INVX1    g08399(.A(new_n8591_), .Y(new_n8592_));
  NAND3X1  g08400(.A(new_n8585_), .B(new_n8565_), .C(new_n3564_), .Y(new_n8593_));
  AOI21X1  g08401(.A0(new_n8593_), .A1(new_n8592_), .B0(new_n8586_), .Y(new_n8594_));
  OR2X1    g08402(.A(new_n8594_), .B(new_n3276_), .Y(new_n8595_));
  AND2X1   g08403(.A(new_n8593_), .B(new_n8592_), .Y(new_n8596_));
  NAND4X1  g08404(.A(\asqrt[28] ), .B(new_n8129_), .C(new_n8127_), .D(new_n8155_), .Y(new_n8597_));
  NAND2X1  g08405(.A(new_n8129_), .B(new_n8155_), .Y(new_n8598_));
  OAI21X1  g08406(.A0(new_n8598_), .A1(new_n8412_), .B0(new_n8128_), .Y(new_n8599_));
  AND2X1   g08407(.A(new_n8599_), .B(new_n8597_), .Y(new_n8600_));
  INVX1    g08408(.A(new_n8600_), .Y(new_n8601_));
  OR2X1    g08409(.A(new_n8586_), .B(\asqrt[42] ), .Y(new_n8602_));
  OAI21X1  g08410(.A0(new_n8602_), .A1(new_n8596_), .B0(new_n8601_), .Y(new_n8603_));
  AOI21X1  g08411(.A0(new_n8603_), .A1(new_n8595_), .B0(new_n3008_), .Y(new_n8604_));
  AND2X1   g08412(.A(new_n8171_), .B(new_n8170_), .Y(new_n8605_));
  NOR3X1   g08413(.A(new_n8605_), .B(new_n8138_), .C(new_n8169_), .Y(new_n8606_));
  NOR3X1   g08414(.A(new_n8412_), .B(new_n8605_), .C(new_n8169_), .Y(new_n8607_));
  NOR2X1   g08415(.A(new_n8607_), .B(new_n8137_), .Y(new_n8608_));
  AOI21X1  g08416(.A0(new_n8606_), .A1(\asqrt[28] ), .B0(new_n8608_), .Y(new_n8609_));
  OR2X1    g08417(.A(new_n8583_), .B(new_n4165_), .Y(new_n8610_));
  NOR2X1   g08418(.A(new_n8555_), .B(new_n8554_), .Y(new_n8611_));
  INVX1    g08419(.A(new_n8562_), .Y(new_n8612_));
  NAND2X1  g08420(.A(new_n8549_), .B(new_n4165_), .Y(new_n8613_));
  OAI21X1  g08421(.A0(new_n8613_), .A1(new_n8611_), .B0(new_n8612_), .Y(new_n8614_));
  AOI21X1  g08422(.A0(new_n8614_), .A1(new_n8610_), .B0(new_n3863_), .Y(new_n8615_));
  AOI21X1  g08423(.A0(new_n8556_), .A1(\asqrt[39] ), .B0(\asqrt[40] ), .Y(new_n8616_));
  AOI21X1  g08424(.A0(new_n8616_), .A1(new_n8614_), .B0(new_n8570_), .Y(new_n8617_));
  OAI21X1  g08425(.A0(new_n8617_), .A1(new_n8615_), .B0(\asqrt[41] ), .Y(new_n8618_));
  NOR3X1   g08426(.A(new_n8617_), .B(new_n8615_), .C(\asqrt[41] ), .Y(new_n8619_));
  OAI21X1  g08427(.A0(new_n8619_), .A1(new_n8591_), .B0(new_n8618_), .Y(new_n8620_));
  AOI21X1  g08428(.A0(new_n8620_), .A1(\asqrt[42] ), .B0(\asqrt[43] ), .Y(new_n8621_));
  AOI21X1  g08429(.A0(new_n8621_), .A1(new_n8603_), .B0(new_n8609_), .Y(new_n8622_));
  OAI21X1  g08430(.A0(new_n8622_), .A1(new_n8604_), .B0(\asqrt[44] ), .Y(new_n8623_));
  AND2X1   g08431(.A(new_n8158_), .B(new_n8140_), .Y(new_n8624_));
  NOR3X1   g08432(.A(new_n8624_), .B(new_n8174_), .C(new_n8141_), .Y(new_n8625_));
  NOR3X1   g08433(.A(new_n8412_), .B(new_n8624_), .C(new_n8141_), .Y(new_n8626_));
  NOR2X1   g08434(.A(new_n8626_), .B(new_n8146_), .Y(new_n8627_));
  AOI21X1  g08435(.A0(new_n8625_), .A1(\asqrt[28] ), .B0(new_n8627_), .Y(new_n8628_));
  NOR3X1   g08436(.A(new_n8622_), .B(new_n8604_), .C(\asqrt[44] ), .Y(new_n8629_));
  OAI21X1  g08437(.A0(new_n8629_), .A1(new_n8628_), .B0(new_n8623_), .Y(new_n8630_));
  AND2X1   g08438(.A(new_n8630_), .B(\asqrt[45] ), .Y(new_n8631_));
  INVX1    g08439(.A(new_n8628_), .Y(new_n8632_));
  AND2X1   g08440(.A(new_n8620_), .B(\asqrt[42] ), .Y(new_n8633_));
  NAND2X1  g08441(.A(new_n8593_), .B(new_n8592_), .Y(new_n8634_));
  NOR2X1   g08442(.A(new_n8586_), .B(\asqrt[42] ), .Y(new_n8635_));
  AOI21X1  g08443(.A0(new_n8635_), .A1(new_n8634_), .B0(new_n8600_), .Y(new_n8636_));
  OAI21X1  g08444(.A0(new_n8636_), .A1(new_n8633_), .B0(\asqrt[43] ), .Y(new_n8637_));
  INVX1    g08445(.A(new_n8609_), .Y(new_n8638_));
  OAI21X1  g08446(.A0(new_n8594_), .A1(new_n3276_), .B0(new_n3008_), .Y(new_n8639_));
  OAI21X1  g08447(.A0(new_n8639_), .A1(new_n8636_), .B0(new_n8638_), .Y(new_n8640_));
  NAND3X1  g08448(.A(new_n8640_), .B(new_n8637_), .C(new_n2769_), .Y(new_n8641_));
  NAND2X1  g08449(.A(new_n8641_), .B(new_n8632_), .Y(new_n8642_));
  NAND4X1  g08450(.A(\asqrt[28] ), .B(new_n8177_), .C(new_n8164_), .D(new_n8160_), .Y(new_n8643_));
  NAND2X1  g08451(.A(new_n8177_), .B(new_n8160_), .Y(new_n8644_));
  OAI21X1  g08452(.A0(new_n8644_), .A1(new_n8412_), .B0(new_n8168_), .Y(new_n8645_));
  AND2X1   g08453(.A(new_n8645_), .B(new_n8643_), .Y(new_n8646_));
  AOI21X1  g08454(.A0(new_n8640_), .A1(new_n8637_), .B0(new_n2769_), .Y(new_n8647_));
  NOR2X1   g08455(.A(new_n8647_), .B(\asqrt[45] ), .Y(new_n8648_));
  AOI21X1  g08456(.A0(new_n8648_), .A1(new_n8642_), .B0(new_n8646_), .Y(new_n8649_));
  OAI21X1  g08457(.A0(new_n8649_), .A1(new_n8631_), .B0(\asqrt[46] ), .Y(new_n8650_));
  AOI21X1  g08458(.A0(new_n8185_), .A1(new_n8178_), .B0(new_n8221_), .Y(new_n8651_));
  AND2X1   g08459(.A(new_n8651_), .B(new_n8219_), .Y(new_n8652_));
  AOI22X1  g08460(.A0(new_n8185_), .A1(new_n8178_), .B0(new_n8166_), .B1(\asqrt[45] ), .Y(new_n8653_));
  AOI21X1  g08461(.A0(new_n8653_), .A1(\asqrt[28] ), .B0(new_n8183_), .Y(new_n8654_));
  AOI21X1  g08462(.A0(new_n8652_), .A1(\asqrt[28] ), .B0(new_n8654_), .Y(new_n8655_));
  INVX1    g08463(.A(new_n8655_), .Y(new_n8656_));
  AOI21X1  g08464(.A0(new_n8641_), .A1(new_n8632_), .B0(new_n8647_), .Y(new_n8657_));
  OAI21X1  g08465(.A0(new_n8657_), .A1(new_n2570_), .B0(new_n2263_), .Y(new_n8658_));
  OAI21X1  g08466(.A0(new_n8658_), .A1(new_n8649_), .B0(new_n8656_), .Y(new_n8659_));
  AOI21X1  g08467(.A0(new_n8659_), .A1(new_n8650_), .B0(new_n2040_), .Y(new_n8660_));
  AND2X1   g08468(.A(new_n8225_), .B(new_n8223_), .Y(new_n8661_));
  NOR3X1   g08469(.A(new_n8661_), .B(new_n8193_), .C(new_n8224_), .Y(new_n8662_));
  NOR3X1   g08470(.A(new_n8412_), .B(new_n8661_), .C(new_n8224_), .Y(new_n8663_));
  NOR2X1   g08471(.A(new_n8663_), .B(new_n8192_), .Y(new_n8664_));
  AOI21X1  g08472(.A0(new_n8662_), .A1(\asqrt[28] ), .B0(new_n8664_), .Y(new_n8665_));
  INVX1    g08473(.A(new_n8665_), .Y(new_n8666_));
  NAND3X1  g08474(.A(new_n8659_), .B(new_n8650_), .C(new_n2040_), .Y(new_n8667_));
  AOI21X1  g08475(.A0(new_n8667_), .A1(new_n8666_), .B0(new_n8660_), .Y(new_n8668_));
  OR2X1    g08476(.A(new_n8668_), .B(new_n1834_), .Y(new_n8669_));
  AND2X1   g08477(.A(new_n8667_), .B(new_n8666_), .Y(new_n8670_));
  OR4X1    g08478(.A(new_n8412_), .B(new_n8229_), .C(new_n8200_), .D(new_n8197_), .Y(new_n8671_));
  NAND2X1  g08479(.A(new_n8201_), .B(new_n8227_), .Y(new_n8672_));
  OAI21X1  g08480(.A0(new_n8672_), .A1(new_n8412_), .B0(new_n8200_), .Y(new_n8673_));
  AND2X1   g08481(.A(new_n8673_), .B(new_n8671_), .Y(new_n8674_));
  INVX1    g08482(.A(new_n8674_), .Y(new_n8675_));
  OR2X1    g08483(.A(new_n8660_), .B(\asqrt[48] ), .Y(new_n8676_));
  OAI21X1  g08484(.A0(new_n8676_), .A1(new_n8670_), .B0(new_n8675_), .Y(new_n8677_));
  AOI21X1  g08485(.A0(new_n8677_), .A1(new_n8669_), .B0(new_n1632_), .Y(new_n8678_));
  AND2X1   g08486(.A(new_n8244_), .B(new_n8243_), .Y(new_n8679_));
  NOR3X1   g08487(.A(new_n8679_), .B(new_n8210_), .C(new_n8242_), .Y(new_n8680_));
  NOR3X1   g08488(.A(new_n8412_), .B(new_n8679_), .C(new_n8242_), .Y(new_n8681_));
  NOR2X1   g08489(.A(new_n8681_), .B(new_n8209_), .Y(new_n8682_));
  AOI21X1  g08490(.A0(new_n8680_), .A1(\asqrt[28] ), .B0(new_n8682_), .Y(new_n8683_));
  OR2X1    g08491(.A(new_n8657_), .B(new_n2570_), .Y(new_n8684_));
  AND2X1   g08492(.A(new_n8641_), .B(new_n8632_), .Y(new_n8685_));
  INVX1    g08493(.A(new_n8646_), .Y(new_n8686_));
  OR2X1    g08494(.A(new_n8647_), .B(\asqrt[45] ), .Y(new_n8687_));
  OAI21X1  g08495(.A0(new_n8687_), .A1(new_n8685_), .B0(new_n8686_), .Y(new_n8688_));
  AOI21X1  g08496(.A0(new_n8688_), .A1(new_n8684_), .B0(new_n2263_), .Y(new_n8689_));
  AOI21X1  g08497(.A0(new_n8630_), .A1(\asqrt[45] ), .B0(\asqrt[46] ), .Y(new_n8690_));
  AOI21X1  g08498(.A0(new_n8690_), .A1(new_n8688_), .B0(new_n8655_), .Y(new_n8691_));
  OAI21X1  g08499(.A0(new_n8691_), .A1(new_n8689_), .B0(\asqrt[47] ), .Y(new_n8692_));
  NOR3X1   g08500(.A(new_n8691_), .B(new_n8689_), .C(\asqrt[47] ), .Y(new_n8693_));
  OAI21X1  g08501(.A0(new_n8693_), .A1(new_n8665_), .B0(new_n8692_), .Y(new_n8694_));
  AOI21X1  g08502(.A0(new_n8694_), .A1(\asqrt[48] ), .B0(\asqrt[49] ), .Y(new_n8695_));
  AOI21X1  g08503(.A0(new_n8695_), .A1(new_n8677_), .B0(new_n8683_), .Y(new_n8696_));
  OAI21X1  g08504(.A0(new_n8696_), .A1(new_n8678_), .B0(\asqrt[50] ), .Y(new_n8697_));
  AND2X1   g08505(.A(new_n8231_), .B(new_n8212_), .Y(new_n8698_));
  NOR3X1   g08506(.A(new_n8698_), .B(new_n8247_), .C(new_n8213_), .Y(new_n8699_));
  NOR3X1   g08507(.A(new_n8412_), .B(new_n8698_), .C(new_n8213_), .Y(new_n8700_));
  NOR2X1   g08508(.A(new_n8700_), .B(new_n8218_), .Y(new_n8701_));
  AOI21X1  g08509(.A0(new_n8699_), .A1(\asqrt[28] ), .B0(new_n8701_), .Y(new_n8702_));
  NOR3X1   g08510(.A(new_n8696_), .B(new_n8678_), .C(\asqrt[50] ), .Y(new_n8703_));
  OAI21X1  g08511(.A0(new_n8703_), .A1(new_n8702_), .B0(new_n8697_), .Y(new_n8704_));
  AND2X1   g08512(.A(new_n8704_), .B(\asqrt[51] ), .Y(new_n8705_));
  INVX1    g08513(.A(new_n8702_), .Y(new_n8706_));
  AND2X1   g08514(.A(new_n8694_), .B(\asqrt[48] ), .Y(new_n8707_));
  NAND2X1  g08515(.A(new_n8667_), .B(new_n8666_), .Y(new_n8708_));
  NOR2X1   g08516(.A(new_n8660_), .B(\asqrt[48] ), .Y(new_n8709_));
  AOI21X1  g08517(.A0(new_n8709_), .A1(new_n8708_), .B0(new_n8674_), .Y(new_n8710_));
  OAI21X1  g08518(.A0(new_n8710_), .A1(new_n8707_), .B0(\asqrt[49] ), .Y(new_n8711_));
  INVX1    g08519(.A(new_n8683_), .Y(new_n8712_));
  OAI21X1  g08520(.A0(new_n8668_), .A1(new_n1834_), .B0(new_n1632_), .Y(new_n8713_));
  OAI21X1  g08521(.A0(new_n8713_), .A1(new_n8710_), .B0(new_n8712_), .Y(new_n8714_));
  NAND3X1  g08522(.A(new_n8714_), .B(new_n8711_), .C(new_n1469_), .Y(new_n8715_));
  NAND2X1  g08523(.A(new_n8715_), .B(new_n8706_), .Y(new_n8716_));
  NAND4X1  g08524(.A(\asqrt[28] ), .B(new_n8250_), .C(new_n8237_), .D(new_n8233_), .Y(new_n8717_));
  NAND2X1  g08525(.A(new_n8250_), .B(new_n8233_), .Y(new_n8718_));
  OAI21X1  g08526(.A0(new_n8718_), .A1(new_n8412_), .B0(new_n8241_), .Y(new_n8719_));
  AND2X1   g08527(.A(new_n8719_), .B(new_n8717_), .Y(new_n8720_));
  AOI21X1  g08528(.A0(new_n8714_), .A1(new_n8711_), .B0(new_n1469_), .Y(new_n8721_));
  NOR2X1   g08529(.A(new_n8721_), .B(\asqrt[51] ), .Y(new_n8722_));
  AOI21X1  g08530(.A0(new_n8722_), .A1(new_n8716_), .B0(new_n8720_), .Y(new_n8723_));
  OAI21X1  g08531(.A0(new_n8723_), .A1(new_n8705_), .B0(\asqrt[52] ), .Y(new_n8724_));
  AOI21X1  g08532(.A0(new_n8258_), .A1(new_n8251_), .B0(new_n8281_), .Y(new_n8725_));
  AND2X1   g08533(.A(new_n8725_), .B(new_n8279_), .Y(new_n8726_));
  AOI22X1  g08534(.A0(new_n8258_), .A1(new_n8251_), .B0(new_n8239_), .B1(\asqrt[51] ), .Y(new_n8727_));
  AOI21X1  g08535(.A0(new_n8727_), .A1(\asqrt[28] ), .B0(new_n8256_), .Y(new_n8728_));
  AOI21X1  g08536(.A0(new_n8726_), .A1(\asqrt[28] ), .B0(new_n8728_), .Y(new_n8729_));
  INVX1    g08537(.A(new_n8729_), .Y(new_n8730_));
  AOI21X1  g08538(.A0(new_n8715_), .A1(new_n8706_), .B0(new_n8721_), .Y(new_n8731_));
  OAI21X1  g08539(.A0(new_n8731_), .A1(new_n1277_), .B0(new_n1111_), .Y(new_n8732_));
  OAI21X1  g08540(.A0(new_n8732_), .A1(new_n8723_), .B0(new_n8730_), .Y(new_n8733_));
  AOI21X1  g08541(.A0(new_n8733_), .A1(new_n8724_), .B0(new_n968_), .Y(new_n8734_));
  AND2X1   g08542(.A(new_n8285_), .B(new_n8283_), .Y(new_n8735_));
  NOR3X1   g08543(.A(new_n8735_), .B(new_n8266_), .C(new_n8284_), .Y(new_n8736_));
  NOR3X1   g08544(.A(new_n8412_), .B(new_n8735_), .C(new_n8284_), .Y(new_n8737_));
  NOR2X1   g08545(.A(new_n8737_), .B(new_n8265_), .Y(new_n8738_));
  AOI21X1  g08546(.A0(new_n8736_), .A1(\asqrt[28] ), .B0(new_n8738_), .Y(new_n8739_));
  INVX1    g08547(.A(new_n8739_), .Y(new_n8740_));
  NAND3X1  g08548(.A(new_n8733_), .B(new_n8724_), .C(new_n968_), .Y(new_n8741_));
  AOI21X1  g08549(.A0(new_n8741_), .A1(new_n8740_), .B0(new_n8734_), .Y(new_n8742_));
  OR2X1    g08550(.A(new_n8742_), .B(new_n902_), .Y(new_n8743_));
  OR2X1    g08551(.A(new_n8731_), .B(new_n1277_), .Y(new_n8744_));
  AND2X1   g08552(.A(new_n8715_), .B(new_n8706_), .Y(new_n8745_));
  INVX1    g08553(.A(new_n8720_), .Y(new_n8746_));
  OR2X1    g08554(.A(new_n8721_), .B(\asqrt[51] ), .Y(new_n8747_));
  OAI21X1  g08555(.A0(new_n8747_), .A1(new_n8745_), .B0(new_n8746_), .Y(new_n8748_));
  AOI21X1  g08556(.A0(new_n8748_), .A1(new_n8744_), .B0(new_n1111_), .Y(new_n8749_));
  AOI21X1  g08557(.A0(new_n8704_), .A1(\asqrt[51] ), .B0(\asqrt[52] ), .Y(new_n8750_));
  AOI21X1  g08558(.A0(new_n8750_), .A1(new_n8748_), .B0(new_n8729_), .Y(new_n8751_));
  NOR3X1   g08559(.A(new_n8751_), .B(new_n8749_), .C(\asqrt[53] ), .Y(new_n8752_));
  NOR2X1   g08560(.A(new_n8752_), .B(new_n8739_), .Y(new_n8753_));
  OR4X1    g08561(.A(new_n8412_), .B(new_n8287_), .C(new_n8275_), .D(new_n8270_), .Y(new_n8754_));
  OR2X1    g08562(.A(new_n8287_), .B(new_n8270_), .Y(new_n8755_));
  OAI21X1  g08563(.A0(new_n8755_), .A1(new_n8412_), .B0(new_n8275_), .Y(new_n8756_));
  AND2X1   g08564(.A(new_n8756_), .B(new_n8754_), .Y(new_n8757_));
  INVX1    g08565(.A(new_n8757_), .Y(new_n8758_));
  OAI21X1  g08566(.A0(new_n8751_), .A1(new_n8749_), .B0(\asqrt[53] ), .Y(new_n8759_));
  NAND2X1  g08567(.A(new_n8759_), .B(new_n902_), .Y(new_n8760_));
  OAI21X1  g08568(.A0(new_n8760_), .A1(new_n8753_), .B0(new_n8758_), .Y(new_n8761_));
  AOI21X1  g08569(.A0(new_n8761_), .A1(new_n8743_), .B0(new_n697_), .Y(new_n8762_));
  AND2X1   g08570(.A(new_n8317_), .B(new_n8316_), .Y(new_n8763_));
  NOR3X1   g08571(.A(new_n8763_), .B(new_n8294_), .C(new_n8315_), .Y(new_n8764_));
  NOR3X1   g08572(.A(new_n8412_), .B(new_n8763_), .C(new_n8315_), .Y(new_n8765_));
  NOR2X1   g08573(.A(new_n8765_), .B(new_n8293_), .Y(new_n8766_));
  AOI21X1  g08574(.A0(new_n8764_), .A1(\asqrt[28] ), .B0(new_n8766_), .Y(new_n8767_));
  OAI21X1  g08575(.A0(new_n8752_), .A1(new_n8739_), .B0(new_n8759_), .Y(new_n8768_));
  AOI21X1  g08576(.A0(new_n8768_), .A1(\asqrt[54] ), .B0(\asqrt[55] ), .Y(new_n8769_));
  AOI21X1  g08577(.A0(new_n8769_), .A1(new_n8761_), .B0(new_n8767_), .Y(new_n8770_));
  OAI21X1  g08578(.A0(new_n8770_), .A1(new_n8762_), .B0(\asqrt[56] ), .Y(new_n8771_));
  AND2X1   g08579(.A(new_n8305_), .B(new_n8297_), .Y(new_n8772_));
  NOR3X1   g08580(.A(new_n8772_), .B(new_n8320_), .C(new_n8298_), .Y(new_n8773_));
  NOR3X1   g08581(.A(new_n8412_), .B(new_n8772_), .C(new_n8298_), .Y(new_n8774_));
  NOR2X1   g08582(.A(new_n8774_), .B(new_n8303_), .Y(new_n8775_));
  AOI21X1  g08583(.A0(new_n8773_), .A1(\asqrt[28] ), .B0(new_n8775_), .Y(new_n8776_));
  NOR3X1   g08584(.A(new_n8770_), .B(new_n8762_), .C(\asqrt[56] ), .Y(new_n8777_));
  OAI21X1  g08585(.A0(new_n8777_), .A1(new_n8776_), .B0(new_n8771_), .Y(new_n8778_));
  AND2X1   g08586(.A(new_n8778_), .B(\asqrt[57] ), .Y(new_n8779_));
  OR2X1    g08587(.A(new_n8777_), .B(new_n8776_), .Y(new_n8780_));
  OR4X1    g08588(.A(new_n8412_), .B(new_n8312_), .C(new_n8310_), .D(new_n8339_), .Y(new_n8781_));
  OR2X1    g08589(.A(new_n8312_), .B(new_n8339_), .Y(new_n8782_));
  OAI21X1  g08590(.A0(new_n8782_), .A1(new_n8412_), .B0(new_n8310_), .Y(new_n8783_));
  AND2X1   g08591(.A(new_n8783_), .B(new_n8781_), .Y(new_n8784_));
  AND2X1   g08592(.A(new_n8771_), .B(new_n481_), .Y(new_n8785_));
  AOI21X1  g08593(.A0(new_n8785_), .A1(new_n8780_), .B0(new_n8784_), .Y(new_n8786_));
  OAI21X1  g08594(.A0(new_n8786_), .A1(new_n8779_), .B0(\asqrt[58] ), .Y(new_n8787_));
  AOI21X1  g08595(.A0(new_n8330_), .A1(new_n8324_), .B0(new_n8354_), .Y(new_n8788_));
  AND2X1   g08596(.A(new_n8788_), .B(new_n8352_), .Y(new_n8789_));
  AOI22X1  g08597(.A0(new_n8330_), .A1(new_n8324_), .B0(new_n8313_), .B1(\asqrt[57] ), .Y(new_n8790_));
  AOI21X1  g08598(.A0(new_n8790_), .A1(\asqrt[28] ), .B0(new_n8329_), .Y(new_n8791_));
  AOI21X1  g08599(.A0(new_n8789_), .A1(\asqrt[28] ), .B0(new_n8791_), .Y(new_n8792_));
  INVX1    g08600(.A(new_n8792_), .Y(new_n8793_));
  AND2X1   g08601(.A(new_n8768_), .B(\asqrt[54] ), .Y(new_n8794_));
  OR2X1    g08602(.A(new_n8752_), .B(new_n8739_), .Y(new_n8795_));
  AND2X1   g08603(.A(new_n8759_), .B(new_n902_), .Y(new_n8796_));
  AOI21X1  g08604(.A0(new_n8796_), .A1(new_n8795_), .B0(new_n8757_), .Y(new_n8797_));
  OAI21X1  g08605(.A0(new_n8797_), .A1(new_n8794_), .B0(\asqrt[55] ), .Y(new_n8798_));
  INVX1    g08606(.A(new_n8767_), .Y(new_n8799_));
  OAI21X1  g08607(.A0(new_n8742_), .A1(new_n902_), .B0(new_n697_), .Y(new_n8800_));
  OAI21X1  g08608(.A0(new_n8800_), .A1(new_n8797_), .B0(new_n8799_), .Y(new_n8801_));
  AOI21X1  g08609(.A0(new_n8801_), .A1(new_n8798_), .B0(new_n582_), .Y(new_n8802_));
  INVX1    g08610(.A(new_n8776_), .Y(new_n8803_));
  NAND3X1  g08611(.A(new_n8801_), .B(new_n8798_), .C(new_n582_), .Y(new_n8804_));
  AOI21X1  g08612(.A0(new_n8804_), .A1(new_n8803_), .B0(new_n8802_), .Y(new_n8805_));
  OAI21X1  g08613(.A0(new_n8805_), .A1(new_n481_), .B0(new_n399_), .Y(new_n8806_));
  OAI21X1  g08614(.A0(new_n8806_), .A1(new_n8786_), .B0(new_n8793_), .Y(new_n8807_));
  AOI21X1  g08615(.A0(new_n8807_), .A1(new_n8787_), .B0(new_n328_), .Y(new_n8808_));
  AND2X1   g08616(.A(new_n8358_), .B(new_n8356_), .Y(new_n8809_));
  NOR3X1   g08617(.A(new_n8809_), .B(new_n8338_), .C(new_n8357_), .Y(new_n8810_));
  NOR3X1   g08618(.A(new_n8412_), .B(new_n8809_), .C(new_n8357_), .Y(new_n8811_));
  NOR2X1   g08619(.A(new_n8811_), .B(new_n8337_), .Y(new_n8812_));
  AOI21X1  g08620(.A0(new_n8810_), .A1(\asqrt[28] ), .B0(new_n8812_), .Y(new_n8813_));
  INVX1    g08621(.A(new_n8813_), .Y(new_n8814_));
  NAND3X1  g08622(.A(new_n8807_), .B(new_n8787_), .C(new_n328_), .Y(new_n8815_));
  AOI21X1  g08623(.A0(new_n8815_), .A1(new_n8814_), .B0(new_n8808_), .Y(new_n8816_));
  OR2X1    g08624(.A(new_n8816_), .B(new_n292_), .Y(new_n8817_));
  OR2X1    g08625(.A(new_n8805_), .B(new_n481_), .Y(new_n8818_));
  NOR2X1   g08626(.A(new_n8777_), .B(new_n8776_), .Y(new_n8819_));
  INVX1    g08627(.A(new_n8784_), .Y(new_n8820_));
  NAND2X1  g08628(.A(new_n8771_), .B(new_n481_), .Y(new_n8821_));
  OAI21X1  g08629(.A0(new_n8821_), .A1(new_n8819_), .B0(new_n8820_), .Y(new_n8822_));
  AOI21X1  g08630(.A0(new_n8822_), .A1(new_n8818_), .B0(new_n399_), .Y(new_n8823_));
  AOI21X1  g08631(.A0(new_n8778_), .A1(\asqrt[57] ), .B0(\asqrt[58] ), .Y(new_n8824_));
  AOI21X1  g08632(.A0(new_n8824_), .A1(new_n8822_), .B0(new_n8792_), .Y(new_n8825_));
  NOR3X1   g08633(.A(new_n8825_), .B(new_n8823_), .C(\asqrt[59] ), .Y(new_n8826_));
  NOR2X1   g08634(.A(new_n8826_), .B(new_n8813_), .Y(new_n8827_));
  OR4X1    g08635(.A(new_n8412_), .B(new_n8360_), .C(new_n8348_), .D(new_n8343_), .Y(new_n8828_));
  OR2X1    g08636(.A(new_n8360_), .B(new_n8343_), .Y(new_n8829_));
  OAI21X1  g08637(.A0(new_n8829_), .A1(new_n8412_), .B0(new_n8348_), .Y(new_n8830_));
  AND2X1   g08638(.A(new_n8830_), .B(new_n8828_), .Y(new_n8831_));
  INVX1    g08639(.A(new_n8831_), .Y(new_n8832_));
  OAI21X1  g08640(.A0(new_n8825_), .A1(new_n8823_), .B0(\asqrt[59] ), .Y(new_n8833_));
  NAND2X1  g08641(.A(new_n8833_), .B(new_n292_), .Y(new_n8834_));
  OAI21X1  g08642(.A0(new_n8834_), .A1(new_n8827_), .B0(new_n8832_), .Y(new_n8835_));
  AOI21X1  g08643(.A0(new_n8835_), .A1(new_n8817_), .B0(new_n217_), .Y(new_n8836_));
  AND2X1   g08644(.A(new_n8421_), .B(new_n8420_), .Y(new_n8837_));
  NOR3X1   g08645(.A(new_n8837_), .B(new_n8367_), .C(new_n8419_), .Y(new_n8838_));
  NOR3X1   g08646(.A(new_n8412_), .B(new_n8837_), .C(new_n8419_), .Y(new_n8839_));
  NOR2X1   g08647(.A(new_n8839_), .B(new_n8366_), .Y(new_n8840_));
  AOI21X1  g08648(.A0(new_n8838_), .A1(\asqrt[28] ), .B0(new_n8840_), .Y(new_n8841_));
  OAI21X1  g08649(.A0(new_n8826_), .A1(new_n8813_), .B0(new_n8833_), .Y(new_n8842_));
  AOI21X1  g08650(.A0(new_n8842_), .A1(\asqrt[60] ), .B0(\asqrt[61] ), .Y(new_n8843_));
  AOI21X1  g08651(.A0(new_n8843_), .A1(new_n8835_), .B0(new_n8841_), .Y(new_n8844_));
  OAI21X1  g08652(.A0(new_n8844_), .A1(new_n8836_), .B0(\asqrt[62] ), .Y(new_n8845_));
  AND2X1   g08653(.A(new_n8378_), .B(new_n8370_), .Y(new_n8846_));
  NOR3X1   g08654(.A(new_n8846_), .B(new_n8424_), .C(new_n8371_), .Y(new_n8847_));
  NOR3X1   g08655(.A(new_n8412_), .B(new_n8846_), .C(new_n8371_), .Y(new_n8848_));
  NOR2X1   g08656(.A(new_n8848_), .B(new_n8376_), .Y(new_n8849_));
  AOI21X1  g08657(.A0(new_n8847_), .A1(\asqrt[28] ), .B0(new_n8849_), .Y(new_n8850_));
  NOR3X1   g08658(.A(new_n8844_), .B(new_n8836_), .C(\asqrt[62] ), .Y(new_n8851_));
  OAI21X1  g08659(.A0(new_n8851_), .A1(new_n8850_), .B0(new_n8845_), .Y(new_n8852_));
  NOR4X1   g08660(.A(new_n8412_), .B(new_n8385_), .C(new_n8428_), .D(new_n8427_), .Y(new_n8853_));
  NOR3X1   g08661(.A(new_n8412_), .B(new_n8385_), .C(new_n8427_), .Y(new_n8854_));
  NOR2X1   g08662(.A(new_n8854_), .B(new_n8384_), .Y(new_n8855_));
  NOR2X1   g08663(.A(new_n8855_), .B(new_n8853_), .Y(new_n8856_));
  INVX1    g08664(.A(new_n8856_), .Y(new_n8857_));
  AND2X1   g08665(.A(new_n8393_), .B(new_n8386_), .Y(new_n8858_));
  AOI21X1  g08666(.A0(new_n8858_), .A1(\asqrt[28] ), .B0(new_n8448_), .Y(new_n8859_));
  AND2X1   g08667(.A(new_n8859_), .B(new_n8857_), .Y(new_n8860_));
  AOI21X1  g08668(.A0(new_n8860_), .A1(new_n8852_), .B0(\asqrt[63] ), .Y(new_n8861_));
  NOR2X1   g08669(.A(new_n8851_), .B(new_n8850_), .Y(new_n8862_));
  NAND2X1  g08670(.A(new_n8856_), .B(new_n8845_), .Y(new_n8863_));
  AOI21X1  g08671(.A0(new_n8436_), .A1(new_n8432_), .B0(new_n8392_), .Y(new_n8864_));
  AOI21X1  g08672(.A0(new_n8393_), .A1(new_n8386_), .B0(new_n193_), .Y(new_n8865_));
  OAI21X1  g08673(.A0(new_n8864_), .A1(new_n8386_), .B0(new_n8865_), .Y(new_n8866_));
  INVX1    g08674(.A(new_n8391_), .Y(new_n8867_));
  NOR4X1   g08675(.A(new_n8409_), .B(new_n8403_), .C(new_n8867_), .D(new_n8388_), .Y(new_n8868_));
  OAI21X1  g08676(.A0(new_n8400_), .A1(new_n8399_), .B0(new_n8868_), .Y(new_n8869_));
  NOR2X1   g08677(.A(new_n8869_), .B(new_n8398_), .Y(new_n8870_));
  INVX1    g08678(.A(new_n8870_), .Y(new_n8871_));
  AND2X1   g08679(.A(new_n8871_), .B(new_n8866_), .Y(new_n8872_));
  OAI21X1  g08680(.A0(new_n8863_), .A1(new_n8862_), .B0(new_n8872_), .Y(new_n8873_));
  NOR2X1   g08681(.A(new_n8873_), .B(new_n8861_), .Y(new_n8874_));
  INVX1    g08682(.A(\a[54] ), .Y(new_n8875_));
  AND2X1   g08683(.A(new_n8842_), .B(\asqrt[60] ), .Y(new_n8876_));
  OR2X1    g08684(.A(new_n8826_), .B(new_n8813_), .Y(new_n8877_));
  AND2X1   g08685(.A(new_n8833_), .B(new_n292_), .Y(new_n8878_));
  AOI21X1  g08686(.A0(new_n8878_), .A1(new_n8877_), .B0(new_n8831_), .Y(new_n8879_));
  OAI21X1  g08687(.A0(new_n8879_), .A1(new_n8876_), .B0(\asqrt[61] ), .Y(new_n8880_));
  INVX1    g08688(.A(new_n8841_), .Y(new_n8881_));
  OAI21X1  g08689(.A0(new_n8816_), .A1(new_n292_), .B0(new_n217_), .Y(new_n8882_));
  OAI21X1  g08690(.A0(new_n8882_), .A1(new_n8879_), .B0(new_n8881_), .Y(new_n8883_));
  AOI21X1  g08691(.A0(new_n8883_), .A1(new_n8880_), .B0(new_n199_), .Y(new_n8884_));
  INVX1    g08692(.A(new_n8850_), .Y(new_n8885_));
  NAND3X1  g08693(.A(new_n8883_), .B(new_n8880_), .C(new_n199_), .Y(new_n8886_));
  AOI21X1  g08694(.A0(new_n8886_), .A1(new_n8885_), .B0(new_n8884_), .Y(new_n8887_));
  INVX1    g08695(.A(new_n8860_), .Y(new_n8888_));
  OAI21X1  g08696(.A0(new_n8888_), .A1(new_n8887_), .B0(new_n193_), .Y(new_n8889_));
  OR2X1    g08697(.A(new_n8851_), .B(new_n8850_), .Y(new_n8890_));
  AND2X1   g08698(.A(new_n8856_), .B(new_n8845_), .Y(new_n8891_));
  INVX1    g08699(.A(new_n8872_), .Y(new_n8892_));
  AOI21X1  g08700(.A0(new_n8891_), .A1(new_n8890_), .B0(new_n8892_), .Y(new_n8893_));
  AOI21X1  g08701(.A0(new_n8893_), .A1(new_n8889_), .B0(new_n8875_), .Y(new_n8894_));
  NOR3X1   g08702(.A(\a[54] ), .B(\a[53] ), .C(\a[52] ), .Y(new_n8895_));
  OR2X1    g08703(.A(new_n8895_), .B(new_n8894_), .Y(new_n8896_));
  OR2X1    g08704(.A(new_n8895_), .B(new_n8409_), .Y(new_n8897_));
  NOR4X1   g08705(.A(new_n8897_), .B(new_n8403_), .C(new_n8448_), .D(new_n8398_), .Y(new_n8898_));
  INVX1    g08706(.A(new_n8898_), .Y(new_n8899_));
  OR2X1    g08707(.A(new_n8899_), .B(new_n8894_), .Y(new_n8900_));
  OAI21X1  g08708(.A0(new_n8873_), .A1(new_n8861_), .B0(new_n8875_), .Y(new_n8901_));
  INVX1    g08709(.A(new_n8416_), .Y(new_n8902_));
  AOI21X1  g08710(.A0(new_n8893_), .A1(new_n8889_), .B0(new_n8902_), .Y(new_n8903_));
  AOI21X1  g08711(.A0(new_n8901_), .A1(\a[55] ), .B0(new_n8903_), .Y(new_n8904_));
  AOI22X1  g08712(.A0(new_n8904_), .A1(new_n8900_), .B0(new_n8896_), .B1(\asqrt[28] ), .Y(new_n8905_));
  OR2X1    g08713(.A(new_n8905_), .B(new_n7970_), .Y(new_n8906_));
  AND2X1   g08714(.A(new_n8904_), .B(new_n8900_), .Y(new_n8907_));
  OAI21X1  g08715(.A0(new_n8895_), .A1(new_n8894_), .B0(\asqrt[28] ), .Y(new_n8908_));
  NAND2X1  g08716(.A(new_n8908_), .B(new_n7970_), .Y(new_n8909_));
  OAI21X1  g08717(.A0(new_n8873_), .A1(new_n8861_), .B0(new_n8416_), .Y(new_n8910_));
  INVX1    g08718(.A(new_n8866_), .Y(new_n8911_));
  NOR3X1   g08719(.A(new_n8870_), .B(new_n8911_), .C(new_n8412_), .Y(new_n8912_));
  OAI21X1  g08720(.A0(new_n8863_), .A1(new_n8862_), .B0(new_n8912_), .Y(new_n8913_));
  OR2X1    g08721(.A(new_n8913_), .B(new_n8861_), .Y(new_n8914_));
  AOI21X1  g08722(.A0(new_n8914_), .A1(new_n8910_), .B0(new_n8415_), .Y(new_n8915_));
  OAI21X1  g08723(.A0(new_n8913_), .A1(new_n8861_), .B0(new_n8415_), .Y(new_n8916_));
  NOR2X1   g08724(.A(new_n8916_), .B(new_n8903_), .Y(new_n8917_));
  OR2X1    g08725(.A(new_n8917_), .B(new_n8915_), .Y(new_n8918_));
  OAI21X1  g08726(.A0(new_n8909_), .A1(new_n8907_), .B0(new_n8918_), .Y(new_n8919_));
  AOI21X1  g08727(.A0(new_n8919_), .A1(new_n8906_), .B0(new_n7527_), .Y(new_n8920_));
  NOR3X1   g08728(.A(new_n8442_), .B(new_n8464_), .C(new_n8418_), .Y(new_n8921_));
  OAI21X1  g08729(.A0(new_n8873_), .A1(new_n8861_), .B0(new_n8921_), .Y(new_n8922_));
  NOR2X1   g08730(.A(new_n8464_), .B(new_n8418_), .Y(new_n8923_));
  OAI21X1  g08731(.A0(new_n8873_), .A1(new_n8861_), .B0(new_n8923_), .Y(new_n8924_));
  NAND2X1  g08732(.A(new_n8924_), .B(new_n8442_), .Y(new_n8925_));
  AND2X1   g08733(.A(new_n8925_), .B(new_n8922_), .Y(new_n8926_));
  NOR2X1   g08734(.A(new_n8899_), .B(new_n8894_), .Y(new_n8927_));
  INVX1    g08735(.A(\a[55] ), .Y(new_n8928_));
  AOI21X1  g08736(.A0(new_n8893_), .A1(new_n8889_), .B0(\a[54] ), .Y(new_n8929_));
  OAI21X1  g08737(.A0(new_n8929_), .A1(new_n8928_), .B0(new_n8910_), .Y(new_n8930_));
  OAI21X1  g08738(.A0(new_n8930_), .A1(new_n8927_), .B0(new_n8908_), .Y(new_n8931_));
  AOI21X1  g08739(.A0(new_n8931_), .A1(\asqrt[29] ), .B0(\asqrt[30] ), .Y(new_n8932_));
  AOI21X1  g08740(.A0(new_n8932_), .A1(new_n8919_), .B0(new_n8926_), .Y(new_n8933_));
  OAI21X1  g08741(.A0(new_n8933_), .A1(new_n8920_), .B0(\asqrt[31] ), .Y(new_n8934_));
  AOI21X1  g08742(.A0(new_n8490_), .A1(new_n8489_), .B0(new_n8454_), .Y(new_n8935_));
  AND2X1   g08743(.A(new_n8935_), .B(new_n8444_), .Y(new_n8936_));
  OAI21X1  g08744(.A0(new_n8873_), .A1(new_n8861_), .B0(new_n8936_), .Y(new_n8937_));
  AOI22X1  g08745(.A0(new_n8490_), .A1(new_n8489_), .B0(new_n8468_), .B1(\asqrt[30] ), .Y(new_n8938_));
  OAI21X1  g08746(.A0(new_n8873_), .A1(new_n8861_), .B0(new_n8938_), .Y(new_n8939_));
  NAND2X1  g08747(.A(new_n8939_), .B(new_n8454_), .Y(new_n8940_));
  AND2X1   g08748(.A(new_n8940_), .B(new_n8937_), .Y(new_n8941_));
  NOR3X1   g08749(.A(new_n8933_), .B(new_n8920_), .C(\asqrt[31] ), .Y(new_n8942_));
  OAI21X1  g08750(.A0(new_n8942_), .A1(new_n8941_), .B0(new_n8934_), .Y(new_n8943_));
  AND2X1   g08751(.A(new_n8943_), .B(\asqrt[32] ), .Y(new_n8944_));
  OR2X1    g08752(.A(new_n8942_), .B(new_n8941_), .Y(new_n8945_));
  INVX1    g08753(.A(new_n8874_), .Y(\asqrt[27] ));
  AND2X1   g08754(.A(new_n8469_), .B(new_n8455_), .Y(new_n8947_));
  NOR3X1   g08755(.A(new_n8947_), .B(new_n8494_), .C(new_n8456_), .Y(new_n8948_));
  NOR2X1   g08756(.A(new_n8947_), .B(new_n8456_), .Y(new_n8949_));
  OAI21X1  g08757(.A0(new_n8873_), .A1(new_n8861_), .B0(new_n8949_), .Y(new_n8950_));
  AOI22X1  g08758(.A0(new_n8950_), .A1(new_n8494_), .B0(new_n8948_), .B1(\asqrt[27] ), .Y(new_n8951_));
  AND2X1   g08759(.A(new_n8934_), .B(new_n6699_), .Y(new_n8952_));
  AOI21X1  g08760(.A0(new_n8952_), .A1(new_n8945_), .B0(new_n8951_), .Y(new_n8953_));
  OAI21X1  g08761(.A0(new_n8953_), .A1(new_n8944_), .B0(\asqrt[33] ), .Y(new_n8954_));
  NAND4X1  g08762(.A(\asqrt[27] ), .B(new_n8508_), .C(new_n8478_), .D(new_n8471_), .Y(new_n8955_));
  NOR3X1   g08763(.A(new_n8874_), .B(new_n8479_), .C(new_n8497_), .Y(new_n8956_));
  OAI21X1  g08764(.A0(new_n8956_), .A1(new_n8478_), .B0(new_n8955_), .Y(new_n8957_));
  AND2X1   g08765(.A(new_n8931_), .B(\asqrt[29] ), .Y(new_n8958_));
  OR2X1    g08766(.A(new_n8930_), .B(new_n8927_), .Y(new_n8959_));
  AND2X1   g08767(.A(new_n8908_), .B(new_n7970_), .Y(new_n8960_));
  NOR2X1   g08768(.A(new_n8917_), .B(new_n8915_), .Y(new_n8961_));
  AOI21X1  g08769(.A0(new_n8960_), .A1(new_n8959_), .B0(new_n8961_), .Y(new_n8962_));
  OAI21X1  g08770(.A0(new_n8962_), .A1(new_n8958_), .B0(\asqrt[30] ), .Y(new_n8963_));
  NAND2X1  g08771(.A(new_n8925_), .B(new_n8922_), .Y(new_n8964_));
  OAI21X1  g08772(.A0(new_n8905_), .A1(new_n7970_), .B0(new_n7527_), .Y(new_n8965_));
  OAI21X1  g08773(.A0(new_n8965_), .A1(new_n8962_), .B0(new_n8964_), .Y(new_n8966_));
  AOI21X1  g08774(.A0(new_n8966_), .A1(new_n8963_), .B0(new_n7103_), .Y(new_n8967_));
  INVX1    g08775(.A(new_n8941_), .Y(new_n8968_));
  NAND3X1  g08776(.A(new_n8966_), .B(new_n8963_), .C(new_n7103_), .Y(new_n8969_));
  AOI21X1  g08777(.A0(new_n8969_), .A1(new_n8968_), .B0(new_n8967_), .Y(new_n8970_));
  OAI21X1  g08778(.A0(new_n8970_), .A1(new_n6699_), .B0(new_n6294_), .Y(new_n8971_));
  OAI21X1  g08779(.A0(new_n8971_), .A1(new_n8953_), .B0(new_n8957_), .Y(new_n8972_));
  AOI21X1  g08780(.A0(new_n8972_), .A1(new_n8954_), .B0(new_n5941_), .Y(new_n8973_));
  AND2X1   g08781(.A(new_n8498_), .B(new_n8482_), .Y(new_n8974_));
  NOR3X1   g08782(.A(new_n8974_), .B(new_n8524_), .C(new_n8481_), .Y(new_n8975_));
  NOR3X1   g08783(.A(new_n8874_), .B(new_n8974_), .C(new_n8481_), .Y(new_n8976_));
  NOR2X1   g08784(.A(new_n8976_), .B(new_n8487_), .Y(new_n8977_));
  AOI21X1  g08785(.A0(new_n8975_), .A1(\asqrt[27] ), .B0(new_n8977_), .Y(new_n8978_));
  INVX1    g08786(.A(new_n8978_), .Y(new_n8979_));
  NAND3X1  g08787(.A(new_n8972_), .B(new_n8954_), .C(new_n5941_), .Y(new_n8980_));
  AOI21X1  g08788(.A0(new_n8980_), .A1(new_n8979_), .B0(new_n8973_), .Y(new_n8981_));
  OR2X1    g08789(.A(new_n8981_), .B(new_n5541_), .Y(new_n8982_));
  AND2X1   g08790(.A(new_n8980_), .B(new_n8979_), .Y(new_n8983_));
  AND2X1   g08791(.A(new_n8528_), .B(new_n8526_), .Y(new_n8984_));
  NOR3X1   g08792(.A(new_n8984_), .B(new_n8506_), .C(new_n8527_), .Y(new_n8985_));
  NOR3X1   g08793(.A(new_n8874_), .B(new_n8984_), .C(new_n8527_), .Y(new_n8986_));
  NOR2X1   g08794(.A(new_n8986_), .B(new_n8505_), .Y(new_n8987_));
  AOI21X1  g08795(.A0(new_n8985_), .A1(\asqrt[27] ), .B0(new_n8987_), .Y(new_n8988_));
  INVX1    g08796(.A(new_n8988_), .Y(new_n8989_));
  OR2X1    g08797(.A(new_n8970_), .B(new_n6699_), .Y(new_n8990_));
  NOR2X1   g08798(.A(new_n8942_), .B(new_n8941_), .Y(new_n8991_));
  INVX1    g08799(.A(new_n8951_), .Y(new_n8992_));
  NAND2X1  g08800(.A(new_n8934_), .B(new_n6699_), .Y(new_n8993_));
  OAI21X1  g08801(.A0(new_n8993_), .A1(new_n8991_), .B0(new_n8992_), .Y(new_n8994_));
  AOI21X1  g08802(.A0(new_n8994_), .A1(new_n8990_), .B0(new_n6294_), .Y(new_n8995_));
  INVX1    g08803(.A(new_n8957_), .Y(new_n8996_));
  AOI21X1  g08804(.A0(new_n8943_), .A1(\asqrt[32] ), .B0(\asqrt[33] ), .Y(new_n8997_));
  AOI21X1  g08805(.A0(new_n8997_), .A1(new_n8994_), .B0(new_n8996_), .Y(new_n8998_));
  OAI21X1  g08806(.A0(new_n8998_), .A1(new_n8995_), .B0(\asqrt[34] ), .Y(new_n8999_));
  NAND2X1  g08807(.A(new_n8999_), .B(new_n5541_), .Y(new_n9000_));
  OAI21X1  g08808(.A0(new_n9000_), .A1(new_n8983_), .B0(new_n8989_), .Y(new_n9001_));
  AOI21X1  g08809(.A0(new_n9001_), .A1(new_n8982_), .B0(new_n5176_), .Y(new_n9002_));
  OR4X1    g08810(.A(new_n8874_), .B(new_n8530_), .C(new_n8518_), .D(new_n8512_), .Y(new_n9003_));
  OR2X1    g08811(.A(new_n8530_), .B(new_n8512_), .Y(new_n9004_));
  OAI21X1  g08812(.A0(new_n9004_), .A1(new_n8874_), .B0(new_n8518_), .Y(new_n9005_));
  AND2X1   g08813(.A(new_n9005_), .B(new_n9003_), .Y(new_n9006_));
  NOR3X1   g08814(.A(new_n8998_), .B(new_n8995_), .C(\asqrt[34] ), .Y(new_n9007_));
  OAI21X1  g08815(.A0(new_n9007_), .A1(new_n8978_), .B0(new_n8999_), .Y(new_n9008_));
  AOI21X1  g08816(.A0(new_n9008_), .A1(\asqrt[35] ), .B0(\asqrt[36] ), .Y(new_n9009_));
  AOI21X1  g08817(.A0(new_n9009_), .A1(new_n9001_), .B0(new_n9006_), .Y(new_n9010_));
  OAI21X1  g08818(.A0(new_n9010_), .A1(new_n9002_), .B0(\asqrt[37] ), .Y(new_n9011_));
  AOI21X1  g08819(.A0(new_n8574_), .A1(new_n8573_), .B0(new_n8536_), .Y(new_n9012_));
  AND2X1   g08820(.A(new_n9012_), .B(new_n8521_), .Y(new_n9013_));
  AOI22X1  g08821(.A0(new_n8574_), .A1(new_n8573_), .B0(new_n8541_), .B1(\asqrt[36] ), .Y(new_n9014_));
  AOI21X1  g08822(.A0(new_n9014_), .A1(\asqrt[27] ), .B0(new_n8535_), .Y(new_n9015_));
  AOI21X1  g08823(.A0(new_n9013_), .A1(\asqrt[27] ), .B0(new_n9015_), .Y(new_n9016_));
  NOR3X1   g08824(.A(new_n9010_), .B(new_n9002_), .C(\asqrt[37] ), .Y(new_n9017_));
  OAI21X1  g08825(.A0(new_n9017_), .A1(new_n9016_), .B0(new_n9011_), .Y(new_n9018_));
  AND2X1   g08826(.A(new_n9018_), .B(\asqrt[38] ), .Y(new_n9019_));
  INVX1    g08827(.A(new_n9016_), .Y(new_n9020_));
  AND2X1   g08828(.A(new_n9008_), .B(\asqrt[35] ), .Y(new_n9021_));
  NAND2X1  g08829(.A(new_n8980_), .B(new_n8979_), .Y(new_n9022_));
  AND2X1   g08830(.A(new_n8999_), .B(new_n5541_), .Y(new_n9023_));
  AOI21X1  g08831(.A0(new_n9023_), .A1(new_n9022_), .B0(new_n8988_), .Y(new_n9024_));
  OAI21X1  g08832(.A0(new_n9024_), .A1(new_n9021_), .B0(\asqrt[36] ), .Y(new_n9025_));
  INVX1    g08833(.A(new_n9006_), .Y(new_n9026_));
  OAI21X1  g08834(.A0(new_n8981_), .A1(new_n5541_), .B0(new_n5176_), .Y(new_n9027_));
  OAI21X1  g08835(.A0(new_n9027_), .A1(new_n9024_), .B0(new_n9026_), .Y(new_n9028_));
  NAND3X1  g08836(.A(new_n9028_), .B(new_n9025_), .C(new_n4826_), .Y(new_n9029_));
  NAND2X1  g08837(.A(new_n9029_), .B(new_n9020_), .Y(new_n9030_));
  AND2X1   g08838(.A(new_n9011_), .B(new_n4493_), .Y(new_n9031_));
  AND2X1   g08839(.A(new_n8542_), .B(new_n8539_), .Y(new_n9032_));
  NOR3X1   g08840(.A(new_n8578_), .B(new_n9032_), .C(new_n8540_), .Y(new_n9033_));
  NOR3X1   g08841(.A(new_n8874_), .B(new_n9032_), .C(new_n8540_), .Y(new_n9034_));
  NOR2X1   g08842(.A(new_n9034_), .B(new_n8547_), .Y(new_n9035_));
  AOI21X1  g08843(.A0(new_n9033_), .A1(\asqrt[27] ), .B0(new_n9035_), .Y(new_n9036_));
  AOI21X1  g08844(.A0(new_n9031_), .A1(new_n9030_), .B0(new_n9036_), .Y(new_n9037_));
  OAI21X1  g08845(.A0(new_n9037_), .A1(new_n9019_), .B0(\asqrt[39] ), .Y(new_n9038_));
  NAND4X1  g08846(.A(\asqrt[27] ), .B(new_n8582_), .C(new_n8554_), .D(new_n8549_), .Y(new_n9039_));
  OR2X1    g08847(.A(new_n8555_), .B(new_n8580_), .Y(new_n9040_));
  OAI21X1  g08848(.A0(new_n9040_), .A1(new_n8874_), .B0(new_n8581_), .Y(new_n9041_));
  AND2X1   g08849(.A(new_n9041_), .B(new_n9039_), .Y(new_n9042_));
  INVX1    g08850(.A(new_n9042_), .Y(new_n9043_));
  AOI21X1  g08851(.A0(new_n9028_), .A1(new_n9025_), .B0(new_n4826_), .Y(new_n9044_));
  AOI21X1  g08852(.A0(new_n9029_), .A1(new_n9020_), .B0(new_n9044_), .Y(new_n9045_));
  OAI21X1  g08853(.A0(new_n9045_), .A1(new_n4493_), .B0(new_n4165_), .Y(new_n9046_));
  OAI21X1  g08854(.A0(new_n9046_), .A1(new_n9037_), .B0(new_n9043_), .Y(new_n9047_));
  AOI21X1  g08855(.A0(new_n9047_), .A1(new_n9038_), .B0(new_n3863_), .Y(new_n9048_));
  AND2X1   g08856(.A(new_n8563_), .B(new_n8558_), .Y(new_n9049_));
  NOR3X1   g08857(.A(new_n9049_), .B(new_n8612_), .C(new_n8557_), .Y(new_n9050_));
  NOR3X1   g08858(.A(new_n8874_), .B(new_n9049_), .C(new_n8557_), .Y(new_n9051_));
  NOR2X1   g08859(.A(new_n9051_), .B(new_n8562_), .Y(new_n9052_));
  AOI21X1  g08860(.A0(new_n9050_), .A1(\asqrt[27] ), .B0(new_n9052_), .Y(new_n9053_));
  INVX1    g08861(.A(new_n9053_), .Y(new_n9054_));
  NAND3X1  g08862(.A(new_n9047_), .B(new_n9038_), .C(new_n3863_), .Y(new_n9055_));
  AOI21X1  g08863(.A0(new_n9055_), .A1(new_n9054_), .B0(new_n9048_), .Y(new_n9056_));
  OR2X1    g08864(.A(new_n9056_), .B(new_n3564_), .Y(new_n9057_));
  AND2X1   g08865(.A(new_n9055_), .B(new_n9054_), .Y(new_n9058_));
  AND2X1   g08866(.A(new_n8616_), .B(new_n8614_), .Y(new_n9059_));
  NOR3X1   g08867(.A(new_n9059_), .B(new_n8571_), .C(new_n8615_), .Y(new_n9060_));
  NOR3X1   g08868(.A(new_n8874_), .B(new_n9059_), .C(new_n8615_), .Y(new_n9061_));
  NOR2X1   g08869(.A(new_n9061_), .B(new_n8570_), .Y(new_n9062_));
  AOI21X1  g08870(.A0(new_n9060_), .A1(\asqrt[27] ), .B0(new_n9062_), .Y(new_n9063_));
  INVX1    g08871(.A(new_n9063_), .Y(new_n9064_));
  OR2X1    g08872(.A(new_n9045_), .B(new_n4493_), .Y(new_n9065_));
  AND2X1   g08873(.A(new_n9029_), .B(new_n9020_), .Y(new_n9066_));
  NAND2X1  g08874(.A(new_n9011_), .B(new_n4493_), .Y(new_n9067_));
  INVX1    g08875(.A(new_n9036_), .Y(new_n9068_));
  OAI21X1  g08876(.A0(new_n9067_), .A1(new_n9066_), .B0(new_n9068_), .Y(new_n9069_));
  AOI21X1  g08877(.A0(new_n9069_), .A1(new_n9065_), .B0(new_n4165_), .Y(new_n9070_));
  AOI21X1  g08878(.A0(new_n9018_), .A1(\asqrt[38] ), .B0(\asqrt[39] ), .Y(new_n9071_));
  AOI21X1  g08879(.A0(new_n9071_), .A1(new_n9069_), .B0(new_n9042_), .Y(new_n9072_));
  OAI21X1  g08880(.A0(new_n9072_), .A1(new_n9070_), .B0(\asqrt[40] ), .Y(new_n9073_));
  NAND2X1  g08881(.A(new_n9073_), .B(new_n3564_), .Y(new_n9074_));
  OAI21X1  g08882(.A0(new_n9074_), .A1(new_n9058_), .B0(new_n9064_), .Y(new_n9075_));
  AOI21X1  g08883(.A0(new_n9075_), .A1(new_n9057_), .B0(new_n3276_), .Y(new_n9076_));
  NAND4X1  g08884(.A(\asqrt[27] ), .B(new_n8593_), .C(new_n8591_), .D(new_n8618_), .Y(new_n9077_));
  NAND2X1  g08885(.A(new_n8593_), .B(new_n8618_), .Y(new_n9078_));
  OAI21X1  g08886(.A0(new_n9078_), .A1(new_n8874_), .B0(new_n8592_), .Y(new_n9079_));
  AND2X1   g08887(.A(new_n9079_), .B(new_n9077_), .Y(new_n9080_));
  NOR3X1   g08888(.A(new_n9072_), .B(new_n9070_), .C(\asqrt[40] ), .Y(new_n9081_));
  OAI21X1  g08889(.A0(new_n9081_), .A1(new_n9053_), .B0(new_n9073_), .Y(new_n9082_));
  AOI21X1  g08890(.A0(new_n9082_), .A1(\asqrt[41] ), .B0(\asqrt[42] ), .Y(new_n9083_));
  AOI21X1  g08891(.A0(new_n9083_), .A1(new_n9075_), .B0(new_n9080_), .Y(new_n9084_));
  OAI21X1  g08892(.A0(new_n9084_), .A1(new_n9076_), .B0(\asqrt[43] ), .Y(new_n9085_));
  AOI21X1  g08893(.A0(new_n8635_), .A1(new_n8634_), .B0(new_n8601_), .Y(new_n9086_));
  AND2X1   g08894(.A(new_n9086_), .B(new_n8595_), .Y(new_n9087_));
  AOI22X1  g08895(.A0(new_n8635_), .A1(new_n8634_), .B0(new_n8620_), .B1(\asqrt[42] ), .Y(new_n9088_));
  AOI21X1  g08896(.A0(new_n9088_), .A1(\asqrt[27] ), .B0(new_n8600_), .Y(new_n9089_));
  AOI21X1  g08897(.A0(new_n9087_), .A1(\asqrt[27] ), .B0(new_n9089_), .Y(new_n9090_));
  NOR3X1   g08898(.A(new_n9084_), .B(new_n9076_), .C(\asqrt[43] ), .Y(new_n9091_));
  OAI21X1  g08899(.A0(new_n9091_), .A1(new_n9090_), .B0(new_n9085_), .Y(new_n9092_));
  AND2X1   g08900(.A(new_n9092_), .B(\asqrt[44] ), .Y(new_n9093_));
  INVX1    g08901(.A(new_n9090_), .Y(new_n9094_));
  AND2X1   g08902(.A(new_n9082_), .B(\asqrt[41] ), .Y(new_n9095_));
  NAND2X1  g08903(.A(new_n9055_), .B(new_n9054_), .Y(new_n9096_));
  AND2X1   g08904(.A(new_n9073_), .B(new_n3564_), .Y(new_n9097_));
  AOI21X1  g08905(.A0(new_n9097_), .A1(new_n9096_), .B0(new_n9063_), .Y(new_n9098_));
  OAI21X1  g08906(.A0(new_n9098_), .A1(new_n9095_), .B0(\asqrt[42] ), .Y(new_n9099_));
  INVX1    g08907(.A(new_n9080_), .Y(new_n9100_));
  OAI21X1  g08908(.A0(new_n9056_), .A1(new_n3564_), .B0(new_n3276_), .Y(new_n9101_));
  OAI21X1  g08909(.A0(new_n9101_), .A1(new_n9098_), .B0(new_n9100_), .Y(new_n9102_));
  NAND3X1  g08910(.A(new_n9102_), .B(new_n9099_), .C(new_n3008_), .Y(new_n9103_));
  NAND2X1  g08911(.A(new_n9103_), .B(new_n9094_), .Y(new_n9104_));
  AND2X1   g08912(.A(new_n8621_), .B(new_n8603_), .Y(new_n9105_));
  NOR3X1   g08913(.A(new_n9105_), .B(new_n8638_), .C(new_n8604_), .Y(new_n9106_));
  NOR3X1   g08914(.A(new_n8874_), .B(new_n9105_), .C(new_n8604_), .Y(new_n9107_));
  NOR2X1   g08915(.A(new_n9107_), .B(new_n8609_), .Y(new_n9108_));
  AOI21X1  g08916(.A0(new_n9106_), .A1(\asqrt[27] ), .B0(new_n9108_), .Y(new_n9109_));
  AND2X1   g08917(.A(new_n9085_), .B(new_n2769_), .Y(new_n9110_));
  AOI21X1  g08918(.A0(new_n9110_), .A1(new_n9104_), .B0(new_n9109_), .Y(new_n9111_));
  OAI21X1  g08919(.A0(new_n9111_), .A1(new_n9093_), .B0(\asqrt[45] ), .Y(new_n9112_));
  NAND4X1  g08920(.A(\asqrt[27] ), .B(new_n8641_), .C(new_n8628_), .D(new_n8623_), .Y(new_n9113_));
  NAND2X1  g08921(.A(new_n8641_), .B(new_n8623_), .Y(new_n9114_));
  OAI21X1  g08922(.A0(new_n9114_), .A1(new_n8874_), .B0(new_n8632_), .Y(new_n9115_));
  AND2X1   g08923(.A(new_n9115_), .B(new_n9113_), .Y(new_n9116_));
  INVX1    g08924(.A(new_n9116_), .Y(new_n9117_));
  AOI21X1  g08925(.A0(new_n9102_), .A1(new_n9099_), .B0(new_n3008_), .Y(new_n9118_));
  AOI21X1  g08926(.A0(new_n9103_), .A1(new_n9094_), .B0(new_n9118_), .Y(new_n9119_));
  OAI21X1  g08927(.A0(new_n9119_), .A1(new_n2769_), .B0(new_n2570_), .Y(new_n9120_));
  OAI21X1  g08928(.A0(new_n9120_), .A1(new_n9111_), .B0(new_n9117_), .Y(new_n9121_));
  AOI21X1  g08929(.A0(new_n9121_), .A1(new_n9112_), .B0(new_n2263_), .Y(new_n9122_));
  AND2X1   g08930(.A(new_n8648_), .B(new_n8642_), .Y(new_n9123_));
  NOR3X1   g08931(.A(new_n9123_), .B(new_n8686_), .C(new_n8631_), .Y(new_n9124_));
  NOR3X1   g08932(.A(new_n8874_), .B(new_n9123_), .C(new_n8631_), .Y(new_n9125_));
  NOR2X1   g08933(.A(new_n9125_), .B(new_n8646_), .Y(new_n9126_));
  AOI21X1  g08934(.A0(new_n9124_), .A1(\asqrt[27] ), .B0(new_n9126_), .Y(new_n9127_));
  INVX1    g08935(.A(new_n9127_), .Y(new_n9128_));
  NAND3X1  g08936(.A(new_n9121_), .B(new_n9112_), .C(new_n2263_), .Y(new_n9129_));
  AOI21X1  g08937(.A0(new_n9129_), .A1(new_n9128_), .B0(new_n9122_), .Y(new_n9130_));
  OR2X1    g08938(.A(new_n9130_), .B(new_n2040_), .Y(new_n9131_));
  AND2X1   g08939(.A(new_n9129_), .B(new_n9128_), .Y(new_n9132_));
  AND2X1   g08940(.A(new_n8690_), .B(new_n8688_), .Y(new_n9133_));
  NOR3X1   g08941(.A(new_n9133_), .B(new_n8656_), .C(new_n8689_), .Y(new_n9134_));
  NOR3X1   g08942(.A(new_n8874_), .B(new_n9133_), .C(new_n8689_), .Y(new_n9135_));
  NOR2X1   g08943(.A(new_n9135_), .B(new_n8655_), .Y(new_n9136_));
  AOI21X1  g08944(.A0(new_n9134_), .A1(\asqrt[27] ), .B0(new_n9136_), .Y(new_n9137_));
  INVX1    g08945(.A(new_n9137_), .Y(new_n9138_));
  OR2X1    g08946(.A(new_n9119_), .B(new_n2769_), .Y(new_n9139_));
  AND2X1   g08947(.A(new_n9103_), .B(new_n9094_), .Y(new_n9140_));
  INVX1    g08948(.A(new_n9109_), .Y(new_n9141_));
  NAND2X1  g08949(.A(new_n9085_), .B(new_n2769_), .Y(new_n9142_));
  OAI21X1  g08950(.A0(new_n9142_), .A1(new_n9140_), .B0(new_n9141_), .Y(new_n9143_));
  AOI21X1  g08951(.A0(new_n9143_), .A1(new_n9139_), .B0(new_n2570_), .Y(new_n9144_));
  AOI21X1  g08952(.A0(new_n9092_), .A1(\asqrt[44] ), .B0(\asqrt[45] ), .Y(new_n9145_));
  AOI21X1  g08953(.A0(new_n9145_), .A1(new_n9143_), .B0(new_n9116_), .Y(new_n9146_));
  OAI21X1  g08954(.A0(new_n9146_), .A1(new_n9144_), .B0(\asqrt[46] ), .Y(new_n9147_));
  NAND2X1  g08955(.A(new_n9147_), .B(new_n2040_), .Y(new_n9148_));
  OAI21X1  g08956(.A0(new_n9148_), .A1(new_n9132_), .B0(new_n9138_), .Y(new_n9149_));
  AOI21X1  g08957(.A0(new_n9149_), .A1(new_n9131_), .B0(new_n1834_), .Y(new_n9150_));
  NAND4X1  g08958(.A(\asqrt[27] ), .B(new_n8667_), .C(new_n8665_), .D(new_n8692_), .Y(new_n9151_));
  NAND2X1  g08959(.A(new_n8667_), .B(new_n8692_), .Y(new_n9152_));
  OAI21X1  g08960(.A0(new_n9152_), .A1(new_n8874_), .B0(new_n8666_), .Y(new_n9153_));
  AND2X1   g08961(.A(new_n9153_), .B(new_n9151_), .Y(new_n9154_));
  NOR3X1   g08962(.A(new_n9146_), .B(new_n9144_), .C(\asqrt[46] ), .Y(new_n9155_));
  OAI21X1  g08963(.A0(new_n9155_), .A1(new_n9127_), .B0(new_n9147_), .Y(new_n9156_));
  AOI21X1  g08964(.A0(new_n9156_), .A1(\asqrt[47] ), .B0(\asqrt[48] ), .Y(new_n9157_));
  AOI21X1  g08965(.A0(new_n9157_), .A1(new_n9149_), .B0(new_n9154_), .Y(new_n9158_));
  OAI21X1  g08966(.A0(new_n9158_), .A1(new_n9150_), .B0(\asqrt[49] ), .Y(new_n9159_));
  AOI21X1  g08967(.A0(new_n8709_), .A1(new_n8708_), .B0(new_n8675_), .Y(new_n9160_));
  AND2X1   g08968(.A(new_n9160_), .B(new_n8669_), .Y(new_n9161_));
  AOI22X1  g08969(.A0(new_n8709_), .A1(new_n8708_), .B0(new_n8694_), .B1(\asqrt[48] ), .Y(new_n9162_));
  AOI21X1  g08970(.A0(new_n9162_), .A1(\asqrt[27] ), .B0(new_n8674_), .Y(new_n9163_));
  AOI21X1  g08971(.A0(new_n9161_), .A1(\asqrt[27] ), .B0(new_n9163_), .Y(new_n9164_));
  NOR3X1   g08972(.A(new_n9158_), .B(new_n9150_), .C(\asqrt[49] ), .Y(new_n9165_));
  OAI21X1  g08973(.A0(new_n9165_), .A1(new_n9164_), .B0(new_n9159_), .Y(new_n9166_));
  AND2X1   g08974(.A(new_n9166_), .B(\asqrt[50] ), .Y(new_n9167_));
  INVX1    g08975(.A(new_n9164_), .Y(new_n9168_));
  AND2X1   g08976(.A(new_n9156_), .B(\asqrt[47] ), .Y(new_n9169_));
  NAND2X1  g08977(.A(new_n9129_), .B(new_n9128_), .Y(new_n9170_));
  AND2X1   g08978(.A(new_n9147_), .B(new_n2040_), .Y(new_n9171_));
  AOI21X1  g08979(.A0(new_n9171_), .A1(new_n9170_), .B0(new_n9137_), .Y(new_n9172_));
  OAI21X1  g08980(.A0(new_n9172_), .A1(new_n9169_), .B0(\asqrt[48] ), .Y(new_n9173_));
  INVX1    g08981(.A(new_n9154_), .Y(new_n9174_));
  OAI21X1  g08982(.A0(new_n9130_), .A1(new_n2040_), .B0(new_n1834_), .Y(new_n9175_));
  OAI21X1  g08983(.A0(new_n9175_), .A1(new_n9172_), .B0(new_n9174_), .Y(new_n9176_));
  NAND3X1  g08984(.A(new_n9176_), .B(new_n9173_), .C(new_n1632_), .Y(new_n9177_));
  NAND2X1  g08985(.A(new_n9177_), .B(new_n9168_), .Y(new_n9178_));
  AND2X1   g08986(.A(new_n8695_), .B(new_n8677_), .Y(new_n9179_));
  NOR3X1   g08987(.A(new_n9179_), .B(new_n8712_), .C(new_n8678_), .Y(new_n9180_));
  NOR3X1   g08988(.A(new_n8874_), .B(new_n9179_), .C(new_n8678_), .Y(new_n9181_));
  NOR2X1   g08989(.A(new_n9181_), .B(new_n8683_), .Y(new_n9182_));
  AOI21X1  g08990(.A0(new_n9180_), .A1(\asqrt[27] ), .B0(new_n9182_), .Y(new_n9183_));
  AND2X1   g08991(.A(new_n9159_), .B(new_n1469_), .Y(new_n9184_));
  AOI21X1  g08992(.A0(new_n9184_), .A1(new_n9178_), .B0(new_n9183_), .Y(new_n9185_));
  OAI21X1  g08993(.A0(new_n9185_), .A1(new_n9167_), .B0(\asqrt[51] ), .Y(new_n9186_));
  NAND4X1  g08994(.A(\asqrt[27] ), .B(new_n8715_), .C(new_n8702_), .D(new_n8697_), .Y(new_n9187_));
  NAND2X1  g08995(.A(new_n8715_), .B(new_n8697_), .Y(new_n9188_));
  OAI21X1  g08996(.A0(new_n9188_), .A1(new_n8874_), .B0(new_n8706_), .Y(new_n9189_));
  AND2X1   g08997(.A(new_n9189_), .B(new_n9187_), .Y(new_n9190_));
  INVX1    g08998(.A(new_n9190_), .Y(new_n9191_));
  AOI21X1  g08999(.A0(new_n9176_), .A1(new_n9173_), .B0(new_n1632_), .Y(new_n9192_));
  AOI21X1  g09000(.A0(new_n9177_), .A1(new_n9168_), .B0(new_n9192_), .Y(new_n9193_));
  OAI21X1  g09001(.A0(new_n9193_), .A1(new_n1469_), .B0(new_n1277_), .Y(new_n9194_));
  OAI21X1  g09002(.A0(new_n9194_), .A1(new_n9185_), .B0(new_n9191_), .Y(new_n9195_));
  AOI21X1  g09003(.A0(new_n9195_), .A1(new_n9186_), .B0(new_n1111_), .Y(new_n9196_));
  AND2X1   g09004(.A(new_n8722_), .B(new_n8716_), .Y(new_n9197_));
  NOR3X1   g09005(.A(new_n9197_), .B(new_n8746_), .C(new_n8705_), .Y(new_n9198_));
  NOR3X1   g09006(.A(new_n8874_), .B(new_n9197_), .C(new_n8705_), .Y(new_n9199_));
  NOR2X1   g09007(.A(new_n9199_), .B(new_n8720_), .Y(new_n9200_));
  AOI21X1  g09008(.A0(new_n9198_), .A1(\asqrt[27] ), .B0(new_n9200_), .Y(new_n9201_));
  INVX1    g09009(.A(new_n9201_), .Y(new_n9202_));
  NAND3X1  g09010(.A(new_n9195_), .B(new_n9186_), .C(new_n1111_), .Y(new_n9203_));
  AOI21X1  g09011(.A0(new_n9203_), .A1(new_n9202_), .B0(new_n9196_), .Y(new_n9204_));
  OR2X1    g09012(.A(new_n9204_), .B(new_n968_), .Y(new_n9205_));
  AND2X1   g09013(.A(new_n9203_), .B(new_n9202_), .Y(new_n9206_));
  AND2X1   g09014(.A(new_n8750_), .B(new_n8748_), .Y(new_n9207_));
  NOR3X1   g09015(.A(new_n9207_), .B(new_n8730_), .C(new_n8749_), .Y(new_n9208_));
  NOR3X1   g09016(.A(new_n8874_), .B(new_n9207_), .C(new_n8749_), .Y(new_n9209_));
  NOR2X1   g09017(.A(new_n9209_), .B(new_n8729_), .Y(new_n9210_));
  AOI21X1  g09018(.A0(new_n9208_), .A1(\asqrt[27] ), .B0(new_n9210_), .Y(new_n9211_));
  INVX1    g09019(.A(new_n9211_), .Y(new_n9212_));
  OR2X1    g09020(.A(new_n9193_), .B(new_n1469_), .Y(new_n9213_));
  AND2X1   g09021(.A(new_n9177_), .B(new_n9168_), .Y(new_n9214_));
  INVX1    g09022(.A(new_n9183_), .Y(new_n9215_));
  NAND2X1  g09023(.A(new_n9159_), .B(new_n1469_), .Y(new_n9216_));
  OAI21X1  g09024(.A0(new_n9216_), .A1(new_n9214_), .B0(new_n9215_), .Y(new_n9217_));
  AOI21X1  g09025(.A0(new_n9217_), .A1(new_n9213_), .B0(new_n1277_), .Y(new_n9218_));
  AOI21X1  g09026(.A0(new_n9166_), .A1(\asqrt[50] ), .B0(\asqrt[51] ), .Y(new_n9219_));
  AOI21X1  g09027(.A0(new_n9219_), .A1(new_n9217_), .B0(new_n9190_), .Y(new_n9220_));
  OAI21X1  g09028(.A0(new_n9220_), .A1(new_n9218_), .B0(\asqrt[52] ), .Y(new_n9221_));
  NAND2X1  g09029(.A(new_n9221_), .B(new_n968_), .Y(new_n9222_));
  OAI21X1  g09030(.A0(new_n9222_), .A1(new_n9206_), .B0(new_n9212_), .Y(new_n9223_));
  AOI21X1  g09031(.A0(new_n9223_), .A1(new_n9205_), .B0(new_n902_), .Y(new_n9224_));
  OR4X1    g09032(.A(new_n8874_), .B(new_n8752_), .C(new_n8740_), .D(new_n8734_), .Y(new_n9225_));
  OR2X1    g09033(.A(new_n8752_), .B(new_n8734_), .Y(new_n9226_));
  OAI21X1  g09034(.A0(new_n9226_), .A1(new_n8874_), .B0(new_n8740_), .Y(new_n9227_));
  AND2X1   g09035(.A(new_n9227_), .B(new_n9225_), .Y(new_n9228_));
  NOR3X1   g09036(.A(new_n9220_), .B(new_n9218_), .C(\asqrt[52] ), .Y(new_n9229_));
  OAI21X1  g09037(.A0(new_n9229_), .A1(new_n9201_), .B0(new_n9221_), .Y(new_n9230_));
  AOI21X1  g09038(.A0(new_n9230_), .A1(\asqrt[53] ), .B0(\asqrt[54] ), .Y(new_n9231_));
  AOI21X1  g09039(.A0(new_n9231_), .A1(new_n9223_), .B0(new_n9228_), .Y(new_n9232_));
  OAI21X1  g09040(.A0(new_n9232_), .A1(new_n9224_), .B0(\asqrt[55] ), .Y(new_n9233_));
  AOI21X1  g09041(.A0(new_n8796_), .A1(new_n8795_), .B0(new_n8758_), .Y(new_n9234_));
  AND2X1   g09042(.A(new_n9234_), .B(new_n8743_), .Y(new_n9235_));
  AOI22X1  g09043(.A0(new_n8796_), .A1(new_n8795_), .B0(new_n8768_), .B1(\asqrt[54] ), .Y(new_n9236_));
  AOI21X1  g09044(.A0(new_n9236_), .A1(\asqrt[27] ), .B0(new_n8757_), .Y(new_n9237_));
  AOI21X1  g09045(.A0(new_n9235_), .A1(\asqrt[27] ), .B0(new_n9237_), .Y(new_n9238_));
  NOR3X1   g09046(.A(new_n9232_), .B(new_n9224_), .C(\asqrt[55] ), .Y(new_n9239_));
  OAI21X1  g09047(.A0(new_n9239_), .A1(new_n9238_), .B0(new_n9233_), .Y(new_n9240_));
  AND2X1   g09048(.A(new_n9240_), .B(\asqrt[56] ), .Y(new_n9241_));
  OR2X1    g09049(.A(new_n9239_), .B(new_n9238_), .Y(new_n9242_));
  AND2X1   g09050(.A(new_n8769_), .B(new_n8761_), .Y(new_n9243_));
  NOR3X1   g09051(.A(new_n9243_), .B(new_n8799_), .C(new_n8762_), .Y(new_n9244_));
  NOR3X1   g09052(.A(new_n8874_), .B(new_n9243_), .C(new_n8762_), .Y(new_n9245_));
  NOR2X1   g09053(.A(new_n9245_), .B(new_n8767_), .Y(new_n9246_));
  AOI21X1  g09054(.A0(new_n9244_), .A1(\asqrt[27] ), .B0(new_n9246_), .Y(new_n9247_));
  AND2X1   g09055(.A(new_n9233_), .B(new_n582_), .Y(new_n9248_));
  AOI21X1  g09056(.A0(new_n9248_), .A1(new_n9242_), .B0(new_n9247_), .Y(new_n9249_));
  OAI21X1  g09057(.A0(new_n9249_), .A1(new_n9241_), .B0(\asqrt[57] ), .Y(new_n9250_));
  OR4X1    g09058(.A(new_n8874_), .B(new_n8777_), .C(new_n8803_), .D(new_n8802_), .Y(new_n9251_));
  OR2X1    g09059(.A(new_n8777_), .B(new_n8802_), .Y(new_n9252_));
  OAI21X1  g09060(.A0(new_n9252_), .A1(new_n8874_), .B0(new_n8803_), .Y(new_n9253_));
  AND2X1   g09061(.A(new_n9253_), .B(new_n9251_), .Y(new_n9254_));
  INVX1    g09062(.A(new_n9254_), .Y(new_n9255_));
  AND2X1   g09063(.A(new_n9230_), .B(\asqrt[53] ), .Y(new_n9256_));
  NAND2X1  g09064(.A(new_n9203_), .B(new_n9202_), .Y(new_n9257_));
  AND2X1   g09065(.A(new_n9221_), .B(new_n968_), .Y(new_n9258_));
  AOI21X1  g09066(.A0(new_n9258_), .A1(new_n9257_), .B0(new_n9211_), .Y(new_n9259_));
  OAI21X1  g09067(.A0(new_n9259_), .A1(new_n9256_), .B0(\asqrt[54] ), .Y(new_n9260_));
  INVX1    g09068(.A(new_n9228_), .Y(new_n9261_));
  OAI21X1  g09069(.A0(new_n9204_), .A1(new_n968_), .B0(new_n902_), .Y(new_n9262_));
  OAI21X1  g09070(.A0(new_n9262_), .A1(new_n9259_), .B0(new_n9261_), .Y(new_n9263_));
  AOI21X1  g09071(.A0(new_n9263_), .A1(new_n9260_), .B0(new_n697_), .Y(new_n9264_));
  INVX1    g09072(.A(new_n9238_), .Y(new_n9265_));
  NAND3X1  g09073(.A(new_n9263_), .B(new_n9260_), .C(new_n697_), .Y(new_n9266_));
  AOI21X1  g09074(.A0(new_n9266_), .A1(new_n9265_), .B0(new_n9264_), .Y(new_n9267_));
  OAI21X1  g09075(.A0(new_n9267_), .A1(new_n582_), .B0(new_n481_), .Y(new_n9268_));
  OAI21X1  g09076(.A0(new_n9268_), .A1(new_n9249_), .B0(new_n9255_), .Y(new_n9269_));
  AOI21X1  g09077(.A0(new_n9269_), .A1(new_n9250_), .B0(new_n399_), .Y(new_n9270_));
  AND2X1   g09078(.A(new_n8785_), .B(new_n8780_), .Y(new_n9271_));
  NOR3X1   g09079(.A(new_n9271_), .B(new_n8820_), .C(new_n8779_), .Y(new_n9272_));
  NOR3X1   g09080(.A(new_n8874_), .B(new_n9271_), .C(new_n8779_), .Y(new_n9273_));
  NOR2X1   g09081(.A(new_n9273_), .B(new_n8784_), .Y(new_n9274_));
  AOI21X1  g09082(.A0(new_n9272_), .A1(\asqrt[27] ), .B0(new_n9274_), .Y(new_n9275_));
  INVX1    g09083(.A(new_n9275_), .Y(new_n9276_));
  NAND3X1  g09084(.A(new_n9269_), .B(new_n9250_), .C(new_n399_), .Y(new_n9277_));
  AOI21X1  g09085(.A0(new_n9277_), .A1(new_n9276_), .B0(new_n9270_), .Y(new_n9278_));
  OR2X1    g09086(.A(new_n9278_), .B(new_n328_), .Y(new_n9279_));
  AND2X1   g09087(.A(new_n9277_), .B(new_n9276_), .Y(new_n9280_));
  AND2X1   g09088(.A(new_n8824_), .B(new_n8822_), .Y(new_n9281_));
  NOR3X1   g09089(.A(new_n9281_), .B(new_n8793_), .C(new_n8823_), .Y(new_n9282_));
  NOR3X1   g09090(.A(new_n8874_), .B(new_n9281_), .C(new_n8823_), .Y(new_n9283_));
  NOR2X1   g09091(.A(new_n9283_), .B(new_n8792_), .Y(new_n9284_));
  AOI21X1  g09092(.A0(new_n9282_), .A1(\asqrt[27] ), .B0(new_n9284_), .Y(new_n9285_));
  INVX1    g09093(.A(new_n9285_), .Y(new_n9286_));
  OR2X1    g09094(.A(new_n9267_), .B(new_n582_), .Y(new_n9287_));
  NOR2X1   g09095(.A(new_n9239_), .B(new_n9238_), .Y(new_n9288_));
  INVX1    g09096(.A(new_n9247_), .Y(new_n9289_));
  NAND2X1  g09097(.A(new_n9233_), .B(new_n582_), .Y(new_n9290_));
  OAI21X1  g09098(.A0(new_n9290_), .A1(new_n9288_), .B0(new_n9289_), .Y(new_n9291_));
  AOI21X1  g09099(.A0(new_n9291_), .A1(new_n9287_), .B0(new_n481_), .Y(new_n9292_));
  AOI21X1  g09100(.A0(new_n9240_), .A1(\asqrt[56] ), .B0(\asqrt[57] ), .Y(new_n9293_));
  AOI21X1  g09101(.A0(new_n9293_), .A1(new_n9291_), .B0(new_n9254_), .Y(new_n9294_));
  OAI21X1  g09102(.A0(new_n9294_), .A1(new_n9292_), .B0(\asqrt[58] ), .Y(new_n9295_));
  NAND2X1  g09103(.A(new_n9295_), .B(new_n328_), .Y(new_n9296_));
  OAI21X1  g09104(.A0(new_n9296_), .A1(new_n9280_), .B0(new_n9286_), .Y(new_n9297_));
  AOI21X1  g09105(.A0(new_n9297_), .A1(new_n9279_), .B0(new_n292_), .Y(new_n9298_));
  OR4X1    g09106(.A(new_n8874_), .B(new_n8826_), .C(new_n8814_), .D(new_n8808_), .Y(new_n9299_));
  OR2X1    g09107(.A(new_n8826_), .B(new_n8808_), .Y(new_n9300_));
  OAI21X1  g09108(.A0(new_n9300_), .A1(new_n8874_), .B0(new_n8814_), .Y(new_n9301_));
  AND2X1   g09109(.A(new_n9301_), .B(new_n9299_), .Y(new_n9302_));
  NOR3X1   g09110(.A(new_n9294_), .B(new_n9292_), .C(\asqrt[58] ), .Y(new_n9303_));
  OAI21X1  g09111(.A0(new_n9303_), .A1(new_n9275_), .B0(new_n9295_), .Y(new_n9304_));
  AOI21X1  g09112(.A0(new_n9304_), .A1(\asqrt[59] ), .B0(\asqrt[60] ), .Y(new_n9305_));
  AOI21X1  g09113(.A0(new_n9305_), .A1(new_n9297_), .B0(new_n9302_), .Y(new_n9306_));
  OAI21X1  g09114(.A0(new_n9306_), .A1(new_n9298_), .B0(\asqrt[61] ), .Y(new_n9307_));
  AOI21X1  g09115(.A0(new_n8878_), .A1(new_n8877_), .B0(new_n8832_), .Y(new_n9308_));
  AND2X1   g09116(.A(new_n9308_), .B(new_n8817_), .Y(new_n9309_));
  AOI22X1  g09117(.A0(new_n8878_), .A1(new_n8877_), .B0(new_n8842_), .B1(\asqrt[60] ), .Y(new_n9310_));
  AOI21X1  g09118(.A0(new_n9310_), .A1(\asqrt[27] ), .B0(new_n8831_), .Y(new_n9311_));
  AOI21X1  g09119(.A0(new_n9309_), .A1(\asqrt[27] ), .B0(new_n9311_), .Y(new_n9312_));
  NOR3X1   g09120(.A(new_n9306_), .B(new_n9298_), .C(\asqrt[61] ), .Y(new_n9313_));
  OAI21X1  g09121(.A0(new_n9313_), .A1(new_n9312_), .B0(new_n9307_), .Y(new_n9314_));
  AND2X1   g09122(.A(new_n9314_), .B(\asqrt[62] ), .Y(new_n9315_));
  OR2X1    g09123(.A(new_n9313_), .B(new_n9312_), .Y(new_n9316_));
  AND2X1   g09124(.A(new_n8843_), .B(new_n8835_), .Y(new_n9317_));
  NOR3X1   g09125(.A(new_n9317_), .B(new_n8881_), .C(new_n8836_), .Y(new_n9318_));
  NOR3X1   g09126(.A(new_n8874_), .B(new_n9317_), .C(new_n8836_), .Y(new_n9319_));
  NOR2X1   g09127(.A(new_n9319_), .B(new_n8841_), .Y(new_n9320_));
  AOI21X1  g09128(.A0(new_n9318_), .A1(\asqrt[27] ), .B0(new_n9320_), .Y(new_n9321_));
  AND2X1   g09129(.A(new_n9307_), .B(new_n199_), .Y(new_n9322_));
  AOI21X1  g09130(.A0(new_n9322_), .A1(new_n9316_), .B0(new_n9321_), .Y(new_n9323_));
  NOR4X1   g09131(.A(new_n8874_), .B(new_n8851_), .C(new_n8885_), .D(new_n8884_), .Y(new_n9324_));
  NAND3X1  g09132(.A(\asqrt[27] ), .B(new_n8886_), .C(new_n8845_), .Y(new_n9325_));
  AOI21X1  g09133(.A0(new_n9325_), .A1(new_n8885_), .B0(new_n9324_), .Y(new_n9326_));
  INVX1    g09134(.A(new_n9326_), .Y(new_n9327_));
  NOR3X1   g09135(.A(new_n8874_), .B(new_n8856_), .C(new_n8887_), .Y(new_n9328_));
  AOI21X1  g09136(.A0(new_n8891_), .A1(new_n8890_), .B0(new_n9328_), .Y(new_n9329_));
  AND2X1   g09137(.A(new_n9329_), .B(new_n9327_), .Y(new_n9330_));
  OAI21X1  g09138(.A0(new_n9323_), .A1(new_n9315_), .B0(new_n9330_), .Y(new_n9331_));
  AND2X1   g09139(.A(new_n9304_), .B(\asqrt[59] ), .Y(new_n9332_));
  NAND2X1  g09140(.A(new_n9277_), .B(new_n9276_), .Y(new_n9333_));
  AND2X1   g09141(.A(new_n9295_), .B(new_n328_), .Y(new_n9334_));
  AOI21X1  g09142(.A0(new_n9334_), .A1(new_n9333_), .B0(new_n9285_), .Y(new_n9335_));
  OAI21X1  g09143(.A0(new_n9335_), .A1(new_n9332_), .B0(\asqrt[60] ), .Y(new_n9336_));
  INVX1    g09144(.A(new_n9302_), .Y(new_n9337_));
  OAI21X1  g09145(.A0(new_n9278_), .A1(new_n328_), .B0(new_n292_), .Y(new_n9338_));
  OAI21X1  g09146(.A0(new_n9338_), .A1(new_n9335_), .B0(new_n9337_), .Y(new_n9339_));
  AOI21X1  g09147(.A0(new_n9339_), .A1(new_n9336_), .B0(new_n217_), .Y(new_n9340_));
  INVX1    g09148(.A(new_n9312_), .Y(new_n9341_));
  NAND3X1  g09149(.A(new_n9339_), .B(new_n9336_), .C(new_n217_), .Y(new_n9342_));
  AOI21X1  g09150(.A0(new_n9342_), .A1(new_n9341_), .B0(new_n9340_), .Y(new_n9343_));
  OAI21X1  g09151(.A0(new_n9343_), .A1(new_n199_), .B0(new_n9326_), .Y(new_n9344_));
  AOI21X1  g09152(.A0(new_n8893_), .A1(new_n8889_), .B0(new_n8856_), .Y(new_n9345_));
  AOI21X1  g09153(.A0(new_n8857_), .A1(new_n8852_), .B0(new_n193_), .Y(new_n9346_));
  OAI21X1  g09154(.A0(new_n9345_), .A1(new_n8852_), .B0(new_n9346_), .Y(new_n9347_));
  OR2X1    g09155(.A(new_n8863_), .B(new_n8862_), .Y(new_n9348_));
  NOR4X1   g09156(.A(new_n8870_), .B(new_n8911_), .C(new_n8855_), .D(new_n8853_), .Y(new_n9349_));
  NAND3X1  g09157(.A(new_n9349_), .B(new_n9348_), .C(new_n8889_), .Y(new_n9350_));
  AND2X1   g09158(.A(new_n9350_), .B(new_n9347_), .Y(new_n9351_));
  OAI21X1  g09159(.A0(new_n9344_), .A1(new_n9323_), .B0(new_n9351_), .Y(new_n9352_));
  AOI21X1  g09160(.A0(new_n9331_), .A1(new_n193_), .B0(new_n9352_), .Y(new_n9353_));
  OR2X1    g09161(.A(new_n9343_), .B(new_n199_), .Y(new_n9354_));
  NOR2X1   g09162(.A(new_n9313_), .B(new_n9312_), .Y(new_n9355_));
  INVX1    g09163(.A(new_n9321_), .Y(new_n9356_));
  NAND2X1  g09164(.A(new_n9307_), .B(new_n199_), .Y(new_n9357_));
  OAI21X1  g09165(.A0(new_n9357_), .A1(new_n9355_), .B0(new_n9356_), .Y(new_n9358_));
  INVX1    g09166(.A(new_n9330_), .Y(new_n9359_));
  AOI21X1  g09167(.A0(new_n9358_), .A1(new_n9354_), .B0(new_n9359_), .Y(new_n9360_));
  AOI21X1  g09168(.A0(new_n9314_), .A1(\asqrt[62] ), .B0(new_n9327_), .Y(new_n9361_));
  INVX1    g09169(.A(new_n9351_), .Y(new_n9362_));
  AOI21X1  g09170(.A0(new_n9361_), .A1(new_n9358_), .B0(new_n9362_), .Y(new_n9363_));
  OAI21X1  g09171(.A0(new_n9360_), .A1(\asqrt[63] ), .B0(new_n9363_), .Y(\asqrt[26] ));
  NOR2X1   g09172(.A(\a[51] ), .B(\a[50] ), .Y(new_n9365_));
  MX2X1    g09173(.A(new_n9365_), .B(\asqrt[26] ), .S0(\a[52] ), .Y(new_n9366_));
  AND2X1   g09174(.A(new_n9366_), .B(\asqrt[27] ), .Y(new_n9367_));
  NOR3X1   g09175(.A(\a[52] ), .B(\a[51] ), .C(\a[50] ), .Y(new_n9368_));
  NOR3X1   g09176(.A(new_n9368_), .B(new_n8870_), .C(new_n8911_), .Y(new_n9369_));
  NAND3X1  g09177(.A(new_n9369_), .B(new_n9348_), .C(new_n8889_), .Y(new_n9370_));
  AOI21X1  g09178(.A0(\asqrt[26] ), .A1(\a[52] ), .B0(new_n9370_), .Y(new_n9371_));
  INVX1    g09179(.A(\a[52] ), .Y(new_n9372_));
  INVX1    g09180(.A(\a[53] ), .Y(new_n9373_));
  AOI21X1  g09181(.A0(\asqrt[26] ), .A1(new_n9372_), .B0(new_n9373_), .Y(new_n9374_));
  NOR2X1   g09182(.A(\a[53] ), .B(\a[52] ), .Y(new_n9375_));
  AND2X1   g09183(.A(\asqrt[26] ), .B(new_n9375_), .Y(new_n9376_));
  NOR3X1   g09184(.A(new_n9376_), .B(new_n9374_), .C(new_n9371_), .Y(new_n9377_));
  OAI21X1  g09185(.A0(new_n9377_), .A1(new_n9367_), .B0(\asqrt[28] ), .Y(new_n9378_));
  INVX1    g09186(.A(new_n9365_), .Y(new_n9379_));
  MX2X1    g09187(.A(new_n9379_), .B(new_n9353_), .S0(\a[52] ), .Y(new_n9380_));
  OAI21X1  g09188(.A0(new_n9380_), .A1(new_n8874_), .B0(new_n8412_), .Y(new_n9381_));
  NAND3X1  g09189(.A(new_n9350_), .B(new_n9347_), .C(\asqrt[27] ), .Y(new_n9382_));
  INVX1    g09190(.A(new_n9382_), .Y(new_n9383_));
  OAI21X1  g09191(.A0(new_n9344_), .A1(new_n9323_), .B0(new_n9383_), .Y(new_n9384_));
  AOI21X1  g09192(.A0(new_n9331_), .A1(new_n193_), .B0(new_n9384_), .Y(new_n9385_));
  AOI21X1  g09193(.A0(\asqrt[26] ), .A1(new_n9375_), .B0(new_n9385_), .Y(new_n9386_));
  OR2X1    g09194(.A(new_n9385_), .B(\a[54] ), .Y(new_n9387_));
  OAI22X1  g09195(.A0(new_n9387_), .A1(new_n9376_), .B0(new_n9386_), .B1(new_n8875_), .Y(new_n9388_));
  OAI21X1  g09196(.A0(new_n9381_), .A1(new_n9377_), .B0(new_n9388_), .Y(new_n9389_));
  AOI21X1  g09197(.A0(new_n9389_), .A1(new_n9378_), .B0(new_n7970_), .Y(new_n9390_));
  AND2X1   g09198(.A(new_n8900_), .B(new_n8908_), .Y(new_n9391_));
  NAND3X1  g09199(.A(new_n9391_), .B(\asqrt[26] ), .C(new_n8930_), .Y(new_n9392_));
  INVX1    g09200(.A(new_n9391_), .Y(new_n9393_));
  OAI21X1  g09201(.A0(new_n9393_), .A1(new_n9353_), .B0(new_n8904_), .Y(new_n9394_));
  AND2X1   g09202(.A(new_n9394_), .B(new_n9392_), .Y(new_n9395_));
  INVX1    g09203(.A(new_n9395_), .Y(new_n9396_));
  NAND3X1  g09204(.A(new_n9389_), .B(new_n9378_), .C(new_n7970_), .Y(new_n9397_));
  AOI21X1  g09205(.A0(new_n9397_), .A1(new_n9396_), .B0(new_n9390_), .Y(new_n9398_));
  OR2X1    g09206(.A(new_n9398_), .B(new_n7527_), .Y(new_n9399_));
  AND2X1   g09207(.A(new_n9397_), .B(new_n9396_), .Y(new_n9400_));
  AOI21X1  g09208(.A0(new_n8960_), .A1(new_n8959_), .B0(new_n8918_), .Y(new_n9401_));
  NAND3X1  g09209(.A(new_n9401_), .B(\asqrt[26] ), .C(new_n8906_), .Y(new_n9402_));
  OAI22X1  g09210(.A0(new_n8909_), .A1(new_n8907_), .B0(new_n8905_), .B1(new_n7970_), .Y(new_n9403_));
  OAI21X1  g09211(.A0(new_n9403_), .A1(new_n9353_), .B0(new_n8918_), .Y(new_n9404_));
  AND2X1   g09212(.A(new_n9404_), .B(new_n9402_), .Y(new_n9405_));
  INVX1    g09213(.A(new_n9405_), .Y(new_n9406_));
  OR2X1    g09214(.A(new_n9390_), .B(\asqrt[30] ), .Y(new_n9407_));
  OAI21X1  g09215(.A0(new_n9407_), .A1(new_n9400_), .B0(new_n9406_), .Y(new_n9408_));
  AOI21X1  g09216(.A0(new_n9408_), .A1(new_n9399_), .B0(new_n7103_), .Y(new_n9409_));
  AND2X1   g09217(.A(new_n8932_), .B(new_n8919_), .Y(new_n9410_));
  OR4X1    g09218(.A(new_n9353_), .B(new_n9410_), .C(new_n8964_), .D(new_n8920_), .Y(new_n9411_));
  OR2X1    g09219(.A(new_n9410_), .B(new_n8920_), .Y(new_n9412_));
  OAI21X1  g09220(.A0(new_n9412_), .A1(new_n9353_), .B0(new_n8964_), .Y(new_n9413_));
  AND2X1   g09221(.A(new_n9413_), .B(new_n9411_), .Y(new_n9414_));
  OR2X1    g09222(.A(new_n9380_), .B(new_n8874_), .Y(new_n9415_));
  INVX1    g09223(.A(new_n9370_), .Y(new_n9416_));
  OAI21X1  g09224(.A0(new_n9353_), .A1(new_n9372_), .B0(new_n9416_), .Y(new_n9417_));
  OAI21X1  g09225(.A0(new_n9353_), .A1(\a[52] ), .B0(\a[53] ), .Y(new_n9418_));
  INVX1    g09226(.A(new_n9375_), .Y(new_n9419_));
  OR2X1    g09227(.A(new_n9353_), .B(new_n9419_), .Y(new_n9420_));
  NAND3X1  g09228(.A(new_n9420_), .B(new_n9418_), .C(new_n9417_), .Y(new_n9421_));
  AOI21X1  g09229(.A0(new_n9421_), .A1(new_n9415_), .B0(new_n8412_), .Y(new_n9422_));
  AOI21X1  g09230(.A0(new_n9366_), .A1(\asqrt[27] ), .B0(\asqrt[28] ), .Y(new_n9423_));
  OR2X1    g09231(.A(new_n9386_), .B(new_n8875_), .Y(new_n9424_));
  OR2X1    g09232(.A(new_n9387_), .B(new_n9376_), .Y(new_n9425_));
  AOI22X1  g09233(.A0(new_n9425_), .A1(new_n9424_), .B0(new_n9423_), .B1(new_n9421_), .Y(new_n9426_));
  OAI21X1  g09234(.A0(new_n9426_), .A1(new_n9422_), .B0(\asqrt[29] ), .Y(new_n9427_));
  NOR3X1   g09235(.A(new_n9426_), .B(new_n9422_), .C(\asqrt[29] ), .Y(new_n9428_));
  OAI21X1  g09236(.A0(new_n9428_), .A1(new_n9395_), .B0(new_n9427_), .Y(new_n9429_));
  AOI21X1  g09237(.A0(new_n9429_), .A1(\asqrt[30] ), .B0(\asqrt[31] ), .Y(new_n9430_));
  AOI21X1  g09238(.A0(new_n9430_), .A1(new_n9408_), .B0(new_n9414_), .Y(new_n9431_));
  OAI21X1  g09239(.A0(new_n9431_), .A1(new_n9409_), .B0(\asqrt[32] ), .Y(new_n9432_));
  OR4X1    g09240(.A(new_n9353_), .B(new_n8942_), .C(new_n8968_), .D(new_n8967_), .Y(new_n9433_));
  NAND2X1  g09241(.A(new_n8969_), .B(new_n8934_), .Y(new_n9434_));
  OAI21X1  g09242(.A0(new_n9434_), .A1(new_n9353_), .B0(new_n8968_), .Y(new_n9435_));
  AND2X1   g09243(.A(new_n9435_), .B(new_n9433_), .Y(new_n9436_));
  NOR3X1   g09244(.A(new_n9431_), .B(new_n9409_), .C(\asqrt[32] ), .Y(new_n9437_));
  OAI21X1  g09245(.A0(new_n9437_), .A1(new_n9436_), .B0(new_n9432_), .Y(new_n9438_));
  AND2X1   g09246(.A(new_n9438_), .B(\asqrt[33] ), .Y(new_n9439_));
  INVX1    g09247(.A(new_n9436_), .Y(new_n9440_));
  AND2X1   g09248(.A(new_n9429_), .B(\asqrt[30] ), .Y(new_n9441_));
  NAND2X1  g09249(.A(new_n9397_), .B(new_n9396_), .Y(new_n9442_));
  NOR2X1   g09250(.A(new_n9390_), .B(\asqrt[30] ), .Y(new_n9443_));
  AOI21X1  g09251(.A0(new_n9443_), .A1(new_n9442_), .B0(new_n9405_), .Y(new_n9444_));
  OAI21X1  g09252(.A0(new_n9444_), .A1(new_n9441_), .B0(\asqrt[31] ), .Y(new_n9445_));
  INVX1    g09253(.A(new_n9414_), .Y(new_n9446_));
  OAI21X1  g09254(.A0(new_n9398_), .A1(new_n7527_), .B0(new_n7103_), .Y(new_n9447_));
  OAI21X1  g09255(.A0(new_n9447_), .A1(new_n9444_), .B0(new_n9446_), .Y(new_n9448_));
  NAND3X1  g09256(.A(new_n9448_), .B(new_n9445_), .C(new_n6699_), .Y(new_n9449_));
  NAND2X1  g09257(.A(new_n9449_), .B(new_n9440_), .Y(new_n9450_));
  AND2X1   g09258(.A(new_n8952_), .B(new_n8945_), .Y(new_n9451_));
  NOR4X1   g09259(.A(new_n9353_), .B(new_n9451_), .C(new_n8992_), .D(new_n8944_), .Y(new_n9452_));
  AOI22X1  g09260(.A0(new_n8952_), .A1(new_n8945_), .B0(new_n8943_), .B1(\asqrt[32] ), .Y(new_n9453_));
  AOI21X1  g09261(.A0(new_n9453_), .A1(\asqrt[26] ), .B0(new_n8951_), .Y(new_n9454_));
  NOR2X1   g09262(.A(new_n9454_), .B(new_n9452_), .Y(new_n9455_));
  AOI21X1  g09263(.A0(new_n9448_), .A1(new_n9445_), .B0(new_n6699_), .Y(new_n9456_));
  NOR2X1   g09264(.A(new_n9456_), .B(\asqrt[33] ), .Y(new_n9457_));
  AOI21X1  g09265(.A0(new_n9457_), .A1(new_n9450_), .B0(new_n9455_), .Y(new_n9458_));
  OAI21X1  g09266(.A0(new_n9458_), .A1(new_n9439_), .B0(\asqrt[34] ), .Y(new_n9459_));
  AND2X1   g09267(.A(new_n8997_), .B(new_n8994_), .Y(new_n9460_));
  OR4X1    g09268(.A(new_n9353_), .B(new_n9460_), .C(new_n8957_), .D(new_n8995_), .Y(new_n9461_));
  OR2X1    g09269(.A(new_n9460_), .B(new_n8995_), .Y(new_n9462_));
  OAI21X1  g09270(.A0(new_n9462_), .A1(new_n9353_), .B0(new_n8957_), .Y(new_n9463_));
  AND2X1   g09271(.A(new_n9463_), .B(new_n9461_), .Y(new_n9464_));
  INVX1    g09272(.A(new_n9464_), .Y(new_n9465_));
  AOI21X1  g09273(.A0(new_n9449_), .A1(new_n9440_), .B0(new_n9456_), .Y(new_n9466_));
  OAI21X1  g09274(.A0(new_n9466_), .A1(new_n6294_), .B0(new_n5941_), .Y(new_n9467_));
  OAI21X1  g09275(.A0(new_n9467_), .A1(new_n9458_), .B0(new_n9465_), .Y(new_n9468_));
  AOI21X1  g09276(.A0(new_n9468_), .A1(new_n9459_), .B0(new_n5541_), .Y(new_n9469_));
  OR4X1    g09277(.A(new_n9353_), .B(new_n9007_), .C(new_n8979_), .D(new_n8973_), .Y(new_n9470_));
  NAND2X1  g09278(.A(new_n8980_), .B(new_n8999_), .Y(new_n9471_));
  OAI21X1  g09279(.A0(new_n9471_), .A1(new_n9353_), .B0(new_n8979_), .Y(new_n9472_));
  AND2X1   g09280(.A(new_n9472_), .B(new_n9470_), .Y(new_n9473_));
  INVX1    g09281(.A(new_n9473_), .Y(new_n9474_));
  NAND3X1  g09282(.A(new_n9468_), .B(new_n9459_), .C(new_n5541_), .Y(new_n9475_));
  AOI21X1  g09283(.A0(new_n9475_), .A1(new_n9474_), .B0(new_n9469_), .Y(new_n9476_));
  OR2X1    g09284(.A(new_n9476_), .B(new_n5176_), .Y(new_n9477_));
  AND2X1   g09285(.A(new_n9475_), .B(new_n9474_), .Y(new_n9478_));
  OAI21X1  g09286(.A0(new_n9000_), .A1(new_n8983_), .B0(new_n8988_), .Y(new_n9479_));
  NOR3X1   g09287(.A(new_n9479_), .B(new_n9353_), .C(new_n9021_), .Y(new_n9480_));
  AOI22X1  g09288(.A0(new_n9023_), .A1(new_n9022_), .B0(new_n9008_), .B1(\asqrt[35] ), .Y(new_n9481_));
  AOI21X1  g09289(.A0(new_n9481_), .A1(\asqrt[26] ), .B0(new_n8988_), .Y(new_n9482_));
  NOR2X1   g09290(.A(new_n9482_), .B(new_n9480_), .Y(new_n9483_));
  INVX1    g09291(.A(new_n9483_), .Y(new_n9484_));
  OR2X1    g09292(.A(new_n9469_), .B(\asqrt[36] ), .Y(new_n9485_));
  OAI21X1  g09293(.A0(new_n9485_), .A1(new_n9478_), .B0(new_n9484_), .Y(new_n9486_));
  AOI21X1  g09294(.A0(new_n9486_), .A1(new_n9477_), .B0(new_n4826_), .Y(new_n9487_));
  AND2X1   g09295(.A(new_n9009_), .B(new_n9001_), .Y(new_n9488_));
  NOR4X1   g09296(.A(new_n9353_), .B(new_n9488_), .C(new_n9026_), .D(new_n9002_), .Y(new_n9489_));
  NOR2X1   g09297(.A(new_n9488_), .B(new_n9002_), .Y(new_n9490_));
  AOI21X1  g09298(.A0(new_n9490_), .A1(\asqrt[26] ), .B0(new_n9006_), .Y(new_n9491_));
  NOR2X1   g09299(.A(new_n9491_), .B(new_n9489_), .Y(new_n9492_));
  OR2X1    g09300(.A(new_n9466_), .B(new_n6294_), .Y(new_n9493_));
  AND2X1   g09301(.A(new_n9449_), .B(new_n9440_), .Y(new_n9494_));
  INVX1    g09302(.A(new_n9455_), .Y(new_n9495_));
  OR2X1    g09303(.A(new_n9456_), .B(\asqrt[33] ), .Y(new_n9496_));
  OAI21X1  g09304(.A0(new_n9496_), .A1(new_n9494_), .B0(new_n9495_), .Y(new_n9497_));
  AOI21X1  g09305(.A0(new_n9497_), .A1(new_n9493_), .B0(new_n5941_), .Y(new_n9498_));
  AOI21X1  g09306(.A0(new_n9438_), .A1(\asqrt[33] ), .B0(\asqrt[34] ), .Y(new_n9499_));
  AOI21X1  g09307(.A0(new_n9499_), .A1(new_n9497_), .B0(new_n9464_), .Y(new_n9500_));
  OAI21X1  g09308(.A0(new_n9500_), .A1(new_n9498_), .B0(\asqrt[35] ), .Y(new_n9501_));
  NOR3X1   g09309(.A(new_n9500_), .B(new_n9498_), .C(\asqrt[35] ), .Y(new_n9502_));
  OAI21X1  g09310(.A0(new_n9502_), .A1(new_n9473_), .B0(new_n9501_), .Y(new_n9503_));
  AOI21X1  g09311(.A0(new_n9503_), .A1(\asqrt[36] ), .B0(\asqrt[37] ), .Y(new_n9504_));
  AOI21X1  g09312(.A0(new_n9504_), .A1(new_n9486_), .B0(new_n9492_), .Y(new_n9505_));
  OAI21X1  g09313(.A0(new_n9505_), .A1(new_n9487_), .B0(\asqrt[38] ), .Y(new_n9506_));
  OR4X1    g09314(.A(new_n9353_), .B(new_n9017_), .C(new_n9020_), .D(new_n9044_), .Y(new_n9507_));
  NAND2X1  g09315(.A(new_n9029_), .B(new_n9011_), .Y(new_n9508_));
  OAI21X1  g09316(.A0(new_n9508_), .A1(new_n9353_), .B0(new_n9020_), .Y(new_n9509_));
  AND2X1   g09317(.A(new_n9509_), .B(new_n9507_), .Y(new_n9510_));
  NOR3X1   g09318(.A(new_n9505_), .B(new_n9487_), .C(\asqrt[38] ), .Y(new_n9511_));
  OAI21X1  g09319(.A0(new_n9511_), .A1(new_n9510_), .B0(new_n9506_), .Y(new_n9512_));
  AND2X1   g09320(.A(new_n9512_), .B(\asqrt[39] ), .Y(new_n9513_));
  INVX1    g09321(.A(new_n9510_), .Y(new_n9514_));
  AND2X1   g09322(.A(new_n9503_), .B(\asqrt[36] ), .Y(new_n9515_));
  NAND2X1  g09323(.A(new_n9475_), .B(new_n9474_), .Y(new_n9516_));
  NOR2X1   g09324(.A(new_n9469_), .B(\asqrt[36] ), .Y(new_n9517_));
  AOI21X1  g09325(.A0(new_n9517_), .A1(new_n9516_), .B0(new_n9483_), .Y(new_n9518_));
  OAI21X1  g09326(.A0(new_n9518_), .A1(new_n9515_), .B0(\asqrt[37] ), .Y(new_n9519_));
  INVX1    g09327(.A(new_n9492_), .Y(new_n9520_));
  OAI21X1  g09328(.A0(new_n9476_), .A1(new_n5176_), .B0(new_n4826_), .Y(new_n9521_));
  OAI21X1  g09329(.A0(new_n9521_), .A1(new_n9518_), .B0(new_n9520_), .Y(new_n9522_));
  NAND3X1  g09330(.A(new_n9522_), .B(new_n9519_), .C(new_n4493_), .Y(new_n9523_));
  NAND2X1  g09331(.A(new_n9523_), .B(new_n9514_), .Y(new_n9524_));
  AOI21X1  g09332(.A0(new_n9522_), .A1(new_n9519_), .B0(new_n4493_), .Y(new_n9525_));
  NOR2X1   g09333(.A(new_n9525_), .B(\asqrt[39] ), .Y(new_n9526_));
  AND2X1   g09334(.A(new_n9031_), .B(new_n9030_), .Y(new_n9527_));
  NOR4X1   g09335(.A(new_n9353_), .B(new_n9068_), .C(new_n9527_), .D(new_n9019_), .Y(new_n9528_));
  AOI22X1  g09336(.A0(new_n9031_), .A1(new_n9030_), .B0(new_n9018_), .B1(\asqrt[38] ), .Y(new_n9529_));
  AOI21X1  g09337(.A0(new_n9529_), .A1(\asqrt[26] ), .B0(new_n9036_), .Y(new_n9530_));
  NOR2X1   g09338(.A(new_n9530_), .B(new_n9528_), .Y(new_n9531_));
  AOI21X1  g09339(.A0(new_n9526_), .A1(new_n9524_), .B0(new_n9531_), .Y(new_n9532_));
  OAI21X1  g09340(.A0(new_n9532_), .A1(new_n9513_), .B0(\asqrt[40] ), .Y(new_n9533_));
  AND2X1   g09341(.A(new_n9071_), .B(new_n9069_), .Y(new_n9534_));
  OR4X1    g09342(.A(new_n9353_), .B(new_n9534_), .C(new_n9043_), .D(new_n9070_), .Y(new_n9535_));
  OR2X1    g09343(.A(new_n9534_), .B(new_n9070_), .Y(new_n9536_));
  OAI21X1  g09344(.A0(new_n9536_), .A1(new_n9353_), .B0(new_n9043_), .Y(new_n9537_));
  AND2X1   g09345(.A(new_n9537_), .B(new_n9535_), .Y(new_n9538_));
  INVX1    g09346(.A(new_n9538_), .Y(new_n9539_));
  AOI21X1  g09347(.A0(new_n9523_), .A1(new_n9514_), .B0(new_n9525_), .Y(new_n9540_));
  OAI21X1  g09348(.A0(new_n9540_), .A1(new_n4165_), .B0(new_n3863_), .Y(new_n9541_));
  OAI21X1  g09349(.A0(new_n9541_), .A1(new_n9532_), .B0(new_n9539_), .Y(new_n9542_));
  AOI21X1  g09350(.A0(new_n9542_), .A1(new_n9533_), .B0(new_n3564_), .Y(new_n9543_));
  OR4X1    g09351(.A(new_n9353_), .B(new_n9081_), .C(new_n9054_), .D(new_n9048_), .Y(new_n9544_));
  NAND2X1  g09352(.A(new_n9055_), .B(new_n9073_), .Y(new_n9545_));
  OAI21X1  g09353(.A0(new_n9545_), .A1(new_n9353_), .B0(new_n9054_), .Y(new_n9546_));
  AND2X1   g09354(.A(new_n9546_), .B(new_n9544_), .Y(new_n9547_));
  INVX1    g09355(.A(new_n9547_), .Y(new_n9548_));
  NAND3X1  g09356(.A(new_n9542_), .B(new_n9533_), .C(new_n3564_), .Y(new_n9549_));
  AOI21X1  g09357(.A0(new_n9549_), .A1(new_n9548_), .B0(new_n9543_), .Y(new_n9550_));
  OR2X1    g09358(.A(new_n9550_), .B(new_n3276_), .Y(new_n9551_));
  AND2X1   g09359(.A(new_n9549_), .B(new_n9548_), .Y(new_n9552_));
  OAI21X1  g09360(.A0(new_n9074_), .A1(new_n9058_), .B0(new_n9063_), .Y(new_n9553_));
  NOR3X1   g09361(.A(new_n9553_), .B(new_n9353_), .C(new_n9095_), .Y(new_n9554_));
  AOI22X1  g09362(.A0(new_n9097_), .A1(new_n9096_), .B0(new_n9082_), .B1(\asqrt[41] ), .Y(new_n9555_));
  AOI21X1  g09363(.A0(new_n9555_), .A1(\asqrt[26] ), .B0(new_n9063_), .Y(new_n9556_));
  NOR2X1   g09364(.A(new_n9556_), .B(new_n9554_), .Y(new_n9557_));
  INVX1    g09365(.A(new_n9557_), .Y(new_n9558_));
  OR2X1    g09366(.A(new_n9543_), .B(\asqrt[42] ), .Y(new_n9559_));
  OAI21X1  g09367(.A0(new_n9559_), .A1(new_n9552_), .B0(new_n9558_), .Y(new_n9560_));
  AOI21X1  g09368(.A0(new_n9560_), .A1(new_n9551_), .B0(new_n3008_), .Y(new_n9561_));
  AND2X1   g09369(.A(new_n9083_), .B(new_n9075_), .Y(new_n9562_));
  OR2X1    g09370(.A(new_n9100_), .B(new_n9076_), .Y(new_n9563_));
  OR2X1    g09371(.A(new_n9563_), .B(new_n9562_), .Y(new_n9564_));
  NOR3X1   g09372(.A(new_n9353_), .B(new_n9562_), .C(new_n9076_), .Y(new_n9565_));
  OAI22X1  g09373(.A0(new_n9565_), .A1(new_n9080_), .B0(new_n9564_), .B1(new_n9353_), .Y(new_n9566_));
  INVX1    g09374(.A(new_n9566_), .Y(new_n9567_));
  OR2X1    g09375(.A(new_n9540_), .B(new_n4165_), .Y(new_n9568_));
  AND2X1   g09376(.A(new_n9523_), .B(new_n9514_), .Y(new_n9569_));
  OR2X1    g09377(.A(new_n9525_), .B(\asqrt[39] ), .Y(new_n9570_));
  INVX1    g09378(.A(new_n9531_), .Y(new_n9571_));
  OAI21X1  g09379(.A0(new_n9570_), .A1(new_n9569_), .B0(new_n9571_), .Y(new_n9572_));
  AOI21X1  g09380(.A0(new_n9572_), .A1(new_n9568_), .B0(new_n3863_), .Y(new_n9573_));
  AOI21X1  g09381(.A0(new_n9512_), .A1(\asqrt[39] ), .B0(\asqrt[40] ), .Y(new_n9574_));
  AOI21X1  g09382(.A0(new_n9574_), .A1(new_n9572_), .B0(new_n9538_), .Y(new_n9575_));
  OAI21X1  g09383(.A0(new_n9575_), .A1(new_n9573_), .B0(\asqrt[41] ), .Y(new_n9576_));
  NOR3X1   g09384(.A(new_n9575_), .B(new_n9573_), .C(\asqrt[41] ), .Y(new_n9577_));
  OAI21X1  g09385(.A0(new_n9577_), .A1(new_n9547_), .B0(new_n9576_), .Y(new_n9578_));
  AOI21X1  g09386(.A0(new_n9578_), .A1(\asqrt[42] ), .B0(\asqrt[43] ), .Y(new_n9579_));
  AOI21X1  g09387(.A0(new_n9579_), .A1(new_n9560_), .B0(new_n9567_), .Y(new_n9580_));
  OAI21X1  g09388(.A0(new_n9580_), .A1(new_n9561_), .B0(\asqrt[44] ), .Y(new_n9581_));
  OR4X1    g09389(.A(new_n9353_), .B(new_n9091_), .C(new_n9094_), .D(new_n9118_), .Y(new_n9582_));
  NAND2X1  g09390(.A(new_n9103_), .B(new_n9085_), .Y(new_n9583_));
  OAI21X1  g09391(.A0(new_n9583_), .A1(new_n9353_), .B0(new_n9094_), .Y(new_n9584_));
  AND2X1   g09392(.A(new_n9584_), .B(new_n9582_), .Y(new_n9585_));
  NOR3X1   g09393(.A(new_n9580_), .B(new_n9561_), .C(\asqrt[44] ), .Y(new_n9586_));
  OAI21X1  g09394(.A0(new_n9586_), .A1(new_n9585_), .B0(new_n9581_), .Y(new_n9587_));
  AND2X1   g09395(.A(new_n9587_), .B(\asqrt[45] ), .Y(new_n9588_));
  INVX1    g09396(.A(new_n9585_), .Y(new_n9589_));
  AND2X1   g09397(.A(new_n9578_), .B(\asqrt[42] ), .Y(new_n9590_));
  NAND2X1  g09398(.A(new_n9549_), .B(new_n9548_), .Y(new_n9591_));
  NOR2X1   g09399(.A(new_n9543_), .B(\asqrt[42] ), .Y(new_n9592_));
  AOI21X1  g09400(.A0(new_n9592_), .A1(new_n9591_), .B0(new_n9557_), .Y(new_n9593_));
  OAI21X1  g09401(.A0(new_n9593_), .A1(new_n9590_), .B0(\asqrt[43] ), .Y(new_n9594_));
  OAI21X1  g09402(.A0(new_n9550_), .A1(new_n3276_), .B0(new_n3008_), .Y(new_n9595_));
  OAI21X1  g09403(.A0(new_n9595_), .A1(new_n9593_), .B0(new_n9566_), .Y(new_n9596_));
  NAND3X1  g09404(.A(new_n9596_), .B(new_n9594_), .C(new_n2769_), .Y(new_n9597_));
  NAND2X1  g09405(.A(new_n9597_), .B(new_n9589_), .Y(new_n9598_));
  AND2X1   g09406(.A(new_n9110_), .B(new_n9104_), .Y(new_n9599_));
  NOR4X1   g09407(.A(new_n9353_), .B(new_n9599_), .C(new_n9141_), .D(new_n9093_), .Y(new_n9600_));
  AOI22X1  g09408(.A0(new_n9110_), .A1(new_n9104_), .B0(new_n9092_), .B1(\asqrt[44] ), .Y(new_n9601_));
  AOI21X1  g09409(.A0(new_n9601_), .A1(\asqrt[26] ), .B0(new_n9109_), .Y(new_n9602_));
  NOR2X1   g09410(.A(new_n9602_), .B(new_n9600_), .Y(new_n9603_));
  AOI21X1  g09411(.A0(new_n9596_), .A1(new_n9594_), .B0(new_n2769_), .Y(new_n9604_));
  NOR2X1   g09412(.A(new_n9604_), .B(\asqrt[45] ), .Y(new_n9605_));
  AOI21X1  g09413(.A0(new_n9605_), .A1(new_n9598_), .B0(new_n9603_), .Y(new_n9606_));
  OAI21X1  g09414(.A0(new_n9606_), .A1(new_n9588_), .B0(\asqrt[46] ), .Y(new_n9607_));
  OAI21X1  g09415(.A0(new_n9120_), .A1(new_n9111_), .B0(new_n9116_), .Y(new_n9608_));
  OR2X1    g09416(.A(new_n9608_), .B(new_n9144_), .Y(new_n9609_));
  AND2X1   g09417(.A(new_n9145_), .B(new_n9143_), .Y(new_n9610_));
  NOR3X1   g09418(.A(new_n9353_), .B(new_n9610_), .C(new_n9144_), .Y(new_n9611_));
  OAI22X1  g09419(.A0(new_n9611_), .A1(new_n9116_), .B0(new_n9609_), .B1(new_n9353_), .Y(new_n9612_));
  AOI21X1  g09420(.A0(new_n9597_), .A1(new_n9589_), .B0(new_n9604_), .Y(new_n9613_));
  OAI21X1  g09421(.A0(new_n9613_), .A1(new_n2570_), .B0(new_n2263_), .Y(new_n9614_));
  OAI21X1  g09422(.A0(new_n9614_), .A1(new_n9606_), .B0(new_n9612_), .Y(new_n9615_));
  AOI21X1  g09423(.A0(new_n9615_), .A1(new_n9607_), .B0(new_n2040_), .Y(new_n9616_));
  OR4X1    g09424(.A(new_n9353_), .B(new_n9155_), .C(new_n9128_), .D(new_n9122_), .Y(new_n9617_));
  NAND2X1  g09425(.A(new_n9129_), .B(new_n9147_), .Y(new_n9618_));
  OAI21X1  g09426(.A0(new_n9618_), .A1(new_n9353_), .B0(new_n9128_), .Y(new_n9619_));
  AND2X1   g09427(.A(new_n9619_), .B(new_n9617_), .Y(new_n9620_));
  INVX1    g09428(.A(new_n9620_), .Y(new_n9621_));
  NAND3X1  g09429(.A(new_n9615_), .B(new_n9607_), .C(new_n2040_), .Y(new_n9622_));
  AOI21X1  g09430(.A0(new_n9622_), .A1(new_n9621_), .B0(new_n9616_), .Y(new_n9623_));
  OR2X1    g09431(.A(new_n9623_), .B(new_n1834_), .Y(new_n9624_));
  AND2X1   g09432(.A(new_n9622_), .B(new_n9621_), .Y(new_n9625_));
  OAI21X1  g09433(.A0(new_n9148_), .A1(new_n9132_), .B0(new_n9137_), .Y(new_n9626_));
  NOR3X1   g09434(.A(new_n9626_), .B(new_n9353_), .C(new_n9169_), .Y(new_n9627_));
  AOI22X1  g09435(.A0(new_n9171_), .A1(new_n9170_), .B0(new_n9156_), .B1(\asqrt[47] ), .Y(new_n9628_));
  AOI21X1  g09436(.A0(new_n9628_), .A1(\asqrt[26] ), .B0(new_n9137_), .Y(new_n9629_));
  NOR2X1   g09437(.A(new_n9629_), .B(new_n9627_), .Y(new_n9630_));
  INVX1    g09438(.A(new_n9630_), .Y(new_n9631_));
  OR2X1    g09439(.A(new_n9616_), .B(\asqrt[48] ), .Y(new_n9632_));
  OAI21X1  g09440(.A0(new_n9632_), .A1(new_n9625_), .B0(new_n9631_), .Y(new_n9633_));
  AOI21X1  g09441(.A0(new_n9633_), .A1(new_n9624_), .B0(new_n1632_), .Y(new_n9634_));
  AND2X1   g09442(.A(new_n9157_), .B(new_n9149_), .Y(new_n9635_));
  OR4X1    g09443(.A(new_n9353_), .B(new_n9635_), .C(new_n9174_), .D(new_n9150_), .Y(new_n9636_));
  OR2X1    g09444(.A(new_n9635_), .B(new_n9150_), .Y(new_n9637_));
  OAI21X1  g09445(.A0(new_n9637_), .A1(new_n9353_), .B0(new_n9174_), .Y(new_n9638_));
  AND2X1   g09446(.A(new_n9638_), .B(new_n9636_), .Y(new_n9639_));
  OR2X1    g09447(.A(new_n9613_), .B(new_n2570_), .Y(new_n9640_));
  AND2X1   g09448(.A(new_n9597_), .B(new_n9589_), .Y(new_n9641_));
  INVX1    g09449(.A(new_n9603_), .Y(new_n9642_));
  OR2X1    g09450(.A(new_n9604_), .B(\asqrt[45] ), .Y(new_n9643_));
  OAI21X1  g09451(.A0(new_n9643_), .A1(new_n9641_), .B0(new_n9642_), .Y(new_n9644_));
  AOI21X1  g09452(.A0(new_n9644_), .A1(new_n9640_), .B0(new_n2263_), .Y(new_n9645_));
  INVX1    g09453(.A(new_n9612_), .Y(new_n9646_));
  AOI21X1  g09454(.A0(new_n9587_), .A1(\asqrt[45] ), .B0(\asqrt[46] ), .Y(new_n9647_));
  AOI21X1  g09455(.A0(new_n9647_), .A1(new_n9644_), .B0(new_n9646_), .Y(new_n9648_));
  OAI21X1  g09456(.A0(new_n9648_), .A1(new_n9645_), .B0(\asqrt[47] ), .Y(new_n9649_));
  NOR3X1   g09457(.A(new_n9648_), .B(new_n9645_), .C(\asqrt[47] ), .Y(new_n9650_));
  OAI21X1  g09458(.A0(new_n9650_), .A1(new_n9620_), .B0(new_n9649_), .Y(new_n9651_));
  AOI21X1  g09459(.A0(new_n9651_), .A1(\asqrt[48] ), .B0(\asqrt[49] ), .Y(new_n9652_));
  AOI21X1  g09460(.A0(new_n9652_), .A1(new_n9633_), .B0(new_n9639_), .Y(new_n9653_));
  OAI21X1  g09461(.A0(new_n9653_), .A1(new_n9634_), .B0(\asqrt[50] ), .Y(new_n9654_));
  OR4X1    g09462(.A(new_n9353_), .B(new_n9165_), .C(new_n9168_), .D(new_n9192_), .Y(new_n9655_));
  NAND2X1  g09463(.A(new_n9177_), .B(new_n9159_), .Y(new_n9656_));
  OAI21X1  g09464(.A0(new_n9656_), .A1(new_n9353_), .B0(new_n9168_), .Y(new_n9657_));
  AND2X1   g09465(.A(new_n9657_), .B(new_n9655_), .Y(new_n9658_));
  NOR3X1   g09466(.A(new_n9653_), .B(new_n9634_), .C(\asqrt[50] ), .Y(new_n9659_));
  OAI21X1  g09467(.A0(new_n9659_), .A1(new_n9658_), .B0(new_n9654_), .Y(new_n9660_));
  AND2X1   g09468(.A(new_n9660_), .B(\asqrt[51] ), .Y(new_n9661_));
  OR2X1    g09469(.A(new_n9659_), .B(new_n9658_), .Y(new_n9662_));
  AND2X1   g09470(.A(new_n9184_), .B(new_n9178_), .Y(new_n9663_));
  NOR4X1   g09471(.A(new_n9353_), .B(new_n9663_), .C(new_n9215_), .D(new_n9167_), .Y(new_n9664_));
  AOI22X1  g09472(.A0(new_n9184_), .A1(new_n9178_), .B0(new_n9166_), .B1(\asqrt[50] ), .Y(new_n9665_));
  AOI21X1  g09473(.A0(new_n9665_), .A1(\asqrt[26] ), .B0(new_n9183_), .Y(new_n9666_));
  NOR2X1   g09474(.A(new_n9666_), .B(new_n9664_), .Y(new_n9667_));
  AND2X1   g09475(.A(new_n9654_), .B(new_n1277_), .Y(new_n9668_));
  AOI21X1  g09476(.A0(new_n9668_), .A1(new_n9662_), .B0(new_n9667_), .Y(new_n9669_));
  OAI21X1  g09477(.A0(new_n9669_), .A1(new_n9661_), .B0(\asqrt[52] ), .Y(new_n9670_));
  AND2X1   g09478(.A(new_n9219_), .B(new_n9217_), .Y(new_n9671_));
  OR4X1    g09479(.A(new_n9353_), .B(new_n9671_), .C(new_n9191_), .D(new_n9218_), .Y(new_n9672_));
  OR2X1    g09480(.A(new_n9671_), .B(new_n9218_), .Y(new_n9673_));
  OAI21X1  g09481(.A0(new_n9673_), .A1(new_n9353_), .B0(new_n9191_), .Y(new_n9674_));
  AND2X1   g09482(.A(new_n9674_), .B(new_n9672_), .Y(new_n9675_));
  INVX1    g09483(.A(new_n9675_), .Y(new_n9676_));
  AND2X1   g09484(.A(new_n9651_), .B(\asqrt[48] ), .Y(new_n9677_));
  NAND2X1  g09485(.A(new_n9622_), .B(new_n9621_), .Y(new_n9678_));
  NOR2X1   g09486(.A(new_n9616_), .B(\asqrt[48] ), .Y(new_n9679_));
  AOI21X1  g09487(.A0(new_n9679_), .A1(new_n9678_), .B0(new_n9630_), .Y(new_n9680_));
  OAI21X1  g09488(.A0(new_n9680_), .A1(new_n9677_), .B0(\asqrt[49] ), .Y(new_n9681_));
  INVX1    g09489(.A(new_n9639_), .Y(new_n9682_));
  OAI21X1  g09490(.A0(new_n9623_), .A1(new_n1834_), .B0(new_n1632_), .Y(new_n9683_));
  OAI21X1  g09491(.A0(new_n9683_), .A1(new_n9680_), .B0(new_n9682_), .Y(new_n9684_));
  AOI21X1  g09492(.A0(new_n9684_), .A1(new_n9681_), .B0(new_n1469_), .Y(new_n9685_));
  INVX1    g09493(.A(new_n9658_), .Y(new_n9686_));
  NAND3X1  g09494(.A(new_n9684_), .B(new_n9681_), .C(new_n1469_), .Y(new_n9687_));
  AOI21X1  g09495(.A0(new_n9687_), .A1(new_n9686_), .B0(new_n9685_), .Y(new_n9688_));
  OAI21X1  g09496(.A0(new_n9688_), .A1(new_n1277_), .B0(new_n1111_), .Y(new_n9689_));
  OAI21X1  g09497(.A0(new_n9689_), .A1(new_n9669_), .B0(new_n9676_), .Y(new_n9690_));
  AOI21X1  g09498(.A0(new_n9690_), .A1(new_n9670_), .B0(new_n968_), .Y(new_n9691_));
  NAND3X1  g09499(.A(new_n9203_), .B(new_n9201_), .C(new_n9221_), .Y(new_n9692_));
  NOR3X1   g09500(.A(new_n9353_), .B(new_n9229_), .C(new_n9196_), .Y(new_n9693_));
  OAI22X1  g09501(.A0(new_n9693_), .A1(new_n9201_), .B0(new_n9692_), .B1(new_n9353_), .Y(new_n9694_));
  NAND3X1  g09502(.A(new_n9690_), .B(new_n9670_), .C(new_n968_), .Y(new_n9695_));
  AOI21X1  g09503(.A0(new_n9695_), .A1(new_n9694_), .B0(new_n9691_), .Y(new_n9696_));
  OR2X1    g09504(.A(new_n9696_), .B(new_n902_), .Y(new_n9697_));
  AND2X1   g09505(.A(new_n9695_), .B(new_n9694_), .Y(new_n9698_));
  OAI21X1  g09506(.A0(new_n9222_), .A1(new_n9206_), .B0(new_n9211_), .Y(new_n9699_));
  NOR3X1   g09507(.A(new_n9699_), .B(new_n9353_), .C(new_n9256_), .Y(new_n9700_));
  AOI22X1  g09508(.A0(new_n9258_), .A1(new_n9257_), .B0(new_n9230_), .B1(\asqrt[53] ), .Y(new_n9701_));
  AOI21X1  g09509(.A0(new_n9701_), .A1(\asqrt[26] ), .B0(new_n9211_), .Y(new_n9702_));
  NOR2X1   g09510(.A(new_n9702_), .B(new_n9700_), .Y(new_n9703_));
  INVX1    g09511(.A(new_n9703_), .Y(new_n9704_));
  OR2X1    g09512(.A(new_n9688_), .B(new_n1277_), .Y(new_n9705_));
  NOR2X1   g09513(.A(new_n9659_), .B(new_n9658_), .Y(new_n9706_));
  INVX1    g09514(.A(new_n9667_), .Y(new_n9707_));
  NAND2X1  g09515(.A(new_n9654_), .B(new_n1277_), .Y(new_n9708_));
  OAI21X1  g09516(.A0(new_n9708_), .A1(new_n9706_), .B0(new_n9707_), .Y(new_n9709_));
  AOI21X1  g09517(.A0(new_n9709_), .A1(new_n9705_), .B0(new_n1111_), .Y(new_n9710_));
  AOI21X1  g09518(.A0(new_n9660_), .A1(\asqrt[51] ), .B0(\asqrt[52] ), .Y(new_n9711_));
  AOI21X1  g09519(.A0(new_n9711_), .A1(new_n9709_), .B0(new_n9675_), .Y(new_n9712_));
  OAI21X1  g09520(.A0(new_n9712_), .A1(new_n9710_), .B0(\asqrt[53] ), .Y(new_n9713_));
  NAND2X1  g09521(.A(new_n9713_), .B(new_n902_), .Y(new_n9714_));
  OAI21X1  g09522(.A0(new_n9714_), .A1(new_n9698_), .B0(new_n9704_), .Y(new_n9715_));
  AOI21X1  g09523(.A0(new_n9715_), .A1(new_n9697_), .B0(new_n697_), .Y(new_n9716_));
  AND2X1   g09524(.A(new_n9231_), .B(new_n9223_), .Y(new_n9717_));
  OR4X1    g09525(.A(new_n9353_), .B(new_n9717_), .C(new_n9261_), .D(new_n9224_), .Y(new_n9718_));
  OR2X1    g09526(.A(new_n9717_), .B(new_n9224_), .Y(new_n9719_));
  OAI21X1  g09527(.A0(new_n9719_), .A1(new_n9353_), .B0(new_n9261_), .Y(new_n9720_));
  AND2X1   g09528(.A(new_n9720_), .B(new_n9718_), .Y(new_n9721_));
  INVX1    g09529(.A(new_n9694_), .Y(new_n9722_));
  NOR3X1   g09530(.A(new_n9712_), .B(new_n9710_), .C(\asqrt[53] ), .Y(new_n9723_));
  OAI21X1  g09531(.A0(new_n9723_), .A1(new_n9722_), .B0(new_n9713_), .Y(new_n9724_));
  AOI21X1  g09532(.A0(new_n9724_), .A1(\asqrt[54] ), .B0(\asqrt[55] ), .Y(new_n9725_));
  AOI21X1  g09533(.A0(new_n9725_), .A1(new_n9715_), .B0(new_n9721_), .Y(new_n9726_));
  OAI21X1  g09534(.A0(new_n9726_), .A1(new_n9716_), .B0(\asqrt[56] ), .Y(new_n9727_));
  OR4X1    g09535(.A(new_n9353_), .B(new_n9239_), .C(new_n9265_), .D(new_n9264_), .Y(new_n9728_));
  OR2X1    g09536(.A(new_n9239_), .B(new_n9264_), .Y(new_n9729_));
  OAI21X1  g09537(.A0(new_n9729_), .A1(new_n9353_), .B0(new_n9265_), .Y(new_n9730_));
  AND2X1   g09538(.A(new_n9730_), .B(new_n9728_), .Y(new_n9731_));
  NOR3X1   g09539(.A(new_n9726_), .B(new_n9716_), .C(\asqrt[56] ), .Y(new_n9732_));
  OAI21X1  g09540(.A0(new_n9732_), .A1(new_n9731_), .B0(new_n9727_), .Y(new_n9733_));
  AND2X1   g09541(.A(new_n9733_), .B(\asqrt[57] ), .Y(new_n9734_));
  OR2X1    g09542(.A(new_n9732_), .B(new_n9731_), .Y(new_n9735_));
  AND2X1   g09543(.A(new_n9248_), .B(new_n9242_), .Y(new_n9736_));
  NOR4X1   g09544(.A(new_n9353_), .B(new_n9736_), .C(new_n9289_), .D(new_n9241_), .Y(new_n9737_));
  AOI22X1  g09545(.A0(new_n9248_), .A1(new_n9242_), .B0(new_n9240_), .B1(\asqrt[56] ), .Y(new_n9738_));
  AOI21X1  g09546(.A0(new_n9738_), .A1(\asqrt[26] ), .B0(new_n9247_), .Y(new_n9739_));
  NOR2X1   g09547(.A(new_n9739_), .B(new_n9737_), .Y(new_n9740_));
  AND2X1   g09548(.A(new_n9727_), .B(new_n481_), .Y(new_n9741_));
  AOI21X1  g09549(.A0(new_n9741_), .A1(new_n9735_), .B0(new_n9740_), .Y(new_n9742_));
  OAI21X1  g09550(.A0(new_n9742_), .A1(new_n9734_), .B0(\asqrt[58] ), .Y(new_n9743_));
  AND2X1   g09551(.A(new_n9293_), .B(new_n9291_), .Y(new_n9744_));
  OR4X1    g09552(.A(new_n9353_), .B(new_n9744_), .C(new_n9255_), .D(new_n9292_), .Y(new_n9745_));
  OR2X1    g09553(.A(new_n9744_), .B(new_n9292_), .Y(new_n9746_));
  OAI21X1  g09554(.A0(new_n9746_), .A1(new_n9353_), .B0(new_n9255_), .Y(new_n9747_));
  AND2X1   g09555(.A(new_n9747_), .B(new_n9745_), .Y(new_n9748_));
  INVX1    g09556(.A(new_n9748_), .Y(new_n9749_));
  AND2X1   g09557(.A(new_n9724_), .B(\asqrt[54] ), .Y(new_n9750_));
  NAND2X1  g09558(.A(new_n9695_), .B(new_n9694_), .Y(new_n9751_));
  AND2X1   g09559(.A(new_n9713_), .B(new_n902_), .Y(new_n9752_));
  AOI21X1  g09560(.A0(new_n9752_), .A1(new_n9751_), .B0(new_n9703_), .Y(new_n9753_));
  OAI21X1  g09561(.A0(new_n9753_), .A1(new_n9750_), .B0(\asqrt[55] ), .Y(new_n9754_));
  INVX1    g09562(.A(new_n9721_), .Y(new_n9755_));
  OAI21X1  g09563(.A0(new_n9696_), .A1(new_n902_), .B0(new_n697_), .Y(new_n9756_));
  OAI21X1  g09564(.A0(new_n9756_), .A1(new_n9753_), .B0(new_n9755_), .Y(new_n9757_));
  AOI21X1  g09565(.A0(new_n9757_), .A1(new_n9754_), .B0(new_n582_), .Y(new_n9758_));
  INVX1    g09566(.A(new_n9731_), .Y(new_n9759_));
  NAND3X1  g09567(.A(new_n9757_), .B(new_n9754_), .C(new_n582_), .Y(new_n9760_));
  AOI21X1  g09568(.A0(new_n9760_), .A1(new_n9759_), .B0(new_n9758_), .Y(new_n9761_));
  OAI21X1  g09569(.A0(new_n9761_), .A1(new_n481_), .B0(new_n399_), .Y(new_n9762_));
  OAI21X1  g09570(.A0(new_n9762_), .A1(new_n9742_), .B0(new_n9749_), .Y(new_n9763_));
  AOI21X1  g09571(.A0(new_n9763_), .A1(new_n9743_), .B0(new_n328_), .Y(new_n9764_));
  OR4X1    g09572(.A(new_n9353_), .B(new_n9303_), .C(new_n9276_), .D(new_n9270_), .Y(new_n9765_));
  OR2X1    g09573(.A(new_n9303_), .B(new_n9270_), .Y(new_n9766_));
  OAI21X1  g09574(.A0(new_n9766_), .A1(new_n9353_), .B0(new_n9276_), .Y(new_n9767_));
  AND2X1   g09575(.A(new_n9767_), .B(new_n9765_), .Y(new_n9768_));
  INVX1    g09576(.A(new_n9768_), .Y(new_n9769_));
  NAND3X1  g09577(.A(new_n9763_), .B(new_n9743_), .C(new_n328_), .Y(new_n9770_));
  AOI21X1  g09578(.A0(new_n9770_), .A1(new_n9769_), .B0(new_n9764_), .Y(new_n9771_));
  OR2X1    g09579(.A(new_n9771_), .B(new_n292_), .Y(new_n9772_));
  OR2X1    g09580(.A(new_n9761_), .B(new_n481_), .Y(new_n9773_));
  NOR2X1   g09581(.A(new_n9732_), .B(new_n9731_), .Y(new_n9774_));
  INVX1    g09582(.A(new_n9740_), .Y(new_n9775_));
  NAND2X1  g09583(.A(new_n9727_), .B(new_n481_), .Y(new_n9776_));
  OAI21X1  g09584(.A0(new_n9776_), .A1(new_n9774_), .B0(new_n9775_), .Y(new_n9777_));
  AOI21X1  g09585(.A0(new_n9777_), .A1(new_n9773_), .B0(new_n399_), .Y(new_n9778_));
  AOI21X1  g09586(.A0(new_n9733_), .A1(\asqrt[57] ), .B0(\asqrt[58] ), .Y(new_n9779_));
  AOI21X1  g09587(.A0(new_n9779_), .A1(new_n9777_), .B0(new_n9748_), .Y(new_n9780_));
  NOR3X1   g09588(.A(new_n9780_), .B(new_n9778_), .C(\asqrt[59] ), .Y(new_n9781_));
  NOR2X1   g09589(.A(new_n9781_), .B(new_n9768_), .Y(new_n9782_));
  OAI21X1  g09590(.A0(new_n9296_), .A1(new_n9280_), .B0(new_n9285_), .Y(new_n9783_));
  NOR3X1   g09591(.A(new_n9783_), .B(new_n9353_), .C(new_n9332_), .Y(new_n9784_));
  AOI22X1  g09592(.A0(new_n9334_), .A1(new_n9333_), .B0(new_n9304_), .B1(\asqrt[59] ), .Y(new_n9785_));
  AOI21X1  g09593(.A0(new_n9785_), .A1(\asqrt[26] ), .B0(new_n9285_), .Y(new_n9786_));
  NOR2X1   g09594(.A(new_n9786_), .B(new_n9784_), .Y(new_n9787_));
  INVX1    g09595(.A(new_n9787_), .Y(new_n9788_));
  OAI21X1  g09596(.A0(new_n9780_), .A1(new_n9778_), .B0(\asqrt[59] ), .Y(new_n9789_));
  NAND2X1  g09597(.A(new_n9789_), .B(new_n292_), .Y(new_n9790_));
  OAI21X1  g09598(.A0(new_n9790_), .A1(new_n9782_), .B0(new_n9788_), .Y(new_n9791_));
  AOI21X1  g09599(.A0(new_n9791_), .A1(new_n9772_), .B0(new_n217_), .Y(new_n9792_));
  AND2X1   g09600(.A(new_n9305_), .B(new_n9297_), .Y(new_n9793_));
  OR4X1    g09601(.A(new_n9353_), .B(new_n9793_), .C(new_n9337_), .D(new_n9298_), .Y(new_n9794_));
  OR2X1    g09602(.A(new_n9793_), .B(new_n9298_), .Y(new_n9795_));
  OAI21X1  g09603(.A0(new_n9795_), .A1(new_n9353_), .B0(new_n9337_), .Y(new_n9796_));
  AND2X1   g09604(.A(new_n9796_), .B(new_n9794_), .Y(new_n9797_));
  OAI21X1  g09605(.A0(new_n9781_), .A1(new_n9768_), .B0(new_n9789_), .Y(new_n9798_));
  AOI21X1  g09606(.A0(new_n9798_), .A1(\asqrt[60] ), .B0(\asqrt[61] ), .Y(new_n9799_));
  AOI21X1  g09607(.A0(new_n9799_), .A1(new_n9791_), .B0(new_n9797_), .Y(new_n9800_));
  OAI21X1  g09608(.A0(new_n9800_), .A1(new_n9792_), .B0(\asqrt[62] ), .Y(new_n9801_));
  OR4X1    g09609(.A(new_n9353_), .B(new_n9313_), .C(new_n9341_), .D(new_n9340_), .Y(new_n9802_));
  OR2X1    g09610(.A(new_n9313_), .B(new_n9340_), .Y(new_n9803_));
  OAI21X1  g09611(.A0(new_n9803_), .A1(new_n9353_), .B0(new_n9341_), .Y(new_n9804_));
  AND2X1   g09612(.A(new_n9804_), .B(new_n9802_), .Y(new_n9805_));
  NOR3X1   g09613(.A(new_n9800_), .B(new_n9792_), .C(\asqrt[62] ), .Y(new_n9806_));
  OAI21X1  g09614(.A0(new_n9806_), .A1(new_n9805_), .B0(new_n9801_), .Y(new_n9807_));
  AND2X1   g09615(.A(new_n9322_), .B(new_n9316_), .Y(new_n9808_));
  NOR4X1   g09616(.A(new_n9353_), .B(new_n9808_), .C(new_n9356_), .D(new_n9315_), .Y(new_n9809_));
  INVX1    g09617(.A(new_n9809_), .Y(new_n9810_));
  OAI22X1  g09618(.A0(new_n9357_), .A1(new_n9355_), .B0(new_n9343_), .B1(new_n199_), .Y(new_n9811_));
  OAI21X1  g09619(.A0(new_n9811_), .A1(new_n9353_), .B0(new_n9356_), .Y(new_n9812_));
  AND2X1   g09620(.A(new_n9812_), .B(new_n9810_), .Y(new_n9813_));
  INVX1    g09621(.A(new_n9813_), .Y(new_n9814_));
  AND2X1   g09622(.A(new_n9361_), .B(new_n9358_), .Y(new_n9815_));
  AOI21X1  g09623(.A0(new_n9358_), .A1(new_n9354_), .B0(new_n9326_), .Y(new_n9816_));
  AOI21X1  g09624(.A0(new_n9816_), .A1(\asqrt[26] ), .B0(new_n9815_), .Y(new_n9817_));
  AND2X1   g09625(.A(new_n9817_), .B(new_n9814_), .Y(new_n9818_));
  AOI21X1  g09626(.A0(new_n9818_), .A1(new_n9807_), .B0(\asqrt[63] ), .Y(new_n9819_));
  NOR2X1   g09627(.A(new_n9806_), .B(new_n9805_), .Y(new_n9820_));
  NAND2X1  g09628(.A(new_n9813_), .B(new_n9801_), .Y(new_n9821_));
  NAND2X1  g09629(.A(new_n9358_), .B(new_n9354_), .Y(new_n9822_));
  AOI21X1  g09630(.A0(\asqrt[26] ), .A1(new_n9327_), .B0(new_n9822_), .Y(new_n9823_));
  NOR3X1   g09631(.A(new_n9823_), .B(new_n9816_), .C(new_n193_), .Y(new_n9824_));
  AND2X1   g09632(.A(new_n9331_), .B(new_n193_), .Y(new_n9825_));
  INVX1    g09633(.A(new_n9350_), .Y(new_n9826_));
  OR2X1    g09634(.A(new_n9826_), .B(new_n9324_), .Y(new_n9827_));
  AOI21X1  g09635(.A0(new_n9325_), .A1(new_n8885_), .B0(new_n9827_), .Y(new_n9828_));
  NAND2X1  g09636(.A(new_n9828_), .B(new_n9347_), .Y(new_n9829_));
  NOR3X1   g09637(.A(new_n9829_), .B(new_n9815_), .C(new_n9825_), .Y(new_n9830_));
  NOR2X1   g09638(.A(new_n9830_), .B(new_n9824_), .Y(new_n9831_));
  OAI21X1  g09639(.A0(new_n9821_), .A1(new_n9820_), .B0(new_n9831_), .Y(new_n9832_));
  NOR2X1   g09640(.A(new_n9832_), .B(new_n9819_), .Y(new_n9833_));
  INVX1    g09641(.A(new_n9833_), .Y(\asqrt[25] ));
  OAI21X1  g09642(.A0(new_n9832_), .A1(new_n9819_), .B0(\a[50] ), .Y(new_n9835_));
  INVX1    g09643(.A(\a[50] ), .Y(new_n9836_));
  NOR2X1   g09644(.A(\a[49] ), .B(\a[48] ), .Y(new_n9837_));
  NAND2X1  g09645(.A(new_n9837_), .B(new_n9836_), .Y(new_n9838_));
  AND2X1   g09646(.A(new_n9838_), .B(new_n9835_), .Y(new_n9839_));
  AND2X1   g09647(.A(new_n9798_), .B(\asqrt[60] ), .Y(new_n9840_));
  OR2X1    g09648(.A(new_n9781_), .B(new_n9768_), .Y(new_n9841_));
  AND2X1   g09649(.A(new_n9789_), .B(new_n292_), .Y(new_n9842_));
  AOI21X1  g09650(.A0(new_n9842_), .A1(new_n9841_), .B0(new_n9787_), .Y(new_n9843_));
  OAI21X1  g09651(.A0(new_n9843_), .A1(new_n9840_), .B0(\asqrt[61] ), .Y(new_n9844_));
  INVX1    g09652(.A(new_n9797_), .Y(new_n9845_));
  OAI21X1  g09653(.A0(new_n9771_), .A1(new_n292_), .B0(new_n217_), .Y(new_n9846_));
  OAI21X1  g09654(.A0(new_n9846_), .A1(new_n9843_), .B0(new_n9845_), .Y(new_n9847_));
  AOI21X1  g09655(.A0(new_n9847_), .A1(new_n9844_), .B0(new_n199_), .Y(new_n9848_));
  INVX1    g09656(.A(new_n9805_), .Y(new_n9849_));
  NAND3X1  g09657(.A(new_n9847_), .B(new_n9844_), .C(new_n199_), .Y(new_n9850_));
  AOI21X1  g09658(.A0(new_n9850_), .A1(new_n9849_), .B0(new_n9848_), .Y(new_n9851_));
  INVX1    g09659(.A(new_n9818_), .Y(new_n9852_));
  OAI21X1  g09660(.A0(new_n9852_), .A1(new_n9851_), .B0(new_n193_), .Y(new_n9853_));
  OR2X1    g09661(.A(new_n9806_), .B(new_n9805_), .Y(new_n9854_));
  AND2X1   g09662(.A(new_n9813_), .B(new_n9801_), .Y(new_n9855_));
  INVX1    g09663(.A(new_n9831_), .Y(new_n9856_));
  AOI21X1  g09664(.A0(new_n9855_), .A1(new_n9854_), .B0(new_n9856_), .Y(new_n9857_));
  AOI21X1  g09665(.A0(new_n9857_), .A1(new_n9853_), .B0(new_n9836_), .Y(new_n9858_));
  NAND3X1  g09666(.A(new_n9838_), .B(new_n9350_), .C(new_n9347_), .Y(new_n9859_));
  NOR4X1   g09667(.A(new_n9859_), .B(new_n9858_), .C(new_n9815_), .D(new_n9825_), .Y(new_n9860_));
  INVX1    g09668(.A(\a[51] ), .Y(new_n9861_));
  AOI21X1  g09669(.A0(new_n9857_), .A1(new_n9853_), .B0(\a[50] ), .Y(new_n9862_));
  OAI21X1  g09670(.A0(new_n9832_), .A1(new_n9819_), .B0(new_n9365_), .Y(new_n9863_));
  OAI21X1  g09671(.A0(new_n9862_), .A1(new_n9861_), .B0(new_n9863_), .Y(new_n9864_));
  OAI22X1  g09672(.A0(new_n9864_), .A1(new_n9860_), .B0(new_n9839_), .B1(new_n9353_), .Y(new_n9865_));
  AND2X1   g09673(.A(new_n9865_), .B(\asqrt[27] ), .Y(new_n9866_));
  OR4X1    g09674(.A(new_n9859_), .B(new_n9858_), .C(new_n9815_), .D(new_n9825_), .Y(new_n9867_));
  OAI21X1  g09675(.A0(new_n9832_), .A1(new_n9819_), .B0(new_n9836_), .Y(new_n9868_));
  AOI21X1  g09676(.A0(new_n9857_), .A1(new_n9853_), .B0(new_n9379_), .Y(new_n9869_));
  AOI21X1  g09677(.A0(new_n9868_), .A1(\a[51] ), .B0(new_n9869_), .Y(new_n9870_));
  NAND2X1  g09678(.A(new_n9870_), .B(new_n9867_), .Y(new_n9871_));
  AOI21X1  g09679(.A0(new_n9838_), .A1(new_n9835_), .B0(new_n9353_), .Y(new_n9872_));
  NOR2X1   g09680(.A(new_n9872_), .B(\asqrt[27] ), .Y(new_n9873_));
  AND2X1   g09681(.A(new_n9855_), .B(new_n9854_), .Y(new_n9874_));
  OR2X1    g09682(.A(new_n9830_), .B(new_n9353_), .Y(new_n9875_));
  OR4X1    g09683(.A(new_n9875_), .B(new_n9824_), .C(new_n9874_), .D(new_n9819_), .Y(new_n9876_));
  AOI21X1  g09684(.A0(new_n9876_), .A1(new_n9863_), .B0(new_n9372_), .Y(new_n9877_));
  NOR4X1   g09685(.A(new_n9875_), .B(new_n9824_), .C(new_n9874_), .D(new_n9819_), .Y(new_n9878_));
  NOR3X1   g09686(.A(new_n9878_), .B(new_n9869_), .C(\a[52] ), .Y(new_n9879_));
  NOR2X1   g09687(.A(new_n9879_), .B(new_n9877_), .Y(new_n9880_));
  AOI21X1  g09688(.A0(new_n9873_), .A1(new_n9871_), .B0(new_n9880_), .Y(new_n9881_));
  OAI21X1  g09689(.A0(new_n9881_), .A1(new_n9866_), .B0(\asqrt[28] ), .Y(new_n9882_));
  AND2X1   g09690(.A(new_n9420_), .B(new_n9418_), .Y(new_n9883_));
  NOR3X1   g09691(.A(new_n9883_), .B(new_n9371_), .C(new_n9367_), .Y(new_n9884_));
  OAI21X1  g09692(.A0(new_n9832_), .A1(new_n9819_), .B0(new_n9884_), .Y(new_n9885_));
  AOI21X1  g09693(.A0(new_n9366_), .A1(\asqrt[27] ), .B0(new_n9371_), .Y(new_n9886_));
  OAI21X1  g09694(.A0(new_n9832_), .A1(new_n9819_), .B0(new_n9886_), .Y(new_n9887_));
  NAND2X1  g09695(.A(new_n9887_), .B(new_n9883_), .Y(new_n9888_));
  NAND2X1  g09696(.A(new_n9888_), .B(new_n9885_), .Y(new_n9889_));
  AOI21X1  g09697(.A0(new_n9870_), .A1(new_n9867_), .B0(new_n9872_), .Y(new_n9890_));
  OAI21X1  g09698(.A0(new_n9890_), .A1(new_n8874_), .B0(new_n8412_), .Y(new_n9891_));
  OAI21X1  g09699(.A0(new_n9891_), .A1(new_n9881_), .B0(new_n9889_), .Y(new_n9892_));
  AOI21X1  g09700(.A0(new_n9892_), .A1(new_n9882_), .B0(new_n7970_), .Y(new_n9893_));
  AND2X1   g09701(.A(new_n9423_), .B(new_n9421_), .Y(new_n9894_));
  NOR3X1   g09702(.A(new_n9388_), .B(new_n9894_), .C(new_n9422_), .Y(new_n9895_));
  OAI21X1  g09703(.A0(new_n9832_), .A1(new_n9819_), .B0(new_n9895_), .Y(new_n9896_));
  NOR2X1   g09704(.A(new_n9894_), .B(new_n9422_), .Y(new_n9897_));
  OAI21X1  g09705(.A0(new_n9832_), .A1(new_n9819_), .B0(new_n9897_), .Y(new_n9898_));
  NAND2X1  g09706(.A(new_n9898_), .B(new_n9388_), .Y(new_n9899_));
  AND2X1   g09707(.A(new_n9899_), .B(new_n9896_), .Y(new_n9900_));
  INVX1    g09708(.A(new_n9900_), .Y(new_n9901_));
  NAND3X1  g09709(.A(new_n9892_), .B(new_n9882_), .C(new_n7970_), .Y(new_n9902_));
  AOI21X1  g09710(.A0(new_n9902_), .A1(new_n9901_), .B0(new_n9893_), .Y(new_n9903_));
  OR2X1    g09711(.A(new_n9903_), .B(new_n7527_), .Y(new_n9904_));
  OR2X1    g09712(.A(new_n9890_), .B(new_n8874_), .Y(new_n9905_));
  AND2X1   g09713(.A(new_n9870_), .B(new_n9867_), .Y(new_n9906_));
  OR2X1    g09714(.A(new_n9872_), .B(\asqrt[27] ), .Y(new_n9907_));
  OR2X1    g09715(.A(new_n9879_), .B(new_n9877_), .Y(new_n9908_));
  OAI21X1  g09716(.A0(new_n9907_), .A1(new_n9906_), .B0(new_n9908_), .Y(new_n9909_));
  AOI21X1  g09717(.A0(new_n9909_), .A1(new_n9905_), .B0(new_n8412_), .Y(new_n9910_));
  AOI21X1  g09718(.A0(new_n9865_), .A1(\asqrt[27] ), .B0(\asqrt[28] ), .Y(new_n9911_));
  AOI22X1  g09719(.A0(new_n9911_), .A1(new_n9909_), .B0(new_n9888_), .B1(new_n9885_), .Y(new_n9912_));
  NOR3X1   g09720(.A(new_n9912_), .B(new_n9910_), .C(\asqrt[29] ), .Y(new_n9913_));
  NOR2X1   g09721(.A(new_n9913_), .B(new_n9900_), .Y(new_n9914_));
  NOR3X1   g09722(.A(new_n9428_), .B(new_n9396_), .C(new_n9390_), .Y(new_n9915_));
  OAI21X1  g09723(.A0(new_n9832_), .A1(new_n9819_), .B0(new_n9915_), .Y(new_n9916_));
  NOR3X1   g09724(.A(new_n9833_), .B(new_n9428_), .C(new_n9390_), .Y(new_n9917_));
  OR2X1    g09725(.A(new_n9917_), .B(new_n9395_), .Y(new_n9918_));
  AND2X1   g09726(.A(new_n9918_), .B(new_n9916_), .Y(new_n9919_));
  INVX1    g09727(.A(new_n9919_), .Y(new_n9920_));
  OR2X1    g09728(.A(new_n9893_), .B(\asqrt[30] ), .Y(new_n9921_));
  OAI21X1  g09729(.A0(new_n9921_), .A1(new_n9914_), .B0(new_n9920_), .Y(new_n9922_));
  AOI21X1  g09730(.A0(new_n9922_), .A1(new_n9904_), .B0(new_n7103_), .Y(new_n9923_));
  AOI21X1  g09731(.A0(new_n9443_), .A1(new_n9442_), .B0(new_n9406_), .Y(new_n9924_));
  AND2X1   g09732(.A(new_n9924_), .B(new_n9399_), .Y(new_n9925_));
  AOI22X1  g09733(.A0(new_n9443_), .A1(new_n9442_), .B0(new_n9429_), .B1(\asqrt[30] ), .Y(new_n9926_));
  AOI21X1  g09734(.A0(new_n9926_), .A1(\asqrt[25] ), .B0(new_n9405_), .Y(new_n9927_));
  AOI21X1  g09735(.A0(new_n9925_), .A1(\asqrt[25] ), .B0(new_n9927_), .Y(new_n9928_));
  OAI21X1  g09736(.A0(new_n9912_), .A1(new_n9910_), .B0(\asqrt[29] ), .Y(new_n9929_));
  OAI21X1  g09737(.A0(new_n9913_), .A1(new_n9900_), .B0(new_n9929_), .Y(new_n9930_));
  AOI21X1  g09738(.A0(new_n9930_), .A1(\asqrt[30] ), .B0(\asqrt[31] ), .Y(new_n9931_));
  AOI21X1  g09739(.A0(new_n9931_), .A1(new_n9922_), .B0(new_n9928_), .Y(new_n9932_));
  OAI21X1  g09740(.A0(new_n9932_), .A1(new_n9923_), .B0(\asqrt[32] ), .Y(new_n9933_));
  AND2X1   g09741(.A(new_n9430_), .B(new_n9408_), .Y(new_n9934_));
  NOR3X1   g09742(.A(new_n9934_), .B(new_n9446_), .C(new_n9409_), .Y(new_n9935_));
  NOR3X1   g09743(.A(new_n9833_), .B(new_n9934_), .C(new_n9409_), .Y(new_n9936_));
  NOR2X1   g09744(.A(new_n9936_), .B(new_n9414_), .Y(new_n9937_));
  AOI21X1  g09745(.A0(new_n9935_), .A1(\asqrt[25] ), .B0(new_n9937_), .Y(new_n9938_));
  NOR3X1   g09746(.A(new_n9932_), .B(new_n9923_), .C(\asqrt[32] ), .Y(new_n9939_));
  OAI21X1  g09747(.A0(new_n9939_), .A1(new_n9938_), .B0(new_n9933_), .Y(new_n9940_));
  AND2X1   g09748(.A(new_n9940_), .B(\asqrt[33] ), .Y(new_n9941_));
  OR2X1    g09749(.A(new_n9939_), .B(new_n9938_), .Y(new_n9942_));
  NAND4X1  g09750(.A(\asqrt[25] ), .B(new_n9449_), .C(new_n9436_), .D(new_n9432_), .Y(new_n9943_));
  NAND2X1  g09751(.A(new_n9449_), .B(new_n9432_), .Y(new_n9944_));
  OAI21X1  g09752(.A0(new_n9944_), .A1(new_n9833_), .B0(new_n9440_), .Y(new_n9945_));
  AND2X1   g09753(.A(new_n9945_), .B(new_n9943_), .Y(new_n9946_));
  AND2X1   g09754(.A(new_n9933_), .B(new_n6294_), .Y(new_n9947_));
  AOI21X1  g09755(.A0(new_n9947_), .A1(new_n9942_), .B0(new_n9946_), .Y(new_n9948_));
  OAI21X1  g09756(.A0(new_n9948_), .A1(new_n9941_), .B0(\asqrt[34] ), .Y(new_n9949_));
  AND2X1   g09757(.A(new_n9457_), .B(new_n9450_), .Y(new_n9950_));
  NOR3X1   g09758(.A(new_n9950_), .B(new_n9495_), .C(new_n9439_), .Y(new_n9951_));
  NOR3X1   g09759(.A(new_n9833_), .B(new_n9950_), .C(new_n9439_), .Y(new_n9952_));
  NOR2X1   g09760(.A(new_n9952_), .B(new_n9455_), .Y(new_n9953_));
  AOI21X1  g09761(.A0(new_n9951_), .A1(\asqrt[25] ), .B0(new_n9953_), .Y(new_n9954_));
  INVX1    g09762(.A(new_n9954_), .Y(new_n9955_));
  AND2X1   g09763(.A(new_n9930_), .B(\asqrt[30] ), .Y(new_n9956_));
  OR2X1    g09764(.A(new_n9913_), .B(new_n9900_), .Y(new_n9957_));
  NOR2X1   g09765(.A(new_n9893_), .B(\asqrt[30] ), .Y(new_n9958_));
  AOI21X1  g09766(.A0(new_n9958_), .A1(new_n9957_), .B0(new_n9919_), .Y(new_n9959_));
  OAI21X1  g09767(.A0(new_n9959_), .A1(new_n9956_), .B0(\asqrt[31] ), .Y(new_n9960_));
  INVX1    g09768(.A(new_n9928_), .Y(new_n9961_));
  OAI21X1  g09769(.A0(new_n9903_), .A1(new_n7527_), .B0(new_n7103_), .Y(new_n9962_));
  OAI21X1  g09770(.A0(new_n9962_), .A1(new_n9959_), .B0(new_n9961_), .Y(new_n9963_));
  AOI21X1  g09771(.A0(new_n9963_), .A1(new_n9960_), .B0(new_n6699_), .Y(new_n9964_));
  INVX1    g09772(.A(new_n9938_), .Y(new_n9965_));
  NAND3X1  g09773(.A(new_n9963_), .B(new_n9960_), .C(new_n6699_), .Y(new_n9966_));
  AOI21X1  g09774(.A0(new_n9966_), .A1(new_n9965_), .B0(new_n9964_), .Y(new_n9967_));
  OAI21X1  g09775(.A0(new_n9967_), .A1(new_n6294_), .B0(new_n5941_), .Y(new_n9968_));
  OAI21X1  g09776(.A0(new_n9968_), .A1(new_n9948_), .B0(new_n9955_), .Y(new_n9969_));
  AOI21X1  g09777(.A0(new_n9969_), .A1(new_n9949_), .B0(new_n5541_), .Y(new_n9970_));
  AND2X1   g09778(.A(new_n9499_), .B(new_n9497_), .Y(new_n9971_));
  NOR3X1   g09779(.A(new_n9971_), .B(new_n9465_), .C(new_n9498_), .Y(new_n9972_));
  NOR3X1   g09780(.A(new_n9833_), .B(new_n9971_), .C(new_n9498_), .Y(new_n9973_));
  NOR2X1   g09781(.A(new_n9973_), .B(new_n9464_), .Y(new_n9974_));
  AOI21X1  g09782(.A0(new_n9972_), .A1(\asqrt[25] ), .B0(new_n9974_), .Y(new_n9975_));
  INVX1    g09783(.A(new_n9975_), .Y(new_n9976_));
  NAND3X1  g09784(.A(new_n9969_), .B(new_n9949_), .C(new_n5541_), .Y(new_n9977_));
  AOI21X1  g09785(.A0(new_n9977_), .A1(new_n9976_), .B0(new_n9970_), .Y(new_n9978_));
  OR2X1    g09786(.A(new_n9978_), .B(new_n5176_), .Y(new_n9979_));
  OR2X1    g09787(.A(new_n9967_), .B(new_n6294_), .Y(new_n9980_));
  NOR2X1   g09788(.A(new_n9939_), .B(new_n9938_), .Y(new_n9981_));
  INVX1    g09789(.A(new_n9946_), .Y(new_n9982_));
  NAND2X1  g09790(.A(new_n9933_), .B(new_n6294_), .Y(new_n9983_));
  OAI21X1  g09791(.A0(new_n9983_), .A1(new_n9981_), .B0(new_n9982_), .Y(new_n9984_));
  AOI21X1  g09792(.A0(new_n9984_), .A1(new_n9980_), .B0(new_n5941_), .Y(new_n9985_));
  AOI21X1  g09793(.A0(new_n9940_), .A1(\asqrt[33] ), .B0(\asqrt[34] ), .Y(new_n9986_));
  AOI21X1  g09794(.A0(new_n9986_), .A1(new_n9984_), .B0(new_n9954_), .Y(new_n9987_));
  NOR3X1   g09795(.A(new_n9987_), .B(new_n9985_), .C(\asqrt[35] ), .Y(new_n9988_));
  NOR2X1   g09796(.A(new_n9988_), .B(new_n9975_), .Y(new_n9989_));
  NAND4X1  g09797(.A(\asqrt[25] ), .B(new_n9475_), .C(new_n9473_), .D(new_n9501_), .Y(new_n9990_));
  NAND2X1  g09798(.A(new_n9475_), .B(new_n9501_), .Y(new_n9991_));
  OAI21X1  g09799(.A0(new_n9991_), .A1(new_n9833_), .B0(new_n9474_), .Y(new_n9992_));
  AND2X1   g09800(.A(new_n9992_), .B(new_n9990_), .Y(new_n9993_));
  INVX1    g09801(.A(new_n9993_), .Y(new_n9994_));
  OAI21X1  g09802(.A0(new_n9987_), .A1(new_n9985_), .B0(\asqrt[35] ), .Y(new_n9995_));
  NAND2X1  g09803(.A(new_n9995_), .B(new_n5176_), .Y(new_n9996_));
  OAI21X1  g09804(.A0(new_n9996_), .A1(new_n9989_), .B0(new_n9994_), .Y(new_n9997_));
  AOI21X1  g09805(.A0(new_n9997_), .A1(new_n9979_), .B0(new_n4826_), .Y(new_n9998_));
  AOI21X1  g09806(.A0(new_n9517_), .A1(new_n9516_), .B0(new_n9484_), .Y(new_n9999_));
  AND2X1   g09807(.A(new_n9999_), .B(new_n9477_), .Y(new_n10000_));
  AOI22X1  g09808(.A0(new_n9517_), .A1(new_n9516_), .B0(new_n9503_), .B1(\asqrt[36] ), .Y(new_n10001_));
  AOI21X1  g09809(.A0(new_n10001_), .A1(\asqrt[25] ), .B0(new_n9483_), .Y(new_n10002_));
  AOI21X1  g09810(.A0(new_n10000_), .A1(\asqrt[25] ), .B0(new_n10002_), .Y(new_n10003_));
  OAI21X1  g09811(.A0(new_n9988_), .A1(new_n9975_), .B0(new_n9995_), .Y(new_n10004_));
  AOI21X1  g09812(.A0(new_n10004_), .A1(\asqrt[36] ), .B0(\asqrt[37] ), .Y(new_n10005_));
  AOI21X1  g09813(.A0(new_n10005_), .A1(new_n9997_), .B0(new_n10003_), .Y(new_n10006_));
  OAI21X1  g09814(.A0(new_n10006_), .A1(new_n9998_), .B0(\asqrt[38] ), .Y(new_n10007_));
  AND2X1   g09815(.A(new_n9504_), .B(new_n9486_), .Y(new_n10008_));
  NOR3X1   g09816(.A(new_n10008_), .B(new_n9520_), .C(new_n9487_), .Y(new_n10009_));
  NOR3X1   g09817(.A(new_n9833_), .B(new_n10008_), .C(new_n9487_), .Y(new_n10010_));
  NOR2X1   g09818(.A(new_n10010_), .B(new_n9492_), .Y(new_n10011_));
  AOI21X1  g09819(.A0(new_n10009_), .A1(\asqrt[25] ), .B0(new_n10011_), .Y(new_n10012_));
  NOR3X1   g09820(.A(new_n10006_), .B(new_n9998_), .C(\asqrt[38] ), .Y(new_n10013_));
  OAI21X1  g09821(.A0(new_n10013_), .A1(new_n10012_), .B0(new_n10007_), .Y(new_n10014_));
  AND2X1   g09822(.A(new_n10014_), .B(\asqrt[39] ), .Y(new_n10015_));
  OR2X1    g09823(.A(new_n10013_), .B(new_n10012_), .Y(new_n10016_));
  NAND4X1  g09824(.A(\asqrt[25] ), .B(new_n9523_), .C(new_n9510_), .D(new_n9506_), .Y(new_n10017_));
  NAND2X1  g09825(.A(new_n9523_), .B(new_n9506_), .Y(new_n10018_));
  OAI21X1  g09826(.A0(new_n10018_), .A1(new_n9833_), .B0(new_n9514_), .Y(new_n10019_));
  AND2X1   g09827(.A(new_n10019_), .B(new_n10017_), .Y(new_n10020_));
  AND2X1   g09828(.A(new_n10004_), .B(\asqrt[36] ), .Y(new_n10021_));
  OR2X1    g09829(.A(new_n9988_), .B(new_n9975_), .Y(new_n10022_));
  AND2X1   g09830(.A(new_n9995_), .B(new_n5176_), .Y(new_n10023_));
  AOI21X1  g09831(.A0(new_n10023_), .A1(new_n10022_), .B0(new_n9993_), .Y(new_n10024_));
  OAI21X1  g09832(.A0(new_n10024_), .A1(new_n10021_), .B0(\asqrt[37] ), .Y(new_n10025_));
  INVX1    g09833(.A(new_n10003_), .Y(new_n10026_));
  OAI21X1  g09834(.A0(new_n9978_), .A1(new_n5176_), .B0(new_n4826_), .Y(new_n10027_));
  OAI21X1  g09835(.A0(new_n10027_), .A1(new_n10024_), .B0(new_n10026_), .Y(new_n10028_));
  AOI21X1  g09836(.A0(new_n10028_), .A1(new_n10025_), .B0(new_n4493_), .Y(new_n10029_));
  NOR2X1   g09837(.A(new_n10029_), .B(\asqrt[39] ), .Y(new_n10030_));
  AOI21X1  g09838(.A0(new_n10030_), .A1(new_n10016_), .B0(new_n10020_), .Y(new_n10031_));
  OAI21X1  g09839(.A0(new_n10031_), .A1(new_n10015_), .B0(\asqrt[40] ), .Y(new_n10032_));
  INVX1    g09840(.A(new_n10012_), .Y(new_n10033_));
  NAND3X1  g09841(.A(new_n10028_), .B(new_n10025_), .C(new_n4493_), .Y(new_n10034_));
  AOI21X1  g09842(.A0(new_n10034_), .A1(new_n10033_), .B0(new_n10029_), .Y(new_n10035_));
  OAI21X1  g09843(.A0(new_n10035_), .A1(new_n4165_), .B0(new_n3863_), .Y(new_n10036_));
  AND2X1   g09844(.A(new_n9526_), .B(new_n9524_), .Y(new_n10037_));
  NOR3X1   g09845(.A(new_n9571_), .B(new_n10037_), .C(new_n9513_), .Y(new_n10038_));
  NOR3X1   g09846(.A(new_n9833_), .B(new_n10037_), .C(new_n9513_), .Y(new_n10039_));
  NOR2X1   g09847(.A(new_n10039_), .B(new_n9531_), .Y(new_n10040_));
  AOI21X1  g09848(.A0(new_n10038_), .A1(\asqrt[25] ), .B0(new_n10040_), .Y(new_n10041_));
  INVX1    g09849(.A(new_n10041_), .Y(new_n10042_));
  OAI21X1  g09850(.A0(new_n10036_), .A1(new_n10031_), .B0(new_n10042_), .Y(new_n10043_));
  AOI21X1  g09851(.A0(new_n10043_), .A1(new_n10032_), .B0(new_n3564_), .Y(new_n10044_));
  AND2X1   g09852(.A(new_n9574_), .B(new_n9572_), .Y(new_n10045_));
  NOR3X1   g09853(.A(new_n10045_), .B(new_n9539_), .C(new_n9573_), .Y(new_n10046_));
  NOR3X1   g09854(.A(new_n9833_), .B(new_n10045_), .C(new_n9573_), .Y(new_n10047_));
  NOR2X1   g09855(.A(new_n10047_), .B(new_n9538_), .Y(new_n10048_));
  AOI21X1  g09856(.A0(new_n10046_), .A1(\asqrt[25] ), .B0(new_n10048_), .Y(new_n10049_));
  INVX1    g09857(.A(new_n10049_), .Y(new_n10050_));
  NAND3X1  g09858(.A(new_n10043_), .B(new_n10032_), .C(new_n3564_), .Y(new_n10051_));
  AOI21X1  g09859(.A0(new_n10051_), .A1(new_n10050_), .B0(new_n10044_), .Y(new_n10052_));
  OR2X1    g09860(.A(new_n10052_), .B(new_n3276_), .Y(new_n10053_));
  AND2X1   g09861(.A(new_n10051_), .B(new_n10050_), .Y(new_n10054_));
  NAND4X1  g09862(.A(\asqrt[25] ), .B(new_n9549_), .C(new_n9547_), .D(new_n9576_), .Y(new_n10055_));
  NAND2X1  g09863(.A(new_n9549_), .B(new_n9576_), .Y(new_n10056_));
  OAI21X1  g09864(.A0(new_n10056_), .A1(new_n9833_), .B0(new_n9548_), .Y(new_n10057_));
  AND2X1   g09865(.A(new_n10057_), .B(new_n10055_), .Y(new_n10058_));
  INVX1    g09866(.A(new_n10058_), .Y(new_n10059_));
  OR2X1    g09867(.A(new_n10044_), .B(\asqrt[42] ), .Y(new_n10060_));
  OAI21X1  g09868(.A0(new_n10060_), .A1(new_n10054_), .B0(new_n10059_), .Y(new_n10061_));
  AOI21X1  g09869(.A0(new_n10061_), .A1(new_n10053_), .B0(new_n3008_), .Y(new_n10062_));
  AOI21X1  g09870(.A0(new_n9592_), .A1(new_n9591_), .B0(new_n9558_), .Y(new_n10063_));
  AND2X1   g09871(.A(new_n10063_), .B(new_n9551_), .Y(new_n10064_));
  AOI22X1  g09872(.A0(new_n9592_), .A1(new_n9591_), .B0(new_n9578_), .B1(\asqrt[42] ), .Y(new_n10065_));
  AOI21X1  g09873(.A0(new_n10065_), .A1(\asqrt[25] ), .B0(new_n9557_), .Y(new_n10066_));
  AOI21X1  g09874(.A0(new_n10064_), .A1(\asqrt[25] ), .B0(new_n10066_), .Y(new_n10067_));
  OR2X1    g09875(.A(new_n10035_), .B(new_n4165_), .Y(new_n10068_));
  NOR2X1   g09876(.A(new_n10013_), .B(new_n10012_), .Y(new_n10069_));
  INVX1    g09877(.A(new_n10020_), .Y(new_n10070_));
  OR2X1    g09878(.A(new_n10029_), .B(\asqrt[39] ), .Y(new_n10071_));
  OAI21X1  g09879(.A0(new_n10071_), .A1(new_n10069_), .B0(new_n10070_), .Y(new_n10072_));
  AOI21X1  g09880(.A0(new_n10072_), .A1(new_n10068_), .B0(new_n3863_), .Y(new_n10073_));
  AOI21X1  g09881(.A0(new_n10014_), .A1(\asqrt[39] ), .B0(\asqrt[40] ), .Y(new_n10074_));
  AOI21X1  g09882(.A0(new_n10074_), .A1(new_n10072_), .B0(new_n10041_), .Y(new_n10075_));
  OAI21X1  g09883(.A0(new_n10075_), .A1(new_n10073_), .B0(\asqrt[41] ), .Y(new_n10076_));
  NOR3X1   g09884(.A(new_n10075_), .B(new_n10073_), .C(\asqrt[41] ), .Y(new_n10077_));
  OAI21X1  g09885(.A0(new_n10077_), .A1(new_n10049_), .B0(new_n10076_), .Y(new_n10078_));
  AOI21X1  g09886(.A0(new_n10078_), .A1(\asqrt[42] ), .B0(\asqrt[43] ), .Y(new_n10079_));
  AOI21X1  g09887(.A0(new_n10079_), .A1(new_n10061_), .B0(new_n10067_), .Y(new_n10080_));
  OAI21X1  g09888(.A0(new_n10080_), .A1(new_n10062_), .B0(\asqrt[44] ), .Y(new_n10081_));
  AND2X1   g09889(.A(new_n9579_), .B(new_n9560_), .Y(new_n10082_));
  NOR3X1   g09890(.A(new_n10082_), .B(new_n9566_), .C(new_n9561_), .Y(new_n10083_));
  NOR3X1   g09891(.A(new_n9833_), .B(new_n10082_), .C(new_n9561_), .Y(new_n10084_));
  NOR2X1   g09892(.A(new_n10084_), .B(new_n9567_), .Y(new_n10085_));
  AOI21X1  g09893(.A0(new_n10083_), .A1(\asqrt[25] ), .B0(new_n10085_), .Y(new_n10086_));
  NOR3X1   g09894(.A(new_n10080_), .B(new_n10062_), .C(\asqrt[44] ), .Y(new_n10087_));
  OAI21X1  g09895(.A0(new_n10087_), .A1(new_n10086_), .B0(new_n10081_), .Y(new_n10088_));
  AND2X1   g09896(.A(new_n10088_), .B(\asqrt[45] ), .Y(new_n10089_));
  OR2X1    g09897(.A(new_n10087_), .B(new_n10086_), .Y(new_n10090_));
  NAND4X1  g09898(.A(\asqrt[25] ), .B(new_n9597_), .C(new_n9585_), .D(new_n9581_), .Y(new_n10091_));
  NAND2X1  g09899(.A(new_n9597_), .B(new_n9581_), .Y(new_n10092_));
  OAI21X1  g09900(.A0(new_n10092_), .A1(new_n9833_), .B0(new_n9589_), .Y(new_n10093_));
  AND2X1   g09901(.A(new_n10093_), .B(new_n10091_), .Y(new_n10094_));
  AND2X1   g09902(.A(new_n10078_), .B(\asqrt[42] ), .Y(new_n10095_));
  NAND2X1  g09903(.A(new_n10051_), .B(new_n10050_), .Y(new_n10096_));
  NOR2X1   g09904(.A(new_n10044_), .B(\asqrt[42] ), .Y(new_n10097_));
  AOI21X1  g09905(.A0(new_n10097_), .A1(new_n10096_), .B0(new_n10058_), .Y(new_n10098_));
  OAI21X1  g09906(.A0(new_n10098_), .A1(new_n10095_), .B0(\asqrt[43] ), .Y(new_n10099_));
  INVX1    g09907(.A(new_n10067_), .Y(new_n10100_));
  OAI21X1  g09908(.A0(new_n10052_), .A1(new_n3276_), .B0(new_n3008_), .Y(new_n10101_));
  OAI21X1  g09909(.A0(new_n10101_), .A1(new_n10098_), .B0(new_n10100_), .Y(new_n10102_));
  AOI21X1  g09910(.A0(new_n10102_), .A1(new_n10099_), .B0(new_n2769_), .Y(new_n10103_));
  NOR2X1   g09911(.A(new_n10103_), .B(\asqrt[45] ), .Y(new_n10104_));
  AOI21X1  g09912(.A0(new_n10104_), .A1(new_n10090_), .B0(new_n10094_), .Y(new_n10105_));
  OAI21X1  g09913(.A0(new_n10105_), .A1(new_n10089_), .B0(\asqrt[46] ), .Y(new_n10106_));
  AND2X1   g09914(.A(new_n9605_), .B(new_n9598_), .Y(new_n10107_));
  NOR3X1   g09915(.A(new_n10107_), .B(new_n9642_), .C(new_n9588_), .Y(new_n10108_));
  NOR3X1   g09916(.A(new_n9833_), .B(new_n10107_), .C(new_n9588_), .Y(new_n10109_));
  NOR2X1   g09917(.A(new_n10109_), .B(new_n9603_), .Y(new_n10110_));
  AOI21X1  g09918(.A0(new_n10108_), .A1(\asqrt[25] ), .B0(new_n10110_), .Y(new_n10111_));
  INVX1    g09919(.A(new_n10111_), .Y(new_n10112_));
  INVX1    g09920(.A(new_n10086_), .Y(new_n10113_));
  NAND3X1  g09921(.A(new_n10102_), .B(new_n10099_), .C(new_n2769_), .Y(new_n10114_));
  AOI21X1  g09922(.A0(new_n10114_), .A1(new_n10113_), .B0(new_n10103_), .Y(new_n10115_));
  OAI21X1  g09923(.A0(new_n10115_), .A1(new_n2570_), .B0(new_n2263_), .Y(new_n10116_));
  OAI21X1  g09924(.A0(new_n10116_), .A1(new_n10105_), .B0(new_n10112_), .Y(new_n10117_));
  AOI21X1  g09925(.A0(new_n10117_), .A1(new_n10106_), .B0(new_n2040_), .Y(new_n10118_));
  AND2X1   g09926(.A(new_n9647_), .B(new_n9644_), .Y(new_n10119_));
  NOR3X1   g09927(.A(new_n10119_), .B(new_n9612_), .C(new_n9645_), .Y(new_n10120_));
  NOR3X1   g09928(.A(new_n9833_), .B(new_n10119_), .C(new_n9645_), .Y(new_n10121_));
  NOR2X1   g09929(.A(new_n10121_), .B(new_n9646_), .Y(new_n10122_));
  AOI21X1  g09930(.A0(new_n10120_), .A1(\asqrt[25] ), .B0(new_n10122_), .Y(new_n10123_));
  INVX1    g09931(.A(new_n10123_), .Y(new_n10124_));
  NAND3X1  g09932(.A(new_n10117_), .B(new_n10106_), .C(new_n2040_), .Y(new_n10125_));
  AOI21X1  g09933(.A0(new_n10125_), .A1(new_n10124_), .B0(new_n10118_), .Y(new_n10126_));
  OR2X1    g09934(.A(new_n10126_), .B(new_n1834_), .Y(new_n10127_));
  OR2X1    g09935(.A(new_n10115_), .B(new_n2570_), .Y(new_n10128_));
  NOR2X1   g09936(.A(new_n10087_), .B(new_n10086_), .Y(new_n10129_));
  INVX1    g09937(.A(new_n10094_), .Y(new_n10130_));
  OR2X1    g09938(.A(new_n10103_), .B(\asqrt[45] ), .Y(new_n10131_));
  OAI21X1  g09939(.A0(new_n10131_), .A1(new_n10129_), .B0(new_n10130_), .Y(new_n10132_));
  AOI21X1  g09940(.A0(new_n10132_), .A1(new_n10128_), .B0(new_n2263_), .Y(new_n10133_));
  AOI21X1  g09941(.A0(new_n10088_), .A1(\asqrt[45] ), .B0(\asqrt[46] ), .Y(new_n10134_));
  AOI21X1  g09942(.A0(new_n10134_), .A1(new_n10132_), .B0(new_n10111_), .Y(new_n10135_));
  NOR3X1   g09943(.A(new_n10135_), .B(new_n10133_), .C(\asqrt[47] ), .Y(new_n10136_));
  NOR2X1   g09944(.A(new_n10136_), .B(new_n10123_), .Y(new_n10137_));
  NAND4X1  g09945(.A(\asqrt[25] ), .B(new_n9622_), .C(new_n9620_), .D(new_n9649_), .Y(new_n10138_));
  NAND2X1  g09946(.A(new_n9622_), .B(new_n9649_), .Y(new_n10139_));
  OAI21X1  g09947(.A0(new_n10139_), .A1(new_n9833_), .B0(new_n9621_), .Y(new_n10140_));
  AND2X1   g09948(.A(new_n10140_), .B(new_n10138_), .Y(new_n10141_));
  INVX1    g09949(.A(new_n10141_), .Y(new_n10142_));
  OAI21X1  g09950(.A0(new_n10135_), .A1(new_n10133_), .B0(\asqrt[47] ), .Y(new_n10143_));
  NAND2X1  g09951(.A(new_n10143_), .B(new_n1834_), .Y(new_n10144_));
  OAI21X1  g09952(.A0(new_n10144_), .A1(new_n10137_), .B0(new_n10142_), .Y(new_n10145_));
  AOI21X1  g09953(.A0(new_n10145_), .A1(new_n10127_), .B0(new_n1632_), .Y(new_n10146_));
  AOI21X1  g09954(.A0(new_n9679_), .A1(new_n9678_), .B0(new_n9631_), .Y(new_n10147_));
  AND2X1   g09955(.A(new_n10147_), .B(new_n9624_), .Y(new_n10148_));
  AOI22X1  g09956(.A0(new_n9679_), .A1(new_n9678_), .B0(new_n9651_), .B1(\asqrt[48] ), .Y(new_n10149_));
  AOI21X1  g09957(.A0(new_n10149_), .A1(\asqrt[25] ), .B0(new_n9630_), .Y(new_n10150_));
  AOI21X1  g09958(.A0(new_n10148_), .A1(\asqrt[25] ), .B0(new_n10150_), .Y(new_n10151_));
  OAI21X1  g09959(.A0(new_n10136_), .A1(new_n10123_), .B0(new_n10143_), .Y(new_n10152_));
  AOI21X1  g09960(.A0(new_n10152_), .A1(\asqrt[48] ), .B0(\asqrt[49] ), .Y(new_n10153_));
  AOI21X1  g09961(.A0(new_n10153_), .A1(new_n10145_), .B0(new_n10151_), .Y(new_n10154_));
  OAI21X1  g09962(.A0(new_n10154_), .A1(new_n10146_), .B0(\asqrt[50] ), .Y(new_n10155_));
  AND2X1   g09963(.A(new_n9652_), .B(new_n9633_), .Y(new_n10156_));
  NOR3X1   g09964(.A(new_n10156_), .B(new_n9682_), .C(new_n9634_), .Y(new_n10157_));
  NOR3X1   g09965(.A(new_n9833_), .B(new_n10156_), .C(new_n9634_), .Y(new_n10158_));
  NOR2X1   g09966(.A(new_n10158_), .B(new_n9639_), .Y(new_n10159_));
  AOI21X1  g09967(.A0(new_n10157_), .A1(\asqrt[25] ), .B0(new_n10159_), .Y(new_n10160_));
  NOR3X1   g09968(.A(new_n10154_), .B(new_n10146_), .C(\asqrt[50] ), .Y(new_n10161_));
  OAI21X1  g09969(.A0(new_n10161_), .A1(new_n10160_), .B0(new_n10155_), .Y(new_n10162_));
  AND2X1   g09970(.A(new_n10162_), .B(\asqrt[51] ), .Y(new_n10163_));
  OR2X1    g09971(.A(new_n10161_), .B(new_n10160_), .Y(new_n10164_));
  OR4X1    g09972(.A(new_n9833_), .B(new_n9659_), .C(new_n9686_), .D(new_n9685_), .Y(new_n10165_));
  OR2X1    g09973(.A(new_n9659_), .B(new_n9685_), .Y(new_n10166_));
  OAI21X1  g09974(.A0(new_n10166_), .A1(new_n9833_), .B0(new_n9686_), .Y(new_n10167_));
  AND2X1   g09975(.A(new_n10167_), .B(new_n10165_), .Y(new_n10168_));
  AND2X1   g09976(.A(new_n10155_), .B(new_n1277_), .Y(new_n10169_));
  AOI21X1  g09977(.A0(new_n10169_), .A1(new_n10164_), .B0(new_n10168_), .Y(new_n10170_));
  OAI21X1  g09978(.A0(new_n10170_), .A1(new_n10163_), .B0(\asqrt[52] ), .Y(new_n10171_));
  AND2X1   g09979(.A(new_n9668_), .B(new_n9662_), .Y(new_n10172_));
  NOR3X1   g09980(.A(new_n10172_), .B(new_n9707_), .C(new_n9661_), .Y(new_n10173_));
  NOR3X1   g09981(.A(new_n9833_), .B(new_n10172_), .C(new_n9661_), .Y(new_n10174_));
  NOR2X1   g09982(.A(new_n10174_), .B(new_n9667_), .Y(new_n10175_));
  AOI21X1  g09983(.A0(new_n10173_), .A1(\asqrt[25] ), .B0(new_n10175_), .Y(new_n10176_));
  INVX1    g09984(.A(new_n10176_), .Y(new_n10177_));
  AND2X1   g09985(.A(new_n10152_), .B(\asqrt[48] ), .Y(new_n10178_));
  OR2X1    g09986(.A(new_n10136_), .B(new_n10123_), .Y(new_n10179_));
  AND2X1   g09987(.A(new_n10143_), .B(new_n1834_), .Y(new_n10180_));
  AOI21X1  g09988(.A0(new_n10180_), .A1(new_n10179_), .B0(new_n10141_), .Y(new_n10181_));
  OAI21X1  g09989(.A0(new_n10181_), .A1(new_n10178_), .B0(\asqrt[49] ), .Y(new_n10182_));
  INVX1    g09990(.A(new_n10151_), .Y(new_n10183_));
  OAI21X1  g09991(.A0(new_n10126_), .A1(new_n1834_), .B0(new_n1632_), .Y(new_n10184_));
  OAI21X1  g09992(.A0(new_n10184_), .A1(new_n10181_), .B0(new_n10183_), .Y(new_n10185_));
  AOI21X1  g09993(.A0(new_n10185_), .A1(new_n10182_), .B0(new_n1469_), .Y(new_n10186_));
  INVX1    g09994(.A(new_n10160_), .Y(new_n10187_));
  NAND3X1  g09995(.A(new_n10185_), .B(new_n10182_), .C(new_n1469_), .Y(new_n10188_));
  AOI21X1  g09996(.A0(new_n10188_), .A1(new_n10187_), .B0(new_n10186_), .Y(new_n10189_));
  OAI21X1  g09997(.A0(new_n10189_), .A1(new_n1277_), .B0(new_n1111_), .Y(new_n10190_));
  OAI21X1  g09998(.A0(new_n10190_), .A1(new_n10170_), .B0(new_n10177_), .Y(new_n10191_));
  AOI21X1  g09999(.A0(new_n10191_), .A1(new_n10171_), .B0(new_n968_), .Y(new_n10192_));
  AND2X1   g10000(.A(new_n9711_), .B(new_n9709_), .Y(new_n10193_));
  NOR3X1   g10001(.A(new_n10193_), .B(new_n9676_), .C(new_n9710_), .Y(new_n10194_));
  NOR3X1   g10002(.A(new_n9833_), .B(new_n10193_), .C(new_n9710_), .Y(new_n10195_));
  NOR2X1   g10003(.A(new_n10195_), .B(new_n9675_), .Y(new_n10196_));
  AOI21X1  g10004(.A0(new_n10194_), .A1(\asqrt[25] ), .B0(new_n10196_), .Y(new_n10197_));
  INVX1    g10005(.A(new_n10197_), .Y(new_n10198_));
  NAND3X1  g10006(.A(new_n10191_), .B(new_n10171_), .C(new_n968_), .Y(new_n10199_));
  AOI21X1  g10007(.A0(new_n10199_), .A1(new_n10198_), .B0(new_n10192_), .Y(new_n10200_));
  OR2X1    g10008(.A(new_n10200_), .B(new_n902_), .Y(new_n10201_));
  OR2X1    g10009(.A(new_n10189_), .B(new_n1277_), .Y(new_n10202_));
  NOR2X1   g10010(.A(new_n10161_), .B(new_n10160_), .Y(new_n10203_));
  INVX1    g10011(.A(new_n10168_), .Y(new_n10204_));
  NAND2X1  g10012(.A(new_n10155_), .B(new_n1277_), .Y(new_n10205_));
  OAI21X1  g10013(.A0(new_n10205_), .A1(new_n10203_), .B0(new_n10204_), .Y(new_n10206_));
  AOI21X1  g10014(.A0(new_n10206_), .A1(new_n10202_), .B0(new_n1111_), .Y(new_n10207_));
  AOI21X1  g10015(.A0(new_n10162_), .A1(\asqrt[51] ), .B0(\asqrt[52] ), .Y(new_n10208_));
  AOI21X1  g10016(.A0(new_n10208_), .A1(new_n10206_), .B0(new_n10176_), .Y(new_n10209_));
  NOR3X1   g10017(.A(new_n10209_), .B(new_n10207_), .C(\asqrt[53] ), .Y(new_n10210_));
  NOR2X1   g10018(.A(new_n10210_), .B(new_n10197_), .Y(new_n10211_));
  OR4X1    g10019(.A(new_n9833_), .B(new_n9723_), .C(new_n9694_), .D(new_n9691_), .Y(new_n10212_));
  OR2X1    g10020(.A(new_n9723_), .B(new_n9691_), .Y(new_n10213_));
  OAI21X1  g10021(.A0(new_n10213_), .A1(new_n9833_), .B0(new_n9694_), .Y(new_n10214_));
  AND2X1   g10022(.A(new_n10214_), .B(new_n10212_), .Y(new_n10215_));
  INVX1    g10023(.A(new_n10215_), .Y(new_n10216_));
  OAI21X1  g10024(.A0(new_n10209_), .A1(new_n10207_), .B0(\asqrt[53] ), .Y(new_n10217_));
  NAND2X1  g10025(.A(new_n10217_), .B(new_n902_), .Y(new_n10218_));
  OAI21X1  g10026(.A0(new_n10218_), .A1(new_n10211_), .B0(new_n10216_), .Y(new_n10219_));
  AOI21X1  g10027(.A0(new_n10219_), .A1(new_n10201_), .B0(new_n697_), .Y(new_n10220_));
  AOI21X1  g10028(.A0(new_n9752_), .A1(new_n9751_), .B0(new_n9704_), .Y(new_n10221_));
  AND2X1   g10029(.A(new_n10221_), .B(new_n9697_), .Y(new_n10222_));
  AOI22X1  g10030(.A0(new_n9752_), .A1(new_n9751_), .B0(new_n9724_), .B1(\asqrt[54] ), .Y(new_n10223_));
  AOI21X1  g10031(.A0(new_n10223_), .A1(\asqrt[25] ), .B0(new_n9703_), .Y(new_n10224_));
  AOI21X1  g10032(.A0(new_n10222_), .A1(\asqrt[25] ), .B0(new_n10224_), .Y(new_n10225_));
  OAI21X1  g10033(.A0(new_n10210_), .A1(new_n10197_), .B0(new_n10217_), .Y(new_n10226_));
  AOI21X1  g10034(.A0(new_n10226_), .A1(\asqrt[54] ), .B0(\asqrt[55] ), .Y(new_n10227_));
  AOI21X1  g10035(.A0(new_n10227_), .A1(new_n10219_), .B0(new_n10225_), .Y(new_n10228_));
  OAI21X1  g10036(.A0(new_n10228_), .A1(new_n10220_), .B0(\asqrt[56] ), .Y(new_n10229_));
  AND2X1   g10037(.A(new_n9725_), .B(new_n9715_), .Y(new_n10230_));
  NOR3X1   g10038(.A(new_n10230_), .B(new_n9755_), .C(new_n9716_), .Y(new_n10231_));
  NOR3X1   g10039(.A(new_n9833_), .B(new_n10230_), .C(new_n9716_), .Y(new_n10232_));
  NOR2X1   g10040(.A(new_n10232_), .B(new_n9721_), .Y(new_n10233_));
  AOI21X1  g10041(.A0(new_n10231_), .A1(\asqrt[25] ), .B0(new_n10233_), .Y(new_n10234_));
  NOR3X1   g10042(.A(new_n10228_), .B(new_n10220_), .C(\asqrt[56] ), .Y(new_n10235_));
  OAI21X1  g10043(.A0(new_n10235_), .A1(new_n10234_), .B0(new_n10229_), .Y(new_n10236_));
  AND2X1   g10044(.A(new_n10236_), .B(\asqrt[57] ), .Y(new_n10237_));
  OR2X1    g10045(.A(new_n10235_), .B(new_n10234_), .Y(new_n10238_));
  OR4X1    g10046(.A(new_n9833_), .B(new_n9732_), .C(new_n9759_), .D(new_n9758_), .Y(new_n10239_));
  OR2X1    g10047(.A(new_n9732_), .B(new_n9758_), .Y(new_n10240_));
  OAI21X1  g10048(.A0(new_n10240_), .A1(new_n9833_), .B0(new_n9759_), .Y(new_n10241_));
  AND2X1   g10049(.A(new_n10241_), .B(new_n10239_), .Y(new_n10242_));
  AND2X1   g10050(.A(new_n10229_), .B(new_n481_), .Y(new_n10243_));
  AOI21X1  g10051(.A0(new_n10243_), .A1(new_n10238_), .B0(new_n10242_), .Y(new_n10244_));
  OAI21X1  g10052(.A0(new_n10244_), .A1(new_n10237_), .B0(\asqrt[58] ), .Y(new_n10245_));
  AND2X1   g10053(.A(new_n9741_), .B(new_n9735_), .Y(new_n10246_));
  NOR3X1   g10054(.A(new_n10246_), .B(new_n9775_), .C(new_n9734_), .Y(new_n10247_));
  NOR3X1   g10055(.A(new_n9833_), .B(new_n10246_), .C(new_n9734_), .Y(new_n10248_));
  NOR2X1   g10056(.A(new_n10248_), .B(new_n9740_), .Y(new_n10249_));
  AOI21X1  g10057(.A0(new_n10247_), .A1(\asqrt[25] ), .B0(new_n10249_), .Y(new_n10250_));
  INVX1    g10058(.A(new_n10250_), .Y(new_n10251_));
  AND2X1   g10059(.A(new_n10226_), .B(\asqrt[54] ), .Y(new_n10252_));
  OR2X1    g10060(.A(new_n10210_), .B(new_n10197_), .Y(new_n10253_));
  AND2X1   g10061(.A(new_n10217_), .B(new_n902_), .Y(new_n10254_));
  AOI21X1  g10062(.A0(new_n10254_), .A1(new_n10253_), .B0(new_n10215_), .Y(new_n10255_));
  OAI21X1  g10063(.A0(new_n10255_), .A1(new_n10252_), .B0(\asqrt[55] ), .Y(new_n10256_));
  INVX1    g10064(.A(new_n10225_), .Y(new_n10257_));
  OAI21X1  g10065(.A0(new_n10200_), .A1(new_n902_), .B0(new_n697_), .Y(new_n10258_));
  OAI21X1  g10066(.A0(new_n10258_), .A1(new_n10255_), .B0(new_n10257_), .Y(new_n10259_));
  AOI21X1  g10067(.A0(new_n10259_), .A1(new_n10256_), .B0(new_n582_), .Y(new_n10260_));
  INVX1    g10068(.A(new_n10234_), .Y(new_n10261_));
  NAND3X1  g10069(.A(new_n10259_), .B(new_n10256_), .C(new_n582_), .Y(new_n10262_));
  AOI21X1  g10070(.A0(new_n10262_), .A1(new_n10261_), .B0(new_n10260_), .Y(new_n10263_));
  OAI21X1  g10071(.A0(new_n10263_), .A1(new_n481_), .B0(new_n399_), .Y(new_n10264_));
  OAI21X1  g10072(.A0(new_n10264_), .A1(new_n10244_), .B0(new_n10251_), .Y(new_n10265_));
  AOI21X1  g10073(.A0(new_n10265_), .A1(new_n10245_), .B0(new_n328_), .Y(new_n10266_));
  AND2X1   g10074(.A(new_n9779_), .B(new_n9777_), .Y(new_n10267_));
  NOR3X1   g10075(.A(new_n10267_), .B(new_n9749_), .C(new_n9778_), .Y(new_n10268_));
  NOR3X1   g10076(.A(new_n9833_), .B(new_n10267_), .C(new_n9778_), .Y(new_n10269_));
  NOR2X1   g10077(.A(new_n10269_), .B(new_n9748_), .Y(new_n10270_));
  AOI21X1  g10078(.A0(new_n10268_), .A1(\asqrt[25] ), .B0(new_n10270_), .Y(new_n10271_));
  INVX1    g10079(.A(new_n10271_), .Y(new_n10272_));
  NAND3X1  g10080(.A(new_n10265_), .B(new_n10245_), .C(new_n328_), .Y(new_n10273_));
  AOI21X1  g10081(.A0(new_n10273_), .A1(new_n10272_), .B0(new_n10266_), .Y(new_n10274_));
  OR2X1    g10082(.A(new_n10274_), .B(new_n292_), .Y(new_n10275_));
  OR2X1    g10083(.A(new_n10263_), .B(new_n481_), .Y(new_n10276_));
  NOR2X1   g10084(.A(new_n10235_), .B(new_n10234_), .Y(new_n10277_));
  INVX1    g10085(.A(new_n10242_), .Y(new_n10278_));
  NAND2X1  g10086(.A(new_n10229_), .B(new_n481_), .Y(new_n10279_));
  OAI21X1  g10087(.A0(new_n10279_), .A1(new_n10277_), .B0(new_n10278_), .Y(new_n10280_));
  AOI21X1  g10088(.A0(new_n10280_), .A1(new_n10276_), .B0(new_n399_), .Y(new_n10281_));
  AOI21X1  g10089(.A0(new_n10236_), .A1(\asqrt[57] ), .B0(\asqrt[58] ), .Y(new_n10282_));
  AOI21X1  g10090(.A0(new_n10282_), .A1(new_n10280_), .B0(new_n10250_), .Y(new_n10283_));
  NOR3X1   g10091(.A(new_n10283_), .B(new_n10281_), .C(\asqrt[59] ), .Y(new_n10284_));
  NOR2X1   g10092(.A(new_n10284_), .B(new_n10271_), .Y(new_n10285_));
  OR4X1    g10093(.A(new_n9833_), .B(new_n9781_), .C(new_n9769_), .D(new_n9764_), .Y(new_n10286_));
  OR2X1    g10094(.A(new_n9781_), .B(new_n9764_), .Y(new_n10287_));
  OAI21X1  g10095(.A0(new_n10287_), .A1(new_n9833_), .B0(new_n9769_), .Y(new_n10288_));
  AND2X1   g10096(.A(new_n10288_), .B(new_n10286_), .Y(new_n10289_));
  INVX1    g10097(.A(new_n10289_), .Y(new_n10290_));
  OAI21X1  g10098(.A0(new_n10283_), .A1(new_n10281_), .B0(\asqrt[59] ), .Y(new_n10291_));
  NAND2X1  g10099(.A(new_n10291_), .B(new_n292_), .Y(new_n10292_));
  OAI21X1  g10100(.A0(new_n10292_), .A1(new_n10285_), .B0(new_n10290_), .Y(new_n10293_));
  AOI21X1  g10101(.A0(new_n10293_), .A1(new_n10275_), .B0(new_n217_), .Y(new_n10294_));
  AOI21X1  g10102(.A0(new_n9842_), .A1(new_n9841_), .B0(new_n9788_), .Y(new_n10295_));
  AND2X1   g10103(.A(new_n10295_), .B(new_n9772_), .Y(new_n10296_));
  AOI22X1  g10104(.A0(new_n9842_), .A1(new_n9841_), .B0(new_n9798_), .B1(\asqrt[60] ), .Y(new_n10297_));
  AOI21X1  g10105(.A0(new_n10297_), .A1(\asqrt[25] ), .B0(new_n9787_), .Y(new_n10298_));
  AOI21X1  g10106(.A0(new_n10296_), .A1(\asqrt[25] ), .B0(new_n10298_), .Y(new_n10299_));
  OAI21X1  g10107(.A0(new_n10284_), .A1(new_n10271_), .B0(new_n10291_), .Y(new_n10300_));
  AOI21X1  g10108(.A0(new_n10300_), .A1(\asqrt[60] ), .B0(\asqrt[61] ), .Y(new_n10301_));
  AOI21X1  g10109(.A0(new_n10301_), .A1(new_n10293_), .B0(new_n10299_), .Y(new_n10302_));
  OAI21X1  g10110(.A0(new_n10302_), .A1(new_n10294_), .B0(\asqrt[62] ), .Y(new_n10303_));
  AND2X1   g10111(.A(new_n9799_), .B(new_n9791_), .Y(new_n10304_));
  NOR3X1   g10112(.A(new_n10304_), .B(new_n9845_), .C(new_n9792_), .Y(new_n10305_));
  NOR3X1   g10113(.A(new_n9833_), .B(new_n10304_), .C(new_n9792_), .Y(new_n10306_));
  NOR2X1   g10114(.A(new_n10306_), .B(new_n9797_), .Y(new_n10307_));
  AOI21X1  g10115(.A0(new_n10305_), .A1(\asqrt[25] ), .B0(new_n10307_), .Y(new_n10308_));
  NOR3X1   g10116(.A(new_n10302_), .B(new_n10294_), .C(\asqrt[62] ), .Y(new_n10309_));
  OAI21X1  g10117(.A0(new_n10309_), .A1(new_n10308_), .B0(new_n10303_), .Y(new_n10310_));
  NOR4X1   g10118(.A(new_n9833_), .B(new_n9806_), .C(new_n9849_), .D(new_n9848_), .Y(new_n10311_));
  NOR3X1   g10119(.A(new_n9833_), .B(new_n9806_), .C(new_n9848_), .Y(new_n10312_));
  NOR2X1   g10120(.A(new_n10312_), .B(new_n9805_), .Y(new_n10313_));
  NOR2X1   g10121(.A(new_n10313_), .B(new_n10311_), .Y(new_n10314_));
  INVX1    g10122(.A(new_n10314_), .Y(new_n10315_));
  AND2X1   g10123(.A(new_n9814_), .B(new_n9807_), .Y(new_n10316_));
  AOI21X1  g10124(.A0(new_n10316_), .A1(\asqrt[25] ), .B0(new_n9874_), .Y(new_n10317_));
  AND2X1   g10125(.A(new_n10317_), .B(new_n10315_), .Y(new_n10318_));
  AOI21X1  g10126(.A0(new_n10318_), .A1(new_n10310_), .B0(\asqrt[63] ), .Y(new_n10319_));
  NOR2X1   g10127(.A(new_n10309_), .B(new_n10308_), .Y(new_n10320_));
  NAND2X1  g10128(.A(new_n10314_), .B(new_n10303_), .Y(new_n10321_));
  AOI21X1  g10129(.A0(new_n9857_), .A1(new_n9853_), .B0(new_n9813_), .Y(new_n10322_));
  AOI21X1  g10130(.A0(new_n9814_), .A1(new_n9807_), .B0(new_n193_), .Y(new_n10323_));
  OAI21X1  g10131(.A0(new_n10322_), .A1(new_n9807_), .B0(new_n10323_), .Y(new_n10324_));
  INVX1    g10132(.A(new_n9812_), .Y(new_n10325_));
  NOR4X1   g10133(.A(new_n9830_), .B(new_n9824_), .C(new_n10325_), .D(new_n9809_), .Y(new_n10326_));
  OAI21X1  g10134(.A0(new_n9821_), .A1(new_n9820_), .B0(new_n10326_), .Y(new_n10327_));
  NOR2X1   g10135(.A(new_n10327_), .B(new_n9819_), .Y(new_n10328_));
  INVX1    g10136(.A(new_n10328_), .Y(new_n10329_));
  AND2X1   g10137(.A(new_n10329_), .B(new_n10324_), .Y(new_n10330_));
  OAI21X1  g10138(.A0(new_n10321_), .A1(new_n10320_), .B0(new_n10330_), .Y(new_n10331_));
  NOR2X1   g10139(.A(new_n10331_), .B(new_n10319_), .Y(new_n10332_));
  INVX1    g10140(.A(\a[48] ), .Y(new_n10333_));
  AND2X1   g10141(.A(new_n10300_), .B(\asqrt[60] ), .Y(new_n10334_));
  OR2X1    g10142(.A(new_n10284_), .B(new_n10271_), .Y(new_n10335_));
  AND2X1   g10143(.A(new_n10291_), .B(new_n292_), .Y(new_n10336_));
  AOI21X1  g10144(.A0(new_n10336_), .A1(new_n10335_), .B0(new_n10289_), .Y(new_n10337_));
  OAI21X1  g10145(.A0(new_n10337_), .A1(new_n10334_), .B0(\asqrt[61] ), .Y(new_n10338_));
  INVX1    g10146(.A(new_n10299_), .Y(new_n10339_));
  OAI21X1  g10147(.A0(new_n10274_), .A1(new_n292_), .B0(new_n217_), .Y(new_n10340_));
  OAI21X1  g10148(.A0(new_n10340_), .A1(new_n10337_), .B0(new_n10339_), .Y(new_n10341_));
  AOI21X1  g10149(.A0(new_n10341_), .A1(new_n10338_), .B0(new_n199_), .Y(new_n10342_));
  INVX1    g10150(.A(new_n10308_), .Y(new_n10343_));
  NAND3X1  g10151(.A(new_n10341_), .B(new_n10338_), .C(new_n199_), .Y(new_n10344_));
  AOI21X1  g10152(.A0(new_n10344_), .A1(new_n10343_), .B0(new_n10342_), .Y(new_n10345_));
  INVX1    g10153(.A(new_n10318_), .Y(new_n10346_));
  OAI21X1  g10154(.A0(new_n10346_), .A1(new_n10345_), .B0(new_n193_), .Y(new_n10347_));
  OR2X1    g10155(.A(new_n10309_), .B(new_n10308_), .Y(new_n10348_));
  AND2X1   g10156(.A(new_n10314_), .B(new_n10303_), .Y(new_n10349_));
  INVX1    g10157(.A(new_n10330_), .Y(new_n10350_));
  AOI21X1  g10158(.A0(new_n10349_), .A1(new_n10348_), .B0(new_n10350_), .Y(new_n10351_));
  AOI21X1  g10159(.A0(new_n10351_), .A1(new_n10347_), .B0(new_n10333_), .Y(new_n10352_));
  NOR3X1   g10160(.A(\a[48] ), .B(\a[47] ), .C(\a[46] ), .Y(new_n10353_));
  OAI21X1  g10161(.A0(new_n10353_), .A1(new_n10352_), .B0(\asqrt[25] ), .Y(new_n10354_));
  OAI21X1  g10162(.A0(new_n10331_), .A1(new_n10319_), .B0(\a[48] ), .Y(new_n10355_));
  OR2X1    g10163(.A(new_n10353_), .B(new_n9830_), .Y(new_n10356_));
  NOR4X1   g10164(.A(new_n10356_), .B(new_n9824_), .C(new_n9874_), .D(new_n9819_), .Y(new_n10357_));
  AND2X1   g10165(.A(new_n10357_), .B(new_n10355_), .Y(new_n10358_));
  INVX1    g10166(.A(\a[49] ), .Y(new_n10359_));
  AOI21X1  g10167(.A0(new_n10351_), .A1(new_n10347_), .B0(\a[48] ), .Y(new_n10360_));
  OAI21X1  g10168(.A0(new_n10331_), .A1(new_n10319_), .B0(new_n9837_), .Y(new_n10361_));
  OAI21X1  g10169(.A0(new_n10360_), .A1(new_n10359_), .B0(new_n10361_), .Y(new_n10362_));
  OAI21X1  g10170(.A0(new_n10362_), .A1(new_n10358_), .B0(new_n10354_), .Y(new_n10363_));
  AND2X1   g10171(.A(new_n10363_), .B(\asqrt[26] ), .Y(new_n10364_));
  NAND2X1  g10172(.A(new_n10357_), .B(new_n10355_), .Y(new_n10365_));
  OAI21X1  g10173(.A0(new_n10331_), .A1(new_n10319_), .B0(new_n10333_), .Y(new_n10366_));
  INVX1    g10174(.A(new_n9837_), .Y(new_n10367_));
  AOI21X1  g10175(.A0(new_n10351_), .A1(new_n10347_), .B0(new_n10367_), .Y(new_n10368_));
  AOI21X1  g10176(.A0(new_n10366_), .A1(\a[49] ), .B0(new_n10368_), .Y(new_n10369_));
  NAND2X1  g10177(.A(new_n10369_), .B(new_n10365_), .Y(new_n10370_));
  AND2X1   g10178(.A(new_n10354_), .B(new_n9353_), .Y(new_n10371_));
  INVX1    g10179(.A(new_n10324_), .Y(new_n10372_));
  NOR3X1   g10180(.A(new_n10328_), .B(new_n10372_), .C(new_n9833_), .Y(new_n10373_));
  OAI21X1  g10181(.A0(new_n10321_), .A1(new_n10320_), .B0(new_n10373_), .Y(new_n10374_));
  OR2X1    g10182(.A(new_n10374_), .B(new_n10319_), .Y(new_n10375_));
  AOI21X1  g10183(.A0(new_n10375_), .A1(new_n10361_), .B0(new_n9836_), .Y(new_n10376_));
  OAI21X1  g10184(.A0(new_n10374_), .A1(new_n10319_), .B0(new_n9836_), .Y(new_n10377_));
  NOR2X1   g10185(.A(new_n10377_), .B(new_n10368_), .Y(new_n10378_));
  NOR2X1   g10186(.A(new_n10378_), .B(new_n10376_), .Y(new_n10379_));
  AOI21X1  g10187(.A0(new_n10371_), .A1(new_n10370_), .B0(new_n10379_), .Y(new_n10380_));
  OAI21X1  g10188(.A0(new_n10380_), .A1(new_n10364_), .B0(\asqrt[27] ), .Y(new_n10381_));
  NOR3X1   g10189(.A(new_n9870_), .B(new_n9860_), .C(new_n9872_), .Y(new_n10382_));
  OAI21X1  g10190(.A0(new_n10331_), .A1(new_n10319_), .B0(new_n10382_), .Y(new_n10383_));
  NOR2X1   g10191(.A(new_n9860_), .B(new_n9872_), .Y(new_n10384_));
  OAI21X1  g10192(.A0(new_n10331_), .A1(new_n10319_), .B0(new_n10384_), .Y(new_n10385_));
  NAND2X1  g10193(.A(new_n10385_), .B(new_n9870_), .Y(new_n10386_));
  NAND2X1  g10194(.A(new_n10386_), .B(new_n10383_), .Y(new_n10387_));
  INVX1    g10195(.A(new_n10353_), .Y(new_n10388_));
  AOI21X1  g10196(.A0(new_n10388_), .A1(new_n10355_), .B0(new_n9833_), .Y(new_n10389_));
  AOI21X1  g10197(.A0(new_n10369_), .A1(new_n10365_), .B0(new_n10389_), .Y(new_n10390_));
  OAI21X1  g10198(.A0(new_n10390_), .A1(new_n9353_), .B0(new_n8874_), .Y(new_n10391_));
  OAI21X1  g10199(.A0(new_n10391_), .A1(new_n10380_), .B0(new_n10387_), .Y(new_n10392_));
  AOI21X1  g10200(.A0(new_n10392_), .A1(new_n10381_), .B0(new_n8412_), .Y(new_n10393_));
  AOI21X1  g10201(.A0(new_n9873_), .A1(new_n9871_), .B0(new_n9908_), .Y(new_n10394_));
  AND2X1   g10202(.A(new_n10394_), .B(new_n9905_), .Y(new_n10395_));
  OAI21X1  g10203(.A0(new_n10331_), .A1(new_n10319_), .B0(new_n10395_), .Y(new_n10396_));
  AOI22X1  g10204(.A0(new_n9873_), .A1(new_n9871_), .B0(new_n9865_), .B1(\asqrt[27] ), .Y(new_n10397_));
  OAI21X1  g10205(.A0(new_n10331_), .A1(new_n10319_), .B0(new_n10397_), .Y(new_n10398_));
  NAND2X1  g10206(.A(new_n10398_), .B(new_n9908_), .Y(new_n10399_));
  AND2X1   g10207(.A(new_n10399_), .B(new_n10396_), .Y(new_n10400_));
  INVX1    g10208(.A(new_n10400_), .Y(new_n10401_));
  NAND3X1  g10209(.A(new_n10392_), .B(new_n10381_), .C(new_n8412_), .Y(new_n10402_));
  AOI21X1  g10210(.A0(new_n10402_), .A1(new_n10401_), .B0(new_n10393_), .Y(new_n10403_));
  OR2X1    g10211(.A(new_n10403_), .B(new_n7970_), .Y(new_n10404_));
  OR2X1    g10212(.A(new_n10390_), .B(new_n9353_), .Y(new_n10405_));
  AND2X1   g10213(.A(new_n10369_), .B(new_n10365_), .Y(new_n10406_));
  OR2X1    g10214(.A(new_n10389_), .B(\asqrt[26] ), .Y(new_n10407_));
  OR2X1    g10215(.A(new_n10378_), .B(new_n10376_), .Y(new_n10408_));
  OAI21X1  g10216(.A0(new_n10407_), .A1(new_n10406_), .B0(new_n10408_), .Y(new_n10409_));
  AOI21X1  g10217(.A0(new_n10409_), .A1(new_n10405_), .B0(new_n8874_), .Y(new_n10410_));
  AND2X1   g10218(.A(new_n10386_), .B(new_n10383_), .Y(new_n10411_));
  AOI21X1  g10219(.A0(new_n10363_), .A1(\asqrt[26] ), .B0(\asqrt[27] ), .Y(new_n10412_));
  AOI21X1  g10220(.A0(new_n10412_), .A1(new_n10409_), .B0(new_n10411_), .Y(new_n10413_));
  NOR3X1   g10221(.A(new_n10413_), .B(new_n10410_), .C(\asqrt[28] ), .Y(new_n10414_));
  NOR2X1   g10222(.A(new_n10414_), .B(new_n10400_), .Y(new_n10415_));
  INVX1    g10223(.A(new_n10332_), .Y(\asqrt[24] ));
  AND2X1   g10224(.A(new_n9911_), .B(new_n9909_), .Y(new_n10417_));
  NOR3X1   g10225(.A(new_n10417_), .B(new_n9889_), .C(new_n9910_), .Y(new_n10418_));
  NOR2X1   g10226(.A(new_n10417_), .B(new_n9910_), .Y(new_n10419_));
  OAI21X1  g10227(.A0(new_n10331_), .A1(new_n10319_), .B0(new_n10419_), .Y(new_n10420_));
  AOI22X1  g10228(.A0(new_n10420_), .A1(new_n9889_), .B0(new_n10418_), .B1(\asqrt[24] ), .Y(new_n10421_));
  INVX1    g10229(.A(new_n10421_), .Y(new_n10422_));
  OAI21X1  g10230(.A0(new_n10413_), .A1(new_n10410_), .B0(\asqrt[28] ), .Y(new_n10423_));
  NAND2X1  g10231(.A(new_n10423_), .B(new_n7970_), .Y(new_n10424_));
  OAI21X1  g10232(.A0(new_n10424_), .A1(new_n10415_), .B0(new_n10422_), .Y(new_n10425_));
  AOI21X1  g10233(.A0(new_n10425_), .A1(new_n10404_), .B0(new_n7527_), .Y(new_n10426_));
  NAND4X1  g10234(.A(\asqrt[24] ), .B(new_n9902_), .C(new_n9900_), .D(new_n9929_), .Y(new_n10427_));
  NOR3X1   g10235(.A(new_n10332_), .B(new_n9913_), .C(new_n9893_), .Y(new_n10428_));
  OAI21X1  g10236(.A0(new_n10428_), .A1(new_n9900_), .B0(new_n10427_), .Y(new_n10429_));
  INVX1    g10237(.A(new_n10429_), .Y(new_n10430_));
  OAI21X1  g10238(.A0(new_n10414_), .A1(new_n10400_), .B0(new_n10423_), .Y(new_n10431_));
  AOI21X1  g10239(.A0(new_n10431_), .A1(\asqrt[29] ), .B0(\asqrt[30] ), .Y(new_n10432_));
  AOI21X1  g10240(.A0(new_n10432_), .A1(new_n10425_), .B0(new_n10430_), .Y(new_n10433_));
  OAI21X1  g10241(.A0(new_n10433_), .A1(new_n10426_), .B0(\asqrt[31] ), .Y(new_n10434_));
  AND2X1   g10242(.A(new_n9958_), .B(new_n9957_), .Y(new_n10435_));
  NOR3X1   g10243(.A(new_n10435_), .B(new_n9920_), .C(new_n9956_), .Y(new_n10436_));
  NOR3X1   g10244(.A(new_n10332_), .B(new_n10435_), .C(new_n9956_), .Y(new_n10437_));
  NOR2X1   g10245(.A(new_n10437_), .B(new_n9919_), .Y(new_n10438_));
  AOI21X1  g10246(.A0(new_n10436_), .A1(\asqrt[24] ), .B0(new_n10438_), .Y(new_n10439_));
  NOR3X1   g10247(.A(new_n10433_), .B(new_n10426_), .C(\asqrt[31] ), .Y(new_n10440_));
  OAI21X1  g10248(.A0(new_n10440_), .A1(new_n10439_), .B0(new_n10434_), .Y(new_n10441_));
  AND2X1   g10249(.A(new_n10441_), .B(\asqrt[32] ), .Y(new_n10442_));
  INVX1    g10250(.A(new_n10439_), .Y(new_n10443_));
  AND2X1   g10251(.A(new_n10431_), .B(\asqrt[29] ), .Y(new_n10444_));
  OR2X1    g10252(.A(new_n10414_), .B(new_n10400_), .Y(new_n10445_));
  AND2X1   g10253(.A(new_n10423_), .B(new_n7970_), .Y(new_n10446_));
  AOI21X1  g10254(.A0(new_n10446_), .A1(new_n10445_), .B0(new_n10421_), .Y(new_n10447_));
  OAI21X1  g10255(.A0(new_n10447_), .A1(new_n10444_), .B0(\asqrt[30] ), .Y(new_n10448_));
  OAI21X1  g10256(.A0(new_n10403_), .A1(new_n7970_), .B0(new_n7527_), .Y(new_n10449_));
  OAI21X1  g10257(.A0(new_n10449_), .A1(new_n10447_), .B0(new_n10429_), .Y(new_n10450_));
  NAND3X1  g10258(.A(new_n10450_), .B(new_n10448_), .C(new_n7103_), .Y(new_n10451_));
  NAND2X1  g10259(.A(new_n10451_), .B(new_n10443_), .Y(new_n10452_));
  AND2X1   g10260(.A(new_n9931_), .B(new_n9922_), .Y(new_n10453_));
  NOR3X1   g10261(.A(new_n10453_), .B(new_n9961_), .C(new_n9923_), .Y(new_n10454_));
  NOR3X1   g10262(.A(new_n10332_), .B(new_n10453_), .C(new_n9923_), .Y(new_n10455_));
  NOR2X1   g10263(.A(new_n10455_), .B(new_n9928_), .Y(new_n10456_));
  AOI21X1  g10264(.A0(new_n10454_), .A1(\asqrt[24] ), .B0(new_n10456_), .Y(new_n10457_));
  AND2X1   g10265(.A(new_n10434_), .B(new_n6699_), .Y(new_n10458_));
  AOI21X1  g10266(.A0(new_n10458_), .A1(new_n10452_), .B0(new_n10457_), .Y(new_n10459_));
  OAI21X1  g10267(.A0(new_n10459_), .A1(new_n10442_), .B0(\asqrt[33] ), .Y(new_n10460_));
  OR4X1    g10268(.A(new_n10332_), .B(new_n9939_), .C(new_n9965_), .D(new_n9964_), .Y(new_n10461_));
  OR2X1    g10269(.A(new_n9939_), .B(new_n9964_), .Y(new_n10462_));
  OAI21X1  g10270(.A0(new_n10462_), .A1(new_n10332_), .B0(new_n9965_), .Y(new_n10463_));
  AND2X1   g10271(.A(new_n10463_), .B(new_n10461_), .Y(new_n10464_));
  INVX1    g10272(.A(new_n10464_), .Y(new_n10465_));
  AOI21X1  g10273(.A0(new_n10450_), .A1(new_n10448_), .B0(new_n7103_), .Y(new_n10466_));
  AOI21X1  g10274(.A0(new_n10451_), .A1(new_n10443_), .B0(new_n10466_), .Y(new_n10467_));
  OAI21X1  g10275(.A0(new_n10467_), .A1(new_n6699_), .B0(new_n6294_), .Y(new_n10468_));
  OAI21X1  g10276(.A0(new_n10468_), .A1(new_n10459_), .B0(new_n10465_), .Y(new_n10469_));
  AOI21X1  g10277(.A0(new_n10469_), .A1(new_n10460_), .B0(new_n5941_), .Y(new_n10470_));
  AOI21X1  g10278(.A0(new_n9947_), .A1(new_n9942_), .B0(new_n9982_), .Y(new_n10471_));
  AND2X1   g10279(.A(new_n10471_), .B(new_n9980_), .Y(new_n10472_));
  AOI22X1  g10280(.A0(new_n9947_), .A1(new_n9942_), .B0(new_n9940_), .B1(\asqrt[33] ), .Y(new_n10473_));
  AOI21X1  g10281(.A0(new_n10473_), .A1(\asqrt[24] ), .B0(new_n9946_), .Y(new_n10474_));
  AOI21X1  g10282(.A0(new_n10472_), .A1(\asqrt[24] ), .B0(new_n10474_), .Y(new_n10475_));
  INVX1    g10283(.A(new_n10475_), .Y(new_n10476_));
  NAND3X1  g10284(.A(new_n10469_), .B(new_n10460_), .C(new_n5941_), .Y(new_n10477_));
  AOI21X1  g10285(.A0(new_n10477_), .A1(new_n10476_), .B0(new_n10470_), .Y(new_n10478_));
  OR2X1    g10286(.A(new_n10478_), .B(new_n5541_), .Y(new_n10479_));
  AND2X1   g10287(.A(new_n10477_), .B(new_n10476_), .Y(new_n10480_));
  AND2X1   g10288(.A(new_n9986_), .B(new_n9984_), .Y(new_n10481_));
  NOR3X1   g10289(.A(new_n10481_), .B(new_n9955_), .C(new_n9985_), .Y(new_n10482_));
  NOR3X1   g10290(.A(new_n10332_), .B(new_n10481_), .C(new_n9985_), .Y(new_n10483_));
  NOR2X1   g10291(.A(new_n10483_), .B(new_n9954_), .Y(new_n10484_));
  AOI21X1  g10292(.A0(new_n10482_), .A1(\asqrt[24] ), .B0(new_n10484_), .Y(new_n10485_));
  INVX1    g10293(.A(new_n10485_), .Y(new_n10486_));
  OR2X1    g10294(.A(new_n10467_), .B(new_n6699_), .Y(new_n10487_));
  AND2X1   g10295(.A(new_n10451_), .B(new_n10443_), .Y(new_n10488_));
  INVX1    g10296(.A(new_n10457_), .Y(new_n10489_));
  NAND2X1  g10297(.A(new_n10434_), .B(new_n6699_), .Y(new_n10490_));
  OAI21X1  g10298(.A0(new_n10490_), .A1(new_n10488_), .B0(new_n10489_), .Y(new_n10491_));
  AOI21X1  g10299(.A0(new_n10491_), .A1(new_n10487_), .B0(new_n6294_), .Y(new_n10492_));
  AOI21X1  g10300(.A0(new_n10441_), .A1(\asqrt[32] ), .B0(\asqrt[33] ), .Y(new_n10493_));
  AOI21X1  g10301(.A0(new_n10493_), .A1(new_n10491_), .B0(new_n10464_), .Y(new_n10494_));
  OAI21X1  g10302(.A0(new_n10494_), .A1(new_n10492_), .B0(\asqrt[34] ), .Y(new_n10495_));
  NAND2X1  g10303(.A(new_n10495_), .B(new_n5541_), .Y(new_n10496_));
  OAI21X1  g10304(.A0(new_n10496_), .A1(new_n10480_), .B0(new_n10486_), .Y(new_n10497_));
  AOI21X1  g10305(.A0(new_n10497_), .A1(new_n10479_), .B0(new_n5176_), .Y(new_n10498_));
  NAND4X1  g10306(.A(\asqrt[24] ), .B(new_n9977_), .C(new_n9975_), .D(new_n9995_), .Y(new_n10499_));
  OR2X1    g10307(.A(new_n9988_), .B(new_n9970_), .Y(new_n10500_));
  OAI21X1  g10308(.A0(new_n10500_), .A1(new_n10332_), .B0(new_n9976_), .Y(new_n10501_));
  AND2X1   g10309(.A(new_n10501_), .B(new_n10499_), .Y(new_n10502_));
  NOR3X1   g10310(.A(new_n10494_), .B(new_n10492_), .C(\asqrt[34] ), .Y(new_n10503_));
  OAI21X1  g10311(.A0(new_n10503_), .A1(new_n10475_), .B0(new_n10495_), .Y(new_n10504_));
  AOI21X1  g10312(.A0(new_n10504_), .A1(\asqrt[35] ), .B0(\asqrt[36] ), .Y(new_n10505_));
  AOI21X1  g10313(.A0(new_n10505_), .A1(new_n10497_), .B0(new_n10502_), .Y(new_n10506_));
  OAI21X1  g10314(.A0(new_n10506_), .A1(new_n10498_), .B0(\asqrt[37] ), .Y(new_n10507_));
  AND2X1   g10315(.A(new_n10023_), .B(new_n10022_), .Y(new_n10508_));
  NOR3X1   g10316(.A(new_n10508_), .B(new_n9994_), .C(new_n10021_), .Y(new_n10509_));
  NOR3X1   g10317(.A(new_n10332_), .B(new_n10508_), .C(new_n10021_), .Y(new_n10510_));
  NOR2X1   g10318(.A(new_n10510_), .B(new_n9993_), .Y(new_n10511_));
  AOI21X1  g10319(.A0(new_n10509_), .A1(\asqrt[24] ), .B0(new_n10511_), .Y(new_n10512_));
  NOR3X1   g10320(.A(new_n10506_), .B(new_n10498_), .C(\asqrt[37] ), .Y(new_n10513_));
  OAI21X1  g10321(.A0(new_n10513_), .A1(new_n10512_), .B0(new_n10507_), .Y(new_n10514_));
  AND2X1   g10322(.A(new_n10514_), .B(\asqrt[38] ), .Y(new_n10515_));
  INVX1    g10323(.A(new_n10512_), .Y(new_n10516_));
  AND2X1   g10324(.A(new_n10504_), .B(\asqrt[35] ), .Y(new_n10517_));
  NAND2X1  g10325(.A(new_n10477_), .B(new_n10476_), .Y(new_n10518_));
  AND2X1   g10326(.A(new_n10495_), .B(new_n5541_), .Y(new_n10519_));
  AOI21X1  g10327(.A0(new_n10519_), .A1(new_n10518_), .B0(new_n10485_), .Y(new_n10520_));
  OAI21X1  g10328(.A0(new_n10520_), .A1(new_n10517_), .B0(\asqrt[36] ), .Y(new_n10521_));
  INVX1    g10329(.A(new_n10502_), .Y(new_n10522_));
  OAI21X1  g10330(.A0(new_n10478_), .A1(new_n5541_), .B0(new_n5176_), .Y(new_n10523_));
  OAI21X1  g10331(.A0(new_n10523_), .A1(new_n10520_), .B0(new_n10522_), .Y(new_n10524_));
  NAND3X1  g10332(.A(new_n10524_), .B(new_n10521_), .C(new_n4826_), .Y(new_n10525_));
  NAND2X1  g10333(.A(new_n10525_), .B(new_n10516_), .Y(new_n10526_));
  AND2X1   g10334(.A(new_n10005_), .B(new_n9997_), .Y(new_n10527_));
  NOR3X1   g10335(.A(new_n10527_), .B(new_n10026_), .C(new_n9998_), .Y(new_n10528_));
  NOR3X1   g10336(.A(new_n10332_), .B(new_n10527_), .C(new_n9998_), .Y(new_n10529_));
  NOR2X1   g10337(.A(new_n10529_), .B(new_n10003_), .Y(new_n10530_));
  AOI21X1  g10338(.A0(new_n10528_), .A1(\asqrt[24] ), .B0(new_n10530_), .Y(new_n10531_));
  AND2X1   g10339(.A(new_n10507_), .B(new_n4493_), .Y(new_n10532_));
  AOI21X1  g10340(.A0(new_n10532_), .A1(new_n10526_), .B0(new_n10531_), .Y(new_n10533_));
  OAI21X1  g10341(.A0(new_n10533_), .A1(new_n10515_), .B0(\asqrt[39] ), .Y(new_n10534_));
  NAND4X1  g10342(.A(\asqrt[24] ), .B(new_n10034_), .C(new_n10012_), .D(new_n10007_), .Y(new_n10535_));
  NAND2X1  g10343(.A(new_n10034_), .B(new_n10007_), .Y(new_n10536_));
  OAI21X1  g10344(.A0(new_n10536_), .A1(new_n10332_), .B0(new_n10033_), .Y(new_n10537_));
  AND2X1   g10345(.A(new_n10537_), .B(new_n10535_), .Y(new_n10538_));
  INVX1    g10346(.A(new_n10538_), .Y(new_n10539_));
  AOI21X1  g10347(.A0(new_n10524_), .A1(new_n10521_), .B0(new_n4826_), .Y(new_n10540_));
  AOI21X1  g10348(.A0(new_n10525_), .A1(new_n10516_), .B0(new_n10540_), .Y(new_n10541_));
  OAI21X1  g10349(.A0(new_n10541_), .A1(new_n4493_), .B0(new_n4165_), .Y(new_n10542_));
  OAI21X1  g10350(.A0(new_n10542_), .A1(new_n10533_), .B0(new_n10539_), .Y(new_n10543_));
  AOI21X1  g10351(.A0(new_n10543_), .A1(new_n10534_), .B0(new_n3863_), .Y(new_n10544_));
  AOI21X1  g10352(.A0(new_n10030_), .A1(new_n10016_), .B0(new_n10070_), .Y(new_n10545_));
  AND2X1   g10353(.A(new_n10545_), .B(new_n10068_), .Y(new_n10546_));
  AOI22X1  g10354(.A0(new_n10030_), .A1(new_n10016_), .B0(new_n10014_), .B1(\asqrt[39] ), .Y(new_n10547_));
  AOI21X1  g10355(.A0(new_n10547_), .A1(\asqrt[24] ), .B0(new_n10020_), .Y(new_n10548_));
  AOI21X1  g10356(.A0(new_n10546_), .A1(\asqrt[24] ), .B0(new_n10548_), .Y(new_n10549_));
  INVX1    g10357(.A(new_n10549_), .Y(new_n10550_));
  NAND3X1  g10358(.A(new_n10543_), .B(new_n10534_), .C(new_n3863_), .Y(new_n10551_));
  AOI21X1  g10359(.A0(new_n10551_), .A1(new_n10550_), .B0(new_n10544_), .Y(new_n10552_));
  OR2X1    g10360(.A(new_n10552_), .B(new_n3564_), .Y(new_n10553_));
  AND2X1   g10361(.A(new_n10551_), .B(new_n10550_), .Y(new_n10554_));
  OR2X1    g10362(.A(new_n10541_), .B(new_n4493_), .Y(new_n10555_));
  AND2X1   g10363(.A(new_n10525_), .B(new_n10516_), .Y(new_n10556_));
  INVX1    g10364(.A(new_n10531_), .Y(new_n10557_));
  NAND2X1  g10365(.A(new_n10507_), .B(new_n4493_), .Y(new_n10558_));
  OAI21X1  g10366(.A0(new_n10558_), .A1(new_n10556_), .B0(new_n10557_), .Y(new_n10559_));
  AOI21X1  g10367(.A0(new_n10559_), .A1(new_n10555_), .B0(new_n4165_), .Y(new_n10560_));
  AOI21X1  g10368(.A0(new_n10514_), .A1(\asqrt[38] ), .B0(\asqrt[39] ), .Y(new_n10561_));
  AOI21X1  g10369(.A0(new_n10561_), .A1(new_n10559_), .B0(new_n10538_), .Y(new_n10562_));
  OAI21X1  g10370(.A0(new_n10562_), .A1(new_n10560_), .B0(\asqrt[40] ), .Y(new_n10563_));
  NAND2X1  g10371(.A(new_n10563_), .B(new_n3564_), .Y(new_n10564_));
  AND2X1   g10372(.A(new_n10074_), .B(new_n10072_), .Y(new_n10565_));
  NOR3X1   g10373(.A(new_n10042_), .B(new_n10565_), .C(new_n10073_), .Y(new_n10566_));
  NOR3X1   g10374(.A(new_n10332_), .B(new_n10565_), .C(new_n10073_), .Y(new_n10567_));
  NOR2X1   g10375(.A(new_n10567_), .B(new_n10041_), .Y(new_n10568_));
  AOI21X1  g10376(.A0(new_n10566_), .A1(\asqrt[24] ), .B0(new_n10568_), .Y(new_n10569_));
  INVX1    g10377(.A(new_n10569_), .Y(new_n10570_));
  OAI21X1  g10378(.A0(new_n10564_), .A1(new_n10554_), .B0(new_n10570_), .Y(new_n10571_));
  AOI21X1  g10379(.A0(new_n10571_), .A1(new_n10553_), .B0(new_n3276_), .Y(new_n10572_));
  NAND4X1  g10380(.A(\asqrt[24] ), .B(new_n10051_), .C(new_n10049_), .D(new_n10076_), .Y(new_n10573_));
  NAND2X1  g10381(.A(new_n10051_), .B(new_n10076_), .Y(new_n10574_));
  OAI21X1  g10382(.A0(new_n10574_), .A1(new_n10332_), .B0(new_n10050_), .Y(new_n10575_));
  AND2X1   g10383(.A(new_n10575_), .B(new_n10573_), .Y(new_n10576_));
  NOR3X1   g10384(.A(new_n10562_), .B(new_n10560_), .C(\asqrt[40] ), .Y(new_n10577_));
  OAI21X1  g10385(.A0(new_n10577_), .A1(new_n10549_), .B0(new_n10563_), .Y(new_n10578_));
  AOI21X1  g10386(.A0(new_n10578_), .A1(\asqrt[41] ), .B0(\asqrt[42] ), .Y(new_n10579_));
  AOI21X1  g10387(.A0(new_n10579_), .A1(new_n10571_), .B0(new_n10576_), .Y(new_n10580_));
  OAI21X1  g10388(.A0(new_n10580_), .A1(new_n10572_), .B0(\asqrt[43] ), .Y(new_n10581_));
  AND2X1   g10389(.A(new_n10097_), .B(new_n10096_), .Y(new_n10582_));
  NOR3X1   g10390(.A(new_n10582_), .B(new_n10059_), .C(new_n10095_), .Y(new_n10583_));
  NOR3X1   g10391(.A(new_n10332_), .B(new_n10582_), .C(new_n10095_), .Y(new_n10584_));
  NOR2X1   g10392(.A(new_n10584_), .B(new_n10058_), .Y(new_n10585_));
  AOI21X1  g10393(.A0(new_n10583_), .A1(\asqrt[24] ), .B0(new_n10585_), .Y(new_n10586_));
  NOR3X1   g10394(.A(new_n10580_), .B(new_n10572_), .C(\asqrt[43] ), .Y(new_n10587_));
  OAI21X1  g10395(.A0(new_n10587_), .A1(new_n10586_), .B0(new_n10581_), .Y(new_n10588_));
  AND2X1   g10396(.A(new_n10588_), .B(\asqrt[44] ), .Y(new_n10589_));
  INVX1    g10397(.A(new_n10586_), .Y(new_n10590_));
  AND2X1   g10398(.A(new_n10578_), .B(\asqrt[41] ), .Y(new_n10591_));
  NAND2X1  g10399(.A(new_n10551_), .B(new_n10550_), .Y(new_n10592_));
  AND2X1   g10400(.A(new_n10563_), .B(new_n3564_), .Y(new_n10593_));
  AOI21X1  g10401(.A0(new_n10593_), .A1(new_n10592_), .B0(new_n10569_), .Y(new_n10594_));
  OAI21X1  g10402(.A0(new_n10594_), .A1(new_n10591_), .B0(\asqrt[42] ), .Y(new_n10595_));
  INVX1    g10403(.A(new_n10576_), .Y(new_n10596_));
  OAI21X1  g10404(.A0(new_n10552_), .A1(new_n3564_), .B0(new_n3276_), .Y(new_n10597_));
  OAI21X1  g10405(.A0(new_n10597_), .A1(new_n10594_), .B0(new_n10596_), .Y(new_n10598_));
  NAND3X1  g10406(.A(new_n10598_), .B(new_n10595_), .C(new_n3008_), .Y(new_n10599_));
  NAND2X1  g10407(.A(new_n10599_), .B(new_n10590_), .Y(new_n10600_));
  AND2X1   g10408(.A(new_n10079_), .B(new_n10061_), .Y(new_n10601_));
  NOR3X1   g10409(.A(new_n10601_), .B(new_n10100_), .C(new_n10062_), .Y(new_n10602_));
  NOR3X1   g10410(.A(new_n10332_), .B(new_n10601_), .C(new_n10062_), .Y(new_n10603_));
  NOR2X1   g10411(.A(new_n10603_), .B(new_n10067_), .Y(new_n10604_));
  AOI21X1  g10412(.A0(new_n10602_), .A1(\asqrt[24] ), .B0(new_n10604_), .Y(new_n10605_));
  AND2X1   g10413(.A(new_n10581_), .B(new_n2769_), .Y(new_n10606_));
  AOI21X1  g10414(.A0(new_n10606_), .A1(new_n10600_), .B0(new_n10605_), .Y(new_n10607_));
  OAI21X1  g10415(.A0(new_n10607_), .A1(new_n10589_), .B0(\asqrt[45] ), .Y(new_n10608_));
  NAND4X1  g10416(.A(\asqrt[24] ), .B(new_n10114_), .C(new_n10086_), .D(new_n10081_), .Y(new_n10609_));
  NAND2X1  g10417(.A(new_n10114_), .B(new_n10081_), .Y(new_n10610_));
  OAI21X1  g10418(.A0(new_n10610_), .A1(new_n10332_), .B0(new_n10113_), .Y(new_n10611_));
  AND2X1   g10419(.A(new_n10611_), .B(new_n10609_), .Y(new_n10612_));
  INVX1    g10420(.A(new_n10612_), .Y(new_n10613_));
  AOI21X1  g10421(.A0(new_n10598_), .A1(new_n10595_), .B0(new_n3008_), .Y(new_n10614_));
  AOI21X1  g10422(.A0(new_n10599_), .A1(new_n10590_), .B0(new_n10614_), .Y(new_n10615_));
  OAI21X1  g10423(.A0(new_n10615_), .A1(new_n2769_), .B0(new_n2570_), .Y(new_n10616_));
  OAI21X1  g10424(.A0(new_n10616_), .A1(new_n10607_), .B0(new_n10613_), .Y(new_n10617_));
  AOI21X1  g10425(.A0(new_n10617_), .A1(new_n10608_), .B0(new_n2263_), .Y(new_n10618_));
  AOI21X1  g10426(.A0(new_n10104_), .A1(new_n10090_), .B0(new_n10130_), .Y(new_n10619_));
  AND2X1   g10427(.A(new_n10619_), .B(new_n10128_), .Y(new_n10620_));
  AOI22X1  g10428(.A0(new_n10104_), .A1(new_n10090_), .B0(new_n10088_), .B1(\asqrt[45] ), .Y(new_n10621_));
  AOI21X1  g10429(.A0(new_n10621_), .A1(\asqrt[24] ), .B0(new_n10094_), .Y(new_n10622_));
  AOI21X1  g10430(.A0(new_n10620_), .A1(\asqrt[24] ), .B0(new_n10622_), .Y(new_n10623_));
  INVX1    g10431(.A(new_n10623_), .Y(new_n10624_));
  NAND3X1  g10432(.A(new_n10617_), .B(new_n10608_), .C(new_n2263_), .Y(new_n10625_));
  AOI21X1  g10433(.A0(new_n10625_), .A1(new_n10624_), .B0(new_n10618_), .Y(new_n10626_));
  OR2X1    g10434(.A(new_n10626_), .B(new_n2040_), .Y(new_n10627_));
  AND2X1   g10435(.A(new_n10625_), .B(new_n10624_), .Y(new_n10628_));
  AND2X1   g10436(.A(new_n10134_), .B(new_n10132_), .Y(new_n10629_));
  NOR3X1   g10437(.A(new_n10629_), .B(new_n10112_), .C(new_n10133_), .Y(new_n10630_));
  NOR3X1   g10438(.A(new_n10332_), .B(new_n10629_), .C(new_n10133_), .Y(new_n10631_));
  NOR2X1   g10439(.A(new_n10631_), .B(new_n10111_), .Y(new_n10632_));
  AOI21X1  g10440(.A0(new_n10630_), .A1(\asqrt[24] ), .B0(new_n10632_), .Y(new_n10633_));
  INVX1    g10441(.A(new_n10633_), .Y(new_n10634_));
  OR2X1    g10442(.A(new_n10615_), .B(new_n2769_), .Y(new_n10635_));
  AND2X1   g10443(.A(new_n10599_), .B(new_n10590_), .Y(new_n10636_));
  INVX1    g10444(.A(new_n10605_), .Y(new_n10637_));
  NAND2X1  g10445(.A(new_n10581_), .B(new_n2769_), .Y(new_n10638_));
  OAI21X1  g10446(.A0(new_n10638_), .A1(new_n10636_), .B0(new_n10637_), .Y(new_n10639_));
  AOI21X1  g10447(.A0(new_n10639_), .A1(new_n10635_), .B0(new_n2570_), .Y(new_n10640_));
  AOI21X1  g10448(.A0(new_n10588_), .A1(\asqrt[44] ), .B0(\asqrt[45] ), .Y(new_n10641_));
  AOI21X1  g10449(.A0(new_n10641_), .A1(new_n10639_), .B0(new_n10612_), .Y(new_n10642_));
  OAI21X1  g10450(.A0(new_n10642_), .A1(new_n10640_), .B0(\asqrt[46] ), .Y(new_n10643_));
  NAND2X1  g10451(.A(new_n10643_), .B(new_n2040_), .Y(new_n10644_));
  OAI21X1  g10452(.A0(new_n10644_), .A1(new_n10628_), .B0(new_n10634_), .Y(new_n10645_));
  AOI21X1  g10453(.A0(new_n10645_), .A1(new_n10627_), .B0(new_n1834_), .Y(new_n10646_));
  NAND4X1  g10454(.A(\asqrt[24] ), .B(new_n10125_), .C(new_n10123_), .D(new_n10143_), .Y(new_n10647_));
  OR2X1    g10455(.A(new_n10136_), .B(new_n10118_), .Y(new_n10648_));
  OAI21X1  g10456(.A0(new_n10648_), .A1(new_n10332_), .B0(new_n10124_), .Y(new_n10649_));
  AND2X1   g10457(.A(new_n10649_), .B(new_n10647_), .Y(new_n10650_));
  NOR3X1   g10458(.A(new_n10642_), .B(new_n10640_), .C(\asqrt[46] ), .Y(new_n10651_));
  OAI21X1  g10459(.A0(new_n10651_), .A1(new_n10623_), .B0(new_n10643_), .Y(new_n10652_));
  AOI21X1  g10460(.A0(new_n10652_), .A1(\asqrt[47] ), .B0(\asqrt[48] ), .Y(new_n10653_));
  AOI21X1  g10461(.A0(new_n10653_), .A1(new_n10645_), .B0(new_n10650_), .Y(new_n10654_));
  OAI21X1  g10462(.A0(new_n10654_), .A1(new_n10646_), .B0(\asqrt[49] ), .Y(new_n10655_));
  AND2X1   g10463(.A(new_n10180_), .B(new_n10179_), .Y(new_n10656_));
  NOR3X1   g10464(.A(new_n10656_), .B(new_n10142_), .C(new_n10178_), .Y(new_n10657_));
  NOR3X1   g10465(.A(new_n10332_), .B(new_n10656_), .C(new_n10178_), .Y(new_n10658_));
  NOR2X1   g10466(.A(new_n10658_), .B(new_n10141_), .Y(new_n10659_));
  AOI21X1  g10467(.A0(new_n10657_), .A1(\asqrt[24] ), .B0(new_n10659_), .Y(new_n10660_));
  NOR3X1   g10468(.A(new_n10654_), .B(new_n10646_), .C(\asqrt[49] ), .Y(new_n10661_));
  OAI21X1  g10469(.A0(new_n10661_), .A1(new_n10660_), .B0(new_n10655_), .Y(new_n10662_));
  AND2X1   g10470(.A(new_n10662_), .B(\asqrt[50] ), .Y(new_n10663_));
  INVX1    g10471(.A(new_n10660_), .Y(new_n10664_));
  AND2X1   g10472(.A(new_n10652_), .B(\asqrt[47] ), .Y(new_n10665_));
  NAND2X1  g10473(.A(new_n10625_), .B(new_n10624_), .Y(new_n10666_));
  AND2X1   g10474(.A(new_n10643_), .B(new_n2040_), .Y(new_n10667_));
  AOI21X1  g10475(.A0(new_n10667_), .A1(new_n10666_), .B0(new_n10633_), .Y(new_n10668_));
  OAI21X1  g10476(.A0(new_n10668_), .A1(new_n10665_), .B0(\asqrt[48] ), .Y(new_n10669_));
  INVX1    g10477(.A(new_n10650_), .Y(new_n10670_));
  OAI21X1  g10478(.A0(new_n10626_), .A1(new_n2040_), .B0(new_n1834_), .Y(new_n10671_));
  OAI21X1  g10479(.A0(new_n10671_), .A1(new_n10668_), .B0(new_n10670_), .Y(new_n10672_));
  NAND3X1  g10480(.A(new_n10672_), .B(new_n10669_), .C(new_n1632_), .Y(new_n10673_));
  NAND2X1  g10481(.A(new_n10673_), .B(new_n10664_), .Y(new_n10674_));
  AND2X1   g10482(.A(new_n10153_), .B(new_n10145_), .Y(new_n10675_));
  NOR3X1   g10483(.A(new_n10675_), .B(new_n10183_), .C(new_n10146_), .Y(new_n10676_));
  NOR3X1   g10484(.A(new_n10332_), .B(new_n10675_), .C(new_n10146_), .Y(new_n10677_));
  NOR2X1   g10485(.A(new_n10677_), .B(new_n10151_), .Y(new_n10678_));
  AOI21X1  g10486(.A0(new_n10676_), .A1(\asqrt[24] ), .B0(new_n10678_), .Y(new_n10679_));
  AND2X1   g10487(.A(new_n10655_), .B(new_n1469_), .Y(new_n10680_));
  AOI21X1  g10488(.A0(new_n10680_), .A1(new_n10674_), .B0(new_n10679_), .Y(new_n10681_));
  OAI21X1  g10489(.A0(new_n10681_), .A1(new_n10663_), .B0(\asqrt[51] ), .Y(new_n10682_));
  OR4X1    g10490(.A(new_n10332_), .B(new_n10161_), .C(new_n10187_), .D(new_n10186_), .Y(new_n10683_));
  OR2X1    g10491(.A(new_n10161_), .B(new_n10186_), .Y(new_n10684_));
  OAI21X1  g10492(.A0(new_n10684_), .A1(new_n10332_), .B0(new_n10187_), .Y(new_n10685_));
  AND2X1   g10493(.A(new_n10685_), .B(new_n10683_), .Y(new_n10686_));
  INVX1    g10494(.A(new_n10686_), .Y(new_n10687_));
  AOI21X1  g10495(.A0(new_n10672_), .A1(new_n10669_), .B0(new_n1632_), .Y(new_n10688_));
  AOI21X1  g10496(.A0(new_n10673_), .A1(new_n10664_), .B0(new_n10688_), .Y(new_n10689_));
  OAI21X1  g10497(.A0(new_n10689_), .A1(new_n1469_), .B0(new_n1277_), .Y(new_n10690_));
  OAI21X1  g10498(.A0(new_n10690_), .A1(new_n10681_), .B0(new_n10687_), .Y(new_n10691_));
  AOI21X1  g10499(.A0(new_n10691_), .A1(new_n10682_), .B0(new_n1111_), .Y(new_n10692_));
  AOI21X1  g10500(.A0(new_n10169_), .A1(new_n10164_), .B0(new_n10204_), .Y(new_n10693_));
  AND2X1   g10501(.A(new_n10693_), .B(new_n10202_), .Y(new_n10694_));
  AOI22X1  g10502(.A0(new_n10169_), .A1(new_n10164_), .B0(new_n10162_), .B1(\asqrt[51] ), .Y(new_n10695_));
  AOI21X1  g10503(.A0(new_n10695_), .A1(\asqrt[24] ), .B0(new_n10168_), .Y(new_n10696_));
  AOI21X1  g10504(.A0(new_n10694_), .A1(\asqrt[24] ), .B0(new_n10696_), .Y(new_n10697_));
  INVX1    g10505(.A(new_n10697_), .Y(new_n10698_));
  NAND3X1  g10506(.A(new_n10691_), .B(new_n10682_), .C(new_n1111_), .Y(new_n10699_));
  AOI21X1  g10507(.A0(new_n10699_), .A1(new_n10698_), .B0(new_n10692_), .Y(new_n10700_));
  OR2X1    g10508(.A(new_n10700_), .B(new_n968_), .Y(new_n10701_));
  OR2X1    g10509(.A(new_n10689_), .B(new_n1469_), .Y(new_n10702_));
  AND2X1   g10510(.A(new_n10673_), .B(new_n10664_), .Y(new_n10703_));
  INVX1    g10511(.A(new_n10679_), .Y(new_n10704_));
  NAND2X1  g10512(.A(new_n10655_), .B(new_n1469_), .Y(new_n10705_));
  OAI21X1  g10513(.A0(new_n10705_), .A1(new_n10703_), .B0(new_n10704_), .Y(new_n10706_));
  AOI21X1  g10514(.A0(new_n10706_), .A1(new_n10702_), .B0(new_n1277_), .Y(new_n10707_));
  AOI21X1  g10515(.A0(new_n10662_), .A1(\asqrt[50] ), .B0(\asqrt[51] ), .Y(new_n10708_));
  AOI21X1  g10516(.A0(new_n10708_), .A1(new_n10706_), .B0(new_n10686_), .Y(new_n10709_));
  NOR3X1   g10517(.A(new_n10709_), .B(new_n10707_), .C(\asqrt[52] ), .Y(new_n10710_));
  NOR2X1   g10518(.A(new_n10710_), .B(new_n10697_), .Y(new_n10711_));
  AND2X1   g10519(.A(new_n10208_), .B(new_n10206_), .Y(new_n10712_));
  NOR3X1   g10520(.A(new_n10712_), .B(new_n10177_), .C(new_n10207_), .Y(new_n10713_));
  NOR3X1   g10521(.A(new_n10332_), .B(new_n10712_), .C(new_n10207_), .Y(new_n10714_));
  NOR2X1   g10522(.A(new_n10714_), .B(new_n10176_), .Y(new_n10715_));
  AOI21X1  g10523(.A0(new_n10713_), .A1(\asqrt[24] ), .B0(new_n10715_), .Y(new_n10716_));
  INVX1    g10524(.A(new_n10716_), .Y(new_n10717_));
  OAI21X1  g10525(.A0(new_n10709_), .A1(new_n10707_), .B0(\asqrt[52] ), .Y(new_n10718_));
  NAND2X1  g10526(.A(new_n10718_), .B(new_n968_), .Y(new_n10719_));
  OAI21X1  g10527(.A0(new_n10719_), .A1(new_n10711_), .B0(new_n10717_), .Y(new_n10720_));
  AOI21X1  g10528(.A0(new_n10720_), .A1(new_n10701_), .B0(new_n902_), .Y(new_n10721_));
  OR4X1    g10529(.A(new_n10332_), .B(new_n10210_), .C(new_n10198_), .D(new_n10192_), .Y(new_n10722_));
  OR2X1    g10530(.A(new_n10210_), .B(new_n10192_), .Y(new_n10723_));
  OAI21X1  g10531(.A0(new_n10723_), .A1(new_n10332_), .B0(new_n10198_), .Y(new_n10724_));
  AND2X1   g10532(.A(new_n10724_), .B(new_n10722_), .Y(new_n10725_));
  OAI21X1  g10533(.A0(new_n10710_), .A1(new_n10697_), .B0(new_n10718_), .Y(new_n10726_));
  AOI21X1  g10534(.A0(new_n10726_), .A1(\asqrt[53] ), .B0(\asqrt[54] ), .Y(new_n10727_));
  AOI21X1  g10535(.A0(new_n10727_), .A1(new_n10720_), .B0(new_n10725_), .Y(new_n10728_));
  OAI21X1  g10536(.A0(new_n10728_), .A1(new_n10721_), .B0(\asqrt[55] ), .Y(new_n10729_));
  AND2X1   g10537(.A(new_n10254_), .B(new_n10253_), .Y(new_n10730_));
  NOR3X1   g10538(.A(new_n10730_), .B(new_n10216_), .C(new_n10252_), .Y(new_n10731_));
  NOR3X1   g10539(.A(new_n10332_), .B(new_n10730_), .C(new_n10252_), .Y(new_n10732_));
  NOR2X1   g10540(.A(new_n10732_), .B(new_n10215_), .Y(new_n10733_));
  AOI21X1  g10541(.A0(new_n10731_), .A1(\asqrt[24] ), .B0(new_n10733_), .Y(new_n10734_));
  NOR3X1   g10542(.A(new_n10728_), .B(new_n10721_), .C(\asqrt[55] ), .Y(new_n10735_));
  OAI21X1  g10543(.A0(new_n10735_), .A1(new_n10734_), .B0(new_n10729_), .Y(new_n10736_));
  AND2X1   g10544(.A(new_n10736_), .B(\asqrt[56] ), .Y(new_n10737_));
  INVX1    g10545(.A(new_n10734_), .Y(new_n10738_));
  AND2X1   g10546(.A(new_n10726_), .B(\asqrt[53] ), .Y(new_n10739_));
  OR2X1    g10547(.A(new_n10710_), .B(new_n10697_), .Y(new_n10740_));
  AND2X1   g10548(.A(new_n10718_), .B(new_n968_), .Y(new_n10741_));
  AOI21X1  g10549(.A0(new_n10741_), .A1(new_n10740_), .B0(new_n10716_), .Y(new_n10742_));
  OAI21X1  g10550(.A0(new_n10742_), .A1(new_n10739_), .B0(\asqrt[54] ), .Y(new_n10743_));
  INVX1    g10551(.A(new_n10725_), .Y(new_n10744_));
  OAI21X1  g10552(.A0(new_n10700_), .A1(new_n968_), .B0(new_n902_), .Y(new_n10745_));
  OAI21X1  g10553(.A0(new_n10745_), .A1(new_n10742_), .B0(new_n10744_), .Y(new_n10746_));
  NAND3X1  g10554(.A(new_n10746_), .B(new_n10743_), .C(new_n697_), .Y(new_n10747_));
  NAND2X1  g10555(.A(new_n10747_), .B(new_n10738_), .Y(new_n10748_));
  AND2X1   g10556(.A(new_n10227_), .B(new_n10219_), .Y(new_n10749_));
  NOR3X1   g10557(.A(new_n10749_), .B(new_n10257_), .C(new_n10220_), .Y(new_n10750_));
  NOR3X1   g10558(.A(new_n10332_), .B(new_n10749_), .C(new_n10220_), .Y(new_n10751_));
  NOR2X1   g10559(.A(new_n10751_), .B(new_n10225_), .Y(new_n10752_));
  AOI21X1  g10560(.A0(new_n10750_), .A1(\asqrt[24] ), .B0(new_n10752_), .Y(new_n10753_));
  AND2X1   g10561(.A(new_n10729_), .B(new_n582_), .Y(new_n10754_));
  AOI21X1  g10562(.A0(new_n10754_), .A1(new_n10748_), .B0(new_n10753_), .Y(new_n10755_));
  OAI21X1  g10563(.A0(new_n10755_), .A1(new_n10737_), .B0(\asqrt[57] ), .Y(new_n10756_));
  OR4X1    g10564(.A(new_n10332_), .B(new_n10235_), .C(new_n10261_), .D(new_n10260_), .Y(new_n10757_));
  OR2X1    g10565(.A(new_n10235_), .B(new_n10260_), .Y(new_n10758_));
  OAI21X1  g10566(.A0(new_n10758_), .A1(new_n10332_), .B0(new_n10261_), .Y(new_n10759_));
  AND2X1   g10567(.A(new_n10759_), .B(new_n10757_), .Y(new_n10760_));
  INVX1    g10568(.A(new_n10760_), .Y(new_n10761_));
  AOI21X1  g10569(.A0(new_n10746_), .A1(new_n10743_), .B0(new_n697_), .Y(new_n10762_));
  AOI21X1  g10570(.A0(new_n10747_), .A1(new_n10738_), .B0(new_n10762_), .Y(new_n10763_));
  OAI21X1  g10571(.A0(new_n10763_), .A1(new_n582_), .B0(new_n481_), .Y(new_n10764_));
  OAI21X1  g10572(.A0(new_n10764_), .A1(new_n10755_), .B0(new_n10761_), .Y(new_n10765_));
  AOI21X1  g10573(.A0(new_n10765_), .A1(new_n10756_), .B0(new_n399_), .Y(new_n10766_));
  AOI21X1  g10574(.A0(new_n10243_), .A1(new_n10238_), .B0(new_n10278_), .Y(new_n10767_));
  AND2X1   g10575(.A(new_n10767_), .B(new_n10276_), .Y(new_n10768_));
  AOI22X1  g10576(.A0(new_n10243_), .A1(new_n10238_), .B0(new_n10236_), .B1(\asqrt[57] ), .Y(new_n10769_));
  AOI21X1  g10577(.A0(new_n10769_), .A1(\asqrt[24] ), .B0(new_n10242_), .Y(new_n10770_));
  AOI21X1  g10578(.A0(new_n10768_), .A1(\asqrt[24] ), .B0(new_n10770_), .Y(new_n10771_));
  INVX1    g10579(.A(new_n10771_), .Y(new_n10772_));
  NAND3X1  g10580(.A(new_n10765_), .B(new_n10756_), .C(new_n399_), .Y(new_n10773_));
  AOI21X1  g10581(.A0(new_n10773_), .A1(new_n10772_), .B0(new_n10766_), .Y(new_n10774_));
  OR2X1    g10582(.A(new_n10774_), .B(new_n328_), .Y(new_n10775_));
  OR2X1    g10583(.A(new_n10763_), .B(new_n582_), .Y(new_n10776_));
  AND2X1   g10584(.A(new_n10747_), .B(new_n10738_), .Y(new_n10777_));
  INVX1    g10585(.A(new_n10753_), .Y(new_n10778_));
  NAND2X1  g10586(.A(new_n10729_), .B(new_n582_), .Y(new_n10779_));
  OAI21X1  g10587(.A0(new_n10779_), .A1(new_n10777_), .B0(new_n10778_), .Y(new_n10780_));
  AOI21X1  g10588(.A0(new_n10780_), .A1(new_n10776_), .B0(new_n481_), .Y(new_n10781_));
  AOI21X1  g10589(.A0(new_n10736_), .A1(\asqrt[56] ), .B0(\asqrt[57] ), .Y(new_n10782_));
  AOI21X1  g10590(.A0(new_n10782_), .A1(new_n10780_), .B0(new_n10760_), .Y(new_n10783_));
  NOR3X1   g10591(.A(new_n10783_), .B(new_n10781_), .C(\asqrt[58] ), .Y(new_n10784_));
  NOR2X1   g10592(.A(new_n10784_), .B(new_n10771_), .Y(new_n10785_));
  AND2X1   g10593(.A(new_n10282_), .B(new_n10280_), .Y(new_n10786_));
  NOR3X1   g10594(.A(new_n10786_), .B(new_n10251_), .C(new_n10281_), .Y(new_n10787_));
  NOR3X1   g10595(.A(new_n10332_), .B(new_n10786_), .C(new_n10281_), .Y(new_n10788_));
  NOR2X1   g10596(.A(new_n10788_), .B(new_n10250_), .Y(new_n10789_));
  AOI21X1  g10597(.A0(new_n10787_), .A1(\asqrt[24] ), .B0(new_n10789_), .Y(new_n10790_));
  INVX1    g10598(.A(new_n10790_), .Y(new_n10791_));
  OAI21X1  g10599(.A0(new_n10783_), .A1(new_n10781_), .B0(\asqrt[58] ), .Y(new_n10792_));
  NAND2X1  g10600(.A(new_n10792_), .B(new_n328_), .Y(new_n10793_));
  OAI21X1  g10601(.A0(new_n10793_), .A1(new_n10785_), .B0(new_n10791_), .Y(new_n10794_));
  AOI21X1  g10602(.A0(new_n10794_), .A1(new_n10775_), .B0(new_n292_), .Y(new_n10795_));
  OR4X1    g10603(.A(new_n10332_), .B(new_n10284_), .C(new_n10272_), .D(new_n10266_), .Y(new_n10796_));
  OR2X1    g10604(.A(new_n10284_), .B(new_n10266_), .Y(new_n10797_));
  OAI21X1  g10605(.A0(new_n10797_), .A1(new_n10332_), .B0(new_n10272_), .Y(new_n10798_));
  AND2X1   g10606(.A(new_n10798_), .B(new_n10796_), .Y(new_n10799_));
  OAI21X1  g10607(.A0(new_n10784_), .A1(new_n10771_), .B0(new_n10792_), .Y(new_n10800_));
  AOI21X1  g10608(.A0(new_n10800_), .A1(\asqrt[59] ), .B0(\asqrt[60] ), .Y(new_n10801_));
  AOI21X1  g10609(.A0(new_n10801_), .A1(new_n10794_), .B0(new_n10799_), .Y(new_n10802_));
  OAI21X1  g10610(.A0(new_n10802_), .A1(new_n10795_), .B0(\asqrt[61] ), .Y(new_n10803_));
  AND2X1   g10611(.A(new_n10336_), .B(new_n10335_), .Y(new_n10804_));
  NOR3X1   g10612(.A(new_n10804_), .B(new_n10290_), .C(new_n10334_), .Y(new_n10805_));
  NOR3X1   g10613(.A(new_n10332_), .B(new_n10804_), .C(new_n10334_), .Y(new_n10806_));
  NOR2X1   g10614(.A(new_n10806_), .B(new_n10289_), .Y(new_n10807_));
  AOI21X1  g10615(.A0(new_n10805_), .A1(\asqrt[24] ), .B0(new_n10807_), .Y(new_n10808_));
  NOR3X1   g10616(.A(new_n10802_), .B(new_n10795_), .C(\asqrt[61] ), .Y(new_n10809_));
  OAI21X1  g10617(.A0(new_n10809_), .A1(new_n10808_), .B0(new_n10803_), .Y(new_n10810_));
  AND2X1   g10618(.A(new_n10810_), .B(\asqrt[62] ), .Y(new_n10811_));
  OR2X1    g10619(.A(new_n10809_), .B(new_n10808_), .Y(new_n10812_));
  AND2X1   g10620(.A(new_n10301_), .B(new_n10293_), .Y(new_n10813_));
  NOR3X1   g10621(.A(new_n10813_), .B(new_n10339_), .C(new_n10294_), .Y(new_n10814_));
  NOR3X1   g10622(.A(new_n10332_), .B(new_n10813_), .C(new_n10294_), .Y(new_n10815_));
  NOR2X1   g10623(.A(new_n10815_), .B(new_n10299_), .Y(new_n10816_));
  AOI21X1  g10624(.A0(new_n10814_), .A1(\asqrt[24] ), .B0(new_n10816_), .Y(new_n10817_));
  AND2X1   g10625(.A(new_n10803_), .B(new_n199_), .Y(new_n10818_));
  AOI21X1  g10626(.A0(new_n10818_), .A1(new_n10812_), .B0(new_n10817_), .Y(new_n10819_));
  NOR4X1   g10627(.A(new_n10332_), .B(new_n10309_), .C(new_n10343_), .D(new_n10342_), .Y(new_n10820_));
  NAND3X1  g10628(.A(\asqrt[24] ), .B(new_n10344_), .C(new_n10303_), .Y(new_n10821_));
  AOI21X1  g10629(.A0(new_n10821_), .A1(new_n10343_), .B0(new_n10820_), .Y(new_n10822_));
  INVX1    g10630(.A(new_n10822_), .Y(new_n10823_));
  NOR3X1   g10631(.A(new_n10332_), .B(new_n10314_), .C(new_n10345_), .Y(new_n10824_));
  AOI21X1  g10632(.A0(new_n10349_), .A1(new_n10348_), .B0(new_n10824_), .Y(new_n10825_));
  AND2X1   g10633(.A(new_n10825_), .B(new_n10823_), .Y(new_n10826_));
  OAI21X1  g10634(.A0(new_n10819_), .A1(new_n10811_), .B0(new_n10826_), .Y(new_n10827_));
  AND2X1   g10635(.A(new_n10800_), .B(\asqrt[59] ), .Y(new_n10828_));
  OR2X1    g10636(.A(new_n10784_), .B(new_n10771_), .Y(new_n10829_));
  AND2X1   g10637(.A(new_n10792_), .B(new_n328_), .Y(new_n10830_));
  AOI21X1  g10638(.A0(new_n10830_), .A1(new_n10829_), .B0(new_n10790_), .Y(new_n10831_));
  OAI21X1  g10639(.A0(new_n10831_), .A1(new_n10828_), .B0(\asqrt[60] ), .Y(new_n10832_));
  INVX1    g10640(.A(new_n10799_), .Y(new_n10833_));
  OAI21X1  g10641(.A0(new_n10774_), .A1(new_n328_), .B0(new_n292_), .Y(new_n10834_));
  OAI21X1  g10642(.A0(new_n10834_), .A1(new_n10831_), .B0(new_n10833_), .Y(new_n10835_));
  AOI21X1  g10643(.A0(new_n10835_), .A1(new_n10832_), .B0(new_n217_), .Y(new_n10836_));
  INVX1    g10644(.A(new_n10808_), .Y(new_n10837_));
  NAND3X1  g10645(.A(new_n10835_), .B(new_n10832_), .C(new_n217_), .Y(new_n10838_));
  AOI21X1  g10646(.A0(new_n10838_), .A1(new_n10837_), .B0(new_n10836_), .Y(new_n10839_));
  OAI21X1  g10647(.A0(new_n10839_), .A1(new_n199_), .B0(new_n10822_), .Y(new_n10840_));
  AOI21X1  g10648(.A0(new_n10351_), .A1(new_n10347_), .B0(new_n10314_), .Y(new_n10841_));
  AOI21X1  g10649(.A0(new_n10315_), .A1(new_n10310_), .B0(new_n193_), .Y(new_n10842_));
  OAI21X1  g10650(.A0(new_n10841_), .A1(new_n10310_), .B0(new_n10842_), .Y(new_n10843_));
  OR2X1    g10651(.A(new_n10321_), .B(new_n10320_), .Y(new_n10844_));
  NOR4X1   g10652(.A(new_n10328_), .B(new_n10372_), .C(new_n10313_), .D(new_n10311_), .Y(new_n10845_));
  NAND3X1  g10653(.A(new_n10845_), .B(new_n10844_), .C(new_n10347_), .Y(new_n10846_));
  AND2X1   g10654(.A(new_n10846_), .B(new_n10843_), .Y(new_n10847_));
  OAI21X1  g10655(.A0(new_n10840_), .A1(new_n10819_), .B0(new_n10847_), .Y(new_n10848_));
  AOI21X1  g10656(.A0(new_n10827_), .A1(new_n193_), .B0(new_n10848_), .Y(new_n10849_));
  NOR2X1   g10657(.A(\a[45] ), .B(\a[44] ), .Y(new_n10850_));
  INVX1    g10658(.A(new_n10850_), .Y(new_n10851_));
  MX2X1    g10659(.A(new_n10851_), .B(new_n10849_), .S0(\a[46] ), .Y(new_n10852_));
  OR2X1    g10660(.A(new_n10852_), .B(new_n10332_), .Y(new_n10853_));
  INVX1    g10661(.A(\a[46] ), .Y(new_n10854_));
  NOR3X1   g10662(.A(\a[46] ), .B(\a[45] ), .C(\a[44] ), .Y(new_n10855_));
  NOR3X1   g10663(.A(new_n10855_), .B(new_n10328_), .C(new_n10372_), .Y(new_n10856_));
  NAND3X1  g10664(.A(new_n10856_), .B(new_n10844_), .C(new_n10347_), .Y(new_n10857_));
  INVX1    g10665(.A(new_n10857_), .Y(new_n10858_));
  OAI21X1  g10666(.A0(new_n10849_), .A1(new_n10854_), .B0(new_n10858_), .Y(new_n10859_));
  OAI21X1  g10667(.A0(new_n10849_), .A1(\a[46] ), .B0(\a[47] ), .Y(new_n10860_));
  NOR2X1   g10668(.A(\a[47] ), .B(\a[46] ), .Y(new_n10861_));
  INVX1    g10669(.A(new_n10861_), .Y(new_n10862_));
  OR2X1    g10670(.A(new_n10849_), .B(new_n10862_), .Y(new_n10863_));
  NAND3X1  g10671(.A(new_n10863_), .B(new_n10860_), .C(new_n10859_), .Y(new_n10864_));
  AOI21X1  g10672(.A0(new_n10864_), .A1(new_n10853_), .B0(new_n9833_), .Y(new_n10865_));
  OR2X1    g10673(.A(new_n10839_), .B(new_n199_), .Y(new_n10866_));
  NOR2X1   g10674(.A(new_n10809_), .B(new_n10808_), .Y(new_n10867_));
  INVX1    g10675(.A(new_n10817_), .Y(new_n10868_));
  NAND2X1  g10676(.A(new_n10803_), .B(new_n199_), .Y(new_n10869_));
  OAI21X1  g10677(.A0(new_n10869_), .A1(new_n10867_), .B0(new_n10868_), .Y(new_n10870_));
  INVX1    g10678(.A(new_n10826_), .Y(new_n10871_));
  AOI21X1  g10679(.A0(new_n10870_), .A1(new_n10866_), .B0(new_n10871_), .Y(new_n10872_));
  AOI21X1  g10680(.A0(new_n10810_), .A1(\asqrt[62] ), .B0(new_n10823_), .Y(new_n10873_));
  INVX1    g10681(.A(new_n10847_), .Y(new_n10874_));
  AOI21X1  g10682(.A0(new_n10873_), .A1(new_n10870_), .B0(new_n10874_), .Y(new_n10875_));
  OAI21X1  g10683(.A0(new_n10872_), .A1(\asqrt[63] ), .B0(new_n10875_), .Y(\asqrt[23] ));
  MX2X1    g10684(.A(new_n10850_), .B(\asqrt[23] ), .S0(\a[46] ), .Y(new_n10877_));
  AOI21X1  g10685(.A0(new_n10877_), .A1(\asqrt[24] ), .B0(\asqrt[25] ), .Y(new_n10878_));
  NAND3X1  g10686(.A(new_n10846_), .B(new_n10843_), .C(\asqrt[24] ), .Y(new_n10879_));
  INVX1    g10687(.A(new_n10879_), .Y(new_n10880_));
  OAI21X1  g10688(.A0(new_n10840_), .A1(new_n10819_), .B0(new_n10880_), .Y(new_n10881_));
  AOI21X1  g10689(.A0(new_n10827_), .A1(new_n193_), .B0(new_n10881_), .Y(new_n10882_));
  AOI21X1  g10690(.A0(\asqrt[23] ), .A1(new_n10861_), .B0(new_n10882_), .Y(new_n10883_));
  OR2X1    g10691(.A(new_n10883_), .B(new_n10333_), .Y(new_n10884_));
  AND2X1   g10692(.A(\asqrt[23] ), .B(new_n10861_), .Y(new_n10885_));
  OR2X1    g10693(.A(new_n10882_), .B(\a[48] ), .Y(new_n10886_));
  OR2X1    g10694(.A(new_n10886_), .B(new_n10885_), .Y(new_n10887_));
  AOI22X1  g10695(.A0(new_n10887_), .A1(new_n10884_), .B0(new_n10878_), .B1(new_n10864_), .Y(new_n10888_));
  OAI21X1  g10696(.A0(new_n10888_), .A1(new_n10865_), .B0(\asqrt[26] ), .Y(new_n10889_));
  AND2X1   g10697(.A(new_n10365_), .B(new_n10354_), .Y(new_n10890_));
  NAND3X1  g10698(.A(new_n10890_), .B(\asqrt[23] ), .C(new_n10362_), .Y(new_n10891_));
  INVX1    g10699(.A(new_n10890_), .Y(new_n10892_));
  OAI21X1  g10700(.A0(new_n10892_), .A1(new_n10849_), .B0(new_n10369_), .Y(new_n10893_));
  AND2X1   g10701(.A(new_n10893_), .B(new_n10891_), .Y(new_n10894_));
  NOR3X1   g10702(.A(new_n10888_), .B(new_n10865_), .C(\asqrt[26] ), .Y(new_n10895_));
  OAI21X1  g10703(.A0(new_n10895_), .A1(new_n10894_), .B0(new_n10889_), .Y(new_n10896_));
  AND2X1   g10704(.A(new_n10896_), .B(\asqrt[27] ), .Y(new_n10897_));
  INVX1    g10705(.A(new_n10894_), .Y(new_n10898_));
  AND2X1   g10706(.A(new_n10877_), .B(\asqrt[24] ), .Y(new_n10899_));
  AOI21X1  g10707(.A0(\asqrt[23] ), .A1(\a[46] ), .B0(new_n10857_), .Y(new_n10900_));
  INVX1    g10708(.A(\a[47] ), .Y(new_n10901_));
  AOI21X1  g10709(.A0(\asqrt[23] ), .A1(new_n10854_), .B0(new_n10901_), .Y(new_n10902_));
  NOR3X1   g10710(.A(new_n10885_), .B(new_n10902_), .C(new_n10900_), .Y(new_n10903_));
  OAI21X1  g10711(.A0(new_n10903_), .A1(new_n10899_), .B0(\asqrt[25] ), .Y(new_n10904_));
  OAI21X1  g10712(.A0(new_n10852_), .A1(new_n10332_), .B0(new_n9833_), .Y(new_n10905_));
  OAI22X1  g10713(.A0(new_n10886_), .A1(new_n10885_), .B0(new_n10883_), .B1(new_n10333_), .Y(new_n10906_));
  OAI21X1  g10714(.A0(new_n10905_), .A1(new_n10903_), .B0(new_n10906_), .Y(new_n10907_));
  NAND3X1  g10715(.A(new_n10907_), .B(new_n10904_), .C(new_n9353_), .Y(new_n10908_));
  NAND2X1  g10716(.A(new_n10908_), .B(new_n10898_), .Y(new_n10909_));
  AOI21X1  g10717(.A0(new_n10371_), .A1(new_n10370_), .B0(new_n10408_), .Y(new_n10910_));
  NAND3X1  g10718(.A(new_n10910_), .B(\asqrt[23] ), .C(new_n10405_), .Y(new_n10911_));
  OAI22X1  g10719(.A0(new_n10407_), .A1(new_n10406_), .B0(new_n10390_), .B1(new_n9353_), .Y(new_n10912_));
  OAI21X1  g10720(.A0(new_n10912_), .A1(new_n10849_), .B0(new_n10408_), .Y(new_n10913_));
  AND2X1   g10721(.A(new_n10913_), .B(new_n10911_), .Y(new_n10914_));
  AOI21X1  g10722(.A0(new_n10907_), .A1(new_n10904_), .B0(new_n9353_), .Y(new_n10915_));
  NOR2X1   g10723(.A(new_n10915_), .B(\asqrt[27] ), .Y(new_n10916_));
  AOI21X1  g10724(.A0(new_n10916_), .A1(new_n10909_), .B0(new_n10914_), .Y(new_n10917_));
  OAI21X1  g10725(.A0(new_n10917_), .A1(new_n10897_), .B0(\asqrt[28] ), .Y(new_n10918_));
  AND2X1   g10726(.A(new_n10412_), .B(new_n10409_), .Y(new_n10919_));
  OR4X1    g10727(.A(new_n10849_), .B(new_n10919_), .C(new_n10387_), .D(new_n10410_), .Y(new_n10920_));
  OR2X1    g10728(.A(new_n10919_), .B(new_n10410_), .Y(new_n10921_));
  OAI21X1  g10729(.A0(new_n10921_), .A1(new_n10849_), .B0(new_n10387_), .Y(new_n10922_));
  AND2X1   g10730(.A(new_n10922_), .B(new_n10920_), .Y(new_n10923_));
  INVX1    g10731(.A(new_n10923_), .Y(new_n10924_));
  AOI21X1  g10732(.A0(new_n10908_), .A1(new_n10898_), .B0(new_n10915_), .Y(new_n10925_));
  OAI21X1  g10733(.A0(new_n10925_), .A1(new_n8874_), .B0(new_n8412_), .Y(new_n10926_));
  OAI21X1  g10734(.A0(new_n10926_), .A1(new_n10917_), .B0(new_n10924_), .Y(new_n10927_));
  AOI21X1  g10735(.A0(new_n10927_), .A1(new_n10918_), .B0(new_n7970_), .Y(new_n10928_));
  NAND3X1  g10736(.A(new_n10402_), .B(new_n10400_), .C(new_n10423_), .Y(new_n10929_));
  NOR3X1   g10737(.A(new_n10849_), .B(new_n10414_), .C(new_n10393_), .Y(new_n10930_));
  OAI22X1  g10738(.A0(new_n10930_), .A1(new_n10400_), .B0(new_n10929_), .B1(new_n10849_), .Y(new_n10931_));
  NAND3X1  g10739(.A(new_n10927_), .B(new_n10918_), .C(new_n7970_), .Y(new_n10932_));
  AOI21X1  g10740(.A0(new_n10932_), .A1(new_n10931_), .B0(new_n10928_), .Y(new_n10933_));
  OR2X1    g10741(.A(new_n10933_), .B(new_n7527_), .Y(new_n10934_));
  AND2X1   g10742(.A(new_n10932_), .B(new_n10931_), .Y(new_n10935_));
  AND2X1   g10743(.A(new_n10446_), .B(new_n10445_), .Y(new_n10936_));
  NOR4X1   g10744(.A(new_n10849_), .B(new_n10936_), .C(new_n10422_), .D(new_n10444_), .Y(new_n10937_));
  AOI22X1  g10745(.A0(new_n10446_), .A1(new_n10445_), .B0(new_n10431_), .B1(\asqrt[29] ), .Y(new_n10938_));
  AOI21X1  g10746(.A0(new_n10938_), .A1(\asqrt[23] ), .B0(new_n10421_), .Y(new_n10939_));
  NOR2X1   g10747(.A(new_n10939_), .B(new_n10937_), .Y(new_n10940_));
  INVX1    g10748(.A(new_n10940_), .Y(new_n10941_));
  OR2X1    g10749(.A(new_n10928_), .B(\asqrt[30] ), .Y(new_n10942_));
  OAI21X1  g10750(.A0(new_n10942_), .A1(new_n10935_), .B0(new_n10941_), .Y(new_n10943_));
  AOI21X1  g10751(.A0(new_n10943_), .A1(new_n10934_), .B0(new_n7103_), .Y(new_n10944_));
  AND2X1   g10752(.A(new_n10432_), .B(new_n10425_), .Y(new_n10945_));
  NOR3X1   g10753(.A(new_n10945_), .B(new_n10429_), .C(new_n10426_), .Y(new_n10946_));
  NOR2X1   g10754(.A(new_n10945_), .B(new_n10426_), .Y(new_n10947_));
  AOI21X1  g10755(.A0(new_n10947_), .A1(\asqrt[23] ), .B0(new_n10430_), .Y(new_n10948_));
  AOI21X1  g10756(.A0(new_n10946_), .A1(\asqrt[23] ), .B0(new_n10948_), .Y(new_n10949_));
  OR2X1    g10757(.A(new_n10925_), .B(new_n8874_), .Y(new_n10950_));
  AND2X1   g10758(.A(new_n10908_), .B(new_n10898_), .Y(new_n10951_));
  INVX1    g10759(.A(new_n10914_), .Y(new_n10952_));
  OR2X1    g10760(.A(new_n10915_), .B(\asqrt[27] ), .Y(new_n10953_));
  OAI21X1  g10761(.A0(new_n10953_), .A1(new_n10951_), .B0(new_n10952_), .Y(new_n10954_));
  AOI21X1  g10762(.A0(new_n10954_), .A1(new_n10950_), .B0(new_n8412_), .Y(new_n10955_));
  AOI21X1  g10763(.A0(new_n10896_), .A1(\asqrt[27] ), .B0(\asqrt[28] ), .Y(new_n10956_));
  AOI21X1  g10764(.A0(new_n10956_), .A1(new_n10954_), .B0(new_n10923_), .Y(new_n10957_));
  OAI21X1  g10765(.A0(new_n10957_), .A1(new_n10955_), .B0(\asqrt[29] ), .Y(new_n10958_));
  INVX1    g10766(.A(new_n10931_), .Y(new_n10959_));
  NOR3X1   g10767(.A(new_n10957_), .B(new_n10955_), .C(\asqrt[29] ), .Y(new_n10960_));
  OAI21X1  g10768(.A0(new_n10960_), .A1(new_n10959_), .B0(new_n10958_), .Y(new_n10961_));
  AOI21X1  g10769(.A0(new_n10961_), .A1(\asqrt[30] ), .B0(\asqrt[31] ), .Y(new_n10962_));
  AOI21X1  g10770(.A0(new_n10962_), .A1(new_n10943_), .B0(new_n10949_), .Y(new_n10963_));
  OAI21X1  g10771(.A0(new_n10963_), .A1(new_n10944_), .B0(\asqrt[32] ), .Y(new_n10964_));
  OR4X1    g10772(.A(new_n10849_), .B(new_n10440_), .C(new_n10443_), .D(new_n10466_), .Y(new_n10965_));
  NAND2X1  g10773(.A(new_n10451_), .B(new_n10434_), .Y(new_n10966_));
  OAI21X1  g10774(.A0(new_n10966_), .A1(new_n10849_), .B0(new_n10443_), .Y(new_n10967_));
  AND2X1   g10775(.A(new_n10967_), .B(new_n10965_), .Y(new_n10968_));
  NOR3X1   g10776(.A(new_n10963_), .B(new_n10944_), .C(\asqrt[32] ), .Y(new_n10969_));
  OAI21X1  g10777(.A0(new_n10969_), .A1(new_n10968_), .B0(new_n10964_), .Y(new_n10970_));
  AND2X1   g10778(.A(new_n10970_), .B(\asqrt[33] ), .Y(new_n10971_));
  INVX1    g10779(.A(new_n10968_), .Y(new_n10972_));
  AND2X1   g10780(.A(new_n10961_), .B(\asqrt[30] ), .Y(new_n10973_));
  NAND2X1  g10781(.A(new_n10932_), .B(new_n10931_), .Y(new_n10974_));
  NOR2X1   g10782(.A(new_n10928_), .B(\asqrt[30] ), .Y(new_n10975_));
  AOI21X1  g10783(.A0(new_n10975_), .A1(new_n10974_), .B0(new_n10940_), .Y(new_n10976_));
  OAI21X1  g10784(.A0(new_n10976_), .A1(new_n10973_), .B0(\asqrt[31] ), .Y(new_n10977_));
  INVX1    g10785(.A(new_n10949_), .Y(new_n10978_));
  OAI21X1  g10786(.A0(new_n10933_), .A1(new_n7527_), .B0(new_n7103_), .Y(new_n10979_));
  OAI21X1  g10787(.A0(new_n10979_), .A1(new_n10976_), .B0(new_n10978_), .Y(new_n10980_));
  NAND3X1  g10788(.A(new_n10980_), .B(new_n10977_), .C(new_n6699_), .Y(new_n10981_));
  NAND2X1  g10789(.A(new_n10981_), .B(new_n10972_), .Y(new_n10982_));
  AOI21X1  g10790(.A0(new_n10458_), .A1(new_n10452_), .B0(new_n10489_), .Y(new_n10983_));
  AND2X1   g10791(.A(new_n10983_), .B(new_n10487_), .Y(new_n10984_));
  AOI22X1  g10792(.A0(new_n10458_), .A1(new_n10452_), .B0(new_n10441_), .B1(\asqrt[32] ), .Y(new_n10985_));
  AOI21X1  g10793(.A0(new_n10985_), .A1(\asqrt[23] ), .B0(new_n10457_), .Y(new_n10986_));
  AOI21X1  g10794(.A0(new_n10984_), .A1(\asqrt[23] ), .B0(new_n10986_), .Y(new_n10987_));
  AOI21X1  g10795(.A0(new_n10980_), .A1(new_n10977_), .B0(new_n6699_), .Y(new_n10988_));
  NOR2X1   g10796(.A(new_n10988_), .B(\asqrt[33] ), .Y(new_n10989_));
  AOI21X1  g10797(.A0(new_n10989_), .A1(new_n10982_), .B0(new_n10987_), .Y(new_n10990_));
  OAI21X1  g10798(.A0(new_n10990_), .A1(new_n10971_), .B0(\asqrt[34] ), .Y(new_n10991_));
  AND2X1   g10799(.A(new_n10493_), .B(new_n10491_), .Y(new_n10992_));
  OR4X1    g10800(.A(new_n10849_), .B(new_n10992_), .C(new_n10465_), .D(new_n10492_), .Y(new_n10993_));
  OR2X1    g10801(.A(new_n10992_), .B(new_n10492_), .Y(new_n10994_));
  OAI21X1  g10802(.A0(new_n10994_), .A1(new_n10849_), .B0(new_n10465_), .Y(new_n10995_));
  AND2X1   g10803(.A(new_n10995_), .B(new_n10993_), .Y(new_n10996_));
  INVX1    g10804(.A(new_n10996_), .Y(new_n10997_));
  AOI21X1  g10805(.A0(new_n10981_), .A1(new_n10972_), .B0(new_n10988_), .Y(new_n10998_));
  OAI21X1  g10806(.A0(new_n10998_), .A1(new_n6294_), .B0(new_n5941_), .Y(new_n10999_));
  OAI21X1  g10807(.A0(new_n10999_), .A1(new_n10990_), .B0(new_n10997_), .Y(new_n11000_));
  AOI21X1  g10808(.A0(new_n11000_), .A1(new_n10991_), .B0(new_n5541_), .Y(new_n11001_));
  OR4X1    g10809(.A(new_n10849_), .B(new_n10503_), .C(new_n10476_), .D(new_n10470_), .Y(new_n11002_));
  NAND2X1  g10810(.A(new_n10477_), .B(new_n10495_), .Y(new_n11003_));
  OAI21X1  g10811(.A0(new_n11003_), .A1(new_n10849_), .B0(new_n10476_), .Y(new_n11004_));
  AND2X1   g10812(.A(new_n11004_), .B(new_n11002_), .Y(new_n11005_));
  INVX1    g10813(.A(new_n11005_), .Y(new_n11006_));
  NAND3X1  g10814(.A(new_n11000_), .B(new_n10991_), .C(new_n5541_), .Y(new_n11007_));
  AOI21X1  g10815(.A0(new_n11007_), .A1(new_n11006_), .B0(new_n11001_), .Y(new_n11008_));
  OR2X1    g10816(.A(new_n11008_), .B(new_n5176_), .Y(new_n11009_));
  AND2X1   g10817(.A(new_n11007_), .B(new_n11006_), .Y(new_n11010_));
  AND2X1   g10818(.A(new_n10519_), .B(new_n10518_), .Y(new_n11011_));
  NOR4X1   g10819(.A(new_n10849_), .B(new_n11011_), .C(new_n10486_), .D(new_n10517_), .Y(new_n11012_));
  AOI22X1  g10820(.A0(new_n10519_), .A1(new_n10518_), .B0(new_n10504_), .B1(\asqrt[35] ), .Y(new_n11013_));
  AOI21X1  g10821(.A0(new_n11013_), .A1(\asqrt[23] ), .B0(new_n10485_), .Y(new_n11014_));
  NOR2X1   g10822(.A(new_n11014_), .B(new_n11012_), .Y(new_n11015_));
  INVX1    g10823(.A(new_n11015_), .Y(new_n11016_));
  OR2X1    g10824(.A(new_n11001_), .B(\asqrt[36] ), .Y(new_n11017_));
  OAI21X1  g10825(.A0(new_n11017_), .A1(new_n11010_), .B0(new_n11016_), .Y(new_n11018_));
  AOI21X1  g10826(.A0(new_n11018_), .A1(new_n11009_), .B0(new_n4826_), .Y(new_n11019_));
  OAI21X1  g10827(.A0(new_n10523_), .A1(new_n10520_), .B0(new_n10502_), .Y(new_n11020_));
  OR2X1    g10828(.A(new_n11020_), .B(new_n10498_), .Y(new_n11021_));
  AND2X1   g10829(.A(new_n10505_), .B(new_n10497_), .Y(new_n11022_));
  NOR3X1   g10830(.A(new_n10849_), .B(new_n11022_), .C(new_n10498_), .Y(new_n11023_));
  OAI22X1  g10831(.A0(new_n11023_), .A1(new_n10502_), .B0(new_n11021_), .B1(new_n10849_), .Y(new_n11024_));
  INVX1    g10832(.A(new_n11024_), .Y(new_n11025_));
  OR2X1    g10833(.A(new_n10998_), .B(new_n6294_), .Y(new_n11026_));
  AND2X1   g10834(.A(new_n10981_), .B(new_n10972_), .Y(new_n11027_));
  INVX1    g10835(.A(new_n10987_), .Y(new_n11028_));
  OR2X1    g10836(.A(new_n10988_), .B(\asqrt[33] ), .Y(new_n11029_));
  OAI21X1  g10837(.A0(new_n11029_), .A1(new_n11027_), .B0(new_n11028_), .Y(new_n11030_));
  AOI21X1  g10838(.A0(new_n11030_), .A1(new_n11026_), .B0(new_n5941_), .Y(new_n11031_));
  AOI21X1  g10839(.A0(new_n10970_), .A1(\asqrt[33] ), .B0(\asqrt[34] ), .Y(new_n11032_));
  AOI21X1  g10840(.A0(new_n11032_), .A1(new_n11030_), .B0(new_n10996_), .Y(new_n11033_));
  OAI21X1  g10841(.A0(new_n11033_), .A1(new_n11031_), .B0(\asqrt[35] ), .Y(new_n11034_));
  NOR3X1   g10842(.A(new_n11033_), .B(new_n11031_), .C(\asqrt[35] ), .Y(new_n11035_));
  OAI21X1  g10843(.A0(new_n11035_), .A1(new_n11005_), .B0(new_n11034_), .Y(new_n11036_));
  AOI21X1  g10844(.A0(new_n11036_), .A1(\asqrt[36] ), .B0(\asqrt[37] ), .Y(new_n11037_));
  AOI21X1  g10845(.A0(new_n11037_), .A1(new_n11018_), .B0(new_n11025_), .Y(new_n11038_));
  OAI21X1  g10846(.A0(new_n11038_), .A1(new_n11019_), .B0(\asqrt[38] ), .Y(new_n11039_));
  NAND3X1  g10847(.A(new_n10525_), .B(new_n10512_), .C(new_n10507_), .Y(new_n11040_));
  NOR3X1   g10848(.A(new_n10849_), .B(new_n10513_), .C(new_n10540_), .Y(new_n11041_));
  OAI22X1  g10849(.A0(new_n11041_), .A1(new_n10512_), .B0(new_n11040_), .B1(new_n10849_), .Y(new_n11042_));
  INVX1    g10850(.A(new_n11042_), .Y(new_n11043_));
  NOR3X1   g10851(.A(new_n11038_), .B(new_n11019_), .C(\asqrt[38] ), .Y(new_n11044_));
  OAI21X1  g10852(.A0(new_n11044_), .A1(new_n11043_), .B0(new_n11039_), .Y(new_n11045_));
  AND2X1   g10853(.A(new_n11045_), .B(\asqrt[39] ), .Y(new_n11046_));
  AND2X1   g10854(.A(new_n11036_), .B(\asqrt[36] ), .Y(new_n11047_));
  NAND2X1  g10855(.A(new_n11007_), .B(new_n11006_), .Y(new_n11048_));
  NOR2X1   g10856(.A(new_n11001_), .B(\asqrt[36] ), .Y(new_n11049_));
  AOI21X1  g10857(.A0(new_n11049_), .A1(new_n11048_), .B0(new_n11015_), .Y(new_n11050_));
  OAI21X1  g10858(.A0(new_n11050_), .A1(new_n11047_), .B0(\asqrt[37] ), .Y(new_n11051_));
  OAI21X1  g10859(.A0(new_n11008_), .A1(new_n5176_), .B0(new_n4826_), .Y(new_n11052_));
  OAI21X1  g10860(.A0(new_n11052_), .A1(new_n11050_), .B0(new_n11024_), .Y(new_n11053_));
  NAND3X1  g10861(.A(new_n11053_), .B(new_n11051_), .C(new_n4493_), .Y(new_n11054_));
  NAND2X1  g10862(.A(new_n11054_), .B(new_n11042_), .Y(new_n11055_));
  OAI21X1  g10863(.A0(new_n10558_), .A1(new_n10556_), .B0(new_n10531_), .Y(new_n11056_));
  NOR3X1   g10864(.A(new_n11056_), .B(new_n10849_), .C(new_n10515_), .Y(new_n11057_));
  AOI22X1  g10865(.A0(new_n10532_), .A1(new_n10526_), .B0(new_n10514_), .B1(\asqrt[38] ), .Y(new_n11058_));
  AOI21X1  g10866(.A0(new_n11058_), .A1(\asqrt[23] ), .B0(new_n10531_), .Y(new_n11059_));
  NOR2X1   g10867(.A(new_n11059_), .B(new_n11057_), .Y(new_n11060_));
  AOI21X1  g10868(.A0(new_n11053_), .A1(new_n11051_), .B0(new_n4493_), .Y(new_n11061_));
  NOR2X1   g10869(.A(new_n11061_), .B(\asqrt[39] ), .Y(new_n11062_));
  AOI21X1  g10870(.A0(new_n11062_), .A1(new_n11055_), .B0(new_n11060_), .Y(new_n11063_));
  OAI21X1  g10871(.A0(new_n11063_), .A1(new_n11046_), .B0(\asqrt[40] ), .Y(new_n11064_));
  AND2X1   g10872(.A(new_n10561_), .B(new_n10559_), .Y(new_n11065_));
  OR4X1    g10873(.A(new_n10849_), .B(new_n11065_), .C(new_n10539_), .D(new_n10560_), .Y(new_n11066_));
  OR2X1    g10874(.A(new_n11065_), .B(new_n10560_), .Y(new_n11067_));
  OAI21X1  g10875(.A0(new_n11067_), .A1(new_n10849_), .B0(new_n10539_), .Y(new_n11068_));
  AND2X1   g10876(.A(new_n11068_), .B(new_n11066_), .Y(new_n11069_));
  INVX1    g10877(.A(new_n11069_), .Y(new_n11070_));
  AOI21X1  g10878(.A0(new_n11054_), .A1(new_n11042_), .B0(new_n11061_), .Y(new_n11071_));
  OAI21X1  g10879(.A0(new_n11071_), .A1(new_n4165_), .B0(new_n3863_), .Y(new_n11072_));
  OAI21X1  g10880(.A0(new_n11072_), .A1(new_n11063_), .B0(new_n11070_), .Y(new_n11073_));
  AOI21X1  g10881(.A0(new_n11073_), .A1(new_n11064_), .B0(new_n3564_), .Y(new_n11074_));
  OR4X1    g10882(.A(new_n10849_), .B(new_n10577_), .C(new_n10550_), .D(new_n10544_), .Y(new_n11075_));
  NAND2X1  g10883(.A(new_n10551_), .B(new_n10563_), .Y(new_n11076_));
  OAI21X1  g10884(.A0(new_n11076_), .A1(new_n10849_), .B0(new_n10550_), .Y(new_n11077_));
  AND2X1   g10885(.A(new_n11077_), .B(new_n11075_), .Y(new_n11078_));
  INVX1    g10886(.A(new_n11078_), .Y(new_n11079_));
  NAND3X1  g10887(.A(new_n11073_), .B(new_n11064_), .C(new_n3564_), .Y(new_n11080_));
  AOI21X1  g10888(.A0(new_n11080_), .A1(new_n11079_), .B0(new_n11074_), .Y(new_n11081_));
  OR2X1    g10889(.A(new_n11081_), .B(new_n3276_), .Y(new_n11082_));
  AND2X1   g10890(.A(new_n11080_), .B(new_n11079_), .Y(new_n11083_));
  OR2X1    g10891(.A(new_n11074_), .B(\asqrt[42] ), .Y(new_n11084_));
  AND2X1   g10892(.A(new_n10593_), .B(new_n10592_), .Y(new_n11085_));
  NOR4X1   g10893(.A(new_n10849_), .B(new_n10570_), .C(new_n11085_), .D(new_n10591_), .Y(new_n11086_));
  AOI22X1  g10894(.A0(new_n10593_), .A1(new_n10592_), .B0(new_n10578_), .B1(\asqrt[41] ), .Y(new_n11087_));
  AOI21X1  g10895(.A0(new_n11087_), .A1(\asqrt[23] ), .B0(new_n10569_), .Y(new_n11088_));
  NOR2X1   g10896(.A(new_n11088_), .B(new_n11086_), .Y(new_n11089_));
  INVX1    g10897(.A(new_n11089_), .Y(new_n11090_));
  OAI21X1  g10898(.A0(new_n11084_), .A1(new_n11083_), .B0(new_n11090_), .Y(new_n11091_));
  AOI21X1  g10899(.A0(new_n11091_), .A1(new_n11082_), .B0(new_n3008_), .Y(new_n11092_));
  AND2X1   g10900(.A(new_n10579_), .B(new_n10571_), .Y(new_n11093_));
  OR4X1    g10901(.A(new_n10849_), .B(new_n11093_), .C(new_n10596_), .D(new_n10572_), .Y(new_n11094_));
  OR2X1    g10902(.A(new_n11093_), .B(new_n10572_), .Y(new_n11095_));
  OAI21X1  g10903(.A0(new_n11095_), .A1(new_n10849_), .B0(new_n10596_), .Y(new_n11096_));
  AND2X1   g10904(.A(new_n11096_), .B(new_n11094_), .Y(new_n11097_));
  OR2X1    g10905(.A(new_n11071_), .B(new_n4165_), .Y(new_n11098_));
  AND2X1   g10906(.A(new_n11054_), .B(new_n11042_), .Y(new_n11099_));
  INVX1    g10907(.A(new_n11060_), .Y(new_n11100_));
  OR2X1    g10908(.A(new_n11061_), .B(\asqrt[39] ), .Y(new_n11101_));
  OAI21X1  g10909(.A0(new_n11101_), .A1(new_n11099_), .B0(new_n11100_), .Y(new_n11102_));
  AOI21X1  g10910(.A0(new_n11102_), .A1(new_n11098_), .B0(new_n3863_), .Y(new_n11103_));
  AOI21X1  g10911(.A0(new_n11045_), .A1(\asqrt[39] ), .B0(\asqrt[40] ), .Y(new_n11104_));
  AOI21X1  g10912(.A0(new_n11104_), .A1(new_n11102_), .B0(new_n11069_), .Y(new_n11105_));
  OAI21X1  g10913(.A0(new_n11105_), .A1(new_n11103_), .B0(\asqrt[41] ), .Y(new_n11106_));
  NOR3X1   g10914(.A(new_n11105_), .B(new_n11103_), .C(\asqrt[41] ), .Y(new_n11107_));
  OAI21X1  g10915(.A0(new_n11107_), .A1(new_n11078_), .B0(new_n11106_), .Y(new_n11108_));
  AOI21X1  g10916(.A0(new_n11108_), .A1(\asqrt[42] ), .B0(\asqrt[43] ), .Y(new_n11109_));
  AOI21X1  g10917(.A0(new_n11109_), .A1(new_n11091_), .B0(new_n11097_), .Y(new_n11110_));
  OAI21X1  g10918(.A0(new_n11110_), .A1(new_n11092_), .B0(\asqrt[44] ), .Y(new_n11111_));
  NAND3X1  g10919(.A(new_n10599_), .B(new_n10586_), .C(new_n10581_), .Y(new_n11112_));
  NOR3X1   g10920(.A(new_n10849_), .B(new_n10587_), .C(new_n10614_), .Y(new_n11113_));
  OAI22X1  g10921(.A0(new_n11113_), .A1(new_n10586_), .B0(new_n11112_), .B1(new_n10849_), .Y(new_n11114_));
  INVX1    g10922(.A(new_n11114_), .Y(new_n11115_));
  NOR3X1   g10923(.A(new_n11110_), .B(new_n11092_), .C(\asqrt[44] ), .Y(new_n11116_));
  OAI21X1  g10924(.A0(new_n11116_), .A1(new_n11115_), .B0(new_n11111_), .Y(new_n11117_));
  AND2X1   g10925(.A(new_n11117_), .B(\asqrt[45] ), .Y(new_n11118_));
  AND2X1   g10926(.A(new_n11108_), .B(\asqrt[42] ), .Y(new_n11119_));
  NAND2X1  g10927(.A(new_n11080_), .B(new_n11079_), .Y(new_n11120_));
  NOR2X1   g10928(.A(new_n11074_), .B(\asqrt[42] ), .Y(new_n11121_));
  AOI21X1  g10929(.A0(new_n11121_), .A1(new_n11120_), .B0(new_n11089_), .Y(new_n11122_));
  OAI21X1  g10930(.A0(new_n11122_), .A1(new_n11119_), .B0(\asqrt[43] ), .Y(new_n11123_));
  INVX1    g10931(.A(new_n11097_), .Y(new_n11124_));
  OAI21X1  g10932(.A0(new_n11081_), .A1(new_n3276_), .B0(new_n3008_), .Y(new_n11125_));
  OAI21X1  g10933(.A0(new_n11125_), .A1(new_n11122_), .B0(new_n11124_), .Y(new_n11126_));
  NAND3X1  g10934(.A(new_n11126_), .B(new_n11123_), .C(new_n2769_), .Y(new_n11127_));
  NAND2X1  g10935(.A(new_n11127_), .B(new_n11114_), .Y(new_n11128_));
  OAI21X1  g10936(.A0(new_n10638_), .A1(new_n10636_), .B0(new_n10605_), .Y(new_n11129_));
  NOR3X1   g10937(.A(new_n11129_), .B(new_n10849_), .C(new_n10589_), .Y(new_n11130_));
  AOI22X1  g10938(.A0(new_n10606_), .A1(new_n10600_), .B0(new_n10588_), .B1(\asqrt[44] ), .Y(new_n11131_));
  AOI21X1  g10939(.A0(new_n11131_), .A1(\asqrt[23] ), .B0(new_n10605_), .Y(new_n11132_));
  NOR2X1   g10940(.A(new_n11132_), .B(new_n11130_), .Y(new_n11133_));
  AND2X1   g10941(.A(new_n11111_), .B(new_n2570_), .Y(new_n11134_));
  AOI21X1  g10942(.A0(new_n11134_), .A1(new_n11128_), .B0(new_n11133_), .Y(new_n11135_));
  OAI21X1  g10943(.A0(new_n11135_), .A1(new_n11118_), .B0(\asqrt[46] ), .Y(new_n11136_));
  AND2X1   g10944(.A(new_n10641_), .B(new_n10639_), .Y(new_n11137_));
  OR4X1    g10945(.A(new_n10849_), .B(new_n11137_), .C(new_n10613_), .D(new_n10640_), .Y(new_n11138_));
  OR2X1    g10946(.A(new_n11137_), .B(new_n10640_), .Y(new_n11139_));
  OAI21X1  g10947(.A0(new_n11139_), .A1(new_n10849_), .B0(new_n10613_), .Y(new_n11140_));
  AND2X1   g10948(.A(new_n11140_), .B(new_n11138_), .Y(new_n11141_));
  INVX1    g10949(.A(new_n11141_), .Y(new_n11142_));
  AOI21X1  g10950(.A0(new_n11126_), .A1(new_n11123_), .B0(new_n2769_), .Y(new_n11143_));
  AOI21X1  g10951(.A0(new_n11127_), .A1(new_n11114_), .B0(new_n11143_), .Y(new_n11144_));
  OAI21X1  g10952(.A0(new_n11144_), .A1(new_n2570_), .B0(new_n2263_), .Y(new_n11145_));
  OAI21X1  g10953(.A0(new_n11145_), .A1(new_n11135_), .B0(new_n11142_), .Y(new_n11146_));
  AOI21X1  g10954(.A0(new_n11146_), .A1(new_n11136_), .B0(new_n2040_), .Y(new_n11147_));
  NAND3X1  g10955(.A(new_n10625_), .B(new_n10623_), .C(new_n10643_), .Y(new_n11148_));
  NOR3X1   g10956(.A(new_n10849_), .B(new_n10651_), .C(new_n10618_), .Y(new_n11149_));
  OAI22X1  g10957(.A0(new_n11149_), .A1(new_n10623_), .B0(new_n11148_), .B1(new_n10849_), .Y(new_n11150_));
  NAND3X1  g10958(.A(new_n11146_), .B(new_n11136_), .C(new_n2040_), .Y(new_n11151_));
  AOI21X1  g10959(.A0(new_n11151_), .A1(new_n11150_), .B0(new_n11147_), .Y(new_n11152_));
  OR2X1    g10960(.A(new_n11152_), .B(new_n1834_), .Y(new_n11153_));
  AND2X1   g10961(.A(new_n11151_), .B(new_n11150_), .Y(new_n11154_));
  AND2X1   g10962(.A(new_n10667_), .B(new_n10666_), .Y(new_n11155_));
  NOR4X1   g10963(.A(new_n10849_), .B(new_n11155_), .C(new_n10634_), .D(new_n10665_), .Y(new_n11156_));
  AOI22X1  g10964(.A0(new_n10667_), .A1(new_n10666_), .B0(new_n10652_), .B1(\asqrt[47] ), .Y(new_n11157_));
  AOI21X1  g10965(.A0(new_n11157_), .A1(\asqrt[23] ), .B0(new_n10633_), .Y(new_n11158_));
  NOR2X1   g10966(.A(new_n11158_), .B(new_n11156_), .Y(new_n11159_));
  INVX1    g10967(.A(new_n11159_), .Y(new_n11160_));
  OR2X1    g10968(.A(new_n11144_), .B(new_n2570_), .Y(new_n11161_));
  AND2X1   g10969(.A(new_n11127_), .B(new_n11114_), .Y(new_n11162_));
  INVX1    g10970(.A(new_n11133_), .Y(new_n11163_));
  NAND2X1  g10971(.A(new_n11111_), .B(new_n2570_), .Y(new_n11164_));
  OAI21X1  g10972(.A0(new_n11164_), .A1(new_n11162_), .B0(new_n11163_), .Y(new_n11165_));
  AOI21X1  g10973(.A0(new_n11165_), .A1(new_n11161_), .B0(new_n2263_), .Y(new_n11166_));
  AOI21X1  g10974(.A0(new_n11117_), .A1(\asqrt[45] ), .B0(\asqrt[46] ), .Y(new_n11167_));
  AOI21X1  g10975(.A0(new_n11167_), .A1(new_n11165_), .B0(new_n11141_), .Y(new_n11168_));
  OAI21X1  g10976(.A0(new_n11168_), .A1(new_n11166_), .B0(\asqrt[47] ), .Y(new_n11169_));
  NAND2X1  g10977(.A(new_n11169_), .B(new_n1834_), .Y(new_n11170_));
  OAI21X1  g10978(.A0(new_n11170_), .A1(new_n11154_), .B0(new_n11160_), .Y(new_n11171_));
  AOI21X1  g10979(.A0(new_n11171_), .A1(new_n11153_), .B0(new_n1632_), .Y(new_n11172_));
  AND2X1   g10980(.A(new_n10653_), .B(new_n10645_), .Y(new_n11173_));
  OR4X1    g10981(.A(new_n10849_), .B(new_n11173_), .C(new_n10670_), .D(new_n10646_), .Y(new_n11174_));
  OR2X1    g10982(.A(new_n11173_), .B(new_n10646_), .Y(new_n11175_));
  OAI21X1  g10983(.A0(new_n11175_), .A1(new_n10849_), .B0(new_n10670_), .Y(new_n11176_));
  AND2X1   g10984(.A(new_n11176_), .B(new_n11174_), .Y(new_n11177_));
  INVX1    g10985(.A(new_n11150_), .Y(new_n11178_));
  NOR3X1   g10986(.A(new_n11168_), .B(new_n11166_), .C(\asqrt[47] ), .Y(new_n11179_));
  OAI21X1  g10987(.A0(new_n11179_), .A1(new_n11178_), .B0(new_n11169_), .Y(new_n11180_));
  AOI21X1  g10988(.A0(new_n11180_), .A1(\asqrt[48] ), .B0(\asqrt[49] ), .Y(new_n11181_));
  AOI21X1  g10989(.A0(new_n11181_), .A1(new_n11171_), .B0(new_n11177_), .Y(new_n11182_));
  OAI21X1  g10990(.A0(new_n11182_), .A1(new_n11172_), .B0(\asqrt[50] ), .Y(new_n11183_));
  OR4X1    g10991(.A(new_n10849_), .B(new_n10661_), .C(new_n10664_), .D(new_n10688_), .Y(new_n11184_));
  NAND2X1  g10992(.A(new_n10673_), .B(new_n10655_), .Y(new_n11185_));
  OAI21X1  g10993(.A0(new_n11185_), .A1(new_n10849_), .B0(new_n10664_), .Y(new_n11186_));
  AND2X1   g10994(.A(new_n11186_), .B(new_n11184_), .Y(new_n11187_));
  NOR3X1   g10995(.A(new_n11182_), .B(new_n11172_), .C(\asqrt[50] ), .Y(new_n11188_));
  OAI21X1  g10996(.A0(new_n11188_), .A1(new_n11187_), .B0(new_n11183_), .Y(new_n11189_));
  AND2X1   g10997(.A(new_n11189_), .B(\asqrt[51] ), .Y(new_n11190_));
  OR2X1    g10998(.A(new_n11188_), .B(new_n11187_), .Y(new_n11191_));
  OAI21X1  g10999(.A0(new_n10705_), .A1(new_n10703_), .B0(new_n10679_), .Y(new_n11192_));
  NOR3X1   g11000(.A(new_n11192_), .B(new_n10849_), .C(new_n10663_), .Y(new_n11193_));
  AOI22X1  g11001(.A0(new_n10680_), .A1(new_n10674_), .B0(new_n10662_), .B1(\asqrt[50] ), .Y(new_n11194_));
  AOI21X1  g11002(.A0(new_n11194_), .A1(\asqrt[23] ), .B0(new_n10679_), .Y(new_n11195_));
  NOR2X1   g11003(.A(new_n11195_), .B(new_n11193_), .Y(new_n11196_));
  AND2X1   g11004(.A(new_n11183_), .B(new_n1277_), .Y(new_n11197_));
  AOI21X1  g11005(.A0(new_n11197_), .A1(new_n11191_), .B0(new_n11196_), .Y(new_n11198_));
  OAI21X1  g11006(.A0(new_n11198_), .A1(new_n11190_), .B0(\asqrt[52] ), .Y(new_n11199_));
  AND2X1   g11007(.A(new_n10708_), .B(new_n10706_), .Y(new_n11200_));
  OR4X1    g11008(.A(new_n10849_), .B(new_n11200_), .C(new_n10687_), .D(new_n10707_), .Y(new_n11201_));
  OR2X1    g11009(.A(new_n11200_), .B(new_n10707_), .Y(new_n11202_));
  OAI21X1  g11010(.A0(new_n11202_), .A1(new_n10849_), .B0(new_n10687_), .Y(new_n11203_));
  AND2X1   g11011(.A(new_n11203_), .B(new_n11201_), .Y(new_n11204_));
  INVX1    g11012(.A(new_n11204_), .Y(new_n11205_));
  AND2X1   g11013(.A(new_n11180_), .B(\asqrt[48] ), .Y(new_n11206_));
  NAND2X1  g11014(.A(new_n11151_), .B(new_n11150_), .Y(new_n11207_));
  AND2X1   g11015(.A(new_n11169_), .B(new_n1834_), .Y(new_n11208_));
  AOI21X1  g11016(.A0(new_n11208_), .A1(new_n11207_), .B0(new_n11159_), .Y(new_n11209_));
  OAI21X1  g11017(.A0(new_n11209_), .A1(new_n11206_), .B0(\asqrt[49] ), .Y(new_n11210_));
  INVX1    g11018(.A(new_n11177_), .Y(new_n11211_));
  OAI21X1  g11019(.A0(new_n11152_), .A1(new_n1834_), .B0(new_n1632_), .Y(new_n11212_));
  OAI21X1  g11020(.A0(new_n11212_), .A1(new_n11209_), .B0(new_n11211_), .Y(new_n11213_));
  AOI21X1  g11021(.A0(new_n11213_), .A1(new_n11210_), .B0(new_n1469_), .Y(new_n11214_));
  INVX1    g11022(.A(new_n11187_), .Y(new_n11215_));
  NAND3X1  g11023(.A(new_n11213_), .B(new_n11210_), .C(new_n1469_), .Y(new_n11216_));
  AOI21X1  g11024(.A0(new_n11216_), .A1(new_n11215_), .B0(new_n11214_), .Y(new_n11217_));
  OAI21X1  g11025(.A0(new_n11217_), .A1(new_n1277_), .B0(new_n1111_), .Y(new_n11218_));
  OAI21X1  g11026(.A0(new_n11218_), .A1(new_n11198_), .B0(new_n11205_), .Y(new_n11219_));
  AOI21X1  g11027(.A0(new_n11219_), .A1(new_n11199_), .B0(new_n968_), .Y(new_n11220_));
  OR4X1    g11028(.A(new_n10849_), .B(new_n10710_), .C(new_n10698_), .D(new_n10692_), .Y(new_n11221_));
  OR2X1    g11029(.A(new_n10710_), .B(new_n10692_), .Y(new_n11222_));
  OAI21X1  g11030(.A0(new_n11222_), .A1(new_n10849_), .B0(new_n10698_), .Y(new_n11223_));
  AND2X1   g11031(.A(new_n11223_), .B(new_n11221_), .Y(new_n11224_));
  INVX1    g11032(.A(new_n11224_), .Y(new_n11225_));
  NAND3X1  g11033(.A(new_n11219_), .B(new_n11199_), .C(new_n968_), .Y(new_n11226_));
  AOI21X1  g11034(.A0(new_n11226_), .A1(new_n11225_), .B0(new_n11220_), .Y(new_n11227_));
  OR2X1    g11035(.A(new_n11227_), .B(new_n902_), .Y(new_n11228_));
  OR2X1    g11036(.A(new_n11217_), .B(new_n1277_), .Y(new_n11229_));
  NOR2X1   g11037(.A(new_n11188_), .B(new_n11187_), .Y(new_n11230_));
  INVX1    g11038(.A(new_n11196_), .Y(new_n11231_));
  NAND2X1  g11039(.A(new_n11183_), .B(new_n1277_), .Y(new_n11232_));
  OAI21X1  g11040(.A0(new_n11232_), .A1(new_n11230_), .B0(new_n11231_), .Y(new_n11233_));
  AOI21X1  g11041(.A0(new_n11233_), .A1(new_n11229_), .B0(new_n1111_), .Y(new_n11234_));
  AOI21X1  g11042(.A0(new_n11189_), .A1(\asqrt[51] ), .B0(\asqrt[52] ), .Y(new_n11235_));
  AOI21X1  g11043(.A0(new_n11235_), .A1(new_n11233_), .B0(new_n11204_), .Y(new_n11236_));
  NOR3X1   g11044(.A(new_n11236_), .B(new_n11234_), .C(\asqrt[53] ), .Y(new_n11237_));
  NOR2X1   g11045(.A(new_n11237_), .B(new_n11224_), .Y(new_n11238_));
  AND2X1   g11046(.A(new_n10741_), .B(new_n10740_), .Y(new_n11239_));
  NOR4X1   g11047(.A(new_n10849_), .B(new_n11239_), .C(new_n10717_), .D(new_n10739_), .Y(new_n11240_));
  AOI22X1  g11048(.A0(new_n10741_), .A1(new_n10740_), .B0(new_n10726_), .B1(\asqrt[53] ), .Y(new_n11241_));
  AOI21X1  g11049(.A0(new_n11241_), .A1(\asqrt[23] ), .B0(new_n10716_), .Y(new_n11242_));
  NOR2X1   g11050(.A(new_n11242_), .B(new_n11240_), .Y(new_n11243_));
  INVX1    g11051(.A(new_n11243_), .Y(new_n11244_));
  OAI21X1  g11052(.A0(new_n11236_), .A1(new_n11234_), .B0(\asqrt[53] ), .Y(new_n11245_));
  NAND2X1  g11053(.A(new_n11245_), .B(new_n902_), .Y(new_n11246_));
  OAI21X1  g11054(.A0(new_n11246_), .A1(new_n11238_), .B0(new_n11244_), .Y(new_n11247_));
  AOI21X1  g11055(.A0(new_n11247_), .A1(new_n11228_), .B0(new_n697_), .Y(new_n11248_));
  AND2X1   g11056(.A(new_n10727_), .B(new_n10720_), .Y(new_n11249_));
  OR4X1    g11057(.A(new_n10849_), .B(new_n11249_), .C(new_n10744_), .D(new_n10721_), .Y(new_n11250_));
  OR2X1    g11058(.A(new_n11249_), .B(new_n10721_), .Y(new_n11251_));
  OAI21X1  g11059(.A0(new_n11251_), .A1(new_n10849_), .B0(new_n10744_), .Y(new_n11252_));
  AND2X1   g11060(.A(new_n11252_), .B(new_n11250_), .Y(new_n11253_));
  OAI21X1  g11061(.A0(new_n11237_), .A1(new_n11224_), .B0(new_n11245_), .Y(new_n11254_));
  AOI21X1  g11062(.A0(new_n11254_), .A1(\asqrt[54] ), .B0(\asqrt[55] ), .Y(new_n11255_));
  AOI21X1  g11063(.A0(new_n11255_), .A1(new_n11247_), .B0(new_n11253_), .Y(new_n11256_));
  OAI21X1  g11064(.A0(new_n11256_), .A1(new_n11248_), .B0(\asqrt[56] ), .Y(new_n11257_));
  OR4X1    g11065(.A(new_n10849_), .B(new_n10735_), .C(new_n10738_), .D(new_n10762_), .Y(new_n11258_));
  OR2X1    g11066(.A(new_n10735_), .B(new_n10762_), .Y(new_n11259_));
  OAI21X1  g11067(.A0(new_n11259_), .A1(new_n10849_), .B0(new_n10738_), .Y(new_n11260_));
  AND2X1   g11068(.A(new_n11260_), .B(new_n11258_), .Y(new_n11261_));
  NOR3X1   g11069(.A(new_n11256_), .B(new_n11248_), .C(\asqrt[56] ), .Y(new_n11262_));
  OAI21X1  g11070(.A0(new_n11262_), .A1(new_n11261_), .B0(new_n11257_), .Y(new_n11263_));
  AND2X1   g11071(.A(new_n11263_), .B(\asqrt[57] ), .Y(new_n11264_));
  OR2X1    g11072(.A(new_n11262_), .B(new_n11261_), .Y(new_n11265_));
  OAI21X1  g11073(.A0(new_n10779_), .A1(new_n10777_), .B0(new_n10753_), .Y(new_n11266_));
  NOR3X1   g11074(.A(new_n11266_), .B(new_n10849_), .C(new_n10737_), .Y(new_n11267_));
  AOI22X1  g11075(.A0(new_n10754_), .A1(new_n10748_), .B0(new_n10736_), .B1(\asqrt[56] ), .Y(new_n11268_));
  AOI21X1  g11076(.A0(new_n11268_), .A1(\asqrt[23] ), .B0(new_n10753_), .Y(new_n11269_));
  NOR2X1   g11077(.A(new_n11269_), .B(new_n11267_), .Y(new_n11270_));
  AND2X1   g11078(.A(new_n11257_), .B(new_n481_), .Y(new_n11271_));
  AOI21X1  g11079(.A0(new_n11271_), .A1(new_n11265_), .B0(new_n11270_), .Y(new_n11272_));
  OAI21X1  g11080(.A0(new_n11272_), .A1(new_n11264_), .B0(\asqrt[58] ), .Y(new_n11273_));
  AND2X1   g11081(.A(new_n10782_), .B(new_n10780_), .Y(new_n11274_));
  OR4X1    g11082(.A(new_n10849_), .B(new_n11274_), .C(new_n10761_), .D(new_n10781_), .Y(new_n11275_));
  OR2X1    g11083(.A(new_n11274_), .B(new_n10781_), .Y(new_n11276_));
  OAI21X1  g11084(.A0(new_n11276_), .A1(new_n10849_), .B0(new_n10761_), .Y(new_n11277_));
  AND2X1   g11085(.A(new_n11277_), .B(new_n11275_), .Y(new_n11278_));
  INVX1    g11086(.A(new_n11278_), .Y(new_n11279_));
  AND2X1   g11087(.A(new_n11254_), .B(\asqrt[54] ), .Y(new_n11280_));
  OR2X1    g11088(.A(new_n11237_), .B(new_n11224_), .Y(new_n11281_));
  AND2X1   g11089(.A(new_n11245_), .B(new_n902_), .Y(new_n11282_));
  AOI21X1  g11090(.A0(new_n11282_), .A1(new_n11281_), .B0(new_n11243_), .Y(new_n11283_));
  OAI21X1  g11091(.A0(new_n11283_), .A1(new_n11280_), .B0(\asqrt[55] ), .Y(new_n11284_));
  INVX1    g11092(.A(new_n11253_), .Y(new_n11285_));
  OAI21X1  g11093(.A0(new_n11227_), .A1(new_n902_), .B0(new_n697_), .Y(new_n11286_));
  OAI21X1  g11094(.A0(new_n11286_), .A1(new_n11283_), .B0(new_n11285_), .Y(new_n11287_));
  AOI21X1  g11095(.A0(new_n11287_), .A1(new_n11284_), .B0(new_n582_), .Y(new_n11288_));
  INVX1    g11096(.A(new_n11261_), .Y(new_n11289_));
  NAND3X1  g11097(.A(new_n11287_), .B(new_n11284_), .C(new_n582_), .Y(new_n11290_));
  AOI21X1  g11098(.A0(new_n11290_), .A1(new_n11289_), .B0(new_n11288_), .Y(new_n11291_));
  OAI21X1  g11099(.A0(new_n11291_), .A1(new_n481_), .B0(new_n399_), .Y(new_n11292_));
  OAI21X1  g11100(.A0(new_n11292_), .A1(new_n11272_), .B0(new_n11279_), .Y(new_n11293_));
  AOI21X1  g11101(.A0(new_n11293_), .A1(new_n11273_), .B0(new_n328_), .Y(new_n11294_));
  NAND3X1  g11102(.A(new_n10773_), .B(new_n10771_), .C(new_n10792_), .Y(new_n11295_));
  NOR3X1   g11103(.A(new_n10849_), .B(new_n10784_), .C(new_n10766_), .Y(new_n11296_));
  OAI22X1  g11104(.A0(new_n11296_), .A1(new_n10771_), .B0(new_n11295_), .B1(new_n10849_), .Y(new_n11297_));
  NAND3X1  g11105(.A(new_n11293_), .B(new_n11273_), .C(new_n328_), .Y(new_n11298_));
  AOI21X1  g11106(.A0(new_n11298_), .A1(new_n11297_), .B0(new_n11294_), .Y(new_n11299_));
  OR2X1    g11107(.A(new_n11299_), .B(new_n292_), .Y(new_n11300_));
  AND2X1   g11108(.A(new_n11298_), .B(new_n11297_), .Y(new_n11301_));
  AND2X1   g11109(.A(new_n10830_), .B(new_n10829_), .Y(new_n11302_));
  NOR4X1   g11110(.A(new_n10849_), .B(new_n11302_), .C(new_n10791_), .D(new_n10828_), .Y(new_n11303_));
  AOI22X1  g11111(.A0(new_n10830_), .A1(new_n10829_), .B0(new_n10800_), .B1(\asqrt[59] ), .Y(new_n11304_));
  AOI21X1  g11112(.A0(new_n11304_), .A1(\asqrt[23] ), .B0(new_n10790_), .Y(new_n11305_));
  NOR2X1   g11113(.A(new_n11305_), .B(new_n11303_), .Y(new_n11306_));
  INVX1    g11114(.A(new_n11306_), .Y(new_n11307_));
  OR2X1    g11115(.A(new_n11291_), .B(new_n481_), .Y(new_n11308_));
  NOR2X1   g11116(.A(new_n11262_), .B(new_n11261_), .Y(new_n11309_));
  INVX1    g11117(.A(new_n11270_), .Y(new_n11310_));
  NAND2X1  g11118(.A(new_n11257_), .B(new_n481_), .Y(new_n11311_));
  OAI21X1  g11119(.A0(new_n11311_), .A1(new_n11309_), .B0(new_n11310_), .Y(new_n11312_));
  AOI21X1  g11120(.A0(new_n11312_), .A1(new_n11308_), .B0(new_n399_), .Y(new_n11313_));
  AOI21X1  g11121(.A0(new_n11263_), .A1(\asqrt[57] ), .B0(\asqrt[58] ), .Y(new_n11314_));
  AOI21X1  g11122(.A0(new_n11314_), .A1(new_n11312_), .B0(new_n11278_), .Y(new_n11315_));
  OAI21X1  g11123(.A0(new_n11315_), .A1(new_n11313_), .B0(\asqrt[59] ), .Y(new_n11316_));
  NAND2X1  g11124(.A(new_n11316_), .B(new_n292_), .Y(new_n11317_));
  OAI21X1  g11125(.A0(new_n11317_), .A1(new_n11301_), .B0(new_n11307_), .Y(new_n11318_));
  AOI21X1  g11126(.A0(new_n11318_), .A1(new_n11300_), .B0(new_n217_), .Y(new_n11319_));
  AND2X1   g11127(.A(new_n10801_), .B(new_n10794_), .Y(new_n11320_));
  OR4X1    g11128(.A(new_n10849_), .B(new_n11320_), .C(new_n10833_), .D(new_n10795_), .Y(new_n11321_));
  OR2X1    g11129(.A(new_n11320_), .B(new_n10795_), .Y(new_n11322_));
  OAI21X1  g11130(.A0(new_n11322_), .A1(new_n10849_), .B0(new_n10833_), .Y(new_n11323_));
  AND2X1   g11131(.A(new_n11323_), .B(new_n11321_), .Y(new_n11324_));
  INVX1    g11132(.A(new_n11297_), .Y(new_n11325_));
  NOR3X1   g11133(.A(new_n11315_), .B(new_n11313_), .C(\asqrt[59] ), .Y(new_n11326_));
  OAI21X1  g11134(.A0(new_n11326_), .A1(new_n11325_), .B0(new_n11316_), .Y(new_n11327_));
  AOI21X1  g11135(.A0(new_n11327_), .A1(\asqrt[60] ), .B0(\asqrt[61] ), .Y(new_n11328_));
  AOI21X1  g11136(.A0(new_n11328_), .A1(new_n11318_), .B0(new_n11324_), .Y(new_n11329_));
  OAI21X1  g11137(.A0(new_n11329_), .A1(new_n11319_), .B0(\asqrt[62] ), .Y(new_n11330_));
  OR4X1    g11138(.A(new_n10849_), .B(new_n10809_), .C(new_n10837_), .D(new_n10836_), .Y(new_n11331_));
  OR2X1    g11139(.A(new_n10809_), .B(new_n10836_), .Y(new_n11332_));
  OAI21X1  g11140(.A0(new_n11332_), .A1(new_n10849_), .B0(new_n10837_), .Y(new_n11333_));
  AND2X1   g11141(.A(new_n11333_), .B(new_n11331_), .Y(new_n11334_));
  NOR3X1   g11142(.A(new_n11329_), .B(new_n11319_), .C(\asqrt[62] ), .Y(new_n11335_));
  OAI21X1  g11143(.A0(new_n11335_), .A1(new_n11334_), .B0(new_n11330_), .Y(new_n11336_));
  AND2X1   g11144(.A(new_n10818_), .B(new_n10812_), .Y(new_n11337_));
  NOR4X1   g11145(.A(new_n10849_), .B(new_n11337_), .C(new_n10868_), .D(new_n10811_), .Y(new_n11338_));
  INVX1    g11146(.A(new_n11338_), .Y(new_n11339_));
  OAI22X1  g11147(.A0(new_n10869_), .A1(new_n10867_), .B0(new_n10839_), .B1(new_n199_), .Y(new_n11340_));
  OAI21X1  g11148(.A0(new_n11340_), .A1(new_n10849_), .B0(new_n10868_), .Y(new_n11341_));
  AND2X1   g11149(.A(new_n11341_), .B(new_n11339_), .Y(new_n11342_));
  INVX1    g11150(.A(new_n11342_), .Y(new_n11343_));
  AND2X1   g11151(.A(new_n10873_), .B(new_n10870_), .Y(new_n11344_));
  AOI21X1  g11152(.A0(new_n10870_), .A1(new_n10866_), .B0(new_n10822_), .Y(new_n11345_));
  AOI21X1  g11153(.A0(new_n11345_), .A1(\asqrt[23] ), .B0(new_n11344_), .Y(new_n11346_));
  AND2X1   g11154(.A(new_n11346_), .B(new_n11343_), .Y(new_n11347_));
  AOI21X1  g11155(.A0(new_n11347_), .A1(new_n11336_), .B0(\asqrt[63] ), .Y(new_n11348_));
  NOR2X1   g11156(.A(new_n11335_), .B(new_n11334_), .Y(new_n11349_));
  NAND2X1  g11157(.A(new_n11342_), .B(new_n11330_), .Y(new_n11350_));
  NAND2X1  g11158(.A(new_n10870_), .B(new_n10866_), .Y(new_n11351_));
  AOI21X1  g11159(.A0(\asqrt[23] ), .A1(new_n10823_), .B0(new_n11351_), .Y(new_n11352_));
  NOR3X1   g11160(.A(new_n11352_), .B(new_n11345_), .C(new_n193_), .Y(new_n11353_));
  AND2X1   g11161(.A(new_n10827_), .B(new_n193_), .Y(new_n11354_));
  INVX1    g11162(.A(new_n10846_), .Y(new_n11355_));
  OR2X1    g11163(.A(new_n11355_), .B(new_n10820_), .Y(new_n11356_));
  AOI21X1  g11164(.A0(new_n10821_), .A1(new_n10343_), .B0(new_n11356_), .Y(new_n11357_));
  NAND2X1  g11165(.A(new_n11357_), .B(new_n10843_), .Y(new_n11358_));
  NOR3X1   g11166(.A(new_n11358_), .B(new_n11344_), .C(new_n11354_), .Y(new_n11359_));
  NOR2X1   g11167(.A(new_n11359_), .B(new_n11353_), .Y(new_n11360_));
  OAI21X1  g11168(.A0(new_n11350_), .A1(new_n11349_), .B0(new_n11360_), .Y(new_n11361_));
  NOR2X1   g11169(.A(new_n11361_), .B(new_n11348_), .Y(new_n11362_));
  INVX1    g11170(.A(new_n11362_), .Y(\asqrt[22] ));
  OAI21X1  g11171(.A0(new_n11361_), .A1(new_n11348_), .B0(\a[44] ), .Y(new_n11364_));
  INVX1    g11172(.A(\a[44] ), .Y(new_n11365_));
  NOR2X1   g11173(.A(\a[43] ), .B(\a[42] ), .Y(new_n11366_));
  NAND2X1  g11174(.A(new_n11366_), .B(new_n11365_), .Y(new_n11367_));
  AOI21X1  g11175(.A0(new_n11367_), .A1(new_n11364_), .B0(new_n10849_), .Y(new_n11368_));
  AND2X1   g11176(.A(new_n11327_), .B(\asqrt[60] ), .Y(new_n11369_));
  NAND2X1  g11177(.A(new_n11298_), .B(new_n11297_), .Y(new_n11370_));
  AND2X1   g11178(.A(new_n11316_), .B(new_n292_), .Y(new_n11371_));
  AOI21X1  g11179(.A0(new_n11371_), .A1(new_n11370_), .B0(new_n11306_), .Y(new_n11372_));
  OAI21X1  g11180(.A0(new_n11372_), .A1(new_n11369_), .B0(\asqrt[61] ), .Y(new_n11373_));
  INVX1    g11181(.A(new_n11324_), .Y(new_n11374_));
  OAI21X1  g11182(.A0(new_n11299_), .A1(new_n292_), .B0(new_n217_), .Y(new_n11375_));
  OAI21X1  g11183(.A0(new_n11375_), .A1(new_n11372_), .B0(new_n11374_), .Y(new_n11376_));
  AOI21X1  g11184(.A0(new_n11376_), .A1(new_n11373_), .B0(new_n199_), .Y(new_n11377_));
  INVX1    g11185(.A(new_n11334_), .Y(new_n11378_));
  NAND3X1  g11186(.A(new_n11376_), .B(new_n11373_), .C(new_n199_), .Y(new_n11379_));
  AOI21X1  g11187(.A0(new_n11379_), .A1(new_n11378_), .B0(new_n11377_), .Y(new_n11380_));
  INVX1    g11188(.A(new_n11347_), .Y(new_n11381_));
  OAI21X1  g11189(.A0(new_n11381_), .A1(new_n11380_), .B0(new_n193_), .Y(new_n11382_));
  OR2X1    g11190(.A(new_n11335_), .B(new_n11334_), .Y(new_n11383_));
  AND2X1   g11191(.A(new_n11342_), .B(new_n11330_), .Y(new_n11384_));
  INVX1    g11192(.A(new_n11360_), .Y(new_n11385_));
  AOI21X1  g11193(.A0(new_n11384_), .A1(new_n11383_), .B0(new_n11385_), .Y(new_n11386_));
  AOI21X1  g11194(.A0(new_n11386_), .A1(new_n11382_), .B0(new_n11365_), .Y(new_n11387_));
  NAND3X1  g11195(.A(new_n11367_), .B(new_n10846_), .C(new_n10843_), .Y(new_n11388_));
  OR4X1    g11196(.A(new_n11388_), .B(new_n11387_), .C(new_n11344_), .D(new_n11354_), .Y(new_n11389_));
  OAI21X1  g11197(.A0(new_n11361_), .A1(new_n11348_), .B0(new_n11365_), .Y(new_n11390_));
  AOI21X1  g11198(.A0(new_n11386_), .A1(new_n11382_), .B0(new_n10851_), .Y(new_n11391_));
  AOI21X1  g11199(.A0(new_n11390_), .A1(\a[45] ), .B0(new_n11391_), .Y(new_n11392_));
  AOI21X1  g11200(.A0(new_n11392_), .A1(new_n11389_), .B0(new_n11368_), .Y(new_n11393_));
  OR2X1    g11201(.A(new_n11393_), .B(new_n10332_), .Y(new_n11394_));
  AND2X1   g11202(.A(new_n11392_), .B(new_n11389_), .Y(new_n11395_));
  OR2X1    g11203(.A(new_n11368_), .B(\asqrt[24] ), .Y(new_n11396_));
  OAI21X1  g11204(.A0(new_n11361_), .A1(new_n11348_), .B0(new_n10850_), .Y(new_n11397_));
  AND2X1   g11205(.A(new_n11384_), .B(new_n11383_), .Y(new_n11398_));
  OR2X1    g11206(.A(new_n11359_), .B(new_n10849_), .Y(new_n11399_));
  OR4X1    g11207(.A(new_n11399_), .B(new_n11353_), .C(new_n11398_), .D(new_n11348_), .Y(new_n11400_));
  AOI21X1  g11208(.A0(new_n11400_), .A1(new_n11397_), .B0(new_n10854_), .Y(new_n11401_));
  NOR4X1   g11209(.A(new_n11399_), .B(new_n11353_), .C(new_n11398_), .D(new_n11348_), .Y(new_n11402_));
  NOR3X1   g11210(.A(new_n11402_), .B(new_n11391_), .C(\a[46] ), .Y(new_n11403_));
  OR2X1    g11211(.A(new_n11403_), .B(new_n11401_), .Y(new_n11404_));
  OAI21X1  g11212(.A0(new_n11396_), .A1(new_n11395_), .B0(new_n11404_), .Y(new_n11405_));
  AOI21X1  g11213(.A0(new_n11405_), .A1(new_n11394_), .B0(new_n9833_), .Y(new_n11406_));
  AND2X1   g11214(.A(new_n10863_), .B(new_n10860_), .Y(new_n11407_));
  NOR3X1   g11215(.A(new_n11407_), .B(new_n10900_), .C(new_n10899_), .Y(new_n11408_));
  OAI21X1  g11216(.A0(new_n11361_), .A1(new_n11348_), .B0(new_n11408_), .Y(new_n11409_));
  AOI21X1  g11217(.A0(new_n10877_), .A1(\asqrt[24] ), .B0(new_n10900_), .Y(new_n11410_));
  OAI21X1  g11218(.A0(new_n11361_), .A1(new_n11348_), .B0(new_n11410_), .Y(new_n11411_));
  NAND2X1  g11219(.A(new_n11411_), .B(new_n11407_), .Y(new_n11412_));
  AND2X1   g11220(.A(new_n11367_), .B(new_n11364_), .Y(new_n11413_));
  NOR4X1   g11221(.A(new_n11388_), .B(new_n11387_), .C(new_n11344_), .D(new_n11354_), .Y(new_n11414_));
  INVX1    g11222(.A(\a[45] ), .Y(new_n11415_));
  AOI21X1  g11223(.A0(new_n11386_), .A1(new_n11382_), .B0(\a[44] ), .Y(new_n11416_));
  OAI21X1  g11224(.A0(new_n11416_), .A1(new_n11415_), .B0(new_n11397_), .Y(new_n11417_));
  OAI22X1  g11225(.A0(new_n11417_), .A1(new_n11414_), .B0(new_n11413_), .B1(new_n10849_), .Y(new_n11418_));
  AOI21X1  g11226(.A0(new_n11418_), .A1(\asqrt[24] ), .B0(\asqrt[25] ), .Y(new_n11419_));
  AOI22X1  g11227(.A0(new_n11419_), .A1(new_n11405_), .B0(new_n11412_), .B1(new_n11409_), .Y(new_n11420_));
  OAI21X1  g11228(.A0(new_n11420_), .A1(new_n11406_), .B0(\asqrt[26] ), .Y(new_n11421_));
  AND2X1   g11229(.A(new_n10878_), .B(new_n10864_), .Y(new_n11422_));
  NOR3X1   g11230(.A(new_n10906_), .B(new_n11422_), .C(new_n10865_), .Y(new_n11423_));
  OAI21X1  g11231(.A0(new_n11361_), .A1(new_n11348_), .B0(new_n11423_), .Y(new_n11424_));
  NOR2X1   g11232(.A(new_n11422_), .B(new_n10865_), .Y(new_n11425_));
  OAI21X1  g11233(.A0(new_n11361_), .A1(new_n11348_), .B0(new_n11425_), .Y(new_n11426_));
  NAND2X1  g11234(.A(new_n11426_), .B(new_n10906_), .Y(new_n11427_));
  AND2X1   g11235(.A(new_n11427_), .B(new_n11424_), .Y(new_n11428_));
  NOR3X1   g11236(.A(new_n11420_), .B(new_n11406_), .C(\asqrt[26] ), .Y(new_n11429_));
  OAI21X1  g11237(.A0(new_n11429_), .A1(new_n11428_), .B0(new_n11421_), .Y(new_n11430_));
  AND2X1   g11238(.A(new_n11430_), .B(\asqrt[27] ), .Y(new_n11431_));
  OR2X1    g11239(.A(new_n11429_), .B(new_n11428_), .Y(new_n11432_));
  NOR3X1   g11240(.A(new_n10895_), .B(new_n10898_), .C(new_n10915_), .Y(new_n11433_));
  NAND3X1  g11241(.A(\asqrt[22] ), .B(new_n10908_), .C(new_n10889_), .Y(new_n11434_));
  AOI22X1  g11242(.A0(new_n11434_), .A1(new_n10898_), .B0(new_n11433_), .B1(\asqrt[22] ), .Y(new_n11435_));
  AND2X1   g11243(.A(new_n11418_), .B(\asqrt[24] ), .Y(new_n11436_));
  NAND2X1  g11244(.A(new_n11392_), .B(new_n11389_), .Y(new_n11437_));
  NOR2X1   g11245(.A(new_n11368_), .B(\asqrt[24] ), .Y(new_n11438_));
  NOR2X1   g11246(.A(new_n11403_), .B(new_n11401_), .Y(new_n11439_));
  AOI21X1  g11247(.A0(new_n11438_), .A1(new_n11437_), .B0(new_n11439_), .Y(new_n11440_));
  OAI21X1  g11248(.A0(new_n11440_), .A1(new_n11436_), .B0(\asqrt[25] ), .Y(new_n11441_));
  NAND2X1  g11249(.A(new_n11412_), .B(new_n11409_), .Y(new_n11442_));
  OAI21X1  g11250(.A0(new_n11393_), .A1(new_n10332_), .B0(new_n9833_), .Y(new_n11443_));
  OAI21X1  g11251(.A0(new_n11443_), .A1(new_n11440_), .B0(new_n11442_), .Y(new_n11444_));
  AOI21X1  g11252(.A0(new_n11444_), .A1(new_n11441_), .B0(new_n9353_), .Y(new_n11445_));
  NOR2X1   g11253(.A(new_n11445_), .B(\asqrt[27] ), .Y(new_n11446_));
  AOI21X1  g11254(.A0(new_n11446_), .A1(new_n11432_), .B0(new_n11435_), .Y(new_n11447_));
  OAI21X1  g11255(.A0(new_n11447_), .A1(new_n11431_), .B0(\asqrt[28] ), .Y(new_n11448_));
  AOI21X1  g11256(.A0(new_n10916_), .A1(new_n10909_), .B0(new_n10952_), .Y(new_n11449_));
  AND2X1   g11257(.A(new_n11449_), .B(new_n10950_), .Y(new_n11450_));
  AOI22X1  g11258(.A0(new_n10916_), .A1(new_n10909_), .B0(new_n10896_), .B1(\asqrt[27] ), .Y(new_n11451_));
  AOI21X1  g11259(.A0(new_n11451_), .A1(\asqrt[22] ), .B0(new_n10914_), .Y(new_n11452_));
  AOI21X1  g11260(.A0(new_n11450_), .A1(\asqrt[22] ), .B0(new_n11452_), .Y(new_n11453_));
  INVX1    g11261(.A(new_n11453_), .Y(new_n11454_));
  INVX1    g11262(.A(new_n11428_), .Y(new_n11455_));
  NAND3X1  g11263(.A(new_n11444_), .B(new_n11441_), .C(new_n9353_), .Y(new_n11456_));
  AOI21X1  g11264(.A0(new_n11456_), .A1(new_n11455_), .B0(new_n11445_), .Y(new_n11457_));
  OAI21X1  g11265(.A0(new_n11457_), .A1(new_n8874_), .B0(new_n8412_), .Y(new_n11458_));
  OAI21X1  g11266(.A0(new_n11458_), .A1(new_n11447_), .B0(new_n11454_), .Y(new_n11459_));
  AOI21X1  g11267(.A0(new_n11459_), .A1(new_n11448_), .B0(new_n7970_), .Y(new_n11460_));
  AND2X1   g11268(.A(new_n10956_), .B(new_n10954_), .Y(new_n11461_));
  NOR3X1   g11269(.A(new_n11461_), .B(new_n10924_), .C(new_n10955_), .Y(new_n11462_));
  NOR3X1   g11270(.A(new_n11362_), .B(new_n11461_), .C(new_n10955_), .Y(new_n11463_));
  NOR2X1   g11271(.A(new_n11463_), .B(new_n10923_), .Y(new_n11464_));
  AOI21X1  g11272(.A0(new_n11462_), .A1(\asqrt[22] ), .B0(new_n11464_), .Y(new_n11465_));
  INVX1    g11273(.A(new_n11465_), .Y(new_n11466_));
  NAND3X1  g11274(.A(new_n11459_), .B(new_n11448_), .C(new_n7970_), .Y(new_n11467_));
  AOI21X1  g11275(.A0(new_n11467_), .A1(new_n11466_), .B0(new_n11460_), .Y(new_n11468_));
  OR2X1    g11276(.A(new_n11468_), .B(new_n7527_), .Y(new_n11469_));
  OR2X1    g11277(.A(new_n11457_), .B(new_n8874_), .Y(new_n11470_));
  NOR2X1   g11278(.A(new_n11429_), .B(new_n11428_), .Y(new_n11471_));
  INVX1    g11279(.A(new_n11435_), .Y(new_n11472_));
  OR2X1    g11280(.A(new_n11445_), .B(\asqrt[27] ), .Y(new_n11473_));
  OAI21X1  g11281(.A0(new_n11473_), .A1(new_n11471_), .B0(new_n11472_), .Y(new_n11474_));
  AOI21X1  g11282(.A0(new_n11474_), .A1(new_n11470_), .B0(new_n8412_), .Y(new_n11475_));
  AOI21X1  g11283(.A0(new_n11430_), .A1(\asqrt[27] ), .B0(\asqrt[28] ), .Y(new_n11476_));
  AOI21X1  g11284(.A0(new_n11476_), .A1(new_n11474_), .B0(new_n11453_), .Y(new_n11477_));
  NOR3X1   g11285(.A(new_n11477_), .B(new_n11475_), .C(\asqrt[29] ), .Y(new_n11478_));
  NOR2X1   g11286(.A(new_n11478_), .B(new_n11465_), .Y(new_n11479_));
  OR4X1    g11287(.A(new_n11362_), .B(new_n10960_), .C(new_n10931_), .D(new_n10928_), .Y(new_n11480_));
  NAND2X1  g11288(.A(new_n10932_), .B(new_n10958_), .Y(new_n11481_));
  OAI21X1  g11289(.A0(new_n11481_), .A1(new_n11362_), .B0(new_n10931_), .Y(new_n11482_));
  AND2X1   g11290(.A(new_n11482_), .B(new_n11480_), .Y(new_n11483_));
  INVX1    g11291(.A(new_n11483_), .Y(new_n11484_));
  OAI21X1  g11292(.A0(new_n11477_), .A1(new_n11475_), .B0(\asqrt[29] ), .Y(new_n11485_));
  NAND2X1  g11293(.A(new_n11485_), .B(new_n7527_), .Y(new_n11486_));
  OAI21X1  g11294(.A0(new_n11486_), .A1(new_n11479_), .B0(new_n11484_), .Y(new_n11487_));
  AOI21X1  g11295(.A0(new_n11487_), .A1(new_n11469_), .B0(new_n7103_), .Y(new_n11488_));
  AND2X1   g11296(.A(new_n10975_), .B(new_n10974_), .Y(new_n11489_));
  NOR3X1   g11297(.A(new_n11489_), .B(new_n10941_), .C(new_n10973_), .Y(new_n11490_));
  NOR3X1   g11298(.A(new_n11362_), .B(new_n11489_), .C(new_n10973_), .Y(new_n11491_));
  NOR2X1   g11299(.A(new_n11491_), .B(new_n10940_), .Y(new_n11492_));
  AOI21X1  g11300(.A0(new_n11490_), .A1(\asqrt[22] ), .B0(new_n11492_), .Y(new_n11493_));
  OAI21X1  g11301(.A0(new_n11478_), .A1(new_n11465_), .B0(new_n11485_), .Y(new_n11494_));
  AOI21X1  g11302(.A0(new_n11494_), .A1(\asqrt[30] ), .B0(\asqrt[31] ), .Y(new_n11495_));
  AOI21X1  g11303(.A0(new_n11495_), .A1(new_n11487_), .B0(new_n11493_), .Y(new_n11496_));
  OAI21X1  g11304(.A0(new_n11496_), .A1(new_n11488_), .B0(\asqrt[32] ), .Y(new_n11497_));
  AND2X1   g11305(.A(new_n10962_), .B(new_n10943_), .Y(new_n11498_));
  NOR3X1   g11306(.A(new_n11498_), .B(new_n10978_), .C(new_n10944_), .Y(new_n11499_));
  NOR3X1   g11307(.A(new_n11362_), .B(new_n11498_), .C(new_n10944_), .Y(new_n11500_));
  NOR2X1   g11308(.A(new_n11500_), .B(new_n10949_), .Y(new_n11501_));
  AOI21X1  g11309(.A0(new_n11499_), .A1(\asqrt[22] ), .B0(new_n11501_), .Y(new_n11502_));
  NOR3X1   g11310(.A(new_n11496_), .B(new_n11488_), .C(\asqrt[32] ), .Y(new_n11503_));
  OAI21X1  g11311(.A0(new_n11503_), .A1(new_n11502_), .B0(new_n11497_), .Y(new_n11504_));
  AND2X1   g11312(.A(new_n11504_), .B(\asqrt[33] ), .Y(new_n11505_));
  INVX1    g11313(.A(new_n11502_), .Y(new_n11506_));
  AND2X1   g11314(.A(new_n11494_), .B(\asqrt[30] ), .Y(new_n11507_));
  OR2X1    g11315(.A(new_n11478_), .B(new_n11465_), .Y(new_n11508_));
  AND2X1   g11316(.A(new_n11485_), .B(new_n7527_), .Y(new_n11509_));
  AOI21X1  g11317(.A0(new_n11509_), .A1(new_n11508_), .B0(new_n11483_), .Y(new_n11510_));
  OAI21X1  g11318(.A0(new_n11510_), .A1(new_n11507_), .B0(\asqrt[31] ), .Y(new_n11511_));
  INVX1    g11319(.A(new_n11493_), .Y(new_n11512_));
  OAI21X1  g11320(.A0(new_n11468_), .A1(new_n7527_), .B0(new_n7103_), .Y(new_n11513_));
  OAI21X1  g11321(.A0(new_n11513_), .A1(new_n11510_), .B0(new_n11512_), .Y(new_n11514_));
  NAND3X1  g11322(.A(new_n11514_), .B(new_n11511_), .C(new_n6699_), .Y(new_n11515_));
  NAND2X1  g11323(.A(new_n11515_), .B(new_n11506_), .Y(new_n11516_));
  NAND4X1  g11324(.A(\asqrt[22] ), .B(new_n10981_), .C(new_n10968_), .D(new_n10964_), .Y(new_n11517_));
  NAND2X1  g11325(.A(new_n10981_), .B(new_n10964_), .Y(new_n11518_));
  OAI21X1  g11326(.A0(new_n11518_), .A1(new_n11362_), .B0(new_n10972_), .Y(new_n11519_));
  AND2X1   g11327(.A(new_n11519_), .B(new_n11517_), .Y(new_n11520_));
  AOI21X1  g11328(.A0(new_n11514_), .A1(new_n11511_), .B0(new_n6699_), .Y(new_n11521_));
  NOR2X1   g11329(.A(new_n11521_), .B(\asqrt[33] ), .Y(new_n11522_));
  AOI21X1  g11330(.A0(new_n11522_), .A1(new_n11516_), .B0(new_n11520_), .Y(new_n11523_));
  OAI21X1  g11331(.A0(new_n11523_), .A1(new_n11505_), .B0(\asqrt[34] ), .Y(new_n11524_));
  AOI21X1  g11332(.A0(new_n10989_), .A1(new_n10982_), .B0(new_n11028_), .Y(new_n11525_));
  AND2X1   g11333(.A(new_n11525_), .B(new_n11026_), .Y(new_n11526_));
  AOI22X1  g11334(.A0(new_n10989_), .A1(new_n10982_), .B0(new_n10970_), .B1(\asqrt[33] ), .Y(new_n11527_));
  AOI21X1  g11335(.A0(new_n11527_), .A1(\asqrt[22] ), .B0(new_n10987_), .Y(new_n11528_));
  AOI21X1  g11336(.A0(new_n11526_), .A1(\asqrt[22] ), .B0(new_n11528_), .Y(new_n11529_));
  INVX1    g11337(.A(new_n11529_), .Y(new_n11530_));
  AOI21X1  g11338(.A0(new_n11515_), .A1(new_n11506_), .B0(new_n11521_), .Y(new_n11531_));
  OAI21X1  g11339(.A0(new_n11531_), .A1(new_n6294_), .B0(new_n5941_), .Y(new_n11532_));
  OAI21X1  g11340(.A0(new_n11532_), .A1(new_n11523_), .B0(new_n11530_), .Y(new_n11533_));
  AOI21X1  g11341(.A0(new_n11533_), .A1(new_n11524_), .B0(new_n5541_), .Y(new_n11534_));
  AND2X1   g11342(.A(new_n11032_), .B(new_n11030_), .Y(new_n11535_));
  NOR3X1   g11343(.A(new_n11535_), .B(new_n10997_), .C(new_n11031_), .Y(new_n11536_));
  NOR3X1   g11344(.A(new_n11362_), .B(new_n11535_), .C(new_n11031_), .Y(new_n11537_));
  NOR2X1   g11345(.A(new_n11537_), .B(new_n10996_), .Y(new_n11538_));
  AOI21X1  g11346(.A0(new_n11536_), .A1(\asqrt[22] ), .B0(new_n11538_), .Y(new_n11539_));
  INVX1    g11347(.A(new_n11539_), .Y(new_n11540_));
  NAND3X1  g11348(.A(new_n11533_), .B(new_n11524_), .C(new_n5541_), .Y(new_n11541_));
  AOI21X1  g11349(.A0(new_n11541_), .A1(new_n11540_), .B0(new_n11534_), .Y(new_n11542_));
  OR2X1    g11350(.A(new_n11542_), .B(new_n5176_), .Y(new_n11543_));
  AND2X1   g11351(.A(new_n11541_), .B(new_n11540_), .Y(new_n11544_));
  OR4X1    g11352(.A(new_n11362_), .B(new_n11035_), .C(new_n11006_), .D(new_n11001_), .Y(new_n11545_));
  NAND2X1  g11353(.A(new_n11007_), .B(new_n11034_), .Y(new_n11546_));
  OAI21X1  g11354(.A0(new_n11546_), .A1(new_n11362_), .B0(new_n11006_), .Y(new_n11547_));
  AND2X1   g11355(.A(new_n11547_), .B(new_n11545_), .Y(new_n11548_));
  INVX1    g11356(.A(new_n11548_), .Y(new_n11549_));
  OR2X1    g11357(.A(new_n11534_), .B(\asqrt[36] ), .Y(new_n11550_));
  OAI21X1  g11358(.A0(new_n11550_), .A1(new_n11544_), .B0(new_n11549_), .Y(new_n11551_));
  AOI21X1  g11359(.A0(new_n11551_), .A1(new_n11543_), .B0(new_n4826_), .Y(new_n11552_));
  AND2X1   g11360(.A(new_n11049_), .B(new_n11048_), .Y(new_n11553_));
  NOR3X1   g11361(.A(new_n11553_), .B(new_n11016_), .C(new_n11047_), .Y(new_n11554_));
  NOR3X1   g11362(.A(new_n11362_), .B(new_n11553_), .C(new_n11047_), .Y(new_n11555_));
  NOR2X1   g11363(.A(new_n11555_), .B(new_n11015_), .Y(new_n11556_));
  AOI21X1  g11364(.A0(new_n11554_), .A1(\asqrt[22] ), .B0(new_n11556_), .Y(new_n11557_));
  OR2X1    g11365(.A(new_n11531_), .B(new_n6294_), .Y(new_n11558_));
  AND2X1   g11366(.A(new_n11515_), .B(new_n11506_), .Y(new_n11559_));
  INVX1    g11367(.A(new_n11520_), .Y(new_n11560_));
  OR2X1    g11368(.A(new_n11521_), .B(\asqrt[33] ), .Y(new_n11561_));
  OAI21X1  g11369(.A0(new_n11561_), .A1(new_n11559_), .B0(new_n11560_), .Y(new_n11562_));
  AOI21X1  g11370(.A0(new_n11562_), .A1(new_n11558_), .B0(new_n5941_), .Y(new_n11563_));
  AOI21X1  g11371(.A0(new_n11504_), .A1(\asqrt[33] ), .B0(\asqrt[34] ), .Y(new_n11564_));
  AOI21X1  g11372(.A0(new_n11564_), .A1(new_n11562_), .B0(new_n11529_), .Y(new_n11565_));
  OAI21X1  g11373(.A0(new_n11565_), .A1(new_n11563_), .B0(\asqrt[35] ), .Y(new_n11566_));
  NOR3X1   g11374(.A(new_n11565_), .B(new_n11563_), .C(\asqrt[35] ), .Y(new_n11567_));
  OAI21X1  g11375(.A0(new_n11567_), .A1(new_n11539_), .B0(new_n11566_), .Y(new_n11568_));
  AOI21X1  g11376(.A0(new_n11568_), .A1(\asqrt[36] ), .B0(\asqrt[37] ), .Y(new_n11569_));
  AOI21X1  g11377(.A0(new_n11569_), .A1(new_n11551_), .B0(new_n11557_), .Y(new_n11570_));
  OAI21X1  g11378(.A0(new_n11570_), .A1(new_n11552_), .B0(\asqrt[38] ), .Y(new_n11571_));
  AND2X1   g11379(.A(new_n11037_), .B(new_n11018_), .Y(new_n11572_));
  NOR3X1   g11380(.A(new_n11572_), .B(new_n11024_), .C(new_n11019_), .Y(new_n11573_));
  NOR3X1   g11381(.A(new_n11362_), .B(new_n11572_), .C(new_n11019_), .Y(new_n11574_));
  NOR2X1   g11382(.A(new_n11574_), .B(new_n11025_), .Y(new_n11575_));
  AOI21X1  g11383(.A0(new_n11573_), .A1(\asqrt[22] ), .B0(new_n11575_), .Y(new_n11576_));
  NOR3X1   g11384(.A(new_n11570_), .B(new_n11552_), .C(\asqrt[38] ), .Y(new_n11577_));
  OAI21X1  g11385(.A0(new_n11577_), .A1(new_n11576_), .B0(new_n11571_), .Y(new_n11578_));
  AND2X1   g11386(.A(new_n11578_), .B(\asqrt[39] ), .Y(new_n11579_));
  OR2X1    g11387(.A(new_n11577_), .B(new_n11576_), .Y(new_n11580_));
  OR4X1    g11388(.A(new_n11362_), .B(new_n11044_), .C(new_n11042_), .D(new_n11061_), .Y(new_n11581_));
  NAND2X1  g11389(.A(new_n11054_), .B(new_n11039_), .Y(new_n11582_));
  OAI21X1  g11390(.A0(new_n11582_), .A1(new_n11362_), .B0(new_n11042_), .Y(new_n11583_));
  AND2X1   g11391(.A(new_n11583_), .B(new_n11581_), .Y(new_n11584_));
  AND2X1   g11392(.A(new_n11568_), .B(\asqrt[36] ), .Y(new_n11585_));
  NAND2X1  g11393(.A(new_n11541_), .B(new_n11540_), .Y(new_n11586_));
  NOR2X1   g11394(.A(new_n11534_), .B(\asqrt[36] ), .Y(new_n11587_));
  AOI21X1  g11395(.A0(new_n11587_), .A1(new_n11586_), .B0(new_n11548_), .Y(new_n11588_));
  OAI21X1  g11396(.A0(new_n11588_), .A1(new_n11585_), .B0(\asqrt[37] ), .Y(new_n11589_));
  INVX1    g11397(.A(new_n11557_), .Y(new_n11590_));
  OAI21X1  g11398(.A0(new_n11542_), .A1(new_n5176_), .B0(new_n4826_), .Y(new_n11591_));
  OAI21X1  g11399(.A0(new_n11591_), .A1(new_n11588_), .B0(new_n11590_), .Y(new_n11592_));
  AOI21X1  g11400(.A0(new_n11592_), .A1(new_n11589_), .B0(new_n4493_), .Y(new_n11593_));
  NOR2X1   g11401(.A(new_n11593_), .B(\asqrt[39] ), .Y(new_n11594_));
  AOI21X1  g11402(.A0(new_n11594_), .A1(new_n11580_), .B0(new_n11584_), .Y(new_n11595_));
  OAI21X1  g11403(.A0(new_n11595_), .A1(new_n11579_), .B0(\asqrt[40] ), .Y(new_n11596_));
  AOI21X1  g11404(.A0(new_n11062_), .A1(new_n11055_), .B0(new_n11100_), .Y(new_n11597_));
  AND2X1   g11405(.A(new_n11597_), .B(new_n11098_), .Y(new_n11598_));
  AOI22X1  g11406(.A0(new_n11062_), .A1(new_n11055_), .B0(new_n11045_), .B1(\asqrt[39] ), .Y(new_n11599_));
  AOI21X1  g11407(.A0(new_n11599_), .A1(\asqrt[22] ), .B0(new_n11060_), .Y(new_n11600_));
  AOI21X1  g11408(.A0(new_n11598_), .A1(\asqrt[22] ), .B0(new_n11600_), .Y(new_n11601_));
  INVX1    g11409(.A(new_n11601_), .Y(new_n11602_));
  INVX1    g11410(.A(new_n11576_), .Y(new_n11603_));
  NAND3X1  g11411(.A(new_n11592_), .B(new_n11589_), .C(new_n4493_), .Y(new_n11604_));
  AOI21X1  g11412(.A0(new_n11604_), .A1(new_n11603_), .B0(new_n11593_), .Y(new_n11605_));
  OAI21X1  g11413(.A0(new_n11605_), .A1(new_n4165_), .B0(new_n3863_), .Y(new_n11606_));
  OAI21X1  g11414(.A0(new_n11606_), .A1(new_n11595_), .B0(new_n11602_), .Y(new_n11607_));
  AOI21X1  g11415(.A0(new_n11607_), .A1(new_n11596_), .B0(new_n3564_), .Y(new_n11608_));
  AND2X1   g11416(.A(new_n11104_), .B(new_n11102_), .Y(new_n11609_));
  NOR3X1   g11417(.A(new_n11609_), .B(new_n11070_), .C(new_n11103_), .Y(new_n11610_));
  NOR3X1   g11418(.A(new_n11362_), .B(new_n11609_), .C(new_n11103_), .Y(new_n11611_));
  NOR2X1   g11419(.A(new_n11611_), .B(new_n11069_), .Y(new_n11612_));
  AOI21X1  g11420(.A0(new_n11610_), .A1(\asqrt[22] ), .B0(new_n11612_), .Y(new_n11613_));
  INVX1    g11421(.A(new_n11613_), .Y(new_n11614_));
  NAND3X1  g11422(.A(new_n11607_), .B(new_n11596_), .C(new_n3564_), .Y(new_n11615_));
  AOI21X1  g11423(.A0(new_n11615_), .A1(new_n11614_), .B0(new_n11608_), .Y(new_n11616_));
  OR2X1    g11424(.A(new_n11616_), .B(new_n3276_), .Y(new_n11617_));
  AND2X1   g11425(.A(new_n11615_), .B(new_n11614_), .Y(new_n11618_));
  NAND4X1  g11426(.A(\asqrt[22] ), .B(new_n11080_), .C(new_n11078_), .D(new_n11106_), .Y(new_n11619_));
  NAND2X1  g11427(.A(new_n11080_), .B(new_n11106_), .Y(new_n11620_));
  OAI21X1  g11428(.A0(new_n11620_), .A1(new_n11362_), .B0(new_n11079_), .Y(new_n11621_));
  AND2X1   g11429(.A(new_n11621_), .B(new_n11619_), .Y(new_n11622_));
  INVX1    g11430(.A(new_n11622_), .Y(new_n11623_));
  OR2X1    g11431(.A(new_n11608_), .B(\asqrt[42] ), .Y(new_n11624_));
  OAI21X1  g11432(.A0(new_n11624_), .A1(new_n11618_), .B0(new_n11623_), .Y(new_n11625_));
  AOI21X1  g11433(.A0(new_n11625_), .A1(new_n11617_), .B0(new_n3008_), .Y(new_n11626_));
  OR2X1    g11434(.A(new_n11605_), .B(new_n4165_), .Y(new_n11627_));
  NOR2X1   g11435(.A(new_n11577_), .B(new_n11576_), .Y(new_n11628_));
  INVX1    g11436(.A(new_n11584_), .Y(new_n11629_));
  OR2X1    g11437(.A(new_n11593_), .B(\asqrt[39] ), .Y(new_n11630_));
  OAI21X1  g11438(.A0(new_n11630_), .A1(new_n11628_), .B0(new_n11629_), .Y(new_n11631_));
  AOI21X1  g11439(.A0(new_n11631_), .A1(new_n11627_), .B0(new_n3863_), .Y(new_n11632_));
  AOI21X1  g11440(.A0(new_n11578_), .A1(\asqrt[39] ), .B0(\asqrt[40] ), .Y(new_n11633_));
  AOI21X1  g11441(.A0(new_n11633_), .A1(new_n11631_), .B0(new_n11601_), .Y(new_n11634_));
  OAI21X1  g11442(.A0(new_n11634_), .A1(new_n11632_), .B0(\asqrt[41] ), .Y(new_n11635_));
  NOR3X1   g11443(.A(new_n11634_), .B(new_n11632_), .C(\asqrt[41] ), .Y(new_n11636_));
  OAI21X1  g11444(.A0(new_n11636_), .A1(new_n11613_), .B0(new_n11635_), .Y(new_n11637_));
  AOI21X1  g11445(.A0(new_n11637_), .A1(\asqrt[42] ), .B0(\asqrt[43] ), .Y(new_n11638_));
  AND2X1   g11446(.A(new_n11121_), .B(new_n11120_), .Y(new_n11639_));
  NOR3X1   g11447(.A(new_n11090_), .B(new_n11639_), .C(new_n11119_), .Y(new_n11640_));
  NOR3X1   g11448(.A(new_n11362_), .B(new_n11639_), .C(new_n11119_), .Y(new_n11641_));
  NOR2X1   g11449(.A(new_n11641_), .B(new_n11089_), .Y(new_n11642_));
  AOI21X1  g11450(.A0(new_n11640_), .A1(\asqrt[22] ), .B0(new_n11642_), .Y(new_n11643_));
  AOI21X1  g11451(.A0(new_n11638_), .A1(new_n11625_), .B0(new_n11643_), .Y(new_n11644_));
  OAI21X1  g11452(.A0(new_n11644_), .A1(new_n11626_), .B0(\asqrt[44] ), .Y(new_n11645_));
  AND2X1   g11453(.A(new_n11109_), .B(new_n11091_), .Y(new_n11646_));
  NOR3X1   g11454(.A(new_n11646_), .B(new_n11124_), .C(new_n11092_), .Y(new_n11647_));
  NOR3X1   g11455(.A(new_n11362_), .B(new_n11646_), .C(new_n11092_), .Y(new_n11648_));
  NOR2X1   g11456(.A(new_n11648_), .B(new_n11097_), .Y(new_n11649_));
  AOI21X1  g11457(.A0(new_n11647_), .A1(\asqrt[22] ), .B0(new_n11649_), .Y(new_n11650_));
  NOR3X1   g11458(.A(new_n11644_), .B(new_n11626_), .C(\asqrt[44] ), .Y(new_n11651_));
  OAI21X1  g11459(.A0(new_n11651_), .A1(new_n11650_), .B0(new_n11645_), .Y(new_n11652_));
  AND2X1   g11460(.A(new_n11652_), .B(\asqrt[45] ), .Y(new_n11653_));
  OR2X1    g11461(.A(new_n11651_), .B(new_n11650_), .Y(new_n11654_));
  OR4X1    g11462(.A(new_n11362_), .B(new_n11116_), .C(new_n11114_), .D(new_n11143_), .Y(new_n11655_));
  OR2X1    g11463(.A(new_n11116_), .B(new_n11143_), .Y(new_n11656_));
  OAI21X1  g11464(.A0(new_n11656_), .A1(new_n11362_), .B0(new_n11114_), .Y(new_n11657_));
  AND2X1   g11465(.A(new_n11657_), .B(new_n11655_), .Y(new_n11658_));
  AND2X1   g11466(.A(new_n11645_), .B(new_n2570_), .Y(new_n11659_));
  AOI21X1  g11467(.A0(new_n11659_), .A1(new_n11654_), .B0(new_n11658_), .Y(new_n11660_));
  OAI21X1  g11468(.A0(new_n11660_), .A1(new_n11653_), .B0(\asqrt[46] ), .Y(new_n11661_));
  AOI21X1  g11469(.A0(new_n11134_), .A1(new_n11128_), .B0(new_n11163_), .Y(new_n11662_));
  AND2X1   g11470(.A(new_n11662_), .B(new_n11161_), .Y(new_n11663_));
  AOI22X1  g11471(.A0(new_n11134_), .A1(new_n11128_), .B0(new_n11117_), .B1(\asqrt[45] ), .Y(new_n11664_));
  AOI21X1  g11472(.A0(new_n11664_), .A1(\asqrt[22] ), .B0(new_n11133_), .Y(new_n11665_));
  AOI21X1  g11473(.A0(new_n11663_), .A1(\asqrt[22] ), .B0(new_n11665_), .Y(new_n11666_));
  INVX1    g11474(.A(new_n11666_), .Y(new_n11667_));
  AND2X1   g11475(.A(new_n11637_), .B(\asqrt[42] ), .Y(new_n11668_));
  NAND2X1  g11476(.A(new_n11615_), .B(new_n11614_), .Y(new_n11669_));
  NOR2X1   g11477(.A(new_n11608_), .B(\asqrt[42] ), .Y(new_n11670_));
  AOI21X1  g11478(.A0(new_n11670_), .A1(new_n11669_), .B0(new_n11622_), .Y(new_n11671_));
  OAI21X1  g11479(.A0(new_n11671_), .A1(new_n11668_), .B0(\asqrt[43] ), .Y(new_n11672_));
  OAI21X1  g11480(.A0(new_n11616_), .A1(new_n3276_), .B0(new_n3008_), .Y(new_n11673_));
  INVX1    g11481(.A(new_n11643_), .Y(new_n11674_));
  OAI21X1  g11482(.A0(new_n11673_), .A1(new_n11671_), .B0(new_n11674_), .Y(new_n11675_));
  AOI21X1  g11483(.A0(new_n11675_), .A1(new_n11672_), .B0(new_n2769_), .Y(new_n11676_));
  INVX1    g11484(.A(new_n11650_), .Y(new_n11677_));
  NAND3X1  g11485(.A(new_n11675_), .B(new_n11672_), .C(new_n2769_), .Y(new_n11678_));
  AOI21X1  g11486(.A0(new_n11678_), .A1(new_n11677_), .B0(new_n11676_), .Y(new_n11679_));
  OAI21X1  g11487(.A0(new_n11679_), .A1(new_n2570_), .B0(new_n2263_), .Y(new_n11680_));
  OAI21X1  g11488(.A0(new_n11680_), .A1(new_n11660_), .B0(new_n11667_), .Y(new_n11681_));
  AOI21X1  g11489(.A0(new_n11681_), .A1(new_n11661_), .B0(new_n2040_), .Y(new_n11682_));
  AND2X1   g11490(.A(new_n11167_), .B(new_n11165_), .Y(new_n11683_));
  NOR3X1   g11491(.A(new_n11683_), .B(new_n11142_), .C(new_n11166_), .Y(new_n11684_));
  NOR3X1   g11492(.A(new_n11362_), .B(new_n11683_), .C(new_n11166_), .Y(new_n11685_));
  NOR2X1   g11493(.A(new_n11685_), .B(new_n11141_), .Y(new_n11686_));
  AOI21X1  g11494(.A0(new_n11684_), .A1(\asqrt[22] ), .B0(new_n11686_), .Y(new_n11687_));
  INVX1    g11495(.A(new_n11687_), .Y(new_n11688_));
  NAND3X1  g11496(.A(new_n11681_), .B(new_n11661_), .C(new_n2040_), .Y(new_n11689_));
  AOI21X1  g11497(.A0(new_n11689_), .A1(new_n11688_), .B0(new_n11682_), .Y(new_n11690_));
  OR2X1    g11498(.A(new_n11690_), .B(new_n1834_), .Y(new_n11691_));
  OR2X1    g11499(.A(new_n11679_), .B(new_n2570_), .Y(new_n11692_));
  NOR2X1   g11500(.A(new_n11651_), .B(new_n11650_), .Y(new_n11693_));
  INVX1    g11501(.A(new_n11658_), .Y(new_n11694_));
  NAND2X1  g11502(.A(new_n11645_), .B(new_n2570_), .Y(new_n11695_));
  OAI21X1  g11503(.A0(new_n11695_), .A1(new_n11693_), .B0(new_n11694_), .Y(new_n11696_));
  AOI21X1  g11504(.A0(new_n11696_), .A1(new_n11692_), .B0(new_n2263_), .Y(new_n11697_));
  AOI21X1  g11505(.A0(new_n11652_), .A1(\asqrt[45] ), .B0(\asqrt[46] ), .Y(new_n11698_));
  AOI21X1  g11506(.A0(new_n11698_), .A1(new_n11696_), .B0(new_n11666_), .Y(new_n11699_));
  NOR3X1   g11507(.A(new_n11699_), .B(new_n11697_), .C(\asqrt[47] ), .Y(new_n11700_));
  NOR2X1   g11508(.A(new_n11700_), .B(new_n11687_), .Y(new_n11701_));
  OR4X1    g11509(.A(new_n11362_), .B(new_n11179_), .C(new_n11150_), .D(new_n11147_), .Y(new_n11702_));
  OR2X1    g11510(.A(new_n11179_), .B(new_n11147_), .Y(new_n11703_));
  OAI21X1  g11511(.A0(new_n11703_), .A1(new_n11362_), .B0(new_n11150_), .Y(new_n11704_));
  AND2X1   g11512(.A(new_n11704_), .B(new_n11702_), .Y(new_n11705_));
  INVX1    g11513(.A(new_n11705_), .Y(new_n11706_));
  OAI21X1  g11514(.A0(new_n11699_), .A1(new_n11697_), .B0(\asqrt[47] ), .Y(new_n11707_));
  NAND2X1  g11515(.A(new_n11707_), .B(new_n1834_), .Y(new_n11708_));
  OAI21X1  g11516(.A0(new_n11708_), .A1(new_n11701_), .B0(new_n11706_), .Y(new_n11709_));
  AOI21X1  g11517(.A0(new_n11709_), .A1(new_n11691_), .B0(new_n1632_), .Y(new_n11710_));
  AND2X1   g11518(.A(new_n11208_), .B(new_n11207_), .Y(new_n11711_));
  NOR3X1   g11519(.A(new_n11711_), .B(new_n11160_), .C(new_n11206_), .Y(new_n11712_));
  NOR3X1   g11520(.A(new_n11362_), .B(new_n11711_), .C(new_n11206_), .Y(new_n11713_));
  NOR2X1   g11521(.A(new_n11713_), .B(new_n11159_), .Y(new_n11714_));
  AOI21X1  g11522(.A0(new_n11712_), .A1(\asqrt[22] ), .B0(new_n11714_), .Y(new_n11715_));
  OAI21X1  g11523(.A0(new_n11700_), .A1(new_n11687_), .B0(new_n11707_), .Y(new_n11716_));
  AOI21X1  g11524(.A0(new_n11716_), .A1(\asqrt[48] ), .B0(\asqrt[49] ), .Y(new_n11717_));
  AOI21X1  g11525(.A0(new_n11717_), .A1(new_n11709_), .B0(new_n11715_), .Y(new_n11718_));
  OAI21X1  g11526(.A0(new_n11718_), .A1(new_n11710_), .B0(\asqrt[50] ), .Y(new_n11719_));
  AND2X1   g11527(.A(new_n11181_), .B(new_n11171_), .Y(new_n11720_));
  NOR3X1   g11528(.A(new_n11720_), .B(new_n11211_), .C(new_n11172_), .Y(new_n11721_));
  NOR3X1   g11529(.A(new_n11362_), .B(new_n11720_), .C(new_n11172_), .Y(new_n11722_));
  NOR2X1   g11530(.A(new_n11722_), .B(new_n11177_), .Y(new_n11723_));
  AOI21X1  g11531(.A0(new_n11721_), .A1(\asqrt[22] ), .B0(new_n11723_), .Y(new_n11724_));
  NOR3X1   g11532(.A(new_n11718_), .B(new_n11710_), .C(\asqrt[50] ), .Y(new_n11725_));
  OAI21X1  g11533(.A0(new_n11725_), .A1(new_n11724_), .B0(new_n11719_), .Y(new_n11726_));
  AND2X1   g11534(.A(new_n11726_), .B(\asqrt[51] ), .Y(new_n11727_));
  OR2X1    g11535(.A(new_n11725_), .B(new_n11724_), .Y(new_n11728_));
  OR4X1    g11536(.A(new_n11362_), .B(new_n11188_), .C(new_n11215_), .D(new_n11214_), .Y(new_n11729_));
  OR2X1    g11537(.A(new_n11188_), .B(new_n11214_), .Y(new_n11730_));
  OAI21X1  g11538(.A0(new_n11730_), .A1(new_n11362_), .B0(new_n11215_), .Y(new_n11731_));
  AND2X1   g11539(.A(new_n11731_), .B(new_n11729_), .Y(new_n11732_));
  AND2X1   g11540(.A(new_n11719_), .B(new_n1277_), .Y(new_n11733_));
  AOI21X1  g11541(.A0(new_n11733_), .A1(new_n11728_), .B0(new_n11732_), .Y(new_n11734_));
  OAI21X1  g11542(.A0(new_n11734_), .A1(new_n11727_), .B0(\asqrt[52] ), .Y(new_n11735_));
  AOI21X1  g11543(.A0(new_n11197_), .A1(new_n11191_), .B0(new_n11231_), .Y(new_n11736_));
  AND2X1   g11544(.A(new_n11736_), .B(new_n11229_), .Y(new_n11737_));
  AOI22X1  g11545(.A0(new_n11197_), .A1(new_n11191_), .B0(new_n11189_), .B1(\asqrt[51] ), .Y(new_n11738_));
  AOI21X1  g11546(.A0(new_n11738_), .A1(\asqrt[22] ), .B0(new_n11196_), .Y(new_n11739_));
  AOI21X1  g11547(.A0(new_n11737_), .A1(\asqrt[22] ), .B0(new_n11739_), .Y(new_n11740_));
  INVX1    g11548(.A(new_n11740_), .Y(new_n11741_));
  AND2X1   g11549(.A(new_n11716_), .B(\asqrt[48] ), .Y(new_n11742_));
  OR2X1    g11550(.A(new_n11700_), .B(new_n11687_), .Y(new_n11743_));
  AND2X1   g11551(.A(new_n11707_), .B(new_n1834_), .Y(new_n11744_));
  AOI21X1  g11552(.A0(new_n11744_), .A1(new_n11743_), .B0(new_n11705_), .Y(new_n11745_));
  OAI21X1  g11553(.A0(new_n11745_), .A1(new_n11742_), .B0(\asqrt[49] ), .Y(new_n11746_));
  INVX1    g11554(.A(new_n11715_), .Y(new_n11747_));
  OAI21X1  g11555(.A0(new_n11690_), .A1(new_n1834_), .B0(new_n1632_), .Y(new_n11748_));
  OAI21X1  g11556(.A0(new_n11748_), .A1(new_n11745_), .B0(new_n11747_), .Y(new_n11749_));
  AOI21X1  g11557(.A0(new_n11749_), .A1(new_n11746_), .B0(new_n1469_), .Y(new_n11750_));
  INVX1    g11558(.A(new_n11724_), .Y(new_n11751_));
  NAND3X1  g11559(.A(new_n11749_), .B(new_n11746_), .C(new_n1469_), .Y(new_n11752_));
  AOI21X1  g11560(.A0(new_n11752_), .A1(new_n11751_), .B0(new_n11750_), .Y(new_n11753_));
  OAI21X1  g11561(.A0(new_n11753_), .A1(new_n1277_), .B0(new_n1111_), .Y(new_n11754_));
  OAI21X1  g11562(.A0(new_n11754_), .A1(new_n11734_), .B0(new_n11741_), .Y(new_n11755_));
  AOI21X1  g11563(.A0(new_n11755_), .A1(new_n11735_), .B0(new_n968_), .Y(new_n11756_));
  AND2X1   g11564(.A(new_n11235_), .B(new_n11233_), .Y(new_n11757_));
  NOR3X1   g11565(.A(new_n11757_), .B(new_n11205_), .C(new_n11234_), .Y(new_n11758_));
  NOR3X1   g11566(.A(new_n11362_), .B(new_n11757_), .C(new_n11234_), .Y(new_n11759_));
  NOR2X1   g11567(.A(new_n11759_), .B(new_n11204_), .Y(new_n11760_));
  AOI21X1  g11568(.A0(new_n11758_), .A1(\asqrt[22] ), .B0(new_n11760_), .Y(new_n11761_));
  INVX1    g11569(.A(new_n11761_), .Y(new_n11762_));
  NAND3X1  g11570(.A(new_n11755_), .B(new_n11735_), .C(new_n968_), .Y(new_n11763_));
  AOI21X1  g11571(.A0(new_n11763_), .A1(new_n11762_), .B0(new_n11756_), .Y(new_n11764_));
  OR2X1    g11572(.A(new_n11764_), .B(new_n902_), .Y(new_n11765_));
  OR2X1    g11573(.A(new_n11753_), .B(new_n1277_), .Y(new_n11766_));
  NOR2X1   g11574(.A(new_n11725_), .B(new_n11724_), .Y(new_n11767_));
  INVX1    g11575(.A(new_n11732_), .Y(new_n11768_));
  NAND2X1  g11576(.A(new_n11719_), .B(new_n1277_), .Y(new_n11769_));
  OAI21X1  g11577(.A0(new_n11769_), .A1(new_n11767_), .B0(new_n11768_), .Y(new_n11770_));
  AOI21X1  g11578(.A0(new_n11770_), .A1(new_n11766_), .B0(new_n1111_), .Y(new_n11771_));
  AOI21X1  g11579(.A0(new_n11726_), .A1(\asqrt[51] ), .B0(\asqrt[52] ), .Y(new_n11772_));
  AOI21X1  g11580(.A0(new_n11772_), .A1(new_n11770_), .B0(new_n11740_), .Y(new_n11773_));
  NOR3X1   g11581(.A(new_n11773_), .B(new_n11771_), .C(\asqrt[53] ), .Y(new_n11774_));
  NOR2X1   g11582(.A(new_n11774_), .B(new_n11761_), .Y(new_n11775_));
  OR4X1    g11583(.A(new_n11362_), .B(new_n11237_), .C(new_n11225_), .D(new_n11220_), .Y(new_n11776_));
  OR2X1    g11584(.A(new_n11237_), .B(new_n11220_), .Y(new_n11777_));
  OAI21X1  g11585(.A0(new_n11777_), .A1(new_n11362_), .B0(new_n11225_), .Y(new_n11778_));
  AND2X1   g11586(.A(new_n11778_), .B(new_n11776_), .Y(new_n11779_));
  INVX1    g11587(.A(new_n11779_), .Y(new_n11780_));
  OAI21X1  g11588(.A0(new_n11773_), .A1(new_n11771_), .B0(\asqrt[53] ), .Y(new_n11781_));
  NAND2X1  g11589(.A(new_n11781_), .B(new_n902_), .Y(new_n11782_));
  OAI21X1  g11590(.A0(new_n11782_), .A1(new_n11775_), .B0(new_n11780_), .Y(new_n11783_));
  AOI21X1  g11591(.A0(new_n11783_), .A1(new_n11765_), .B0(new_n697_), .Y(new_n11784_));
  AND2X1   g11592(.A(new_n11282_), .B(new_n11281_), .Y(new_n11785_));
  NOR3X1   g11593(.A(new_n11785_), .B(new_n11244_), .C(new_n11280_), .Y(new_n11786_));
  NOR3X1   g11594(.A(new_n11362_), .B(new_n11785_), .C(new_n11280_), .Y(new_n11787_));
  NOR2X1   g11595(.A(new_n11787_), .B(new_n11243_), .Y(new_n11788_));
  AOI21X1  g11596(.A0(new_n11786_), .A1(\asqrt[22] ), .B0(new_n11788_), .Y(new_n11789_));
  OAI21X1  g11597(.A0(new_n11774_), .A1(new_n11761_), .B0(new_n11781_), .Y(new_n11790_));
  AOI21X1  g11598(.A0(new_n11790_), .A1(\asqrt[54] ), .B0(\asqrt[55] ), .Y(new_n11791_));
  AOI21X1  g11599(.A0(new_n11791_), .A1(new_n11783_), .B0(new_n11789_), .Y(new_n11792_));
  OAI21X1  g11600(.A0(new_n11792_), .A1(new_n11784_), .B0(\asqrt[56] ), .Y(new_n11793_));
  AND2X1   g11601(.A(new_n11255_), .B(new_n11247_), .Y(new_n11794_));
  NOR3X1   g11602(.A(new_n11794_), .B(new_n11285_), .C(new_n11248_), .Y(new_n11795_));
  NOR3X1   g11603(.A(new_n11362_), .B(new_n11794_), .C(new_n11248_), .Y(new_n11796_));
  NOR2X1   g11604(.A(new_n11796_), .B(new_n11253_), .Y(new_n11797_));
  AOI21X1  g11605(.A0(new_n11795_), .A1(\asqrt[22] ), .B0(new_n11797_), .Y(new_n11798_));
  NOR3X1   g11606(.A(new_n11792_), .B(new_n11784_), .C(\asqrt[56] ), .Y(new_n11799_));
  OAI21X1  g11607(.A0(new_n11799_), .A1(new_n11798_), .B0(new_n11793_), .Y(new_n11800_));
  AND2X1   g11608(.A(new_n11800_), .B(\asqrt[57] ), .Y(new_n11801_));
  OR2X1    g11609(.A(new_n11799_), .B(new_n11798_), .Y(new_n11802_));
  OR4X1    g11610(.A(new_n11362_), .B(new_n11262_), .C(new_n11289_), .D(new_n11288_), .Y(new_n11803_));
  OR2X1    g11611(.A(new_n11262_), .B(new_n11288_), .Y(new_n11804_));
  OAI21X1  g11612(.A0(new_n11804_), .A1(new_n11362_), .B0(new_n11289_), .Y(new_n11805_));
  AND2X1   g11613(.A(new_n11805_), .B(new_n11803_), .Y(new_n11806_));
  AND2X1   g11614(.A(new_n11793_), .B(new_n481_), .Y(new_n11807_));
  AOI21X1  g11615(.A0(new_n11807_), .A1(new_n11802_), .B0(new_n11806_), .Y(new_n11808_));
  OAI21X1  g11616(.A0(new_n11808_), .A1(new_n11801_), .B0(\asqrt[58] ), .Y(new_n11809_));
  AOI21X1  g11617(.A0(new_n11271_), .A1(new_n11265_), .B0(new_n11310_), .Y(new_n11810_));
  AND2X1   g11618(.A(new_n11810_), .B(new_n11308_), .Y(new_n11811_));
  AOI22X1  g11619(.A0(new_n11271_), .A1(new_n11265_), .B0(new_n11263_), .B1(\asqrt[57] ), .Y(new_n11812_));
  AOI21X1  g11620(.A0(new_n11812_), .A1(\asqrt[22] ), .B0(new_n11270_), .Y(new_n11813_));
  AOI21X1  g11621(.A0(new_n11811_), .A1(\asqrt[22] ), .B0(new_n11813_), .Y(new_n11814_));
  INVX1    g11622(.A(new_n11814_), .Y(new_n11815_));
  AND2X1   g11623(.A(new_n11790_), .B(\asqrt[54] ), .Y(new_n11816_));
  OR2X1    g11624(.A(new_n11774_), .B(new_n11761_), .Y(new_n11817_));
  AND2X1   g11625(.A(new_n11781_), .B(new_n902_), .Y(new_n11818_));
  AOI21X1  g11626(.A0(new_n11818_), .A1(new_n11817_), .B0(new_n11779_), .Y(new_n11819_));
  OAI21X1  g11627(.A0(new_n11819_), .A1(new_n11816_), .B0(\asqrt[55] ), .Y(new_n11820_));
  INVX1    g11628(.A(new_n11789_), .Y(new_n11821_));
  OAI21X1  g11629(.A0(new_n11764_), .A1(new_n902_), .B0(new_n697_), .Y(new_n11822_));
  OAI21X1  g11630(.A0(new_n11822_), .A1(new_n11819_), .B0(new_n11821_), .Y(new_n11823_));
  AOI21X1  g11631(.A0(new_n11823_), .A1(new_n11820_), .B0(new_n582_), .Y(new_n11824_));
  INVX1    g11632(.A(new_n11798_), .Y(new_n11825_));
  NAND3X1  g11633(.A(new_n11823_), .B(new_n11820_), .C(new_n582_), .Y(new_n11826_));
  AOI21X1  g11634(.A0(new_n11826_), .A1(new_n11825_), .B0(new_n11824_), .Y(new_n11827_));
  OAI21X1  g11635(.A0(new_n11827_), .A1(new_n481_), .B0(new_n399_), .Y(new_n11828_));
  OAI21X1  g11636(.A0(new_n11828_), .A1(new_n11808_), .B0(new_n11815_), .Y(new_n11829_));
  AOI21X1  g11637(.A0(new_n11829_), .A1(new_n11809_), .B0(new_n328_), .Y(new_n11830_));
  AND2X1   g11638(.A(new_n11314_), .B(new_n11312_), .Y(new_n11831_));
  NOR3X1   g11639(.A(new_n11831_), .B(new_n11279_), .C(new_n11313_), .Y(new_n11832_));
  NOR3X1   g11640(.A(new_n11362_), .B(new_n11831_), .C(new_n11313_), .Y(new_n11833_));
  NOR2X1   g11641(.A(new_n11833_), .B(new_n11278_), .Y(new_n11834_));
  AOI21X1  g11642(.A0(new_n11832_), .A1(\asqrt[22] ), .B0(new_n11834_), .Y(new_n11835_));
  INVX1    g11643(.A(new_n11835_), .Y(new_n11836_));
  NAND3X1  g11644(.A(new_n11829_), .B(new_n11809_), .C(new_n328_), .Y(new_n11837_));
  AOI21X1  g11645(.A0(new_n11837_), .A1(new_n11836_), .B0(new_n11830_), .Y(new_n11838_));
  OR2X1    g11646(.A(new_n11838_), .B(new_n292_), .Y(new_n11839_));
  OR2X1    g11647(.A(new_n11827_), .B(new_n481_), .Y(new_n11840_));
  NOR2X1   g11648(.A(new_n11799_), .B(new_n11798_), .Y(new_n11841_));
  INVX1    g11649(.A(new_n11806_), .Y(new_n11842_));
  NAND2X1  g11650(.A(new_n11793_), .B(new_n481_), .Y(new_n11843_));
  OAI21X1  g11651(.A0(new_n11843_), .A1(new_n11841_), .B0(new_n11842_), .Y(new_n11844_));
  AOI21X1  g11652(.A0(new_n11844_), .A1(new_n11840_), .B0(new_n399_), .Y(new_n11845_));
  AOI21X1  g11653(.A0(new_n11800_), .A1(\asqrt[57] ), .B0(\asqrt[58] ), .Y(new_n11846_));
  AOI21X1  g11654(.A0(new_n11846_), .A1(new_n11844_), .B0(new_n11814_), .Y(new_n11847_));
  NOR3X1   g11655(.A(new_n11847_), .B(new_n11845_), .C(\asqrt[59] ), .Y(new_n11848_));
  NOR2X1   g11656(.A(new_n11848_), .B(new_n11835_), .Y(new_n11849_));
  OR4X1    g11657(.A(new_n11362_), .B(new_n11326_), .C(new_n11297_), .D(new_n11294_), .Y(new_n11850_));
  OR2X1    g11658(.A(new_n11326_), .B(new_n11294_), .Y(new_n11851_));
  OAI21X1  g11659(.A0(new_n11851_), .A1(new_n11362_), .B0(new_n11297_), .Y(new_n11852_));
  AND2X1   g11660(.A(new_n11852_), .B(new_n11850_), .Y(new_n11853_));
  INVX1    g11661(.A(new_n11853_), .Y(new_n11854_));
  OAI21X1  g11662(.A0(new_n11847_), .A1(new_n11845_), .B0(\asqrt[59] ), .Y(new_n11855_));
  NAND2X1  g11663(.A(new_n11855_), .B(new_n292_), .Y(new_n11856_));
  OAI21X1  g11664(.A0(new_n11856_), .A1(new_n11849_), .B0(new_n11854_), .Y(new_n11857_));
  AOI21X1  g11665(.A0(new_n11857_), .A1(new_n11839_), .B0(new_n217_), .Y(new_n11858_));
  AND2X1   g11666(.A(new_n11371_), .B(new_n11370_), .Y(new_n11859_));
  NOR3X1   g11667(.A(new_n11859_), .B(new_n11307_), .C(new_n11369_), .Y(new_n11860_));
  NOR3X1   g11668(.A(new_n11362_), .B(new_n11859_), .C(new_n11369_), .Y(new_n11861_));
  NOR2X1   g11669(.A(new_n11861_), .B(new_n11306_), .Y(new_n11862_));
  AOI21X1  g11670(.A0(new_n11860_), .A1(\asqrt[22] ), .B0(new_n11862_), .Y(new_n11863_));
  OAI21X1  g11671(.A0(new_n11848_), .A1(new_n11835_), .B0(new_n11855_), .Y(new_n11864_));
  AOI21X1  g11672(.A0(new_n11864_), .A1(\asqrt[60] ), .B0(\asqrt[61] ), .Y(new_n11865_));
  AOI21X1  g11673(.A0(new_n11865_), .A1(new_n11857_), .B0(new_n11863_), .Y(new_n11866_));
  OAI21X1  g11674(.A0(new_n11866_), .A1(new_n11858_), .B0(\asqrt[62] ), .Y(new_n11867_));
  AND2X1   g11675(.A(new_n11328_), .B(new_n11318_), .Y(new_n11868_));
  NOR3X1   g11676(.A(new_n11868_), .B(new_n11374_), .C(new_n11319_), .Y(new_n11869_));
  NOR3X1   g11677(.A(new_n11362_), .B(new_n11868_), .C(new_n11319_), .Y(new_n11870_));
  NOR2X1   g11678(.A(new_n11870_), .B(new_n11324_), .Y(new_n11871_));
  AOI21X1  g11679(.A0(new_n11869_), .A1(\asqrt[22] ), .B0(new_n11871_), .Y(new_n11872_));
  NOR3X1   g11680(.A(new_n11866_), .B(new_n11858_), .C(\asqrt[62] ), .Y(new_n11873_));
  OAI21X1  g11681(.A0(new_n11873_), .A1(new_n11872_), .B0(new_n11867_), .Y(new_n11874_));
  NOR4X1   g11682(.A(new_n11362_), .B(new_n11335_), .C(new_n11378_), .D(new_n11377_), .Y(new_n11875_));
  NOR3X1   g11683(.A(new_n11362_), .B(new_n11335_), .C(new_n11377_), .Y(new_n11876_));
  NOR2X1   g11684(.A(new_n11876_), .B(new_n11334_), .Y(new_n11877_));
  NOR2X1   g11685(.A(new_n11877_), .B(new_n11875_), .Y(new_n11878_));
  INVX1    g11686(.A(new_n11878_), .Y(new_n11879_));
  AND2X1   g11687(.A(new_n11343_), .B(new_n11336_), .Y(new_n11880_));
  AOI21X1  g11688(.A0(new_n11880_), .A1(\asqrt[22] ), .B0(new_n11398_), .Y(new_n11881_));
  AND2X1   g11689(.A(new_n11881_), .B(new_n11879_), .Y(new_n11882_));
  AOI21X1  g11690(.A0(new_n11882_), .A1(new_n11874_), .B0(\asqrt[63] ), .Y(new_n11883_));
  NOR2X1   g11691(.A(new_n11873_), .B(new_n11872_), .Y(new_n11884_));
  NAND2X1  g11692(.A(new_n11878_), .B(new_n11867_), .Y(new_n11885_));
  AOI21X1  g11693(.A0(new_n11386_), .A1(new_n11382_), .B0(new_n11342_), .Y(new_n11886_));
  AOI21X1  g11694(.A0(new_n11343_), .A1(new_n11336_), .B0(new_n193_), .Y(new_n11887_));
  OAI21X1  g11695(.A0(new_n11886_), .A1(new_n11336_), .B0(new_n11887_), .Y(new_n11888_));
  INVX1    g11696(.A(new_n11341_), .Y(new_n11889_));
  NOR4X1   g11697(.A(new_n11359_), .B(new_n11353_), .C(new_n11889_), .D(new_n11338_), .Y(new_n11890_));
  OAI21X1  g11698(.A0(new_n11350_), .A1(new_n11349_), .B0(new_n11890_), .Y(new_n11891_));
  NOR2X1   g11699(.A(new_n11891_), .B(new_n11348_), .Y(new_n11892_));
  INVX1    g11700(.A(new_n11892_), .Y(new_n11893_));
  AND2X1   g11701(.A(new_n11893_), .B(new_n11888_), .Y(new_n11894_));
  OAI21X1  g11702(.A0(new_n11885_), .A1(new_n11884_), .B0(new_n11894_), .Y(new_n11895_));
  NOR2X1   g11703(.A(new_n11895_), .B(new_n11883_), .Y(new_n11896_));
  OAI21X1  g11704(.A0(new_n11895_), .A1(new_n11883_), .B0(\a[42] ), .Y(new_n11897_));
  NOR3X1   g11705(.A(\a[42] ), .B(\a[41] ), .C(\a[40] ), .Y(new_n11898_));
  INVX1    g11706(.A(new_n11898_), .Y(new_n11899_));
  AOI21X1  g11707(.A0(new_n11899_), .A1(new_n11897_), .B0(new_n11362_), .Y(new_n11900_));
  OR2X1    g11708(.A(new_n11898_), .B(new_n11359_), .Y(new_n11901_));
  NOR4X1   g11709(.A(new_n11901_), .B(new_n11353_), .C(new_n11398_), .D(new_n11348_), .Y(new_n11902_));
  NAND2X1  g11710(.A(new_n11902_), .B(new_n11897_), .Y(new_n11903_));
  INVX1    g11711(.A(\a[42] ), .Y(new_n11904_));
  OAI21X1  g11712(.A0(new_n11895_), .A1(new_n11883_), .B0(new_n11904_), .Y(new_n11905_));
  INVX1    g11713(.A(new_n11366_), .Y(new_n11906_));
  AND2X1   g11714(.A(new_n11864_), .B(\asqrt[60] ), .Y(new_n11907_));
  OR2X1    g11715(.A(new_n11848_), .B(new_n11835_), .Y(new_n11908_));
  AND2X1   g11716(.A(new_n11855_), .B(new_n292_), .Y(new_n11909_));
  AOI21X1  g11717(.A0(new_n11909_), .A1(new_n11908_), .B0(new_n11853_), .Y(new_n11910_));
  OAI21X1  g11718(.A0(new_n11910_), .A1(new_n11907_), .B0(\asqrt[61] ), .Y(new_n11911_));
  INVX1    g11719(.A(new_n11863_), .Y(new_n11912_));
  OAI21X1  g11720(.A0(new_n11838_), .A1(new_n292_), .B0(new_n217_), .Y(new_n11913_));
  OAI21X1  g11721(.A0(new_n11913_), .A1(new_n11910_), .B0(new_n11912_), .Y(new_n11914_));
  AOI21X1  g11722(.A0(new_n11914_), .A1(new_n11911_), .B0(new_n199_), .Y(new_n11915_));
  INVX1    g11723(.A(new_n11872_), .Y(new_n11916_));
  NAND3X1  g11724(.A(new_n11914_), .B(new_n11911_), .C(new_n199_), .Y(new_n11917_));
  AOI21X1  g11725(.A0(new_n11917_), .A1(new_n11916_), .B0(new_n11915_), .Y(new_n11918_));
  INVX1    g11726(.A(new_n11882_), .Y(new_n11919_));
  OAI21X1  g11727(.A0(new_n11919_), .A1(new_n11918_), .B0(new_n193_), .Y(new_n11920_));
  OR2X1    g11728(.A(new_n11873_), .B(new_n11872_), .Y(new_n11921_));
  AND2X1   g11729(.A(new_n11878_), .B(new_n11867_), .Y(new_n11922_));
  INVX1    g11730(.A(new_n11894_), .Y(new_n11923_));
  AOI21X1  g11731(.A0(new_n11922_), .A1(new_n11921_), .B0(new_n11923_), .Y(new_n11924_));
  AOI21X1  g11732(.A0(new_n11924_), .A1(new_n11920_), .B0(new_n11906_), .Y(new_n11925_));
  AOI21X1  g11733(.A0(new_n11905_), .A1(\a[43] ), .B0(new_n11925_), .Y(new_n11926_));
  AOI21X1  g11734(.A0(new_n11926_), .A1(new_n11903_), .B0(new_n11900_), .Y(new_n11927_));
  OR2X1    g11735(.A(new_n11927_), .B(new_n10849_), .Y(new_n11928_));
  AND2X1   g11736(.A(new_n11926_), .B(new_n11903_), .Y(new_n11929_));
  OR2X1    g11737(.A(new_n11900_), .B(\asqrt[23] ), .Y(new_n11930_));
  OAI21X1  g11738(.A0(new_n11895_), .A1(new_n11883_), .B0(new_n11366_), .Y(new_n11931_));
  INVX1    g11739(.A(new_n11888_), .Y(new_n11932_));
  NOR3X1   g11740(.A(new_n11892_), .B(new_n11932_), .C(new_n11362_), .Y(new_n11933_));
  OAI21X1  g11741(.A0(new_n11885_), .A1(new_n11884_), .B0(new_n11933_), .Y(new_n11934_));
  OR2X1    g11742(.A(new_n11934_), .B(new_n11883_), .Y(new_n11935_));
  AOI21X1  g11743(.A0(new_n11935_), .A1(new_n11931_), .B0(new_n11365_), .Y(new_n11936_));
  OAI21X1  g11744(.A0(new_n11934_), .A1(new_n11883_), .B0(new_n11365_), .Y(new_n11937_));
  NOR2X1   g11745(.A(new_n11937_), .B(new_n11925_), .Y(new_n11938_));
  OR2X1    g11746(.A(new_n11938_), .B(new_n11936_), .Y(new_n11939_));
  OAI21X1  g11747(.A0(new_n11930_), .A1(new_n11929_), .B0(new_n11939_), .Y(new_n11940_));
  AOI21X1  g11748(.A0(new_n11940_), .A1(new_n11928_), .B0(new_n10332_), .Y(new_n11941_));
  OR4X1    g11749(.A(new_n11896_), .B(new_n11392_), .C(new_n11414_), .D(new_n11368_), .Y(new_n11942_));
  NOR3X1   g11750(.A(new_n11896_), .B(new_n11414_), .C(new_n11368_), .Y(new_n11943_));
  OR2X1    g11751(.A(new_n11943_), .B(new_n11417_), .Y(new_n11944_));
  AOI21X1  g11752(.A0(new_n11924_), .A1(new_n11920_), .B0(new_n11904_), .Y(new_n11945_));
  OAI21X1  g11753(.A0(new_n11898_), .A1(new_n11945_), .B0(\asqrt[22] ), .Y(new_n11946_));
  AND2X1   g11754(.A(new_n11902_), .B(new_n11897_), .Y(new_n11947_));
  INVX1    g11755(.A(\a[43] ), .Y(new_n11948_));
  AOI21X1  g11756(.A0(new_n11924_), .A1(new_n11920_), .B0(\a[42] ), .Y(new_n11949_));
  OAI21X1  g11757(.A0(new_n11949_), .A1(new_n11948_), .B0(new_n11931_), .Y(new_n11950_));
  OAI21X1  g11758(.A0(new_n11950_), .A1(new_n11947_), .B0(new_n11946_), .Y(new_n11951_));
  AOI21X1  g11759(.A0(new_n11951_), .A1(\asqrt[23] ), .B0(\asqrt[24] ), .Y(new_n11952_));
  AOI22X1  g11760(.A0(new_n11952_), .A1(new_n11940_), .B0(new_n11944_), .B1(new_n11942_), .Y(new_n11953_));
  OAI21X1  g11761(.A0(new_n11953_), .A1(new_n11941_), .B0(\asqrt[25] ), .Y(new_n11954_));
  AOI21X1  g11762(.A0(new_n11438_), .A1(new_n11437_), .B0(new_n11404_), .Y(new_n11955_));
  AND2X1   g11763(.A(new_n11955_), .B(new_n11394_), .Y(new_n11956_));
  OAI21X1  g11764(.A0(new_n11895_), .A1(new_n11883_), .B0(new_n11956_), .Y(new_n11957_));
  AOI22X1  g11765(.A0(new_n11438_), .A1(new_n11437_), .B0(new_n11418_), .B1(\asqrt[24] ), .Y(new_n11958_));
  OAI21X1  g11766(.A0(new_n11895_), .A1(new_n11883_), .B0(new_n11958_), .Y(new_n11959_));
  NAND2X1  g11767(.A(new_n11959_), .B(new_n11404_), .Y(new_n11960_));
  AND2X1   g11768(.A(new_n11960_), .B(new_n11957_), .Y(new_n11961_));
  NOR3X1   g11769(.A(new_n11953_), .B(new_n11941_), .C(\asqrt[25] ), .Y(new_n11962_));
  OAI21X1  g11770(.A0(new_n11962_), .A1(new_n11961_), .B0(new_n11954_), .Y(new_n11963_));
  AND2X1   g11771(.A(new_n11963_), .B(\asqrt[26] ), .Y(new_n11964_));
  OR2X1    g11772(.A(new_n11962_), .B(new_n11961_), .Y(new_n11965_));
  INVX1    g11773(.A(new_n11896_), .Y(\asqrt[21] ));
  AND2X1   g11774(.A(new_n11419_), .B(new_n11405_), .Y(new_n11967_));
  NOR3X1   g11775(.A(new_n11967_), .B(new_n11442_), .C(new_n11406_), .Y(new_n11968_));
  NOR2X1   g11776(.A(new_n11967_), .B(new_n11406_), .Y(new_n11969_));
  OAI21X1  g11777(.A0(new_n11895_), .A1(new_n11883_), .B0(new_n11969_), .Y(new_n11970_));
  AOI22X1  g11778(.A0(new_n11970_), .A1(new_n11442_), .B0(new_n11968_), .B1(\asqrt[21] ), .Y(new_n11971_));
  AND2X1   g11779(.A(new_n11954_), .B(new_n9353_), .Y(new_n11972_));
  AOI21X1  g11780(.A0(new_n11972_), .A1(new_n11965_), .B0(new_n11971_), .Y(new_n11973_));
  OAI21X1  g11781(.A0(new_n11973_), .A1(new_n11964_), .B0(\asqrt[27] ), .Y(new_n11974_));
  NAND4X1  g11782(.A(\asqrt[21] ), .B(new_n11456_), .C(new_n11428_), .D(new_n11421_), .Y(new_n11975_));
  NOR3X1   g11783(.A(new_n11896_), .B(new_n11429_), .C(new_n11445_), .Y(new_n11976_));
  OAI21X1  g11784(.A0(new_n11976_), .A1(new_n11428_), .B0(new_n11975_), .Y(new_n11977_));
  AND2X1   g11785(.A(new_n11951_), .B(\asqrt[23] ), .Y(new_n11978_));
  NAND2X1  g11786(.A(new_n11926_), .B(new_n11903_), .Y(new_n11979_));
  AND2X1   g11787(.A(new_n11946_), .B(new_n10849_), .Y(new_n11980_));
  NOR2X1   g11788(.A(new_n11938_), .B(new_n11936_), .Y(new_n11981_));
  AOI21X1  g11789(.A0(new_n11980_), .A1(new_n11979_), .B0(new_n11981_), .Y(new_n11982_));
  OAI21X1  g11790(.A0(new_n11982_), .A1(new_n11978_), .B0(\asqrt[24] ), .Y(new_n11983_));
  OAI21X1  g11791(.A0(new_n11943_), .A1(new_n11417_), .B0(new_n11942_), .Y(new_n11984_));
  OAI21X1  g11792(.A0(new_n11927_), .A1(new_n10849_), .B0(new_n10332_), .Y(new_n11985_));
  OAI21X1  g11793(.A0(new_n11985_), .A1(new_n11982_), .B0(new_n11984_), .Y(new_n11986_));
  AOI21X1  g11794(.A0(new_n11986_), .A1(new_n11983_), .B0(new_n9833_), .Y(new_n11987_));
  INVX1    g11795(.A(new_n11961_), .Y(new_n11988_));
  NAND3X1  g11796(.A(new_n11986_), .B(new_n11983_), .C(new_n9833_), .Y(new_n11989_));
  AOI21X1  g11797(.A0(new_n11989_), .A1(new_n11988_), .B0(new_n11987_), .Y(new_n11990_));
  OAI21X1  g11798(.A0(new_n11990_), .A1(new_n9353_), .B0(new_n8874_), .Y(new_n11991_));
  OAI21X1  g11799(.A0(new_n11991_), .A1(new_n11973_), .B0(new_n11977_), .Y(new_n11992_));
  AOI21X1  g11800(.A0(new_n11992_), .A1(new_n11974_), .B0(new_n8412_), .Y(new_n11993_));
  AND2X1   g11801(.A(new_n11446_), .B(new_n11432_), .Y(new_n11994_));
  NOR3X1   g11802(.A(new_n11994_), .B(new_n11472_), .C(new_n11431_), .Y(new_n11995_));
  NOR3X1   g11803(.A(new_n11896_), .B(new_n11994_), .C(new_n11431_), .Y(new_n11996_));
  NOR2X1   g11804(.A(new_n11996_), .B(new_n11435_), .Y(new_n11997_));
  AOI21X1  g11805(.A0(new_n11995_), .A1(\asqrt[21] ), .B0(new_n11997_), .Y(new_n11998_));
  INVX1    g11806(.A(new_n11998_), .Y(new_n11999_));
  NAND3X1  g11807(.A(new_n11992_), .B(new_n11974_), .C(new_n8412_), .Y(new_n12000_));
  AOI21X1  g11808(.A0(new_n12000_), .A1(new_n11999_), .B0(new_n11993_), .Y(new_n12001_));
  OR2X1    g11809(.A(new_n12001_), .B(new_n7970_), .Y(new_n12002_));
  AND2X1   g11810(.A(new_n12000_), .B(new_n11999_), .Y(new_n12003_));
  AND2X1   g11811(.A(new_n11476_), .B(new_n11474_), .Y(new_n12004_));
  NOR3X1   g11812(.A(new_n12004_), .B(new_n11454_), .C(new_n11475_), .Y(new_n12005_));
  NOR3X1   g11813(.A(new_n11896_), .B(new_n12004_), .C(new_n11475_), .Y(new_n12006_));
  NOR2X1   g11814(.A(new_n12006_), .B(new_n11453_), .Y(new_n12007_));
  AOI21X1  g11815(.A0(new_n12005_), .A1(\asqrt[21] ), .B0(new_n12007_), .Y(new_n12008_));
  INVX1    g11816(.A(new_n12008_), .Y(new_n12009_));
  OR2X1    g11817(.A(new_n11990_), .B(new_n9353_), .Y(new_n12010_));
  NOR2X1   g11818(.A(new_n11962_), .B(new_n11961_), .Y(new_n12011_));
  INVX1    g11819(.A(new_n11971_), .Y(new_n12012_));
  NAND2X1  g11820(.A(new_n11954_), .B(new_n9353_), .Y(new_n12013_));
  OAI21X1  g11821(.A0(new_n12013_), .A1(new_n12011_), .B0(new_n12012_), .Y(new_n12014_));
  AOI21X1  g11822(.A0(new_n12014_), .A1(new_n12010_), .B0(new_n8874_), .Y(new_n12015_));
  INVX1    g11823(.A(new_n11977_), .Y(new_n12016_));
  AOI21X1  g11824(.A0(new_n11963_), .A1(\asqrt[26] ), .B0(\asqrt[27] ), .Y(new_n12017_));
  AOI21X1  g11825(.A0(new_n12017_), .A1(new_n12014_), .B0(new_n12016_), .Y(new_n12018_));
  OAI21X1  g11826(.A0(new_n12018_), .A1(new_n12015_), .B0(\asqrt[28] ), .Y(new_n12019_));
  NAND2X1  g11827(.A(new_n12019_), .B(new_n7970_), .Y(new_n12020_));
  OAI21X1  g11828(.A0(new_n12020_), .A1(new_n12003_), .B0(new_n12009_), .Y(new_n12021_));
  AOI21X1  g11829(.A0(new_n12021_), .A1(new_n12002_), .B0(new_n7527_), .Y(new_n12022_));
  OR4X1    g11830(.A(new_n11896_), .B(new_n11478_), .C(new_n11466_), .D(new_n11460_), .Y(new_n12023_));
  OR2X1    g11831(.A(new_n11478_), .B(new_n11460_), .Y(new_n12024_));
  OAI21X1  g11832(.A0(new_n12024_), .A1(new_n11896_), .B0(new_n11466_), .Y(new_n12025_));
  AND2X1   g11833(.A(new_n12025_), .B(new_n12023_), .Y(new_n12026_));
  NOR3X1   g11834(.A(new_n12018_), .B(new_n12015_), .C(\asqrt[28] ), .Y(new_n12027_));
  OAI21X1  g11835(.A0(new_n12027_), .A1(new_n11998_), .B0(new_n12019_), .Y(new_n12028_));
  AOI21X1  g11836(.A0(new_n12028_), .A1(\asqrt[29] ), .B0(\asqrt[30] ), .Y(new_n12029_));
  AOI21X1  g11837(.A0(new_n12029_), .A1(new_n12021_), .B0(new_n12026_), .Y(new_n12030_));
  OAI21X1  g11838(.A0(new_n12030_), .A1(new_n12022_), .B0(\asqrt[31] ), .Y(new_n12031_));
  AOI21X1  g11839(.A0(new_n11509_), .A1(new_n11508_), .B0(new_n11484_), .Y(new_n12032_));
  AND2X1   g11840(.A(new_n12032_), .B(new_n11469_), .Y(new_n12033_));
  AOI22X1  g11841(.A0(new_n11509_), .A1(new_n11508_), .B0(new_n11494_), .B1(\asqrt[30] ), .Y(new_n12034_));
  AOI21X1  g11842(.A0(new_n12034_), .A1(\asqrt[21] ), .B0(new_n11483_), .Y(new_n12035_));
  AOI21X1  g11843(.A0(new_n12033_), .A1(\asqrt[21] ), .B0(new_n12035_), .Y(new_n12036_));
  NOR3X1   g11844(.A(new_n12030_), .B(new_n12022_), .C(\asqrt[31] ), .Y(new_n12037_));
  OAI21X1  g11845(.A0(new_n12037_), .A1(new_n12036_), .B0(new_n12031_), .Y(new_n12038_));
  AND2X1   g11846(.A(new_n12038_), .B(\asqrt[32] ), .Y(new_n12039_));
  INVX1    g11847(.A(new_n12036_), .Y(new_n12040_));
  AND2X1   g11848(.A(new_n12028_), .B(\asqrt[29] ), .Y(new_n12041_));
  NAND2X1  g11849(.A(new_n12000_), .B(new_n11999_), .Y(new_n12042_));
  AND2X1   g11850(.A(new_n12019_), .B(new_n7970_), .Y(new_n12043_));
  AOI21X1  g11851(.A0(new_n12043_), .A1(new_n12042_), .B0(new_n12008_), .Y(new_n12044_));
  OAI21X1  g11852(.A0(new_n12044_), .A1(new_n12041_), .B0(\asqrt[30] ), .Y(new_n12045_));
  INVX1    g11853(.A(new_n12026_), .Y(new_n12046_));
  OAI21X1  g11854(.A0(new_n12001_), .A1(new_n7970_), .B0(new_n7527_), .Y(new_n12047_));
  OAI21X1  g11855(.A0(new_n12047_), .A1(new_n12044_), .B0(new_n12046_), .Y(new_n12048_));
  NAND3X1  g11856(.A(new_n12048_), .B(new_n12045_), .C(new_n7103_), .Y(new_n12049_));
  NAND2X1  g11857(.A(new_n12049_), .B(new_n12040_), .Y(new_n12050_));
  AND2X1   g11858(.A(new_n11495_), .B(new_n11487_), .Y(new_n12051_));
  NOR3X1   g11859(.A(new_n12051_), .B(new_n11512_), .C(new_n11488_), .Y(new_n12052_));
  NOR3X1   g11860(.A(new_n11896_), .B(new_n12051_), .C(new_n11488_), .Y(new_n12053_));
  NOR2X1   g11861(.A(new_n12053_), .B(new_n11493_), .Y(new_n12054_));
  AOI21X1  g11862(.A0(new_n12052_), .A1(\asqrt[21] ), .B0(new_n12054_), .Y(new_n12055_));
  AND2X1   g11863(.A(new_n12031_), .B(new_n6699_), .Y(new_n12056_));
  AOI21X1  g11864(.A0(new_n12056_), .A1(new_n12050_), .B0(new_n12055_), .Y(new_n12057_));
  OAI21X1  g11865(.A0(new_n12057_), .A1(new_n12039_), .B0(\asqrt[33] ), .Y(new_n12058_));
  OR4X1    g11866(.A(new_n11896_), .B(new_n11503_), .C(new_n11506_), .D(new_n11521_), .Y(new_n12059_));
  OR2X1    g11867(.A(new_n11503_), .B(new_n11521_), .Y(new_n12060_));
  OAI21X1  g11868(.A0(new_n12060_), .A1(new_n11896_), .B0(new_n11506_), .Y(new_n12061_));
  AND2X1   g11869(.A(new_n12061_), .B(new_n12059_), .Y(new_n12062_));
  INVX1    g11870(.A(new_n12062_), .Y(new_n12063_));
  AOI21X1  g11871(.A0(new_n12048_), .A1(new_n12045_), .B0(new_n7103_), .Y(new_n12064_));
  AOI21X1  g11872(.A0(new_n12049_), .A1(new_n12040_), .B0(new_n12064_), .Y(new_n12065_));
  OAI21X1  g11873(.A0(new_n12065_), .A1(new_n6699_), .B0(new_n6294_), .Y(new_n12066_));
  OAI21X1  g11874(.A0(new_n12066_), .A1(new_n12057_), .B0(new_n12063_), .Y(new_n12067_));
  AOI21X1  g11875(.A0(new_n12067_), .A1(new_n12058_), .B0(new_n5941_), .Y(new_n12068_));
  AND2X1   g11876(.A(new_n11522_), .B(new_n11516_), .Y(new_n12069_));
  NOR3X1   g11877(.A(new_n12069_), .B(new_n11560_), .C(new_n11505_), .Y(new_n12070_));
  NOR3X1   g11878(.A(new_n11896_), .B(new_n12069_), .C(new_n11505_), .Y(new_n12071_));
  NOR2X1   g11879(.A(new_n12071_), .B(new_n11520_), .Y(new_n12072_));
  AOI21X1  g11880(.A0(new_n12070_), .A1(\asqrt[21] ), .B0(new_n12072_), .Y(new_n12073_));
  INVX1    g11881(.A(new_n12073_), .Y(new_n12074_));
  NAND3X1  g11882(.A(new_n12067_), .B(new_n12058_), .C(new_n5941_), .Y(new_n12075_));
  AOI21X1  g11883(.A0(new_n12075_), .A1(new_n12074_), .B0(new_n12068_), .Y(new_n12076_));
  OR2X1    g11884(.A(new_n12076_), .B(new_n5541_), .Y(new_n12077_));
  AND2X1   g11885(.A(new_n12075_), .B(new_n12074_), .Y(new_n12078_));
  AND2X1   g11886(.A(new_n11564_), .B(new_n11562_), .Y(new_n12079_));
  NOR3X1   g11887(.A(new_n12079_), .B(new_n11530_), .C(new_n11563_), .Y(new_n12080_));
  NOR3X1   g11888(.A(new_n11896_), .B(new_n12079_), .C(new_n11563_), .Y(new_n12081_));
  NOR2X1   g11889(.A(new_n12081_), .B(new_n11529_), .Y(new_n12082_));
  AOI21X1  g11890(.A0(new_n12080_), .A1(\asqrt[21] ), .B0(new_n12082_), .Y(new_n12083_));
  INVX1    g11891(.A(new_n12083_), .Y(new_n12084_));
  OR2X1    g11892(.A(new_n12065_), .B(new_n6699_), .Y(new_n12085_));
  AND2X1   g11893(.A(new_n12049_), .B(new_n12040_), .Y(new_n12086_));
  INVX1    g11894(.A(new_n12055_), .Y(new_n12087_));
  NAND2X1  g11895(.A(new_n12031_), .B(new_n6699_), .Y(new_n12088_));
  OAI21X1  g11896(.A0(new_n12088_), .A1(new_n12086_), .B0(new_n12087_), .Y(new_n12089_));
  AOI21X1  g11897(.A0(new_n12089_), .A1(new_n12085_), .B0(new_n6294_), .Y(new_n12090_));
  AOI21X1  g11898(.A0(new_n12038_), .A1(\asqrt[32] ), .B0(\asqrt[33] ), .Y(new_n12091_));
  AOI21X1  g11899(.A0(new_n12091_), .A1(new_n12089_), .B0(new_n12062_), .Y(new_n12092_));
  OAI21X1  g11900(.A0(new_n12092_), .A1(new_n12090_), .B0(\asqrt[34] ), .Y(new_n12093_));
  NAND2X1  g11901(.A(new_n12093_), .B(new_n5541_), .Y(new_n12094_));
  OAI21X1  g11902(.A0(new_n12094_), .A1(new_n12078_), .B0(new_n12084_), .Y(new_n12095_));
  AOI21X1  g11903(.A0(new_n12095_), .A1(new_n12077_), .B0(new_n5176_), .Y(new_n12096_));
  NAND4X1  g11904(.A(\asqrt[21] ), .B(new_n11541_), .C(new_n11539_), .D(new_n11566_), .Y(new_n12097_));
  NAND2X1  g11905(.A(new_n11541_), .B(new_n11566_), .Y(new_n12098_));
  OAI21X1  g11906(.A0(new_n12098_), .A1(new_n11896_), .B0(new_n11540_), .Y(new_n12099_));
  AND2X1   g11907(.A(new_n12099_), .B(new_n12097_), .Y(new_n12100_));
  NOR3X1   g11908(.A(new_n12092_), .B(new_n12090_), .C(\asqrt[34] ), .Y(new_n12101_));
  OAI21X1  g11909(.A0(new_n12101_), .A1(new_n12073_), .B0(new_n12093_), .Y(new_n12102_));
  AOI21X1  g11910(.A0(new_n12102_), .A1(\asqrt[35] ), .B0(\asqrt[36] ), .Y(new_n12103_));
  AOI21X1  g11911(.A0(new_n12103_), .A1(new_n12095_), .B0(new_n12100_), .Y(new_n12104_));
  OAI21X1  g11912(.A0(new_n12104_), .A1(new_n12096_), .B0(\asqrt[37] ), .Y(new_n12105_));
  AOI21X1  g11913(.A0(new_n11587_), .A1(new_n11586_), .B0(new_n11549_), .Y(new_n12106_));
  AND2X1   g11914(.A(new_n12106_), .B(new_n11543_), .Y(new_n12107_));
  AOI22X1  g11915(.A0(new_n11587_), .A1(new_n11586_), .B0(new_n11568_), .B1(\asqrt[36] ), .Y(new_n12108_));
  AOI21X1  g11916(.A0(new_n12108_), .A1(\asqrt[21] ), .B0(new_n11548_), .Y(new_n12109_));
  AOI21X1  g11917(.A0(new_n12107_), .A1(\asqrt[21] ), .B0(new_n12109_), .Y(new_n12110_));
  NOR3X1   g11918(.A(new_n12104_), .B(new_n12096_), .C(\asqrt[37] ), .Y(new_n12111_));
  OAI21X1  g11919(.A0(new_n12111_), .A1(new_n12110_), .B0(new_n12105_), .Y(new_n12112_));
  AND2X1   g11920(.A(new_n12112_), .B(\asqrt[38] ), .Y(new_n12113_));
  INVX1    g11921(.A(new_n12110_), .Y(new_n12114_));
  AND2X1   g11922(.A(new_n12102_), .B(\asqrt[35] ), .Y(new_n12115_));
  NAND2X1  g11923(.A(new_n12075_), .B(new_n12074_), .Y(new_n12116_));
  AND2X1   g11924(.A(new_n12093_), .B(new_n5541_), .Y(new_n12117_));
  AOI21X1  g11925(.A0(new_n12117_), .A1(new_n12116_), .B0(new_n12083_), .Y(new_n12118_));
  OAI21X1  g11926(.A0(new_n12118_), .A1(new_n12115_), .B0(\asqrt[36] ), .Y(new_n12119_));
  INVX1    g11927(.A(new_n12100_), .Y(new_n12120_));
  OAI21X1  g11928(.A0(new_n12076_), .A1(new_n5541_), .B0(new_n5176_), .Y(new_n12121_));
  OAI21X1  g11929(.A0(new_n12121_), .A1(new_n12118_), .B0(new_n12120_), .Y(new_n12122_));
  NAND3X1  g11930(.A(new_n12122_), .B(new_n12119_), .C(new_n4826_), .Y(new_n12123_));
  NAND2X1  g11931(.A(new_n12123_), .B(new_n12114_), .Y(new_n12124_));
  AND2X1   g11932(.A(new_n11569_), .B(new_n11551_), .Y(new_n12125_));
  NOR3X1   g11933(.A(new_n12125_), .B(new_n11590_), .C(new_n11552_), .Y(new_n12126_));
  NOR3X1   g11934(.A(new_n11896_), .B(new_n12125_), .C(new_n11552_), .Y(new_n12127_));
  NOR2X1   g11935(.A(new_n12127_), .B(new_n11557_), .Y(new_n12128_));
  AOI21X1  g11936(.A0(new_n12126_), .A1(\asqrt[21] ), .B0(new_n12128_), .Y(new_n12129_));
  AND2X1   g11937(.A(new_n12105_), .B(new_n4493_), .Y(new_n12130_));
  AOI21X1  g11938(.A0(new_n12130_), .A1(new_n12124_), .B0(new_n12129_), .Y(new_n12131_));
  OAI21X1  g11939(.A0(new_n12131_), .A1(new_n12113_), .B0(\asqrt[39] ), .Y(new_n12132_));
  NAND4X1  g11940(.A(\asqrt[21] ), .B(new_n11604_), .C(new_n11576_), .D(new_n11571_), .Y(new_n12133_));
  NAND2X1  g11941(.A(new_n11604_), .B(new_n11571_), .Y(new_n12134_));
  OAI21X1  g11942(.A0(new_n12134_), .A1(new_n11896_), .B0(new_n11603_), .Y(new_n12135_));
  AND2X1   g11943(.A(new_n12135_), .B(new_n12133_), .Y(new_n12136_));
  INVX1    g11944(.A(new_n12136_), .Y(new_n12137_));
  AOI21X1  g11945(.A0(new_n12122_), .A1(new_n12119_), .B0(new_n4826_), .Y(new_n12138_));
  AOI21X1  g11946(.A0(new_n12123_), .A1(new_n12114_), .B0(new_n12138_), .Y(new_n12139_));
  OAI21X1  g11947(.A0(new_n12139_), .A1(new_n4493_), .B0(new_n4165_), .Y(new_n12140_));
  OAI21X1  g11948(.A0(new_n12140_), .A1(new_n12131_), .B0(new_n12137_), .Y(new_n12141_));
  AOI21X1  g11949(.A0(new_n12141_), .A1(new_n12132_), .B0(new_n3863_), .Y(new_n12142_));
  AND2X1   g11950(.A(new_n11594_), .B(new_n11580_), .Y(new_n12143_));
  NOR3X1   g11951(.A(new_n12143_), .B(new_n11629_), .C(new_n11579_), .Y(new_n12144_));
  NOR3X1   g11952(.A(new_n11896_), .B(new_n12143_), .C(new_n11579_), .Y(new_n12145_));
  NOR2X1   g11953(.A(new_n12145_), .B(new_n11584_), .Y(new_n12146_));
  AOI21X1  g11954(.A0(new_n12144_), .A1(\asqrt[21] ), .B0(new_n12146_), .Y(new_n12147_));
  INVX1    g11955(.A(new_n12147_), .Y(new_n12148_));
  NAND3X1  g11956(.A(new_n12141_), .B(new_n12132_), .C(new_n3863_), .Y(new_n12149_));
  AOI21X1  g11957(.A0(new_n12149_), .A1(new_n12148_), .B0(new_n12142_), .Y(new_n12150_));
  OR2X1    g11958(.A(new_n12150_), .B(new_n3564_), .Y(new_n12151_));
  AND2X1   g11959(.A(new_n12149_), .B(new_n12148_), .Y(new_n12152_));
  AND2X1   g11960(.A(new_n11633_), .B(new_n11631_), .Y(new_n12153_));
  NOR3X1   g11961(.A(new_n12153_), .B(new_n11602_), .C(new_n11632_), .Y(new_n12154_));
  NOR3X1   g11962(.A(new_n11896_), .B(new_n12153_), .C(new_n11632_), .Y(new_n12155_));
  NOR2X1   g11963(.A(new_n12155_), .B(new_n11601_), .Y(new_n12156_));
  AOI21X1  g11964(.A0(new_n12154_), .A1(\asqrt[21] ), .B0(new_n12156_), .Y(new_n12157_));
  INVX1    g11965(.A(new_n12157_), .Y(new_n12158_));
  OR2X1    g11966(.A(new_n12139_), .B(new_n4493_), .Y(new_n12159_));
  AND2X1   g11967(.A(new_n12123_), .B(new_n12114_), .Y(new_n12160_));
  INVX1    g11968(.A(new_n12129_), .Y(new_n12161_));
  NAND2X1  g11969(.A(new_n12105_), .B(new_n4493_), .Y(new_n12162_));
  OAI21X1  g11970(.A0(new_n12162_), .A1(new_n12160_), .B0(new_n12161_), .Y(new_n12163_));
  AOI21X1  g11971(.A0(new_n12163_), .A1(new_n12159_), .B0(new_n4165_), .Y(new_n12164_));
  AOI21X1  g11972(.A0(new_n12112_), .A1(\asqrt[38] ), .B0(\asqrt[39] ), .Y(new_n12165_));
  AOI21X1  g11973(.A0(new_n12165_), .A1(new_n12163_), .B0(new_n12136_), .Y(new_n12166_));
  OAI21X1  g11974(.A0(new_n12166_), .A1(new_n12164_), .B0(\asqrt[40] ), .Y(new_n12167_));
  NAND2X1  g11975(.A(new_n12167_), .B(new_n3564_), .Y(new_n12168_));
  OAI21X1  g11976(.A0(new_n12168_), .A1(new_n12152_), .B0(new_n12158_), .Y(new_n12169_));
  AOI21X1  g11977(.A0(new_n12169_), .A1(new_n12151_), .B0(new_n3276_), .Y(new_n12170_));
  NAND4X1  g11978(.A(\asqrt[21] ), .B(new_n11615_), .C(new_n11613_), .D(new_n11635_), .Y(new_n12171_));
  NAND2X1  g11979(.A(new_n11615_), .B(new_n11635_), .Y(new_n12172_));
  OAI21X1  g11980(.A0(new_n12172_), .A1(new_n11896_), .B0(new_n11614_), .Y(new_n12173_));
  AND2X1   g11981(.A(new_n12173_), .B(new_n12171_), .Y(new_n12174_));
  NOR3X1   g11982(.A(new_n12166_), .B(new_n12164_), .C(\asqrt[40] ), .Y(new_n12175_));
  OAI21X1  g11983(.A0(new_n12175_), .A1(new_n12147_), .B0(new_n12167_), .Y(new_n12176_));
  AOI21X1  g11984(.A0(new_n12176_), .A1(\asqrt[41] ), .B0(\asqrt[42] ), .Y(new_n12177_));
  AOI21X1  g11985(.A0(new_n12177_), .A1(new_n12169_), .B0(new_n12174_), .Y(new_n12178_));
  OAI21X1  g11986(.A0(new_n12178_), .A1(new_n12170_), .B0(\asqrt[43] ), .Y(new_n12179_));
  AOI21X1  g11987(.A0(new_n11670_), .A1(new_n11669_), .B0(new_n11623_), .Y(new_n12180_));
  AND2X1   g11988(.A(new_n12180_), .B(new_n11617_), .Y(new_n12181_));
  AOI22X1  g11989(.A0(new_n11670_), .A1(new_n11669_), .B0(new_n11637_), .B1(\asqrt[42] ), .Y(new_n12182_));
  AOI21X1  g11990(.A0(new_n12182_), .A1(\asqrt[21] ), .B0(new_n11622_), .Y(new_n12183_));
  AOI21X1  g11991(.A0(new_n12181_), .A1(\asqrt[21] ), .B0(new_n12183_), .Y(new_n12184_));
  NOR3X1   g11992(.A(new_n12178_), .B(new_n12170_), .C(\asqrt[43] ), .Y(new_n12185_));
  OAI21X1  g11993(.A0(new_n12185_), .A1(new_n12184_), .B0(new_n12179_), .Y(new_n12186_));
  AND2X1   g11994(.A(new_n12186_), .B(\asqrt[44] ), .Y(new_n12187_));
  INVX1    g11995(.A(new_n12184_), .Y(new_n12188_));
  AND2X1   g11996(.A(new_n12176_), .B(\asqrt[41] ), .Y(new_n12189_));
  NAND2X1  g11997(.A(new_n12149_), .B(new_n12148_), .Y(new_n12190_));
  AND2X1   g11998(.A(new_n12167_), .B(new_n3564_), .Y(new_n12191_));
  AOI21X1  g11999(.A0(new_n12191_), .A1(new_n12190_), .B0(new_n12157_), .Y(new_n12192_));
  OAI21X1  g12000(.A0(new_n12192_), .A1(new_n12189_), .B0(\asqrt[42] ), .Y(new_n12193_));
  INVX1    g12001(.A(new_n12174_), .Y(new_n12194_));
  OAI21X1  g12002(.A0(new_n12150_), .A1(new_n3564_), .B0(new_n3276_), .Y(new_n12195_));
  OAI21X1  g12003(.A0(new_n12195_), .A1(new_n12192_), .B0(new_n12194_), .Y(new_n12196_));
  NAND3X1  g12004(.A(new_n12196_), .B(new_n12193_), .C(new_n3008_), .Y(new_n12197_));
  NAND2X1  g12005(.A(new_n12197_), .B(new_n12188_), .Y(new_n12198_));
  AND2X1   g12006(.A(new_n12179_), .B(new_n2769_), .Y(new_n12199_));
  AND2X1   g12007(.A(new_n11638_), .B(new_n11625_), .Y(new_n12200_));
  NOR3X1   g12008(.A(new_n11674_), .B(new_n12200_), .C(new_n11626_), .Y(new_n12201_));
  NOR3X1   g12009(.A(new_n11896_), .B(new_n12200_), .C(new_n11626_), .Y(new_n12202_));
  NOR2X1   g12010(.A(new_n12202_), .B(new_n11643_), .Y(new_n12203_));
  AOI21X1  g12011(.A0(new_n12201_), .A1(\asqrt[21] ), .B0(new_n12203_), .Y(new_n12204_));
  AOI21X1  g12012(.A0(new_n12199_), .A1(new_n12198_), .B0(new_n12204_), .Y(new_n12205_));
  OAI21X1  g12013(.A0(new_n12205_), .A1(new_n12187_), .B0(\asqrt[45] ), .Y(new_n12206_));
  NAND4X1  g12014(.A(\asqrt[21] ), .B(new_n11678_), .C(new_n11650_), .D(new_n11645_), .Y(new_n12207_));
  OR2X1    g12015(.A(new_n11651_), .B(new_n11676_), .Y(new_n12208_));
  OAI21X1  g12016(.A0(new_n12208_), .A1(new_n11896_), .B0(new_n11677_), .Y(new_n12209_));
  AND2X1   g12017(.A(new_n12209_), .B(new_n12207_), .Y(new_n12210_));
  INVX1    g12018(.A(new_n12210_), .Y(new_n12211_));
  AOI21X1  g12019(.A0(new_n12196_), .A1(new_n12193_), .B0(new_n3008_), .Y(new_n12212_));
  AOI21X1  g12020(.A0(new_n12197_), .A1(new_n12188_), .B0(new_n12212_), .Y(new_n12213_));
  OAI21X1  g12021(.A0(new_n12213_), .A1(new_n2769_), .B0(new_n2570_), .Y(new_n12214_));
  OAI21X1  g12022(.A0(new_n12214_), .A1(new_n12205_), .B0(new_n12211_), .Y(new_n12215_));
  AOI21X1  g12023(.A0(new_n12215_), .A1(new_n12206_), .B0(new_n2263_), .Y(new_n12216_));
  AND2X1   g12024(.A(new_n11659_), .B(new_n11654_), .Y(new_n12217_));
  NOR3X1   g12025(.A(new_n12217_), .B(new_n11694_), .C(new_n11653_), .Y(new_n12218_));
  NOR3X1   g12026(.A(new_n11896_), .B(new_n12217_), .C(new_n11653_), .Y(new_n12219_));
  NOR2X1   g12027(.A(new_n12219_), .B(new_n11658_), .Y(new_n12220_));
  AOI21X1  g12028(.A0(new_n12218_), .A1(\asqrt[21] ), .B0(new_n12220_), .Y(new_n12221_));
  INVX1    g12029(.A(new_n12221_), .Y(new_n12222_));
  NAND3X1  g12030(.A(new_n12215_), .B(new_n12206_), .C(new_n2263_), .Y(new_n12223_));
  AOI21X1  g12031(.A0(new_n12223_), .A1(new_n12222_), .B0(new_n12216_), .Y(new_n12224_));
  OR2X1    g12032(.A(new_n12224_), .B(new_n2040_), .Y(new_n12225_));
  AND2X1   g12033(.A(new_n12223_), .B(new_n12222_), .Y(new_n12226_));
  AND2X1   g12034(.A(new_n11698_), .B(new_n11696_), .Y(new_n12227_));
  NOR3X1   g12035(.A(new_n12227_), .B(new_n11667_), .C(new_n11697_), .Y(new_n12228_));
  NOR3X1   g12036(.A(new_n11896_), .B(new_n12227_), .C(new_n11697_), .Y(new_n12229_));
  NOR2X1   g12037(.A(new_n12229_), .B(new_n11666_), .Y(new_n12230_));
  AOI21X1  g12038(.A0(new_n12228_), .A1(\asqrt[21] ), .B0(new_n12230_), .Y(new_n12231_));
  INVX1    g12039(.A(new_n12231_), .Y(new_n12232_));
  OR2X1    g12040(.A(new_n12213_), .B(new_n2769_), .Y(new_n12233_));
  AND2X1   g12041(.A(new_n12197_), .B(new_n12188_), .Y(new_n12234_));
  NAND2X1  g12042(.A(new_n12179_), .B(new_n2769_), .Y(new_n12235_));
  INVX1    g12043(.A(new_n12204_), .Y(new_n12236_));
  OAI21X1  g12044(.A0(new_n12235_), .A1(new_n12234_), .B0(new_n12236_), .Y(new_n12237_));
  AOI21X1  g12045(.A0(new_n12237_), .A1(new_n12233_), .B0(new_n2570_), .Y(new_n12238_));
  AOI21X1  g12046(.A0(new_n12186_), .A1(\asqrt[44] ), .B0(\asqrt[45] ), .Y(new_n12239_));
  AOI21X1  g12047(.A0(new_n12239_), .A1(new_n12237_), .B0(new_n12210_), .Y(new_n12240_));
  OAI21X1  g12048(.A0(new_n12240_), .A1(new_n12238_), .B0(\asqrt[46] ), .Y(new_n12241_));
  NAND2X1  g12049(.A(new_n12241_), .B(new_n2040_), .Y(new_n12242_));
  OAI21X1  g12050(.A0(new_n12242_), .A1(new_n12226_), .B0(new_n12232_), .Y(new_n12243_));
  AOI21X1  g12051(.A0(new_n12243_), .A1(new_n12225_), .B0(new_n1834_), .Y(new_n12244_));
  OR4X1    g12052(.A(new_n11896_), .B(new_n11700_), .C(new_n11688_), .D(new_n11682_), .Y(new_n12245_));
  OR2X1    g12053(.A(new_n11700_), .B(new_n11682_), .Y(new_n12246_));
  OAI21X1  g12054(.A0(new_n12246_), .A1(new_n11896_), .B0(new_n11688_), .Y(new_n12247_));
  AND2X1   g12055(.A(new_n12247_), .B(new_n12245_), .Y(new_n12248_));
  NOR3X1   g12056(.A(new_n12240_), .B(new_n12238_), .C(\asqrt[46] ), .Y(new_n12249_));
  OAI21X1  g12057(.A0(new_n12249_), .A1(new_n12221_), .B0(new_n12241_), .Y(new_n12250_));
  AOI21X1  g12058(.A0(new_n12250_), .A1(\asqrt[47] ), .B0(\asqrt[48] ), .Y(new_n12251_));
  AOI21X1  g12059(.A0(new_n12251_), .A1(new_n12243_), .B0(new_n12248_), .Y(new_n12252_));
  OAI21X1  g12060(.A0(new_n12252_), .A1(new_n12244_), .B0(\asqrt[49] ), .Y(new_n12253_));
  AOI21X1  g12061(.A0(new_n11744_), .A1(new_n11743_), .B0(new_n11706_), .Y(new_n12254_));
  AND2X1   g12062(.A(new_n12254_), .B(new_n11691_), .Y(new_n12255_));
  AOI22X1  g12063(.A0(new_n11744_), .A1(new_n11743_), .B0(new_n11716_), .B1(\asqrt[48] ), .Y(new_n12256_));
  AOI21X1  g12064(.A0(new_n12256_), .A1(\asqrt[21] ), .B0(new_n11705_), .Y(new_n12257_));
  AOI21X1  g12065(.A0(new_n12255_), .A1(\asqrt[21] ), .B0(new_n12257_), .Y(new_n12258_));
  NOR3X1   g12066(.A(new_n12252_), .B(new_n12244_), .C(\asqrt[49] ), .Y(new_n12259_));
  OAI21X1  g12067(.A0(new_n12259_), .A1(new_n12258_), .B0(new_n12253_), .Y(new_n12260_));
  AND2X1   g12068(.A(new_n12260_), .B(\asqrt[50] ), .Y(new_n12261_));
  INVX1    g12069(.A(new_n12258_), .Y(new_n12262_));
  AND2X1   g12070(.A(new_n12250_), .B(\asqrt[47] ), .Y(new_n12263_));
  NAND2X1  g12071(.A(new_n12223_), .B(new_n12222_), .Y(new_n12264_));
  AND2X1   g12072(.A(new_n12241_), .B(new_n2040_), .Y(new_n12265_));
  AOI21X1  g12073(.A0(new_n12265_), .A1(new_n12264_), .B0(new_n12231_), .Y(new_n12266_));
  OAI21X1  g12074(.A0(new_n12266_), .A1(new_n12263_), .B0(\asqrt[48] ), .Y(new_n12267_));
  INVX1    g12075(.A(new_n12248_), .Y(new_n12268_));
  OAI21X1  g12076(.A0(new_n12224_), .A1(new_n2040_), .B0(new_n1834_), .Y(new_n12269_));
  OAI21X1  g12077(.A0(new_n12269_), .A1(new_n12266_), .B0(new_n12268_), .Y(new_n12270_));
  NAND3X1  g12078(.A(new_n12270_), .B(new_n12267_), .C(new_n1632_), .Y(new_n12271_));
  NAND2X1  g12079(.A(new_n12271_), .B(new_n12262_), .Y(new_n12272_));
  AND2X1   g12080(.A(new_n11717_), .B(new_n11709_), .Y(new_n12273_));
  NOR3X1   g12081(.A(new_n12273_), .B(new_n11747_), .C(new_n11710_), .Y(new_n12274_));
  NOR3X1   g12082(.A(new_n11896_), .B(new_n12273_), .C(new_n11710_), .Y(new_n12275_));
  NOR2X1   g12083(.A(new_n12275_), .B(new_n11715_), .Y(new_n12276_));
  AOI21X1  g12084(.A0(new_n12274_), .A1(\asqrt[21] ), .B0(new_n12276_), .Y(new_n12277_));
  AND2X1   g12085(.A(new_n12253_), .B(new_n1469_), .Y(new_n12278_));
  AOI21X1  g12086(.A0(new_n12278_), .A1(new_n12272_), .B0(new_n12277_), .Y(new_n12279_));
  OAI21X1  g12087(.A0(new_n12279_), .A1(new_n12261_), .B0(\asqrt[51] ), .Y(new_n12280_));
  OR4X1    g12088(.A(new_n11896_), .B(new_n11725_), .C(new_n11751_), .D(new_n11750_), .Y(new_n12281_));
  OR2X1    g12089(.A(new_n11725_), .B(new_n11750_), .Y(new_n12282_));
  OAI21X1  g12090(.A0(new_n12282_), .A1(new_n11896_), .B0(new_n11751_), .Y(new_n12283_));
  AND2X1   g12091(.A(new_n12283_), .B(new_n12281_), .Y(new_n12284_));
  INVX1    g12092(.A(new_n12284_), .Y(new_n12285_));
  AOI21X1  g12093(.A0(new_n12270_), .A1(new_n12267_), .B0(new_n1632_), .Y(new_n12286_));
  AOI21X1  g12094(.A0(new_n12271_), .A1(new_n12262_), .B0(new_n12286_), .Y(new_n12287_));
  OAI21X1  g12095(.A0(new_n12287_), .A1(new_n1469_), .B0(new_n1277_), .Y(new_n12288_));
  OAI21X1  g12096(.A0(new_n12288_), .A1(new_n12279_), .B0(new_n12285_), .Y(new_n12289_));
  AOI21X1  g12097(.A0(new_n12289_), .A1(new_n12280_), .B0(new_n1111_), .Y(new_n12290_));
  AND2X1   g12098(.A(new_n11733_), .B(new_n11728_), .Y(new_n12291_));
  NOR3X1   g12099(.A(new_n12291_), .B(new_n11768_), .C(new_n11727_), .Y(new_n12292_));
  NOR3X1   g12100(.A(new_n11896_), .B(new_n12291_), .C(new_n11727_), .Y(new_n12293_));
  NOR2X1   g12101(.A(new_n12293_), .B(new_n11732_), .Y(new_n12294_));
  AOI21X1  g12102(.A0(new_n12292_), .A1(\asqrt[21] ), .B0(new_n12294_), .Y(new_n12295_));
  INVX1    g12103(.A(new_n12295_), .Y(new_n12296_));
  NAND3X1  g12104(.A(new_n12289_), .B(new_n12280_), .C(new_n1111_), .Y(new_n12297_));
  AOI21X1  g12105(.A0(new_n12297_), .A1(new_n12296_), .B0(new_n12290_), .Y(new_n12298_));
  OR2X1    g12106(.A(new_n12298_), .B(new_n968_), .Y(new_n12299_));
  OR2X1    g12107(.A(new_n12287_), .B(new_n1469_), .Y(new_n12300_));
  AND2X1   g12108(.A(new_n12271_), .B(new_n12262_), .Y(new_n12301_));
  INVX1    g12109(.A(new_n12277_), .Y(new_n12302_));
  NAND2X1  g12110(.A(new_n12253_), .B(new_n1469_), .Y(new_n12303_));
  OAI21X1  g12111(.A0(new_n12303_), .A1(new_n12301_), .B0(new_n12302_), .Y(new_n12304_));
  AOI21X1  g12112(.A0(new_n12304_), .A1(new_n12300_), .B0(new_n1277_), .Y(new_n12305_));
  AOI21X1  g12113(.A0(new_n12260_), .A1(\asqrt[50] ), .B0(\asqrt[51] ), .Y(new_n12306_));
  AOI21X1  g12114(.A0(new_n12306_), .A1(new_n12304_), .B0(new_n12284_), .Y(new_n12307_));
  NOR3X1   g12115(.A(new_n12307_), .B(new_n12305_), .C(\asqrt[52] ), .Y(new_n12308_));
  NOR2X1   g12116(.A(new_n12308_), .B(new_n12295_), .Y(new_n12309_));
  AND2X1   g12117(.A(new_n11772_), .B(new_n11770_), .Y(new_n12310_));
  NOR3X1   g12118(.A(new_n12310_), .B(new_n11741_), .C(new_n11771_), .Y(new_n12311_));
  NOR3X1   g12119(.A(new_n11896_), .B(new_n12310_), .C(new_n11771_), .Y(new_n12312_));
  NOR2X1   g12120(.A(new_n12312_), .B(new_n11740_), .Y(new_n12313_));
  AOI21X1  g12121(.A0(new_n12311_), .A1(\asqrt[21] ), .B0(new_n12313_), .Y(new_n12314_));
  INVX1    g12122(.A(new_n12314_), .Y(new_n12315_));
  OAI21X1  g12123(.A0(new_n12307_), .A1(new_n12305_), .B0(\asqrt[52] ), .Y(new_n12316_));
  NAND2X1  g12124(.A(new_n12316_), .B(new_n968_), .Y(new_n12317_));
  OAI21X1  g12125(.A0(new_n12317_), .A1(new_n12309_), .B0(new_n12315_), .Y(new_n12318_));
  AOI21X1  g12126(.A0(new_n12318_), .A1(new_n12299_), .B0(new_n902_), .Y(new_n12319_));
  OR4X1    g12127(.A(new_n11896_), .B(new_n11774_), .C(new_n11762_), .D(new_n11756_), .Y(new_n12320_));
  OR2X1    g12128(.A(new_n11774_), .B(new_n11756_), .Y(new_n12321_));
  OAI21X1  g12129(.A0(new_n12321_), .A1(new_n11896_), .B0(new_n11762_), .Y(new_n12322_));
  AND2X1   g12130(.A(new_n12322_), .B(new_n12320_), .Y(new_n12323_));
  OAI21X1  g12131(.A0(new_n12308_), .A1(new_n12295_), .B0(new_n12316_), .Y(new_n12324_));
  AOI21X1  g12132(.A0(new_n12324_), .A1(\asqrt[53] ), .B0(\asqrt[54] ), .Y(new_n12325_));
  AOI21X1  g12133(.A0(new_n12325_), .A1(new_n12318_), .B0(new_n12323_), .Y(new_n12326_));
  OAI21X1  g12134(.A0(new_n12326_), .A1(new_n12319_), .B0(\asqrt[55] ), .Y(new_n12327_));
  AOI21X1  g12135(.A0(new_n11818_), .A1(new_n11817_), .B0(new_n11780_), .Y(new_n12328_));
  AND2X1   g12136(.A(new_n12328_), .B(new_n11765_), .Y(new_n12329_));
  AOI22X1  g12137(.A0(new_n11818_), .A1(new_n11817_), .B0(new_n11790_), .B1(\asqrt[54] ), .Y(new_n12330_));
  AOI21X1  g12138(.A0(new_n12330_), .A1(\asqrt[21] ), .B0(new_n11779_), .Y(new_n12331_));
  AOI21X1  g12139(.A0(new_n12329_), .A1(\asqrt[21] ), .B0(new_n12331_), .Y(new_n12332_));
  NOR3X1   g12140(.A(new_n12326_), .B(new_n12319_), .C(\asqrt[55] ), .Y(new_n12333_));
  OAI21X1  g12141(.A0(new_n12333_), .A1(new_n12332_), .B0(new_n12327_), .Y(new_n12334_));
  AND2X1   g12142(.A(new_n12334_), .B(\asqrt[56] ), .Y(new_n12335_));
  OR2X1    g12143(.A(new_n12333_), .B(new_n12332_), .Y(new_n12336_));
  AND2X1   g12144(.A(new_n11791_), .B(new_n11783_), .Y(new_n12337_));
  NOR3X1   g12145(.A(new_n12337_), .B(new_n11821_), .C(new_n11784_), .Y(new_n12338_));
  NOR3X1   g12146(.A(new_n11896_), .B(new_n12337_), .C(new_n11784_), .Y(new_n12339_));
  NOR2X1   g12147(.A(new_n12339_), .B(new_n11789_), .Y(new_n12340_));
  AOI21X1  g12148(.A0(new_n12338_), .A1(\asqrt[21] ), .B0(new_n12340_), .Y(new_n12341_));
  AND2X1   g12149(.A(new_n12327_), .B(new_n582_), .Y(new_n12342_));
  AOI21X1  g12150(.A0(new_n12342_), .A1(new_n12336_), .B0(new_n12341_), .Y(new_n12343_));
  OAI21X1  g12151(.A0(new_n12343_), .A1(new_n12335_), .B0(\asqrt[57] ), .Y(new_n12344_));
  OR4X1    g12152(.A(new_n11896_), .B(new_n11799_), .C(new_n11825_), .D(new_n11824_), .Y(new_n12345_));
  OR2X1    g12153(.A(new_n11799_), .B(new_n11824_), .Y(new_n12346_));
  OAI21X1  g12154(.A0(new_n12346_), .A1(new_n11896_), .B0(new_n11825_), .Y(new_n12347_));
  AND2X1   g12155(.A(new_n12347_), .B(new_n12345_), .Y(new_n12348_));
  INVX1    g12156(.A(new_n12348_), .Y(new_n12349_));
  AND2X1   g12157(.A(new_n12324_), .B(\asqrt[53] ), .Y(new_n12350_));
  OR2X1    g12158(.A(new_n12308_), .B(new_n12295_), .Y(new_n12351_));
  AND2X1   g12159(.A(new_n12316_), .B(new_n968_), .Y(new_n12352_));
  AOI21X1  g12160(.A0(new_n12352_), .A1(new_n12351_), .B0(new_n12314_), .Y(new_n12353_));
  OAI21X1  g12161(.A0(new_n12353_), .A1(new_n12350_), .B0(\asqrt[54] ), .Y(new_n12354_));
  INVX1    g12162(.A(new_n12323_), .Y(new_n12355_));
  OAI21X1  g12163(.A0(new_n12298_), .A1(new_n968_), .B0(new_n902_), .Y(new_n12356_));
  OAI21X1  g12164(.A0(new_n12356_), .A1(new_n12353_), .B0(new_n12355_), .Y(new_n12357_));
  AOI21X1  g12165(.A0(new_n12357_), .A1(new_n12354_), .B0(new_n697_), .Y(new_n12358_));
  INVX1    g12166(.A(new_n12332_), .Y(new_n12359_));
  NAND3X1  g12167(.A(new_n12357_), .B(new_n12354_), .C(new_n697_), .Y(new_n12360_));
  AOI21X1  g12168(.A0(new_n12360_), .A1(new_n12359_), .B0(new_n12358_), .Y(new_n12361_));
  OAI21X1  g12169(.A0(new_n12361_), .A1(new_n582_), .B0(new_n481_), .Y(new_n12362_));
  OAI21X1  g12170(.A0(new_n12362_), .A1(new_n12343_), .B0(new_n12349_), .Y(new_n12363_));
  AOI21X1  g12171(.A0(new_n12363_), .A1(new_n12344_), .B0(new_n399_), .Y(new_n12364_));
  AND2X1   g12172(.A(new_n11807_), .B(new_n11802_), .Y(new_n12365_));
  NOR3X1   g12173(.A(new_n12365_), .B(new_n11842_), .C(new_n11801_), .Y(new_n12366_));
  NOR3X1   g12174(.A(new_n11896_), .B(new_n12365_), .C(new_n11801_), .Y(new_n12367_));
  NOR2X1   g12175(.A(new_n12367_), .B(new_n11806_), .Y(new_n12368_));
  AOI21X1  g12176(.A0(new_n12366_), .A1(\asqrt[21] ), .B0(new_n12368_), .Y(new_n12369_));
  INVX1    g12177(.A(new_n12369_), .Y(new_n12370_));
  NAND3X1  g12178(.A(new_n12363_), .B(new_n12344_), .C(new_n399_), .Y(new_n12371_));
  AOI21X1  g12179(.A0(new_n12371_), .A1(new_n12370_), .B0(new_n12364_), .Y(new_n12372_));
  OR2X1    g12180(.A(new_n12372_), .B(new_n328_), .Y(new_n12373_));
  OR2X1    g12181(.A(new_n12361_), .B(new_n582_), .Y(new_n12374_));
  NOR2X1   g12182(.A(new_n12333_), .B(new_n12332_), .Y(new_n12375_));
  INVX1    g12183(.A(new_n12341_), .Y(new_n12376_));
  NAND2X1  g12184(.A(new_n12327_), .B(new_n582_), .Y(new_n12377_));
  OAI21X1  g12185(.A0(new_n12377_), .A1(new_n12375_), .B0(new_n12376_), .Y(new_n12378_));
  AOI21X1  g12186(.A0(new_n12378_), .A1(new_n12374_), .B0(new_n481_), .Y(new_n12379_));
  AOI21X1  g12187(.A0(new_n12334_), .A1(\asqrt[56] ), .B0(\asqrt[57] ), .Y(new_n12380_));
  AOI21X1  g12188(.A0(new_n12380_), .A1(new_n12378_), .B0(new_n12348_), .Y(new_n12381_));
  NOR3X1   g12189(.A(new_n12381_), .B(new_n12379_), .C(\asqrt[58] ), .Y(new_n12382_));
  NOR2X1   g12190(.A(new_n12382_), .B(new_n12369_), .Y(new_n12383_));
  AND2X1   g12191(.A(new_n11846_), .B(new_n11844_), .Y(new_n12384_));
  NOR3X1   g12192(.A(new_n12384_), .B(new_n11815_), .C(new_n11845_), .Y(new_n12385_));
  NOR3X1   g12193(.A(new_n11896_), .B(new_n12384_), .C(new_n11845_), .Y(new_n12386_));
  NOR2X1   g12194(.A(new_n12386_), .B(new_n11814_), .Y(new_n12387_));
  AOI21X1  g12195(.A0(new_n12385_), .A1(\asqrt[21] ), .B0(new_n12387_), .Y(new_n12388_));
  INVX1    g12196(.A(new_n12388_), .Y(new_n12389_));
  OAI21X1  g12197(.A0(new_n12381_), .A1(new_n12379_), .B0(\asqrt[58] ), .Y(new_n12390_));
  NAND2X1  g12198(.A(new_n12390_), .B(new_n328_), .Y(new_n12391_));
  OAI21X1  g12199(.A0(new_n12391_), .A1(new_n12383_), .B0(new_n12389_), .Y(new_n12392_));
  AOI21X1  g12200(.A0(new_n12392_), .A1(new_n12373_), .B0(new_n292_), .Y(new_n12393_));
  OR4X1    g12201(.A(new_n11896_), .B(new_n11848_), .C(new_n11836_), .D(new_n11830_), .Y(new_n12394_));
  OR2X1    g12202(.A(new_n11848_), .B(new_n11830_), .Y(new_n12395_));
  OAI21X1  g12203(.A0(new_n12395_), .A1(new_n11896_), .B0(new_n11836_), .Y(new_n12396_));
  AND2X1   g12204(.A(new_n12396_), .B(new_n12394_), .Y(new_n12397_));
  OAI21X1  g12205(.A0(new_n12382_), .A1(new_n12369_), .B0(new_n12390_), .Y(new_n12398_));
  AOI21X1  g12206(.A0(new_n12398_), .A1(\asqrt[59] ), .B0(\asqrt[60] ), .Y(new_n12399_));
  AOI21X1  g12207(.A0(new_n12399_), .A1(new_n12392_), .B0(new_n12397_), .Y(new_n12400_));
  OAI21X1  g12208(.A0(new_n12400_), .A1(new_n12393_), .B0(\asqrt[61] ), .Y(new_n12401_));
  AOI21X1  g12209(.A0(new_n11909_), .A1(new_n11908_), .B0(new_n11854_), .Y(new_n12402_));
  AND2X1   g12210(.A(new_n12402_), .B(new_n11839_), .Y(new_n12403_));
  AOI22X1  g12211(.A0(new_n11909_), .A1(new_n11908_), .B0(new_n11864_), .B1(\asqrt[60] ), .Y(new_n12404_));
  AOI21X1  g12212(.A0(new_n12404_), .A1(\asqrt[21] ), .B0(new_n11853_), .Y(new_n12405_));
  AOI21X1  g12213(.A0(new_n12403_), .A1(\asqrt[21] ), .B0(new_n12405_), .Y(new_n12406_));
  NOR3X1   g12214(.A(new_n12400_), .B(new_n12393_), .C(\asqrt[61] ), .Y(new_n12407_));
  OAI21X1  g12215(.A0(new_n12407_), .A1(new_n12406_), .B0(new_n12401_), .Y(new_n12408_));
  AND2X1   g12216(.A(new_n12408_), .B(\asqrt[62] ), .Y(new_n12409_));
  INVX1    g12217(.A(new_n12406_), .Y(new_n12410_));
  AND2X1   g12218(.A(new_n12398_), .B(\asqrt[59] ), .Y(new_n12411_));
  OR2X1    g12219(.A(new_n12382_), .B(new_n12369_), .Y(new_n12412_));
  AND2X1   g12220(.A(new_n12390_), .B(new_n328_), .Y(new_n12413_));
  AOI21X1  g12221(.A0(new_n12413_), .A1(new_n12412_), .B0(new_n12388_), .Y(new_n12414_));
  OAI21X1  g12222(.A0(new_n12414_), .A1(new_n12411_), .B0(\asqrt[60] ), .Y(new_n12415_));
  INVX1    g12223(.A(new_n12397_), .Y(new_n12416_));
  OAI21X1  g12224(.A0(new_n12372_), .A1(new_n328_), .B0(new_n292_), .Y(new_n12417_));
  OAI21X1  g12225(.A0(new_n12417_), .A1(new_n12414_), .B0(new_n12416_), .Y(new_n12418_));
  NAND3X1  g12226(.A(new_n12418_), .B(new_n12415_), .C(new_n217_), .Y(new_n12419_));
  NAND2X1  g12227(.A(new_n12419_), .B(new_n12410_), .Y(new_n12420_));
  AND2X1   g12228(.A(new_n11865_), .B(new_n11857_), .Y(new_n12421_));
  NOR3X1   g12229(.A(new_n12421_), .B(new_n11912_), .C(new_n11858_), .Y(new_n12422_));
  NOR3X1   g12230(.A(new_n11896_), .B(new_n12421_), .C(new_n11858_), .Y(new_n12423_));
  NOR2X1   g12231(.A(new_n12423_), .B(new_n11863_), .Y(new_n12424_));
  AOI21X1  g12232(.A0(new_n12422_), .A1(\asqrt[21] ), .B0(new_n12424_), .Y(new_n12425_));
  AND2X1   g12233(.A(new_n12401_), .B(new_n199_), .Y(new_n12426_));
  AOI21X1  g12234(.A0(new_n12426_), .A1(new_n12420_), .B0(new_n12425_), .Y(new_n12427_));
  NOR4X1   g12235(.A(new_n11896_), .B(new_n11873_), .C(new_n11916_), .D(new_n11915_), .Y(new_n12428_));
  NAND3X1  g12236(.A(\asqrt[21] ), .B(new_n11917_), .C(new_n11867_), .Y(new_n12429_));
  AOI21X1  g12237(.A0(new_n12429_), .A1(new_n11916_), .B0(new_n12428_), .Y(new_n12430_));
  INVX1    g12238(.A(new_n12430_), .Y(new_n12431_));
  NOR3X1   g12239(.A(new_n11896_), .B(new_n11878_), .C(new_n11918_), .Y(new_n12432_));
  AOI21X1  g12240(.A0(new_n11922_), .A1(new_n11921_), .B0(new_n12432_), .Y(new_n12433_));
  AND2X1   g12241(.A(new_n12433_), .B(new_n12431_), .Y(new_n12434_));
  OAI21X1  g12242(.A0(new_n12427_), .A1(new_n12409_), .B0(new_n12434_), .Y(new_n12435_));
  AOI21X1  g12243(.A0(new_n12418_), .A1(new_n12415_), .B0(new_n217_), .Y(new_n12436_));
  AOI21X1  g12244(.A0(new_n12419_), .A1(new_n12410_), .B0(new_n12436_), .Y(new_n12437_));
  OAI21X1  g12245(.A0(new_n12437_), .A1(new_n199_), .B0(new_n12430_), .Y(new_n12438_));
  AOI21X1  g12246(.A0(new_n11924_), .A1(new_n11920_), .B0(new_n11878_), .Y(new_n12439_));
  AOI21X1  g12247(.A0(new_n11879_), .A1(new_n11874_), .B0(new_n193_), .Y(new_n12440_));
  OAI21X1  g12248(.A0(new_n12439_), .A1(new_n11874_), .B0(new_n12440_), .Y(new_n12441_));
  OR2X1    g12249(.A(new_n11885_), .B(new_n11884_), .Y(new_n12442_));
  NOR4X1   g12250(.A(new_n11892_), .B(new_n11932_), .C(new_n11877_), .D(new_n11875_), .Y(new_n12443_));
  NAND3X1  g12251(.A(new_n12443_), .B(new_n12442_), .C(new_n11920_), .Y(new_n12444_));
  AND2X1   g12252(.A(new_n12444_), .B(new_n12441_), .Y(new_n12445_));
  OAI21X1  g12253(.A0(new_n12438_), .A1(new_n12427_), .B0(new_n12445_), .Y(new_n12446_));
  AOI21X1  g12254(.A0(new_n12435_), .A1(new_n193_), .B0(new_n12446_), .Y(new_n12447_));
  OR2X1    g12255(.A(new_n12437_), .B(new_n199_), .Y(new_n12448_));
  AND2X1   g12256(.A(new_n12419_), .B(new_n12410_), .Y(new_n12449_));
  INVX1    g12257(.A(new_n12425_), .Y(new_n12450_));
  NAND2X1  g12258(.A(new_n12401_), .B(new_n199_), .Y(new_n12451_));
  OAI21X1  g12259(.A0(new_n12451_), .A1(new_n12449_), .B0(new_n12450_), .Y(new_n12452_));
  INVX1    g12260(.A(new_n12434_), .Y(new_n12453_));
  AOI21X1  g12261(.A0(new_n12452_), .A1(new_n12448_), .B0(new_n12453_), .Y(new_n12454_));
  AOI21X1  g12262(.A0(new_n12408_), .A1(\asqrt[62] ), .B0(new_n12431_), .Y(new_n12455_));
  INVX1    g12263(.A(new_n12445_), .Y(new_n12456_));
  AOI21X1  g12264(.A0(new_n12455_), .A1(new_n12452_), .B0(new_n12456_), .Y(new_n12457_));
  OAI21X1  g12265(.A0(new_n12454_), .A1(\asqrt[63] ), .B0(new_n12457_), .Y(\asqrt[20] ));
  NOR2X1   g12266(.A(\a[39] ), .B(\a[38] ), .Y(new_n12459_));
  MX2X1    g12267(.A(new_n12459_), .B(\asqrt[20] ), .S0(\a[40] ), .Y(new_n12460_));
  AND2X1   g12268(.A(new_n12460_), .B(\asqrt[21] ), .Y(new_n12461_));
  NOR3X1   g12269(.A(\a[40] ), .B(\a[39] ), .C(\a[38] ), .Y(new_n12462_));
  NOR3X1   g12270(.A(new_n12462_), .B(new_n11892_), .C(new_n11932_), .Y(new_n12463_));
  NAND3X1  g12271(.A(new_n12463_), .B(new_n12442_), .C(new_n11920_), .Y(new_n12464_));
  AOI21X1  g12272(.A0(\asqrt[20] ), .A1(\a[40] ), .B0(new_n12464_), .Y(new_n12465_));
  INVX1    g12273(.A(\a[40] ), .Y(new_n12466_));
  INVX1    g12274(.A(\a[41] ), .Y(new_n12467_));
  AOI21X1  g12275(.A0(\asqrt[20] ), .A1(new_n12466_), .B0(new_n12467_), .Y(new_n12468_));
  NOR2X1   g12276(.A(\a[41] ), .B(\a[40] ), .Y(new_n12469_));
  AND2X1   g12277(.A(\asqrt[20] ), .B(new_n12469_), .Y(new_n12470_));
  NOR3X1   g12278(.A(new_n12470_), .B(new_n12468_), .C(new_n12465_), .Y(new_n12471_));
  OAI21X1  g12279(.A0(new_n12471_), .A1(new_n12461_), .B0(\asqrt[22] ), .Y(new_n12472_));
  INVX1    g12280(.A(new_n12459_), .Y(new_n12473_));
  MX2X1    g12281(.A(new_n12473_), .B(new_n12447_), .S0(\a[40] ), .Y(new_n12474_));
  OAI21X1  g12282(.A0(new_n12474_), .A1(new_n11896_), .B0(new_n11362_), .Y(new_n12475_));
  NAND3X1  g12283(.A(new_n12444_), .B(new_n12441_), .C(\asqrt[21] ), .Y(new_n12476_));
  INVX1    g12284(.A(new_n12476_), .Y(new_n12477_));
  OAI21X1  g12285(.A0(new_n12438_), .A1(new_n12427_), .B0(new_n12477_), .Y(new_n12478_));
  AOI21X1  g12286(.A0(new_n12435_), .A1(new_n193_), .B0(new_n12478_), .Y(new_n12479_));
  AOI21X1  g12287(.A0(\asqrt[20] ), .A1(new_n12469_), .B0(new_n12479_), .Y(new_n12480_));
  OR2X1    g12288(.A(new_n12479_), .B(\a[42] ), .Y(new_n12481_));
  OAI22X1  g12289(.A0(new_n12481_), .A1(new_n12470_), .B0(new_n12480_), .B1(new_n11904_), .Y(new_n12482_));
  OAI21X1  g12290(.A0(new_n12475_), .A1(new_n12471_), .B0(new_n12482_), .Y(new_n12483_));
  AOI21X1  g12291(.A0(new_n12483_), .A1(new_n12472_), .B0(new_n10849_), .Y(new_n12484_));
  AND2X1   g12292(.A(new_n11903_), .B(new_n11946_), .Y(new_n12485_));
  NAND3X1  g12293(.A(new_n12485_), .B(\asqrt[20] ), .C(new_n11950_), .Y(new_n12486_));
  INVX1    g12294(.A(new_n12485_), .Y(new_n12487_));
  OAI21X1  g12295(.A0(new_n12487_), .A1(new_n12447_), .B0(new_n11926_), .Y(new_n12488_));
  AND2X1   g12296(.A(new_n12488_), .B(new_n12486_), .Y(new_n12489_));
  INVX1    g12297(.A(new_n12489_), .Y(new_n12490_));
  NAND3X1  g12298(.A(new_n12483_), .B(new_n12472_), .C(new_n10849_), .Y(new_n12491_));
  AOI21X1  g12299(.A0(new_n12491_), .A1(new_n12490_), .B0(new_n12484_), .Y(new_n12492_));
  OR2X1    g12300(.A(new_n12492_), .B(new_n10332_), .Y(new_n12493_));
  AND2X1   g12301(.A(new_n12491_), .B(new_n12490_), .Y(new_n12494_));
  AOI21X1  g12302(.A0(new_n11980_), .A1(new_n11979_), .B0(new_n11939_), .Y(new_n12495_));
  NAND3X1  g12303(.A(new_n12495_), .B(\asqrt[20] ), .C(new_n11928_), .Y(new_n12496_));
  OAI22X1  g12304(.A0(new_n11930_), .A1(new_n11929_), .B0(new_n11927_), .B1(new_n10849_), .Y(new_n12497_));
  OAI21X1  g12305(.A0(new_n12497_), .A1(new_n12447_), .B0(new_n11939_), .Y(new_n12498_));
  AND2X1   g12306(.A(new_n12498_), .B(new_n12496_), .Y(new_n12499_));
  INVX1    g12307(.A(new_n12499_), .Y(new_n12500_));
  OR2X1    g12308(.A(new_n12484_), .B(\asqrt[24] ), .Y(new_n12501_));
  OAI21X1  g12309(.A0(new_n12501_), .A1(new_n12494_), .B0(new_n12500_), .Y(new_n12502_));
  AOI21X1  g12310(.A0(new_n12502_), .A1(new_n12493_), .B0(new_n9833_), .Y(new_n12503_));
  AND2X1   g12311(.A(new_n11952_), .B(new_n11940_), .Y(new_n12504_));
  OR4X1    g12312(.A(new_n12447_), .B(new_n12504_), .C(new_n11984_), .D(new_n11941_), .Y(new_n12505_));
  OR2X1    g12313(.A(new_n12504_), .B(new_n11941_), .Y(new_n12506_));
  OAI21X1  g12314(.A0(new_n12506_), .A1(new_n12447_), .B0(new_n11984_), .Y(new_n12507_));
  AND2X1   g12315(.A(new_n12507_), .B(new_n12505_), .Y(new_n12508_));
  OR2X1    g12316(.A(new_n12474_), .B(new_n11896_), .Y(new_n12509_));
  INVX1    g12317(.A(new_n12464_), .Y(new_n12510_));
  OAI21X1  g12318(.A0(new_n12447_), .A1(new_n12466_), .B0(new_n12510_), .Y(new_n12511_));
  OAI21X1  g12319(.A0(new_n12447_), .A1(\a[40] ), .B0(\a[41] ), .Y(new_n12512_));
  INVX1    g12320(.A(new_n12469_), .Y(new_n12513_));
  OR2X1    g12321(.A(new_n12447_), .B(new_n12513_), .Y(new_n12514_));
  NAND3X1  g12322(.A(new_n12514_), .B(new_n12512_), .C(new_n12511_), .Y(new_n12515_));
  AOI21X1  g12323(.A0(new_n12515_), .A1(new_n12509_), .B0(new_n11362_), .Y(new_n12516_));
  AOI21X1  g12324(.A0(new_n12460_), .A1(\asqrt[21] ), .B0(\asqrt[22] ), .Y(new_n12517_));
  OR2X1    g12325(.A(new_n12480_), .B(new_n11904_), .Y(new_n12518_));
  OR2X1    g12326(.A(new_n12481_), .B(new_n12470_), .Y(new_n12519_));
  AOI22X1  g12327(.A0(new_n12519_), .A1(new_n12518_), .B0(new_n12517_), .B1(new_n12515_), .Y(new_n12520_));
  OAI21X1  g12328(.A0(new_n12520_), .A1(new_n12516_), .B0(\asqrt[23] ), .Y(new_n12521_));
  NOR3X1   g12329(.A(new_n12520_), .B(new_n12516_), .C(\asqrt[23] ), .Y(new_n12522_));
  OAI21X1  g12330(.A0(new_n12522_), .A1(new_n12489_), .B0(new_n12521_), .Y(new_n12523_));
  AOI21X1  g12331(.A0(new_n12523_), .A1(\asqrt[24] ), .B0(\asqrt[25] ), .Y(new_n12524_));
  AOI21X1  g12332(.A0(new_n12524_), .A1(new_n12502_), .B0(new_n12508_), .Y(new_n12525_));
  OAI21X1  g12333(.A0(new_n12525_), .A1(new_n12503_), .B0(\asqrt[26] ), .Y(new_n12526_));
  OR4X1    g12334(.A(new_n12447_), .B(new_n11962_), .C(new_n11988_), .D(new_n11987_), .Y(new_n12527_));
  NAND2X1  g12335(.A(new_n11989_), .B(new_n11954_), .Y(new_n12528_));
  OAI21X1  g12336(.A0(new_n12528_), .A1(new_n12447_), .B0(new_n11988_), .Y(new_n12529_));
  AND2X1   g12337(.A(new_n12529_), .B(new_n12527_), .Y(new_n12530_));
  NOR3X1   g12338(.A(new_n12525_), .B(new_n12503_), .C(\asqrt[26] ), .Y(new_n12531_));
  OAI21X1  g12339(.A0(new_n12531_), .A1(new_n12530_), .B0(new_n12526_), .Y(new_n12532_));
  AND2X1   g12340(.A(new_n12532_), .B(\asqrt[27] ), .Y(new_n12533_));
  INVX1    g12341(.A(new_n12530_), .Y(new_n12534_));
  AND2X1   g12342(.A(new_n12523_), .B(\asqrt[24] ), .Y(new_n12535_));
  NAND2X1  g12343(.A(new_n12491_), .B(new_n12490_), .Y(new_n12536_));
  NOR2X1   g12344(.A(new_n12484_), .B(\asqrt[24] ), .Y(new_n12537_));
  AOI21X1  g12345(.A0(new_n12537_), .A1(new_n12536_), .B0(new_n12499_), .Y(new_n12538_));
  OAI21X1  g12346(.A0(new_n12538_), .A1(new_n12535_), .B0(\asqrt[25] ), .Y(new_n12539_));
  INVX1    g12347(.A(new_n12508_), .Y(new_n12540_));
  OAI21X1  g12348(.A0(new_n12492_), .A1(new_n10332_), .B0(new_n9833_), .Y(new_n12541_));
  OAI21X1  g12349(.A0(new_n12541_), .A1(new_n12538_), .B0(new_n12540_), .Y(new_n12542_));
  NAND3X1  g12350(.A(new_n12542_), .B(new_n12539_), .C(new_n9353_), .Y(new_n12543_));
  NAND2X1  g12351(.A(new_n12543_), .B(new_n12534_), .Y(new_n12544_));
  AND2X1   g12352(.A(new_n11972_), .B(new_n11965_), .Y(new_n12545_));
  NOR4X1   g12353(.A(new_n12447_), .B(new_n12545_), .C(new_n12012_), .D(new_n11964_), .Y(new_n12546_));
  AOI22X1  g12354(.A0(new_n11972_), .A1(new_n11965_), .B0(new_n11963_), .B1(\asqrt[26] ), .Y(new_n12547_));
  AOI21X1  g12355(.A0(new_n12547_), .A1(\asqrt[20] ), .B0(new_n11971_), .Y(new_n12548_));
  NOR2X1   g12356(.A(new_n12548_), .B(new_n12546_), .Y(new_n12549_));
  AOI21X1  g12357(.A0(new_n12542_), .A1(new_n12539_), .B0(new_n9353_), .Y(new_n12550_));
  NOR2X1   g12358(.A(new_n12550_), .B(\asqrt[27] ), .Y(new_n12551_));
  AOI21X1  g12359(.A0(new_n12551_), .A1(new_n12544_), .B0(new_n12549_), .Y(new_n12552_));
  OAI21X1  g12360(.A0(new_n12552_), .A1(new_n12533_), .B0(\asqrt[28] ), .Y(new_n12553_));
  AND2X1   g12361(.A(new_n12017_), .B(new_n12014_), .Y(new_n12554_));
  OR4X1    g12362(.A(new_n12447_), .B(new_n12554_), .C(new_n11977_), .D(new_n12015_), .Y(new_n12555_));
  OR2X1    g12363(.A(new_n12554_), .B(new_n12015_), .Y(new_n12556_));
  OAI21X1  g12364(.A0(new_n12556_), .A1(new_n12447_), .B0(new_n11977_), .Y(new_n12557_));
  AND2X1   g12365(.A(new_n12557_), .B(new_n12555_), .Y(new_n12558_));
  INVX1    g12366(.A(new_n12558_), .Y(new_n12559_));
  AOI21X1  g12367(.A0(new_n12543_), .A1(new_n12534_), .B0(new_n12550_), .Y(new_n12560_));
  OAI21X1  g12368(.A0(new_n12560_), .A1(new_n8874_), .B0(new_n8412_), .Y(new_n12561_));
  OAI21X1  g12369(.A0(new_n12561_), .A1(new_n12552_), .B0(new_n12559_), .Y(new_n12562_));
  AOI21X1  g12370(.A0(new_n12562_), .A1(new_n12553_), .B0(new_n7970_), .Y(new_n12563_));
  OR4X1    g12371(.A(new_n12447_), .B(new_n12027_), .C(new_n11999_), .D(new_n11993_), .Y(new_n12564_));
  NAND2X1  g12372(.A(new_n12000_), .B(new_n12019_), .Y(new_n12565_));
  OAI21X1  g12373(.A0(new_n12565_), .A1(new_n12447_), .B0(new_n11999_), .Y(new_n12566_));
  AND2X1   g12374(.A(new_n12566_), .B(new_n12564_), .Y(new_n12567_));
  INVX1    g12375(.A(new_n12567_), .Y(new_n12568_));
  NAND3X1  g12376(.A(new_n12562_), .B(new_n12553_), .C(new_n7970_), .Y(new_n12569_));
  AOI21X1  g12377(.A0(new_n12569_), .A1(new_n12568_), .B0(new_n12563_), .Y(new_n12570_));
  OR2X1    g12378(.A(new_n12570_), .B(new_n7527_), .Y(new_n12571_));
  AND2X1   g12379(.A(new_n12569_), .B(new_n12568_), .Y(new_n12572_));
  OAI21X1  g12380(.A0(new_n12020_), .A1(new_n12003_), .B0(new_n12008_), .Y(new_n12573_));
  NOR3X1   g12381(.A(new_n12573_), .B(new_n12447_), .C(new_n12041_), .Y(new_n12574_));
  AOI22X1  g12382(.A0(new_n12043_), .A1(new_n12042_), .B0(new_n12028_), .B1(\asqrt[29] ), .Y(new_n12575_));
  AOI21X1  g12383(.A0(new_n12575_), .A1(\asqrt[20] ), .B0(new_n12008_), .Y(new_n12576_));
  NOR2X1   g12384(.A(new_n12576_), .B(new_n12574_), .Y(new_n12577_));
  INVX1    g12385(.A(new_n12577_), .Y(new_n12578_));
  OR2X1    g12386(.A(new_n12563_), .B(\asqrt[30] ), .Y(new_n12579_));
  OAI21X1  g12387(.A0(new_n12579_), .A1(new_n12572_), .B0(new_n12578_), .Y(new_n12580_));
  AOI21X1  g12388(.A0(new_n12580_), .A1(new_n12571_), .B0(new_n7103_), .Y(new_n12581_));
  AND2X1   g12389(.A(new_n12029_), .B(new_n12021_), .Y(new_n12582_));
  OR4X1    g12390(.A(new_n12447_), .B(new_n12582_), .C(new_n12046_), .D(new_n12022_), .Y(new_n12583_));
  OR2X1    g12391(.A(new_n12582_), .B(new_n12022_), .Y(new_n12584_));
  OAI21X1  g12392(.A0(new_n12584_), .A1(new_n12447_), .B0(new_n12046_), .Y(new_n12585_));
  AND2X1   g12393(.A(new_n12585_), .B(new_n12583_), .Y(new_n12586_));
  OR2X1    g12394(.A(new_n12560_), .B(new_n8874_), .Y(new_n12587_));
  AND2X1   g12395(.A(new_n12543_), .B(new_n12534_), .Y(new_n12588_));
  INVX1    g12396(.A(new_n12549_), .Y(new_n12589_));
  OR2X1    g12397(.A(new_n12550_), .B(\asqrt[27] ), .Y(new_n12590_));
  OAI21X1  g12398(.A0(new_n12590_), .A1(new_n12588_), .B0(new_n12589_), .Y(new_n12591_));
  AOI21X1  g12399(.A0(new_n12591_), .A1(new_n12587_), .B0(new_n8412_), .Y(new_n12592_));
  AOI21X1  g12400(.A0(new_n12532_), .A1(\asqrt[27] ), .B0(\asqrt[28] ), .Y(new_n12593_));
  AOI21X1  g12401(.A0(new_n12593_), .A1(new_n12591_), .B0(new_n12558_), .Y(new_n12594_));
  OAI21X1  g12402(.A0(new_n12594_), .A1(new_n12592_), .B0(\asqrt[29] ), .Y(new_n12595_));
  NOR3X1   g12403(.A(new_n12594_), .B(new_n12592_), .C(\asqrt[29] ), .Y(new_n12596_));
  OAI21X1  g12404(.A0(new_n12596_), .A1(new_n12567_), .B0(new_n12595_), .Y(new_n12597_));
  AOI21X1  g12405(.A0(new_n12597_), .A1(\asqrt[30] ), .B0(\asqrt[31] ), .Y(new_n12598_));
  AOI21X1  g12406(.A0(new_n12598_), .A1(new_n12580_), .B0(new_n12586_), .Y(new_n12599_));
  OAI21X1  g12407(.A0(new_n12599_), .A1(new_n12581_), .B0(\asqrt[32] ), .Y(new_n12600_));
  OR4X1    g12408(.A(new_n12447_), .B(new_n12037_), .C(new_n12040_), .D(new_n12064_), .Y(new_n12601_));
  NAND2X1  g12409(.A(new_n12049_), .B(new_n12031_), .Y(new_n12602_));
  OAI21X1  g12410(.A0(new_n12602_), .A1(new_n12447_), .B0(new_n12040_), .Y(new_n12603_));
  AND2X1   g12411(.A(new_n12603_), .B(new_n12601_), .Y(new_n12604_));
  NOR3X1   g12412(.A(new_n12599_), .B(new_n12581_), .C(\asqrt[32] ), .Y(new_n12605_));
  OAI21X1  g12413(.A0(new_n12605_), .A1(new_n12604_), .B0(new_n12600_), .Y(new_n12606_));
  AND2X1   g12414(.A(new_n12606_), .B(\asqrt[33] ), .Y(new_n12607_));
  INVX1    g12415(.A(new_n12604_), .Y(new_n12608_));
  AND2X1   g12416(.A(new_n12597_), .B(\asqrt[30] ), .Y(new_n12609_));
  NAND2X1  g12417(.A(new_n12569_), .B(new_n12568_), .Y(new_n12610_));
  NOR2X1   g12418(.A(new_n12563_), .B(\asqrt[30] ), .Y(new_n12611_));
  AOI21X1  g12419(.A0(new_n12611_), .A1(new_n12610_), .B0(new_n12577_), .Y(new_n12612_));
  OAI21X1  g12420(.A0(new_n12612_), .A1(new_n12609_), .B0(\asqrt[31] ), .Y(new_n12613_));
  INVX1    g12421(.A(new_n12586_), .Y(new_n12614_));
  OAI21X1  g12422(.A0(new_n12570_), .A1(new_n7527_), .B0(new_n7103_), .Y(new_n12615_));
  OAI21X1  g12423(.A0(new_n12615_), .A1(new_n12612_), .B0(new_n12614_), .Y(new_n12616_));
  NAND3X1  g12424(.A(new_n12616_), .B(new_n12613_), .C(new_n6699_), .Y(new_n12617_));
  NAND2X1  g12425(.A(new_n12617_), .B(new_n12608_), .Y(new_n12618_));
  AND2X1   g12426(.A(new_n12056_), .B(new_n12050_), .Y(new_n12619_));
  NOR4X1   g12427(.A(new_n12447_), .B(new_n12619_), .C(new_n12087_), .D(new_n12039_), .Y(new_n12620_));
  AOI22X1  g12428(.A0(new_n12056_), .A1(new_n12050_), .B0(new_n12038_), .B1(\asqrt[32] ), .Y(new_n12621_));
  AOI21X1  g12429(.A0(new_n12621_), .A1(\asqrt[20] ), .B0(new_n12055_), .Y(new_n12622_));
  NOR2X1   g12430(.A(new_n12622_), .B(new_n12620_), .Y(new_n12623_));
  AOI21X1  g12431(.A0(new_n12616_), .A1(new_n12613_), .B0(new_n6699_), .Y(new_n12624_));
  NOR2X1   g12432(.A(new_n12624_), .B(\asqrt[33] ), .Y(new_n12625_));
  AOI21X1  g12433(.A0(new_n12625_), .A1(new_n12618_), .B0(new_n12623_), .Y(new_n12626_));
  OAI21X1  g12434(.A0(new_n12626_), .A1(new_n12607_), .B0(\asqrt[34] ), .Y(new_n12627_));
  OR2X1    g12435(.A(new_n12066_), .B(new_n12057_), .Y(new_n12628_));
  NAND4X1  g12436(.A(\asqrt[20] ), .B(new_n12628_), .C(new_n12062_), .D(new_n12058_), .Y(new_n12629_));
  NAND2X1  g12437(.A(new_n12628_), .B(new_n12058_), .Y(new_n12630_));
  OAI21X1  g12438(.A0(new_n12630_), .A1(new_n12447_), .B0(new_n12063_), .Y(new_n12631_));
  AND2X1   g12439(.A(new_n12631_), .B(new_n12629_), .Y(new_n12632_));
  INVX1    g12440(.A(new_n12632_), .Y(new_n12633_));
  AOI21X1  g12441(.A0(new_n12617_), .A1(new_n12608_), .B0(new_n12624_), .Y(new_n12634_));
  OAI21X1  g12442(.A0(new_n12634_), .A1(new_n6294_), .B0(new_n5941_), .Y(new_n12635_));
  OAI21X1  g12443(.A0(new_n12635_), .A1(new_n12626_), .B0(new_n12633_), .Y(new_n12636_));
  AOI21X1  g12444(.A0(new_n12636_), .A1(new_n12627_), .B0(new_n5541_), .Y(new_n12637_));
  OR4X1    g12445(.A(new_n12447_), .B(new_n12101_), .C(new_n12074_), .D(new_n12068_), .Y(new_n12638_));
  NAND2X1  g12446(.A(new_n12075_), .B(new_n12093_), .Y(new_n12639_));
  OAI21X1  g12447(.A0(new_n12639_), .A1(new_n12447_), .B0(new_n12074_), .Y(new_n12640_));
  AND2X1   g12448(.A(new_n12640_), .B(new_n12638_), .Y(new_n12641_));
  INVX1    g12449(.A(new_n12641_), .Y(new_n12642_));
  NAND3X1  g12450(.A(new_n12636_), .B(new_n12627_), .C(new_n5541_), .Y(new_n12643_));
  AOI21X1  g12451(.A0(new_n12643_), .A1(new_n12642_), .B0(new_n12637_), .Y(new_n12644_));
  OR2X1    g12452(.A(new_n12644_), .B(new_n5176_), .Y(new_n12645_));
  AND2X1   g12453(.A(new_n12643_), .B(new_n12642_), .Y(new_n12646_));
  OAI21X1  g12454(.A0(new_n12094_), .A1(new_n12078_), .B0(new_n12083_), .Y(new_n12647_));
  NOR3X1   g12455(.A(new_n12647_), .B(new_n12447_), .C(new_n12115_), .Y(new_n12648_));
  AOI22X1  g12456(.A0(new_n12117_), .A1(new_n12116_), .B0(new_n12102_), .B1(\asqrt[35] ), .Y(new_n12649_));
  AOI21X1  g12457(.A0(new_n12649_), .A1(\asqrt[20] ), .B0(new_n12083_), .Y(new_n12650_));
  NOR2X1   g12458(.A(new_n12650_), .B(new_n12648_), .Y(new_n12651_));
  INVX1    g12459(.A(new_n12651_), .Y(new_n12652_));
  OR2X1    g12460(.A(new_n12637_), .B(\asqrt[36] ), .Y(new_n12653_));
  OAI21X1  g12461(.A0(new_n12653_), .A1(new_n12646_), .B0(new_n12652_), .Y(new_n12654_));
  AOI21X1  g12462(.A0(new_n12654_), .A1(new_n12645_), .B0(new_n4826_), .Y(new_n12655_));
  AND2X1   g12463(.A(new_n12103_), .B(new_n12095_), .Y(new_n12656_));
  OR4X1    g12464(.A(new_n12447_), .B(new_n12656_), .C(new_n12120_), .D(new_n12096_), .Y(new_n12657_));
  OR2X1    g12465(.A(new_n12656_), .B(new_n12096_), .Y(new_n12658_));
  OAI21X1  g12466(.A0(new_n12658_), .A1(new_n12447_), .B0(new_n12120_), .Y(new_n12659_));
  AND2X1   g12467(.A(new_n12659_), .B(new_n12657_), .Y(new_n12660_));
  OR2X1    g12468(.A(new_n12634_), .B(new_n6294_), .Y(new_n12661_));
  AND2X1   g12469(.A(new_n12617_), .B(new_n12608_), .Y(new_n12662_));
  INVX1    g12470(.A(new_n12623_), .Y(new_n12663_));
  OR2X1    g12471(.A(new_n12624_), .B(\asqrt[33] ), .Y(new_n12664_));
  OAI21X1  g12472(.A0(new_n12664_), .A1(new_n12662_), .B0(new_n12663_), .Y(new_n12665_));
  AOI21X1  g12473(.A0(new_n12665_), .A1(new_n12661_), .B0(new_n5941_), .Y(new_n12666_));
  AOI21X1  g12474(.A0(new_n12606_), .A1(\asqrt[33] ), .B0(\asqrt[34] ), .Y(new_n12667_));
  AOI21X1  g12475(.A0(new_n12667_), .A1(new_n12665_), .B0(new_n12632_), .Y(new_n12668_));
  OAI21X1  g12476(.A0(new_n12668_), .A1(new_n12666_), .B0(\asqrt[35] ), .Y(new_n12669_));
  NOR3X1   g12477(.A(new_n12668_), .B(new_n12666_), .C(\asqrt[35] ), .Y(new_n12670_));
  OAI21X1  g12478(.A0(new_n12670_), .A1(new_n12641_), .B0(new_n12669_), .Y(new_n12671_));
  AOI21X1  g12479(.A0(new_n12671_), .A1(\asqrt[36] ), .B0(\asqrt[37] ), .Y(new_n12672_));
  AOI21X1  g12480(.A0(new_n12672_), .A1(new_n12654_), .B0(new_n12660_), .Y(new_n12673_));
  OAI21X1  g12481(.A0(new_n12673_), .A1(new_n12655_), .B0(\asqrt[38] ), .Y(new_n12674_));
  OR4X1    g12482(.A(new_n12447_), .B(new_n12111_), .C(new_n12114_), .D(new_n12138_), .Y(new_n12675_));
  NAND2X1  g12483(.A(new_n12123_), .B(new_n12105_), .Y(new_n12676_));
  OAI21X1  g12484(.A0(new_n12676_), .A1(new_n12447_), .B0(new_n12114_), .Y(new_n12677_));
  AND2X1   g12485(.A(new_n12677_), .B(new_n12675_), .Y(new_n12678_));
  NOR3X1   g12486(.A(new_n12673_), .B(new_n12655_), .C(\asqrt[38] ), .Y(new_n12679_));
  OAI21X1  g12487(.A0(new_n12679_), .A1(new_n12678_), .B0(new_n12674_), .Y(new_n12680_));
  AND2X1   g12488(.A(new_n12680_), .B(\asqrt[39] ), .Y(new_n12681_));
  INVX1    g12489(.A(new_n12678_), .Y(new_n12682_));
  AND2X1   g12490(.A(new_n12671_), .B(\asqrt[36] ), .Y(new_n12683_));
  NAND2X1  g12491(.A(new_n12643_), .B(new_n12642_), .Y(new_n12684_));
  NOR2X1   g12492(.A(new_n12637_), .B(\asqrt[36] ), .Y(new_n12685_));
  AOI21X1  g12493(.A0(new_n12685_), .A1(new_n12684_), .B0(new_n12651_), .Y(new_n12686_));
  OAI21X1  g12494(.A0(new_n12686_), .A1(new_n12683_), .B0(\asqrt[37] ), .Y(new_n12687_));
  INVX1    g12495(.A(new_n12660_), .Y(new_n12688_));
  OAI21X1  g12496(.A0(new_n12644_), .A1(new_n5176_), .B0(new_n4826_), .Y(new_n12689_));
  OAI21X1  g12497(.A0(new_n12689_), .A1(new_n12686_), .B0(new_n12688_), .Y(new_n12690_));
  NAND3X1  g12498(.A(new_n12690_), .B(new_n12687_), .C(new_n4493_), .Y(new_n12691_));
  NAND2X1  g12499(.A(new_n12691_), .B(new_n12682_), .Y(new_n12692_));
  AND2X1   g12500(.A(new_n12130_), .B(new_n12124_), .Y(new_n12693_));
  NOR4X1   g12501(.A(new_n12447_), .B(new_n12693_), .C(new_n12161_), .D(new_n12113_), .Y(new_n12694_));
  AOI22X1  g12502(.A0(new_n12130_), .A1(new_n12124_), .B0(new_n12112_), .B1(\asqrt[38] ), .Y(new_n12695_));
  AOI21X1  g12503(.A0(new_n12695_), .A1(\asqrt[20] ), .B0(new_n12129_), .Y(new_n12696_));
  NOR2X1   g12504(.A(new_n12696_), .B(new_n12694_), .Y(new_n12697_));
  AOI21X1  g12505(.A0(new_n12690_), .A1(new_n12687_), .B0(new_n4493_), .Y(new_n12698_));
  NOR2X1   g12506(.A(new_n12698_), .B(\asqrt[39] ), .Y(new_n12699_));
  AOI21X1  g12507(.A0(new_n12699_), .A1(new_n12692_), .B0(new_n12697_), .Y(new_n12700_));
  OAI21X1  g12508(.A0(new_n12700_), .A1(new_n12681_), .B0(\asqrt[40] ), .Y(new_n12701_));
  AND2X1   g12509(.A(new_n12165_), .B(new_n12163_), .Y(new_n12702_));
  OR4X1    g12510(.A(new_n12447_), .B(new_n12702_), .C(new_n12137_), .D(new_n12164_), .Y(new_n12703_));
  OR2X1    g12511(.A(new_n12702_), .B(new_n12164_), .Y(new_n12704_));
  OAI21X1  g12512(.A0(new_n12704_), .A1(new_n12447_), .B0(new_n12137_), .Y(new_n12705_));
  AND2X1   g12513(.A(new_n12705_), .B(new_n12703_), .Y(new_n12706_));
  INVX1    g12514(.A(new_n12706_), .Y(new_n12707_));
  AOI21X1  g12515(.A0(new_n12691_), .A1(new_n12682_), .B0(new_n12698_), .Y(new_n12708_));
  OAI21X1  g12516(.A0(new_n12708_), .A1(new_n4165_), .B0(new_n3863_), .Y(new_n12709_));
  OAI21X1  g12517(.A0(new_n12709_), .A1(new_n12700_), .B0(new_n12707_), .Y(new_n12710_));
  AOI21X1  g12518(.A0(new_n12710_), .A1(new_n12701_), .B0(new_n3564_), .Y(new_n12711_));
  OR4X1    g12519(.A(new_n12447_), .B(new_n12175_), .C(new_n12148_), .D(new_n12142_), .Y(new_n12712_));
  NAND2X1  g12520(.A(new_n12149_), .B(new_n12167_), .Y(new_n12713_));
  OAI21X1  g12521(.A0(new_n12713_), .A1(new_n12447_), .B0(new_n12148_), .Y(new_n12714_));
  AND2X1   g12522(.A(new_n12714_), .B(new_n12712_), .Y(new_n12715_));
  INVX1    g12523(.A(new_n12715_), .Y(new_n12716_));
  NAND3X1  g12524(.A(new_n12710_), .B(new_n12701_), .C(new_n3564_), .Y(new_n12717_));
  AOI21X1  g12525(.A0(new_n12717_), .A1(new_n12716_), .B0(new_n12711_), .Y(new_n12718_));
  OR2X1    g12526(.A(new_n12718_), .B(new_n3276_), .Y(new_n12719_));
  OR2X1    g12527(.A(new_n12708_), .B(new_n4165_), .Y(new_n12720_));
  AND2X1   g12528(.A(new_n12691_), .B(new_n12682_), .Y(new_n12721_));
  INVX1    g12529(.A(new_n12697_), .Y(new_n12722_));
  OR2X1    g12530(.A(new_n12698_), .B(\asqrt[39] ), .Y(new_n12723_));
  OAI21X1  g12531(.A0(new_n12723_), .A1(new_n12721_), .B0(new_n12722_), .Y(new_n12724_));
  AOI21X1  g12532(.A0(new_n12724_), .A1(new_n12720_), .B0(new_n3863_), .Y(new_n12725_));
  AOI21X1  g12533(.A0(new_n12680_), .A1(\asqrt[39] ), .B0(\asqrt[40] ), .Y(new_n12726_));
  AOI21X1  g12534(.A0(new_n12726_), .A1(new_n12724_), .B0(new_n12706_), .Y(new_n12727_));
  NOR3X1   g12535(.A(new_n12727_), .B(new_n12725_), .C(\asqrt[41] ), .Y(new_n12728_));
  NOR2X1   g12536(.A(new_n12728_), .B(new_n12715_), .Y(new_n12729_));
  OAI21X1  g12537(.A0(new_n12168_), .A1(new_n12152_), .B0(new_n12157_), .Y(new_n12730_));
  NOR3X1   g12538(.A(new_n12730_), .B(new_n12447_), .C(new_n12189_), .Y(new_n12731_));
  AOI22X1  g12539(.A0(new_n12191_), .A1(new_n12190_), .B0(new_n12176_), .B1(\asqrt[41] ), .Y(new_n12732_));
  AOI21X1  g12540(.A0(new_n12732_), .A1(\asqrt[20] ), .B0(new_n12157_), .Y(new_n12733_));
  NOR2X1   g12541(.A(new_n12733_), .B(new_n12731_), .Y(new_n12734_));
  INVX1    g12542(.A(new_n12734_), .Y(new_n12735_));
  OAI21X1  g12543(.A0(new_n12727_), .A1(new_n12725_), .B0(\asqrt[41] ), .Y(new_n12736_));
  NAND2X1  g12544(.A(new_n12736_), .B(new_n3276_), .Y(new_n12737_));
  OAI21X1  g12545(.A0(new_n12737_), .A1(new_n12729_), .B0(new_n12735_), .Y(new_n12738_));
  AOI21X1  g12546(.A0(new_n12738_), .A1(new_n12719_), .B0(new_n3008_), .Y(new_n12739_));
  AND2X1   g12547(.A(new_n12177_), .B(new_n12169_), .Y(new_n12740_));
  OR4X1    g12548(.A(new_n12447_), .B(new_n12740_), .C(new_n12194_), .D(new_n12170_), .Y(new_n12741_));
  OR2X1    g12549(.A(new_n12740_), .B(new_n12170_), .Y(new_n12742_));
  OAI21X1  g12550(.A0(new_n12742_), .A1(new_n12447_), .B0(new_n12194_), .Y(new_n12743_));
  AND2X1   g12551(.A(new_n12743_), .B(new_n12741_), .Y(new_n12744_));
  OAI21X1  g12552(.A0(new_n12728_), .A1(new_n12715_), .B0(new_n12736_), .Y(new_n12745_));
  AOI21X1  g12553(.A0(new_n12745_), .A1(\asqrt[42] ), .B0(\asqrt[43] ), .Y(new_n12746_));
  AOI21X1  g12554(.A0(new_n12746_), .A1(new_n12738_), .B0(new_n12744_), .Y(new_n12747_));
  OAI21X1  g12555(.A0(new_n12747_), .A1(new_n12739_), .B0(\asqrt[44] ), .Y(new_n12748_));
  OR4X1    g12556(.A(new_n12447_), .B(new_n12185_), .C(new_n12188_), .D(new_n12212_), .Y(new_n12749_));
  NAND2X1  g12557(.A(new_n12197_), .B(new_n12179_), .Y(new_n12750_));
  OAI21X1  g12558(.A0(new_n12750_), .A1(new_n12447_), .B0(new_n12188_), .Y(new_n12751_));
  AND2X1   g12559(.A(new_n12751_), .B(new_n12749_), .Y(new_n12752_));
  NOR3X1   g12560(.A(new_n12747_), .B(new_n12739_), .C(\asqrt[44] ), .Y(new_n12753_));
  OAI21X1  g12561(.A0(new_n12753_), .A1(new_n12752_), .B0(new_n12748_), .Y(new_n12754_));
  AND2X1   g12562(.A(new_n12754_), .B(\asqrt[45] ), .Y(new_n12755_));
  OR2X1    g12563(.A(new_n12753_), .B(new_n12752_), .Y(new_n12756_));
  AND2X1   g12564(.A(new_n12748_), .B(new_n2570_), .Y(new_n12757_));
  AND2X1   g12565(.A(new_n12199_), .B(new_n12198_), .Y(new_n12758_));
  NOR4X1   g12566(.A(new_n12447_), .B(new_n12236_), .C(new_n12758_), .D(new_n12187_), .Y(new_n12759_));
  AOI22X1  g12567(.A0(new_n12199_), .A1(new_n12198_), .B0(new_n12186_), .B1(\asqrt[44] ), .Y(new_n12760_));
  AOI21X1  g12568(.A0(new_n12760_), .A1(\asqrt[20] ), .B0(new_n12204_), .Y(new_n12761_));
  NOR2X1   g12569(.A(new_n12761_), .B(new_n12759_), .Y(new_n12762_));
  AOI21X1  g12570(.A0(new_n12757_), .A1(new_n12756_), .B0(new_n12762_), .Y(new_n12763_));
  OAI21X1  g12571(.A0(new_n12763_), .A1(new_n12755_), .B0(\asqrt[46] ), .Y(new_n12764_));
  AND2X1   g12572(.A(new_n12239_), .B(new_n12237_), .Y(new_n12765_));
  OR4X1    g12573(.A(new_n12447_), .B(new_n12765_), .C(new_n12211_), .D(new_n12238_), .Y(new_n12766_));
  OR2X1    g12574(.A(new_n12765_), .B(new_n12238_), .Y(new_n12767_));
  OAI21X1  g12575(.A0(new_n12767_), .A1(new_n12447_), .B0(new_n12211_), .Y(new_n12768_));
  AND2X1   g12576(.A(new_n12768_), .B(new_n12766_), .Y(new_n12769_));
  INVX1    g12577(.A(new_n12769_), .Y(new_n12770_));
  AND2X1   g12578(.A(new_n12745_), .B(\asqrt[42] ), .Y(new_n12771_));
  OR2X1    g12579(.A(new_n12728_), .B(new_n12715_), .Y(new_n12772_));
  AND2X1   g12580(.A(new_n12736_), .B(new_n3276_), .Y(new_n12773_));
  AOI21X1  g12581(.A0(new_n12773_), .A1(new_n12772_), .B0(new_n12734_), .Y(new_n12774_));
  OAI21X1  g12582(.A0(new_n12774_), .A1(new_n12771_), .B0(\asqrt[43] ), .Y(new_n12775_));
  INVX1    g12583(.A(new_n12744_), .Y(new_n12776_));
  OAI21X1  g12584(.A0(new_n12718_), .A1(new_n3276_), .B0(new_n3008_), .Y(new_n12777_));
  OAI21X1  g12585(.A0(new_n12777_), .A1(new_n12774_), .B0(new_n12776_), .Y(new_n12778_));
  AOI21X1  g12586(.A0(new_n12778_), .A1(new_n12775_), .B0(new_n2769_), .Y(new_n12779_));
  INVX1    g12587(.A(new_n12752_), .Y(new_n12780_));
  NAND3X1  g12588(.A(new_n12778_), .B(new_n12775_), .C(new_n2769_), .Y(new_n12781_));
  AOI21X1  g12589(.A0(new_n12781_), .A1(new_n12780_), .B0(new_n12779_), .Y(new_n12782_));
  OAI21X1  g12590(.A0(new_n12782_), .A1(new_n2570_), .B0(new_n2263_), .Y(new_n12783_));
  OAI21X1  g12591(.A0(new_n12783_), .A1(new_n12763_), .B0(new_n12770_), .Y(new_n12784_));
  AOI21X1  g12592(.A0(new_n12784_), .A1(new_n12764_), .B0(new_n2040_), .Y(new_n12785_));
  NAND3X1  g12593(.A(new_n12223_), .B(new_n12221_), .C(new_n12241_), .Y(new_n12786_));
  NOR3X1   g12594(.A(new_n12447_), .B(new_n12249_), .C(new_n12216_), .Y(new_n12787_));
  OAI22X1  g12595(.A0(new_n12787_), .A1(new_n12221_), .B0(new_n12786_), .B1(new_n12447_), .Y(new_n12788_));
  NAND3X1  g12596(.A(new_n12784_), .B(new_n12764_), .C(new_n2040_), .Y(new_n12789_));
  AOI21X1  g12597(.A0(new_n12789_), .A1(new_n12788_), .B0(new_n12785_), .Y(new_n12790_));
  OR2X1    g12598(.A(new_n12790_), .B(new_n1834_), .Y(new_n12791_));
  AND2X1   g12599(.A(new_n12789_), .B(new_n12788_), .Y(new_n12792_));
  OAI21X1  g12600(.A0(new_n12242_), .A1(new_n12226_), .B0(new_n12231_), .Y(new_n12793_));
  NOR3X1   g12601(.A(new_n12793_), .B(new_n12447_), .C(new_n12263_), .Y(new_n12794_));
  AOI22X1  g12602(.A0(new_n12265_), .A1(new_n12264_), .B0(new_n12250_), .B1(\asqrt[47] ), .Y(new_n12795_));
  AOI21X1  g12603(.A0(new_n12795_), .A1(\asqrt[20] ), .B0(new_n12231_), .Y(new_n12796_));
  NOR2X1   g12604(.A(new_n12796_), .B(new_n12794_), .Y(new_n12797_));
  INVX1    g12605(.A(new_n12797_), .Y(new_n12798_));
  OR2X1    g12606(.A(new_n12782_), .B(new_n2570_), .Y(new_n12799_));
  NOR2X1   g12607(.A(new_n12753_), .B(new_n12752_), .Y(new_n12800_));
  NAND2X1  g12608(.A(new_n12748_), .B(new_n2570_), .Y(new_n12801_));
  INVX1    g12609(.A(new_n12762_), .Y(new_n12802_));
  OAI21X1  g12610(.A0(new_n12801_), .A1(new_n12800_), .B0(new_n12802_), .Y(new_n12803_));
  AOI21X1  g12611(.A0(new_n12803_), .A1(new_n12799_), .B0(new_n2263_), .Y(new_n12804_));
  AOI21X1  g12612(.A0(new_n12754_), .A1(\asqrt[45] ), .B0(\asqrt[46] ), .Y(new_n12805_));
  AOI21X1  g12613(.A0(new_n12805_), .A1(new_n12803_), .B0(new_n12769_), .Y(new_n12806_));
  OAI21X1  g12614(.A0(new_n12806_), .A1(new_n12804_), .B0(\asqrt[47] ), .Y(new_n12807_));
  NAND2X1  g12615(.A(new_n12807_), .B(new_n1834_), .Y(new_n12808_));
  OAI21X1  g12616(.A0(new_n12808_), .A1(new_n12792_), .B0(new_n12798_), .Y(new_n12809_));
  AOI21X1  g12617(.A0(new_n12809_), .A1(new_n12791_), .B0(new_n1632_), .Y(new_n12810_));
  AND2X1   g12618(.A(new_n12251_), .B(new_n12243_), .Y(new_n12811_));
  OR4X1    g12619(.A(new_n12447_), .B(new_n12811_), .C(new_n12268_), .D(new_n12244_), .Y(new_n12812_));
  OR2X1    g12620(.A(new_n12811_), .B(new_n12244_), .Y(new_n12813_));
  OAI21X1  g12621(.A0(new_n12813_), .A1(new_n12447_), .B0(new_n12268_), .Y(new_n12814_));
  AND2X1   g12622(.A(new_n12814_), .B(new_n12812_), .Y(new_n12815_));
  INVX1    g12623(.A(new_n12788_), .Y(new_n12816_));
  NOR3X1   g12624(.A(new_n12806_), .B(new_n12804_), .C(\asqrt[47] ), .Y(new_n12817_));
  OAI21X1  g12625(.A0(new_n12817_), .A1(new_n12816_), .B0(new_n12807_), .Y(new_n12818_));
  AOI21X1  g12626(.A0(new_n12818_), .A1(\asqrt[48] ), .B0(\asqrt[49] ), .Y(new_n12819_));
  AOI21X1  g12627(.A0(new_n12819_), .A1(new_n12809_), .B0(new_n12815_), .Y(new_n12820_));
  OAI21X1  g12628(.A0(new_n12820_), .A1(new_n12810_), .B0(\asqrt[50] ), .Y(new_n12821_));
  OR4X1    g12629(.A(new_n12447_), .B(new_n12259_), .C(new_n12262_), .D(new_n12286_), .Y(new_n12822_));
  NAND2X1  g12630(.A(new_n12271_), .B(new_n12253_), .Y(new_n12823_));
  OAI21X1  g12631(.A0(new_n12823_), .A1(new_n12447_), .B0(new_n12262_), .Y(new_n12824_));
  AND2X1   g12632(.A(new_n12824_), .B(new_n12822_), .Y(new_n12825_));
  NOR3X1   g12633(.A(new_n12820_), .B(new_n12810_), .C(\asqrt[50] ), .Y(new_n12826_));
  OAI21X1  g12634(.A0(new_n12826_), .A1(new_n12825_), .B0(new_n12821_), .Y(new_n12827_));
  AND2X1   g12635(.A(new_n12827_), .B(\asqrt[51] ), .Y(new_n12828_));
  OR2X1    g12636(.A(new_n12826_), .B(new_n12825_), .Y(new_n12829_));
  AND2X1   g12637(.A(new_n12278_), .B(new_n12272_), .Y(new_n12830_));
  NOR4X1   g12638(.A(new_n12447_), .B(new_n12830_), .C(new_n12302_), .D(new_n12261_), .Y(new_n12831_));
  AOI22X1  g12639(.A0(new_n12278_), .A1(new_n12272_), .B0(new_n12260_), .B1(\asqrt[50] ), .Y(new_n12832_));
  AOI21X1  g12640(.A0(new_n12832_), .A1(\asqrt[20] ), .B0(new_n12277_), .Y(new_n12833_));
  NOR2X1   g12641(.A(new_n12833_), .B(new_n12831_), .Y(new_n12834_));
  AND2X1   g12642(.A(new_n12821_), .B(new_n1277_), .Y(new_n12835_));
  AOI21X1  g12643(.A0(new_n12835_), .A1(new_n12829_), .B0(new_n12834_), .Y(new_n12836_));
  OAI21X1  g12644(.A0(new_n12836_), .A1(new_n12828_), .B0(\asqrt[52] ), .Y(new_n12837_));
  AND2X1   g12645(.A(new_n12306_), .B(new_n12304_), .Y(new_n12838_));
  OR4X1    g12646(.A(new_n12447_), .B(new_n12838_), .C(new_n12285_), .D(new_n12305_), .Y(new_n12839_));
  OR2X1    g12647(.A(new_n12838_), .B(new_n12305_), .Y(new_n12840_));
  OAI21X1  g12648(.A0(new_n12840_), .A1(new_n12447_), .B0(new_n12285_), .Y(new_n12841_));
  AND2X1   g12649(.A(new_n12841_), .B(new_n12839_), .Y(new_n12842_));
  INVX1    g12650(.A(new_n12842_), .Y(new_n12843_));
  AND2X1   g12651(.A(new_n12818_), .B(\asqrt[48] ), .Y(new_n12844_));
  NAND2X1  g12652(.A(new_n12789_), .B(new_n12788_), .Y(new_n12845_));
  AND2X1   g12653(.A(new_n12807_), .B(new_n1834_), .Y(new_n12846_));
  AOI21X1  g12654(.A0(new_n12846_), .A1(new_n12845_), .B0(new_n12797_), .Y(new_n12847_));
  OAI21X1  g12655(.A0(new_n12847_), .A1(new_n12844_), .B0(\asqrt[49] ), .Y(new_n12848_));
  INVX1    g12656(.A(new_n12815_), .Y(new_n12849_));
  OAI21X1  g12657(.A0(new_n12790_), .A1(new_n1834_), .B0(new_n1632_), .Y(new_n12850_));
  OAI21X1  g12658(.A0(new_n12850_), .A1(new_n12847_), .B0(new_n12849_), .Y(new_n12851_));
  AOI21X1  g12659(.A0(new_n12851_), .A1(new_n12848_), .B0(new_n1469_), .Y(new_n12852_));
  INVX1    g12660(.A(new_n12825_), .Y(new_n12853_));
  NAND3X1  g12661(.A(new_n12851_), .B(new_n12848_), .C(new_n1469_), .Y(new_n12854_));
  AOI21X1  g12662(.A0(new_n12854_), .A1(new_n12853_), .B0(new_n12852_), .Y(new_n12855_));
  OAI21X1  g12663(.A0(new_n12855_), .A1(new_n1277_), .B0(new_n1111_), .Y(new_n12856_));
  OAI21X1  g12664(.A0(new_n12856_), .A1(new_n12836_), .B0(new_n12843_), .Y(new_n12857_));
  AOI21X1  g12665(.A0(new_n12857_), .A1(new_n12837_), .B0(new_n968_), .Y(new_n12858_));
  OR4X1    g12666(.A(new_n12447_), .B(new_n12308_), .C(new_n12296_), .D(new_n12290_), .Y(new_n12859_));
  OR2X1    g12667(.A(new_n12308_), .B(new_n12290_), .Y(new_n12860_));
  OAI21X1  g12668(.A0(new_n12860_), .A1(new_n12447_), .B0(new_n12296_), .Y(new_n12861_));
  AND2X1   g12669(.A(new_n12861_), .B(new_n12859_), .Y(new_n12862_));
  INVX1    g12670(.A(new_n12862_), .Y(new_n12863_));
  NAND3X1  g12671(.A(new_n12857_), .B(new_n12837_), .C(new_n968_), .Y(new_n12864_));
  AOI21X1  g12672(.A0(new_n12864_), .A1(new_n12863_), .B0(new_n12858_), .Y(new_n12865_));
  OR2X1    g12673(.A(new_n12865_), .B(new_n902_), .Y(new_n12866_));
  OR2X1    g12674(.A(new_n12855_), .B(new_n1277_), .Y(new_n12867_));
  NOR2X1   g12675(.A(new_n12826_), .B(new_n12825_), .Y(new_n12868_));
  INVX1    g12676(.A(new_n12834_), .Y(new_n12869_));
  NAND2X1  g12677(.A(new_n12821_), .B(new_n1277_), .Y(new_n12870_));
  OAI21X1  g12678(.A0(new_n12870_), .A1(new_n12868_), .B0(new_n12869_), .Y(new_n12871_));
  AOI21X1  g12679(.A0(new_n12871_), .A1(new_n12867_), .B0(new_n1111_), .Y(new_n12872_));
  AOI21X1  g12680(.A0(new_n12827_), .A1(\asqrt[51] ), .B0(\asqrt[52] ), .Y(new_n12873_));
  AOI21X1  g12681(.A0(new_n12873_), .A1(new_n12871_), .B0(new_n12842_), .Y(new_n12874_));
  NOR3X1   g12682(.A(new_n12874_), .B(new_n12872_), .C(\asqrt[53] ), .Y(new_n12875_));
  NOR2X1   g12683(.A(new_n12875_), .B(new_n12862_), .Y(new_n12876_));
  OAI21X1  g12684(.A0(new_n12317_), .A1(new_n12309_), .B0(new_n12314_), .Y(new_n12877_));
  NOR3X1   g12685(.A(new_n12877_), .B(new_n12447_), .C(new_n12350_), .Y(new_n12878_));
  AOI22X1  g12686(.A0(new_n12352_), .A1(new_n12351_), .B0(new_n12324_), .B1(\asqrt[53] ), .Y(new_n12879_));
  AOI21X1  g12687(.A0(new_n12879_), .A1(\asqrt[20] ), .B0(new_n12314_), .Y(new_n12880_));
  NOR2X1   g12688(.A(new_n12880_), .B(new_n12878_), .Y(new_n12881_));
  INVX1    g12689(.A(new_n12881_), .Y(new_n12882_));
  OAI21X1  g12690(.A0(new_n12874_), .A1(new_n12872_), .B0(\asqrt[53] ), .Y(new_n12883_));
  NAND2X1  g12691(.A(new_n12883_), .B(new_n902_), .Y(new_n12884_));
  OAI21X1  g12692(.A0(new_n12884_), .A1(new_n12876_), .B0(new_n12882_), .Y(new_n12885_));
  AOI21X1  g12693(.A0(new_n12885_), .A1(new_n12866_), .B0(new_n697_), .Y(new_n12886_));
  AND2X1   g12694(.A(new_n12325_), .B(new_n12318_), .Y(new_n12887_));
  OR4X1    g12695(.A(new_n12447_), .B(new_n12887_), .C(new_n12355_), .D(new_n12319_), .Y(new_n12888_));
  OR2X1    g12696(.A(new_n12887_), .B(new_n12319_), .Y(new_n12889_));
  OAI21X1  g12697(.A0(new_n12889_), .A1(new_n12447_), .B0(new_n12355_), .Y(new_n12890_));
  AND2X1   g12698(.A(new_n12890_), .B(new_n12888_), .Y(new_n12891_));
  OAI21X1  g12699(.A0(new_n12875_), .A1(new_n12862_), .B0(new_n12883_), .Y(new_n12892_));
  AOI21X1  g12700(.A0(new_n12892_), .A1(\asqrt[54] ), .B0(\asqrt[55] ), .Y(new_n12893_));
  AOI21X1  g12701(.A0(new_n12893_), .A1(new_n12885_), .B0(new_n12891_), .Y(new_n12894_));
  OAI21X1  g12702(.A0(new_n12894_), .A1(new_n12886_), .B0(\asqrt[56] ), .Y(new_n12895_));
  NAND3X1  g12703(.A(new_n12360_), .B(new_n12332_), .C(new_n12327_), .Y(new_n12896_));
  NOR3X1   g12704(.A(new_n12447_), .B(new_n12333_), .C(new_n12358_), .Y(new_n12897_));
  OAI22X1  g12705(.A0(new_n12897_), .A1(new_n12332_), .B0(new_n12896_), .B1(new_n12447_), .Y(new_n12898_));
  INVX1    g12706(.A(new_n12898_), .Y(new_n12899_));
  NOR3X1   g12707(.A(new_n12894_), .B(new_n12886_), .C(\asqrt[56] ), .Y(new_n12900_));
  OAI21X1  g12708(.A0(new_n12900_), .A1(new_n12899_), .B0(new_n12895_), .Y(new_n12901_));
  AND2X1   g12709(.A(new_n12901_), .B(\asqrt[57] ), .Y(new_n12902_));
  AND2X1   g12710(.A(new_n12892_), .B(\asqrt[54] ), .Y(new_n12903_));
  OR2X1    g12711(.A(new_n12875_), .B(new_n12862_), .Y(new_n12904_));
  AND2X1   g12712(.A(new_n12883_), .B(new_n902_), .Y(new_n12905_));
  AOI21X1  g12713(.A0(new_n12905_), .A1(new_n12904_), .B0(new_n12881_), .Y(new_n12906_));
  OAI21X1  g12714(.A0(new_n12906_), .A1(new_n12903_), .B0(\asqrt[55] ), .Y(new_n12907_));
  INVX1    g12715(.A(new_n12891_), .Y(new_n12908_));
  OAI21X1  g12716(.A0(new_n12865_), .A1(new_n902_), .B0(new_n697_), .Y(new_n12909_));
  OAI21X1  g12717(.A0(new_n12909_), .A1(new_n12906_), .B0(new_n12908_), .Y(new_n12910_));
  NAND3X1  g12718(.A(new_n12910_), .B(new_n12907_), .C(new_n582_), .Y(new_n12911_));
  NAND2X1  g12719(.A(new_n12911_), .B(new_n12898_), .Y(new_n12912_));
  AND2X1   g12720(.A(new_n12342_), .B(new_n12336_), .Y(new_n12913_));
  NOR4X1   g12721(.A(new_n12447_), .B(new_n12913_), .C(new_n12376_), .D(new_n12335_), .Y(new_n12914_));
  AOI22X1  g12722(.A0(new_n12342_), .A1(new_n12336_), .B0(new_n12334_), .B1(\asqrt[56] ), .Y(new_n12915_));
  AOI21X1  g12723(.A0(new_n12915_), .A1(\asqrt[20] ), .B0(new_n12341_), .Y(new_n12916_));
  NOR2X1   g12724(.A(new_n12916_), .B(new_n12914_), .Y(new_n12917_));
  AND2X1   g12725(.A(new_n12895_), .B(new_n481_), .Y(new_n12918_));
  AOI21X1  g12726(.A0(new_n12918_), .A1(new_n12912_), .B0(new_n12917_), .Y(new_n12919_));
  OAI21X1  g12727(.A0(new_n12919_), .A1(new_n12902_), .B0(\asqrt[58] ), .Y(new_n12920_));
  AND2X1   g12728(.A(new_n12380_), .B(new_n12378_), .Y(new_n12921_));
  OR4X1    g12729(.A(new_n12447_), .B(new_n12921_), .C(new_n12349_), .D(new_n12379_), .Y(new_n12922_));
  OR2X1    g12730(.A(new_n12921_), .B(new_n12379_), .Y(new_n12923_));
  OAI21X1  g12731(.A0(new_n12923_), .A1(new_n12447_), .B0(new_n12349_), .Y(new_n12924_));
  AND2X1   g12732(.A(new_n12924_), .B(new_n12922_), .Y(new_n12925_));
  INVX1    g12733(.A(new_n12925_), .Y(new_n12926_));
  AOI21X1  g12734(.A0(new_n12910_), .A1(new_n12907_), .B0(new_n582_), .Y(new_n12927_));
  AOI21X1  g12735(.A0(new_n12911_), .A1(new_n12898_), .B0(new_n12927_), .Y(new_n12928_));
  OAI21X1  g12736(.A0(new_n12928_), .A1(new_n481_), .B0(new_n399_), .Y(new_n12929_));
  OAI21X1  g12737(.A0(new_n12929_), .A1(new_n12919_), .B0(new_n12926_), .Y(new_n12930_));
  AOI21X1  g12738(.A0(new_n12930_), .A1(new_n12920_), .B0(new_n328_), .Y(new_n12931_));
  OR4X1    g12739(.A(new_n12447_), .B(new_n12382_), .C(new_n12370_), .D(new_n12364_), .Y(new_n12932_));
  OR2X1    g12740(.A(new_n12382_), .B(new_n12364_), .Y(new_n12933_));
  OAI21X1  g12741(.A0(new_n12933_), .A1(new_n12447_), .B0(new_n12370_), .Y(new_n12934_));
  AND2X1   g12742(.A(new_n12934_), .B(new_n12932_), .Y(new_n12935_));
  INVX1    g12743(.A(new_n12935_), .Y(new_n12936_));
  NAND3X1  g12744(.A(new_n12930_), .B(new_n12920_), .C(new_n328_), .Y(new_n12937_));
  AOI21X1  g12745(.A0(new_n12937_), .A1(new_n12936_), .B0(new_n12931_), .Y(new_n12938_));
  OR2X1    g12746(.A(new_n12938_), .B(new_n292_), .Y(new_n12939_));
  OR2X1    g12747(.A(new_n12928_), .B(new_n481_), .Y(new_n12940_));
  AND2X1   g12748(.A(new_n12911_), .B(new_n12898_), .Y(new_n12941_));
  INVX1    g12749(.A(new_n12917_), .Y(new_n12942_));
  NAND2X1  g12750(.A(new_n12895_), .B(new_n481_), .Y(new_n12943_));
  OAI21X1  g12751(.A0(new_n12943_), .A1(new_n12941_), .B0(new_n12942_), .Y(new_n12944_));
  AOI21X1  g12752(.A0(new_n12944_), .A1(new_n12940_), .B0(new_n399_), .Y(new_n12945_));
  AOI21X1  g12753(.A0(new_n12901_), .A1(\asqrt[57] ), .B0(\asqrt[58] ), .Y(new_n12946_));
  AOI21X1  g12754(.A0(new_n12946_), .A1(new_n12944_), .B0(new_n12925_), .Y(new_n12947_));
  NOR3X1   g12755(.A(new_n12947_), .B(new_n12945_), .C(\asqrt[59] ), .Y(new_n12948_));
  NOR2X1   g12756(.A(new_n12948_), .B(new_n12935_), .Y(new_n12949_));
  OAI21X1  g12757(.A0(new_n12391_), .A1(new_n12383_), .B0(new_n12388_), .Y(new_n12950_));
  NOR3X1   g12758(.A(new_n12950_), .B(new_n12447_), .C(new_n12411_), .Y(new_n12951_));
  AOI22X1  g12759(.A0(new_n12413_), .A1(new_n12412_), .B0(new_n12398_), .B1(\asqrt[59] ), .Y(new_n12952_));
  AOI21X1  g12760(.A0(new_n12952_), .A1(\asqrt[20] ), .B0(new_n12388_), .Y(new_n12953_));
  NOR2X1   g12761(.A(new_n12953_), .B(new_n12951_), .Y(new_n12954_));
  INVX1    g12762(.A(new_n12954_), .Y(new_n12955_));
  OAI21X1  g12763(.A0(new_n12947_), .A1(new_n12945_), .B0(\asqrt[59] ), .Y(new_n12956_));
  NAND2X1  g12764(.A(new_n12956_), .B(new_n292_), .Y(new_n12957_));
  OAI21X1  g12765(.A0(new_n12957_), .A1(new_n12949_), .B0(new_n12955_), .Y(new_n12958_));
  AOI21X1  g12766(.A0(new_n12958_), .A1(new_n12939_), .B0(new_n217_), .Y(new_n12959_));
  AND2X1   g12767(.A(new_n12399_), .B(new_n12392_), .Y(new_n12960_));
  OR4X1    g12768(.A(new_n12447_), .B(new_n12960_), .C(new_n12416_), .D(new_n12393_), .Y(new_n12961_));
  OR2X1    g12769(.A(new_n12960_), .B(new_n12393_), .Y(new_n12962_));
  OAI21X1  g12770(.A0(new_n12962_), .A1(new_n12447_), .B0(new_n12416_), .Y(new_n12963_));
  AND2X1   g12771(.A(new_n12963_), .B(new_n12961_), .Y(new_n12964_));
  OAI21X1  g12772(.A0(new_n12948_), .A1(new_n12935_), .B0(new_n12956_), .Y(new_n12965_));
  AOI21X1  g12773(.A0(new_n12965_), .A1(\asqrt[60] ), .B0(\asqrt[61] ), .Y(new_n12966_));
  AOI21X1  g12774(.A0(new_n12966_), .A1(new_n12958_), .B0(new_n12964_), .Y(new_n12967_));
  OAI21X1  g12775(.A0(new_n12967_), .A1(new_n12959_), .B0(\asqrt[62] ), .Y(new_n12968_));
  OR4X1    g12776(.A(new_n12447_), .B(new_n12407_), .C(new_n12410_), .D(new_n12436_), .Y(new_n12969_));
  OR2X1    g12777(.A(new_n12407_), .B(new_n12436_), .Y(new_n12970_));
  OAI21X1  g12778(.A0(new_n12970_), .A1(new_n12447_), .B0(new_n12410_), .Y(new_n12971_));
  AND2X1   g12779(.A(new_n12971_), .B(new_n12969_), .Y(new_n12972_));
  NOR3X1   g12780(.A(new_n12967_), .B(new_n12959_), .C(\asqrt[62] ), .Y(new_n12973_));
  OAI21X1  g12781(.A0(new_n12973_), .A1(new_n12972_), .B0(new_n12968_), .Y(new_n12974_));
  AND2X1   g12782(.A(new_n12426_), .B(new_n12420_), .Y(new_n12975_));
  NOR4X1   g12783(.A(new_n12447_), .B(new_n12975_), .C(new_n12450_), .D(new_n12409_), .Y(new_n12976_));
  INVX1    g12784(.A(new_n12976_), .Y(new_n12977_));
  OAI22X1  g12785(.A0(new_n12451_), .A1(new_n12449_), .B0(new_n12437_), .B1(new_n199_), .Y(new_n12978_));
  OAI21X1  g12786(.A0(new_n12978_), .A1(new_n12447_), .B0(new_n12450_), .Y(new_n12979_));
  AND2X1   g12787(.A(new_n12979_), .B(new_n12977_), .Y(new_n12980_));
  INVX1    g12788(.A(new_n12980_), .Y(new_n12981_));
  AND2X1   g12789(.A(new_n12455_), .B(new_n12452_), .Y(new_n12982_));
  AOI21X1  g12790(.A0(new_n12452_), .A1(new_n12448_), .B0(new_n12430_), .Y(new_n12983_));
  AOI21X1  g12791(.A0(new_n12983_), .A1(\asqrt[20] ), .B0(new_n12982_), .Y(new_n12984_));
  AND2X1   g12792(.A(new_n12984_), .B(new_n12981_), .Y(new_n12985_));
  AOI21X1  g12793(.A0(new_n12985_), .A1(new_n12974_), .B0(\asqrt[63] ), .Y(new_n12986_));
  NOR2X1   g12794(.A(new_n12973_), .B(new_n12972_), .Y(new_n12987_));
  NAND2X1  g12795(.A(new_n12980_), .B(new_n12968_), .Y(new_n12988_));
  NAND2X1  g12796(.A(new_n12452_), .B(new_n12448_), .Y(new_n12989_));
  AOI21X1  g12797(.A0(\asqrt[20] ), .A1(new_n12431_), .B0(new_n12989_), .Y(new_n12990_));
  NOR3X1   g12798(.A(new_n12990_), .B(new_n12983_), .C(new_n193_), .Y(new_n12991_));
  AND2X1   g12799(.A(new_n12435_), .B(new_n193_), .Y(new_n12992_));
  INVX1    g12800(.A(new_n12444_), .Y(new_n12993_));
  OR2X1    g12801(.A(new_n12993_), .B(new_n12428_), .Y(new_n12994_));
  AOI21X1  g12802(.A0(new_n12429_), .A1(new_n11916_), .B0(new_n12994_), .Y(new_n12995_));
  NAND2X1  g12803(.A(new_n12995_), .B(new_n12441_), .Y(new_n12996_));
  NOR3X1   g12804(.A(new_n12996_), .B(new_n12982_), .C(new_n12992_), .Y(new_n12997_));
  NOR2X1   g12805(.A(new_n12997_), .B(new_n12991_), .Y(new_n12998_));
  OAI21X1  g12806(.A0(new_n12988_), .A1(new_n12987_), .B0(new_n12998_), .Y(new_n12999_));
  NOR2X1   g12807(.A(new_n12999_), .B(new_n12986_), .Y(new_n13000_));
  INVX1    g12808(.A(new_n13000_), .Y(\asqrt[19] ));
  OAI21X1  g12809(.A0(new_n12999_), .A1(new_n12986_), .B0(\a[38] ), .Y(new_n13002_));
  INVX1    g12810(.A(\a[38] ), .Y(new_n13003_));
  NOR2X1   g12811(.A(\a[37] ), .B(\a[36] ), .Y(new_n13004_));
  NAND2X1  g12812(.A(new_n13004_), .B(new_n13003_), .Y(new_n13005_));
  AND2X1   g12813(.A(new_n13005_), .B(new_n13002_), .Y(new_n13006_));
  AND2X1   g12814(.A(new_n12965_), .B(\asqrt[60] ), .Y(new_n13007_));
  OR2X1    g12815(.A(new_n12948_), .B(new_n12935_), .Y(new_n13008_));
  AND2X1   g12816(.A(new_n12956_), .B(new_n292_), .Y(new_n13009_));
  AOI21X1  g12817(.A0(new_n13009_), .A1(new_n13008_), .B0(new_n12954_), .Y(new_n13010_));
  OAI21X1  g12818(.A0(new_n13010_), .A1(new_n13007_), .B0(\asqrt[61] ), .Y(new_n13011_));
  INVX1    g12819(.A(new_n12964_), .Y(new_n13012_));
  OAI21X1  g12820(.A0(new_n12938_), .A1(new_n292_), .B0(new_n217_), .Y(new_n13013_));
  OAI21X1  g12821(.A0(new_n13013_), .A1(new_n13010_), .B0(new_n13012_), .Y(new_n13014_));
  AOI21X1  g12822(.A0(new_n13014_), .A1(new_n13011_), .B0(new_n199_), .Y(new_n13015_));
  INVX1    g12823(.A(new_n12972_), .Y(new_n13016_));
  NAND3X1  g12824(.A(new_n13014_), .B(new_n13011_), .C(new_n199_), .Y(new_n13017_));
  AOI21X1  g12825(.A0(new_n13017_), .A1(new_n13016_), .B0(new_n13015_), .Y(new_n13018_));
  INVX1    g12826(.A(new_n12985_), .Y(new_n13019_));
  OAI21X1  g12827(.A0(new_n13019_), .A1(new_n13018_), .B0(new_n193_), .Y(new_n13020_));
  OR2X1    g12828(.A(new_n12973_), .B(new_n12972_), .Y(new_n13021_));
  AND2X1   g12829(.A(new_n12980_), .B(new_n12968_), .Y(new_n13022_));
  INVX1    g12830(.A(new_n12998_), .Y(new_n13023_));
  AOI21X1  g12831(.A0(new_n13022_), .A1(new_n13021_), .B0(new_n13023_), .Y(new_n13024_));
  AOI21X1  g12832(.A0(new_n13024_), .A1(new_n13020_), .B0(new_n13003_), .Y(new_n13025_));
  NAND3X1  g12833(.A(new_n13005_), .B(new_n12444_), .C(new_n12441_), .Y(new_n13026_));
  NOR4X1   g12834(.A(new_n13026_), .B(new_n13025_), .C(new_n12982_), .D(new_n12992_), .Y(new_n13027_));
  INVX1    g12835(.A(\a[39] ), .Y(new_n13028_));
  AOI21X1  g12836(.A0(new_n13024_), .A1(new_n13020_), .B0(\a[38] ), .Y(new_n13029_));
  OAI21X1  g12837(.A0(new_n12999_), .A1(new_n12986_), .B0(new_n12459_), .Y(new_n13030_));
  OAI21X1  g12838(.A0(new_n13029_), .A1(new_n13028_), .B0(new_n13030_), .Y(new_n13031_));
  OAI22X1  g12839(.A0(new_n13031_), .A1(new_n13027_), .B0(new_n13006_), .B1(new_n12447_), .Y(new_n13032_));
  AND2X1   g12840(.A(new_n13032_), .B(\asqrt[21] ), .Y(new_n13033_));
  OR4X1    g12841(.A(new_n13026_), .B(new_n13025_), .C(new_n12982_), .D(new_n12992_), .Y(new_n13034_));
  OAI21X1  g12842(.A0(new_n12999_), .A1(new_n12986_), .B0(new_n13003_), .Y(new_n13035_));
  AOI21X1  g12843(.A0(new_n13024_), .A1(new_n13020_), .B0(new_n12473_), .Y(new_n13036_));
  AOI21X1  g12844(.A0(new_n13035_), .A1(\a[39] ), .B0(new_n13036_), .Y(new_n13037_));
  NAND2X1  g12845(.A(new_n13037_), .B(new_n13034_), .Y(new_n13038_));
  AOI21X1  g12846(.A0(new_n13005_), .A1(new_n13002_), .B0(new_n12447_), .Y(new_n13039_));
  NOR2X1   g12847(.A(new_n13039_), .B(\asqrt[21] ), .Y(new_n13040_));
  AND2X1   g12848(.A(new_n13022_), .B(new_n13021_), .Y(new_n13041_));
  OR2X1    g12849(.A(new_n12997_), .B(new_n12447_), .Y(new_n13042_));
  OR4X1    g12850(.A(new_n13042_), .B(new_n12991_), .C(new_n13041_), .D(new_n12986_), .Y(new_n13043_));
  AOI21X1  g12851(.A0(new_n13043_), .A1(new_n13030_), .B0(new_n12466_), .Y(new_n13044_));
  NOR4X1   g12852(.A(new_n13042_), .B(new_n12991_), .C(new_n13041_), .D(new_n12986_), .Y(new_n13045_));
  NOR3X1   g12853(.A(new_n13045_), .B(new_n13036_), .C(\a[40] ), .Y(new_n13046_));
  NOR2X1   g12854(.A(new_n13046_), .B(new_n13044_), .Y(new_n13047_));
  AOI21X1  g12855(.A0(new_n13040_), .A1(new_n13038_), .B0(new_n13047_), .Y(new_n13048_));
  OAI21X1  g12856(.A0(new_n13048_), .A1(new_n13033_), .B0(\asqrt[22] ), .Y(new_n13049_));
  AND2X1   g12857(.A(new_n12514_), .B(new_n12512_), .Y(new_n13050_));
  NOR3X1   g12858(.A(new_n13050_), .B(new_n12465_), .C(new_n12461_), .Y(new_n13051_));
  OAI21X1  g12859(.A0(new_n12999_), .A1(new_n12986_), .B0(new_n13051_), .Y(new_n13052_));
  AOI21X1  g12860(.A0(new_n12460_), .A1(\asqrt[21] ), .B0(new_n12465_), .Y(new_n13053_));
  OAI21X1  g12861(.A0(new_n12999_), .A1(new_n12986_), .B0(new_n13053_), .Y(new_n13054_));
  NAND2X1  g12862(.A(new_n13054_), .B(new_n13050_), .Y(new_n13055_));
  NAND2X1  g12863(.A(new_n13055_), .B(new_n13052_), .Y(new_n13056_));
  AOI21X1  g12864(.A0(new_n13037_), .A1(new_n13034_), .B0(new_n13039_), .Y(new_n13057_));
  OAI21X1  g12865(.A0(new_n13057_), .A1(new_n11896_), .B0(new_n11362_), .Y(new_n13058_));
  OAI21X1  g12866(.A0(new_n13058_), .A1(new_n13048_), .B0(new_n13056_), .Y(new_n13059_));
  AOI21X1  g12867(.A0(new_n13059_), .A1(new_n13049_), .B0(new_n10849_), .Y(new_n13060_));
  AND2X1   g12868(.A(new_n12517_), .B(new_n12515_), .Y(new_n13061_));
  NOR3X1   g12869(.A(new_n12482_), .B(new_n13061_), .C(new_n12516_), .Y(new_n13062_));
  OAI21X1  g12870(.A0(new_n12999_), .A1(new_n12986_), .B0(new_n13062_), .Y(new_n13063_));
  NOR2X1   g12871(.A(new_n13061_), .B(new_n12516_), .Y(new_n13064_));
  OAI21X1  g12872(.A0(new_n12999_), .A1(new_n12986_), .B0(new_n13064_), .Y(new_n13065_));
  NAND2X1  g12873(.A(new_n13065_), .B(new_n12482_), .Y(new_n13066_));
  AND2X1   g12874(.A(new_n13066_), .B(new_n13063_), .Y(new_n13067_));
  INVX1    g12875(.A(new_n13067_), .Y(new_n13068_));
  NAND3X1  g12876(.A(new_n13059_), .B(new_n13049_), .C(new_n10849_), .Y(new_n13069_));
  AOI21X1  g12877(.A0(new_n13069_), .A1(new_n13068_), .B0(new_n13060_), .Y(new_n13070_));
  OR2X1    g12878(.A(new_n13070_), .B(new_n10332_), .Y(new_n13071_));
  OR2X1    g12879(.A(new_n13057_), .B(new_n11896_), .Y(new_n13072_));
  AND2X1   g12880(.A(new_n13037_), .B(new_n13034_), .Y(new_n13073_));
  OR2X1    g12881(.A(new_n13039_), .B(\asqrt[21] ), .Y(new_n13074_));
  OR2X1    g12882(.A(new_n13046_), .B(new_n13044_), .Y(new_n13075_));
  OAI21X1  g12883(.A0(new_n13074_), .A1(new_n13073_), .B0(new_n13075_), .Y(new_n13076_));
  AOI21X1  g12884(.A0(new_n13076_), .A1(new_n13072_), .B0(new_n11362_), .Y(new_n13077_));
  AOI21X1  g12885(.A0(new_n13032_), .A1(\asqrt[21] ), .B0(\asqrt[22] ), .Y(new_n13078_));
  AOI22X1  g12886(.A0(new_n13078_), .A1(new_n13076_), .B0(new_n13055_), .B1(new_n13052_), .Y(new_n13079_));
  NOR3X1   g12887(.A(new_n13079_), .B(new_n13077_), .C(\asqrt[23] ), .Y(new_n13080_));
  NOR2X1   g12888(.A(new_n13080_), .B(new_n13067_), .Y(new_n13081_));
  NOR3X1   g12889(.A(new_n12522_), .B(new_n12490_), .C(new_n12484_), .Y(new_n13082_));
  NAND3X1  g12890(.A(\asqrt[19] ), .B(new_n12491_), .C(new_n12521_), .Y(new_n13083_));
  AOI22X1  g12891(.A0(new_n13083_), .A1(new_n12490_), .B0(new_n13082_), .B1(\asqrt[19] ), .Y(new_n13084_));
  INVX1    g12892(.A(new_n13084_), .Y(new_n13085_));
  OR2X1    g12893(.A(new_n13060_), .B(\asqrt[24] ), .Y(new_n13086_));
  OAI21X1  g12894(.A0(new_n13086_), .A1(new_n13081_), .B0(new_n13085_), .Y(new_n13087_));
  AOI21X1  g12895(.A0(new_n13087_), .A1(new_n13071_), .B0(new_n9833_), .Y(new_n13088_));
  AOI21X1  g12896(.A0(new_n12537_), .A1(new_n12536_), .B0(new_n12500_), .Y(new_n13089_));
  AND2X1   g12897(.A(new_n13089_), .B(new_n12493_), .Y(new_n13090_));
  AOI22X1  g12898(.A0(new_n12537_), .A1(new_n12536_), .B0(new_n12523_), .B1(\asqrt[24] ), .Y(new_n13091_));
  AOI21X1  g12899(.A0(new_n13091_), .A1(\asqrt[19] ), .B0(new_n12499_), .Y(new_n13092_));
  AOI21X1  g12900(.A0(new_n13090_), .A1(\asqrt[19] ), .B0(new_n13092_), .Y(new_n13093_));
  OAI21X1  g12901(.A0(new_n13079_), .A1(new_n13077_), .B0(\asqrt[23] ), .Y(new_n13094_));
  OAI21X1  g12902(.A0(new_n13080_), .A1(new_n13067_), .B0(new_n13094_), .Y(new_n13095_));
  AOI21X1  g12903(.A0(new_n13095_), .A1(\asqrt[24] ), .B0(\asqrt[25] ), .Y(new_n13096_));
  AOI21X1  g12904(.A0(new_n13096_), .A1(new_n13087_), .B0(new_n13093_), .Y(new_n13097_));
  OAI21X1  g12905(.A0(new_n13097_), .A1(new_n13088_), .B0(\asqrt[26] ), .Y(new_n13098_));
  AND2X1   g12906(.A(new_n12524_), .B(new_n12502_), .Y(new_n13099_));
  NOR3X1   g12907(.A(new_n13099_), .B(new_n12540_), .C(new_n12503_), .Y(new_n13100_));
  NOR3X1   g12908(.A(new_n13000_), .B(new_n13099_), .C(new_n12503_), .Y(new_n13101_));
  NOR2X1   g12909(.A(new_n13101_), .B(new_n12508_), .Y(new_n13102_));
  AOI21X1  g12910(.A0(new_n13100_), .A1(\asqrt[19] ), .B0(new_n13102_), .Y(new_n13103_));
  NOR3X1   g12911(.A(new_n13097_), .B(new_n13088_), .C(\asqrt[26] ), .Y(new_n13104_));
  OAI21X1  g12912(.A0(new_n13104_), .A1(new_n13103_), .B0(new_n13098_), .Y(new_n13105_));
  AND2X1   g12913(.A(new_n13105_), .B(\asqrt[27] ), .Y(new_n13106_));
  OR2X1    g12914(.A(new_n13104_), .B(new_n13103_), .Y(new_n13107_));
  NAND4X1  g12915(.A(\asqrt[19] ), .B(new_n12543_), .C(new_n12530_), .D(new_n12526_), .Y(new_n13108_));
  NAND2X1  g12916(.A(new_n12543_), .B(new_n12526_), .Y(new_n13109_));
  OAI21X1  g12917(.A0(new_n13109_), .A1(new_n13000_), .B0(new_n12534_), .Y(new_n13110_));
  AND2X1   g12918(.A(new_n13110_), .B(new_n13108_), .Y(new_n13111_));
  AND2X1   g12919(.A(new_n13098_), .B(new_n8874_), .Y(new_n13112_));
  AOI21X1  g12920(.A0(new_n13112_), .A1(new_n13107_), .B0(new_n13111_), .Y(new_n13113_));
  OAI21X1  g12921(.A0(new_n13113_), .A1(new_n13106_), .B0(\asqrt[28] ), .Y(new_n13114_));
  AND2X1   g12922(.A(new_n12551_), .B(new_n12544_), .Y(new_n13115_));
  NOR3X1   g12923(.A(new_n13115_), .B(new_n12589_), .C(new_n12533_), .Y(new_n13116_));
  NOR3X1   g12924(.A(new_n13000_), .B(new_n13115_), .C(new_n12533_), .Y(new_n13117_));
  NOR2X1   g12925(.A(new_n13117_), .B(new_n12549_), .Y(new_n13118_));
  AOI21X1  g12926(.A0(new_n13116_), .A1(\asqrt[19] ), .B0(new_n13118_), .Y(new_n13119_));
  INVX1    g12927(.A(new_n13119_), .Y(new_n13120_));
  AND2X1   g12928(.A(new_n13095_), .B(\asqrt[24] ), .Y(new_n13121_));
  OR2X1    g12929(.A(new_n13080_), .B(new_n13067_), .Y(new_n13122_));
  NOR2X1   g12930(.A(new_n13060_), .B(\asqrt[24] ), .Y(new_n13123_));
  AOI21X1  g12931(.A0(new_n13123_), .A1(new_n13122_), .B0(new_n13084_), .Y(new_n13124_));
  OAI21X1  g12932(.A0(new_n13124_), .A1(new_n13121_), .B0(\asqrt[25] ), .Y(new_n13125_));
  INVX1    g12933(.A(new_n13093_), .Y(new_n13126_));
  OAI21X1  g12934(.A0(new_n13070_), .A1(new_n10332_), .B0(new_n9833_), .Y(new_n13127_));
  OAI21X1  g12935(.A0(new_n13127_), .A1(new_n13124_), .B0(new_n13126_), .Y(new_n13128_));
  AOI21X1  g12936(.A0(new_n13128_), .A1(new_n13125_), .B0(new_n9353_), .Y(new_n13129_));
  INVX1    g12937(.A(new_n13103_), .Y(new_n13130_));
  NAND3X1  g12938(.A(new_n13128_), .B(new_n13125_), .C(new_n9353_), .Y(new_n13131_));
  AOI21X1  g12939(.A0(new_n13131_), .A1(new_n13130_), .B0(new_n13129_), .Y(new_n13132_));
  OAI21X1  g12940(.A0(new_n13132_), .A1(new_n8874_), .B0(new_n8412_), .Y(new_n13133_));
  OAI21X1  g12941(.A0(new_n13133_), .A1(new_n13113_), .B0(new_n13120_), .Y(new_n13134_));
  AOI21X1  g12942(.A0(new_n13134_), .A1(new_n13114_), .B0(new_n7970_), .Y(new_n13135_));
  AND2X1   g12943(.A(new_n12593_), .B(new_n12591_), .Y(new_n13136_));
  NOR3X1   g12944(.A(new_n13136_), .B(new_n12559_), .C(new_n12592_), .Y(new_n13137_));
  NOR3X1   g12945(.A(new_n13000_), .B(new_n13136_), .C(new_n12592_), .Y(new_n13138_));
  NOR2X1   g12946(.A(new_n13138_), .B(new_n12558_), .Y(new_n13139_));
  AOI21X1  g12947(.A0(new_n13137_), .A1(\asqrt[19] ), .B0(new_n13139_), .Y(new_n13140_));
  INVX1    g12948(.A(new_n13140_), .Y(new_n13141_));
  NAND3X1  g12949(.A(new_n13134_), .B(new_n13114_), .C(new_n7970_), .Y(new_n13142_));
  AOI21X1  g12950(.A0(new_n13142_), .A1(new_n13141_), .B0(new_n13135_), .Y(new_n13143_));
  OR2X1    g12951(.A(new_n13143_), .B(new_n7527_), .Y(new_n13144_));
  OR2X1    g12952(.A(new_n13132_), .B(new_n8874_), .Y(new_n13145_));
  NOR2X1   g12953(.A(new_n13104_), .B(new_n13103_), .Y(new_n13146_));
  INVX1    g12954(.A(new_n13111_), .Y(new_n13147_));
  NAND2X1  g12955(.A(new_n13098_), .B(new_n8874_), .Y(new_n13148_));
  OAI21X1  g12956(.A0(new_n13148_), .A1(new_n13146_), .B0(new_n13147_), .Y(new_n13149_));
  AOI21X1  g12957(.A0(new_n13149_), .A1(new_n13145_), .B0(new_n8412_), .Y(new_n13150_));
  AOI21X1  g12958(.A0(new_n13105_), .A1(\asqrt[27] ), .B0(\asqrt[28] ), .Y(new_n13151_));
  AOI21X1  g12959(.A0(new_n13151_), .A1(new_n13149_), .B0(new_n13119_), .Y(new_n13152_));
  NOR3X1   g12960(.A(new_n13152_), .B(new_n13150_), .C(\asqrt[29] ), .Y(new_n13153_));
  NOR2X1   g12961(.A(new_n13153_), .B(new_n13140_), .Y(new_n13154_));
  NAND4X1  g12962(.A(\asqrt[19] ), .B(new_n12569_), .C(new_n12567_), .D(new_n12595_), .Y(new_n13155_));
  NAND2X1  g12963(.A(new_n12569_), .B(new_n12595_), .Y(new_n13156_));
  OAI21X1  g12964(.A0(new_n13156_), .A1(new_n13000_), .B0(new_n12568_), .Y(new_n13157_));
  AND2X1   g12965(.A(new_n13157_), .B(new_n13155_), .Y(new_n13158_));
  INVX1    g12966(.A(new_n13158_), .Y(new_n13159_));
  OAI21X1  g12967(.A0(new_n13152_), .A1(new_n13150_), .B0(\asqrt[29] ), .Y(new_n13160_));
  NAND2X1  g12968(.A(new_n13160_), .B(new_n7527_), .Y(new_n13161_));
  OAI21X1  g12969(.A0(new_n13161_), .A1(new_n13154_), .B0(new_n13159_), .Y(new_n13162_));
  AOI21X1  g12970(.A0(new_n13162_), .A1(new_n13144_), .B0(new_n7103_), .Y(new_n13163_));
  AOI21X1  g12971(.A0(new_n12611_), .A1(new_n12610_), .B0(new_n12578_), .Y(new_n13164_));
  AND2X1   g12972(.A(new_n13164_), .B(new_n12571_), .Y(new_n13165_));
  AOI22X1  g12973(.A0(new_n12611_), .A1(new_n12610_), .B0(new_n12597_), .B1(\asqrt[30] ), .Y(new_n13166_));
  AOI21X1  g12974(.A0(new_n13166_), .A1(\asqrt[19] ), .B0(new_n12577_), .Y(new_n13167_));
  AOI21X1  g12975(.A0(new_n13165_), .A1(\asqrt[19] ), .B0(new_n13167_), .Y(new_n13168_));
  OAI21X1  g12976(.A0(new_n13153_), .A1(new_n13140_), .B0(new_n13160_), .Y(new_n13169_));
  AOI21X1  g12977(.A0(new_n13169_), .A1(\asqrt[30] ), .B0(\asqrt[31] ), .Y(new_n13170_));
  AOI21X1  g12978(.A0(new_n13170_), .A1(new_n13162_), .B0(new_n13168_), .Y(new_n13171_));
  OAI21X1  g12979(.A0(new_n13171_), .A1(new_n13163_), .B0(\asqrt[32] ), .Y(new_n13172_));
  AND2X1   g12980(.A(new_n12598_), .B(new_n12580_), .Y(new_n13173_));
  NOR3X1   g12981(.A(new_n13173_), .B(new_n12614_), .C(new_n12581_), .Y(new_n13174_));
  NOR3X1   g12982(.A(new_n13000_), .B(new_n13173_), .C(new_n12581_), .Y(new_n13175_));
  NOR2X1   g12983(.A(new_n13175_), .B(new_n12586_), .Y(new_n13176_));
  AOI21X1  g12984(.A0(new_n13174_), .A1(\asqrt[19] ), .B0(new_n13176_), .Y(new_n13177_));
  NOR3X1   g12985(.A(new_n13171_), .B(new_n13163_), .C(\asqrt[32] ), .Y(new_n13178_));
  OAI21X1  g12986(.A0(new_n13178_), .A1(new_n13177_), .B0(new_n13172_), .Y(new_n13179_));
  AND2X1   g12987(.A(new_n13179_), .B(\asqrt[33] ), .Y(new_n13180_));
  INVX1    g12988(.A(new_n13177_), .Y(new_n13181_));
  AND2X1   g12989(.A(new_n13169_), .B(\asqrt[30] ), .Y(new_n13182_));
  OR2X1    g12990(.A(new_n13153_), .B(new_n13140_), .Y(new_n13183_));
  AND2X1   g12991(.A(new_n13160_), .B(new_n7527_), .Y(new_n13184_));
  AOI21X1  g12992(.A0(new_n13184_), .A1(new_n13183_), .B0(new_n13158_), .Y(new_n13185_));
  OAI21X1  g12993(.A0(new_n13185_), .A1(new_n13182_), .B0(\asqrt[31] ), .Y(new_n13186_));
  INVX1    g12994(.A(new_n13168_), .Y(new_n13187_));
  OAI21X1  g12995(.A0(new_n13143_), .A1(new_n7527_), .B0(new_n7103_), .Y(new_n13188_));
  OAI21X1  g12996(.A0(new_n13188_), .A1(new_n13185_), .B0(new_n13187_), .Y(new_n13189_));
  NAND3X1  g12997(.A(new_n13189_), .B(new_n13186_), .C(new_n6699_), .Y(new_n13190_));
  NAND2X1  g12998(.A(new_n13190_), .B(new_n13181_), .Y(new_n13191_));
  NAND4X1  g12999(.A(\asqrt[19] ), .B(new_n12617_), .C(new_n12604_), .D(new_n12600_), .Y(new_n13192_));
  NAND2X1  g13000(.A(new_n12617_), .B(new_n12600_), .Y(new_n13193_));
  OAI21X1  g13001(.A0(new_n13193_), .A1(new_n13000_), .B0(new_n12608_), .Y(new_n13194_));
  AND2X1   g13002(.A(new_n13194_), .B(new_n13192_), .Y(new_n13195_));
  AOI21X1  g13003(.A0(new_n13189_), .A1(new_n13186_), .B0(new_n6699_), .Y(new_n13196_));
  NOR2X1   g13004(.A(new_n13196_), .B(\asqrt[33] ), .Y(new_n13197_));
  AOI21X1  g13005(.A0(new_n13197_), .A1(new_n13191_), .B0(new_n13195_), .Y(new_n13198_));
  OAI21X1  g13006(.A0(new_n13198_), .A1(new_n13180_), .B0(\asqrt[34] ), .Y(new_n13199_));
  AND2X1   g13007(.A(new_n12625_), .B(new_n12618_), .Y(new_n13200_));
  NOR3X1   g13008(.A(new_n13200_), .B(new_n12663_), .C(new_n12607_), .Y(new_n13201_));
  NOR3X1   g13009(.A(new_n13000_), .B(new_n13200_), .C(new_n12607_), .Y(new_n13202_));
  NOR2X1   g13010(.A(new_n13202_), .B(new_n12623_), .Y(new_n13203_));
  AOI21X1  g13011(.A0(new_n13201_), .A1(\asqrt[19] ), .B0(new_n13203_), .Y(new_n13204_));
  INVX1    g13012(.A(new_n13204_), .Y(new_n13205_));
  AOI21X1  g13013(.A0(new_n13190_), .A1(new_n13181_), .B0(new_n13196_), .Y(new_n13206_));
  OAI21X1  g13014(.A0(new_n13206_), .A1(new_n6294_), .B0(new_n5941_), .Y(new_n13207_));
  OAI21X1  g13015(.A0(new_n13207_), .A1(new_n13198_), .B0(new_n13205_), .Y(new_n13208_));
  AOI21X1  g13016(.A0(new_n13208_), .A1(new_n13199_), .B0(new_n5541_), .Y(new_n13209_));
  AND2X1   g13017(.A(new_n12667_), .B(new_n12665_), .Y(new_n13210_));
  NOR3X1   g13018(.A(new_n13210_), .B(new_n12633_), .C(new_n12666_), .Y(new_n13211_));
  NOR3X1   g13019(.A(new_n13000_), .B(new_n13210_), .C(new_n12666_), .Y(new_n13212_));
  NOR2X1   g13020(.A(new_n13212_), .B(new_n12632_), .Y(new_n13213_));
  AOI21X1  g13021(.A0(new_n13211_), .A1(\asqrt[19] ), .B0(new_n13213_), .Y(new_n13214_));
  INVX1    g13022(.A(new_n13214_), .Y(new_n13215_));
  NAND3X1  g13023(.A(new_n13208_), .B(new_n13199_), .C(new_n5541_), .Y(new_n13216_));
  AOI21X1  g13024(.A0(new_n13216_), .A1(new_n13215_), .B0(new_n13209_), .Y(new_n13217_));
  OR2X1    g13025(.A(new_n13217_), .B(new_n5176_), .Y(new_n13218_));
  OR2X1    g13026(.A(new_n13206_), .B(new_n6294_), .Y(new_n13219_));
  AND2X1   g13027(.A(new_n13190_), .B(new_n13181_), .Y(new_n13220_));
  INVX1    g13028(.A(new_n13195_), .Y(new_n13221_));
  OR2X1    g13029(.A(new_n13196_), .B(\asqrt[33] ), .Y(new_n13222_));
  OAI21X1  g13030(.A0(new_n13222_), .A1(new_n13220_), .B0(new_n13221_), .Y(new_n13223_));
  AOI21X1  g13031(.A0(new_n13223_), .A1(new_n13219_), .B0(new_n5941_), .Y(new_n13224_));
  AOI21X1  g13032(.A0(new_n13179_), .A1(\asqrt[33] ), .B0(\asqrt[34] ), .Y(new_n13225_));
  AOI21X1  g13033(.A0(new_n13225_), .A1(new_n13223_), .B0(new_n13204_), .Y(new_n13226_));
  NOR3X1   g13034(.A(new_n13226_), .B(new_n13224_), .C(\asqrt[35] ), .Y(new_n13227_));
  NOR2X1   g13035(.A(new_n13227_), .B(new_n13214_), .Y(new_n13228_));
  NAND4X1  g13036(.A(\asqrt[19] ), .B(new_n12643_), .C(new_n12641_), .D(new_n12669_), .Y(new_n13229_));
  NAND2X1  g13037(.A(new_n12643_), .B(new_n12669_), .Y(new_n13230_));
  OAI21X1  g13038(.A0(new_n13230_), .A1(new_n13000_), .B0(new_n12642_), .Y(new_n13231_));
  AND2X1   g13039(.A(new_n13231_), .B(new_n13229_), .Y(new_n13232_));
  INVX1    g13040(.A(new_n13232_), .Y(new_n13233_));
  OR2X1    g13041(.A(new_n13209_), .B(\asqrt[36] ), .Y(new_n13234_));
  OAI21X1  g13042(.A0(new_n13234_), .A1(new_n13228_), .B0(new_n13233_), .Y(new_n13235_));
  AOI21X1  g13043(.A0(new_n13235_), .A1(new_n13218_), .B0(new_n4826_), .Y(new_n13236_));
  AOI21X1  g13044(.A0(new_n12685_), .A1(new_n12684_), .B0(new_n12652_), .Y(new_n13237_));
  AND2X1   g13045(.A(new_n13237_), .B(new_n12645_), .Y(new_n13238_));
  AOI22X1  g13046(.A0(new_n12685_), .A1(new_n12684_), .B0(new_n12671_), .B1(\asqrt[36] ), .Y(new_n13239_));
  AOI21X1  g13047(.A0(new_n13239_), .A1(\asqrt[19] ), .B0(new_n12651_), .Y(new_n13240_));
  AOI21X1  g13048(.A0(new_n13238_), .A1(\asqrt[19] ), .B0(new_n13240_), .Y(new_n13241_));
  OAI21X1  g13049(.A0(new_n13226_), .A1(new_n13224_), .B0(\asqrt[35] ), .Y(new_n13242_));
  OAI21X1  g13050(.A0(new_n13227_), .A1(new_n13214_), .B0(new_n13242_), .Y(new_n13243_));
  AOI21X1  g13051(.A0(new_n13243_), .A1(\asqrt[36] ), .B0(\asqrt[37] ), .Y(new_n13244_));
  AOI21X1  g13052(.A0(new_n13244_), .A1(new_n13235_), .B0(new_n13241_), .Y(new_n13245_));
  OAI21X1  g13053(.A0(new_n13245_), .A1(new_n13236_), .B0(\asqrt[38] ), .Y(new_n13246_));
  AND2X1   g13054(.A(new_n12672_), .B(new_n12654_), .Y(new_n13247_));
  NOR3X1   g13055(.A(new_n13247_), .B(new_n12688_), .C(new_n12655_), .Y(new_n13248_));
  NOR3X1   g13056(.A(new_n13000_), .B(new_n13247_), .C(new_n12655_), .Y(new_n13249_));
  NOR2X1   g13057(.A(new_n13249_), .B(new_n12660_), .Y(new_n13250_));
  AOI21X1  g13058(.A0(new_n13248_), .A1(\asqrt[19] ), .B0(new_n13250_), .Y(new_n13251_));
  NOR3X1   g13059(.A(new_n13245_), .B(new_n13236_), .C(\asqrt[38] ), .Y(new_n13252_));
  OAI21X1  g13060(.A0(new_n13252_), .A1(new_n13251_), .B0(new_n13246_), .Y(new_n13253_));
  AND2X1   g13061(.A(new_n13253_), .B(\asqrt[39] ), .Y(new_n13254_));
  INVX1    g13062(.A(new_n13251_), .Y(new_n13255_));
  AND2X1   g13063(.A(new_n13243_), .B(\asqrt[36] ), .Y(new_n13256_));
  OR2X1    g13064(.A(new_n13227_), .B(new_n13214_), .Y(new_n13257_));
  NOR2X1   g13065(.A(new_n13209_), .B(\asqrt[36] ), .Y(new_n13258_));
  AOI21X1  g13066(.A0(new_n13258_), .A1(new_n13257_), .B0(new_n13232_), .Y(new_n13259_));
  OAI21X1  g13067(.A0(new_n13259_), .A1(new_n13256_), .B0(\asqrt[37] ), .Y(new_n13260_));
  INVX1    g13068(.A(new_n13241_), .Y(new_n13261_));
  OAI21X1  g13069(.A0(new_n13217_), .A1(new_n5176_), .B0(new_n4826_), .Y(new_n13262_));
  OAI21X1  g13070(.A0(new_n13262_), .A1(new_n13259_), .B0(new_n13261_), .Y(new_n13263_));
  NAND3X1  g13071(.A(new_n13263_), .B(new_n13260_), .C(new_n4493_), .Y(new_n13264_));
  NAND2X1  g13072(.A(new_n13264_), .B(new_n13255_), .Y(new_n13265_));
  NAND4X1  g13073(.A(\asqrt[19] ), .B(new_n12691_), .C(new_n12678_), .D(new_n12674_), .Y(new_n13266_));
  NAND2X1  g13074(.A(new_n12691_), .B(new_n12674_), .Y(new_n13267_));
  OAI21X1  g13075(.A0(new_n13267_), .A1(new_n13000_), .B0(new_n12682_), .Y(new_n13268_));
  AND2X1   g13076(.A(new_n13268_), .B(new_n13266_), .Y(new_n13269_));
  AOI21X1  g13077(.A0(new_n13263_), .A1(new_n13260_), .B0(new_n4493_), .Y(new_n13270_));
  NOR2X1   g13078(.A(new_n13270_), .B(\asqrt[39] ), .Y(new_n13271_));
  AOI21X1  g13079(.A0(new_n13271_), .A1(new_n13265_), .B0(new_n13269_), .Y(new_n13272_));
  OAI21X1  g13080(.A0(new_n13272_), .A1(new_n13254_), .B0(\asqrt[40] ), .Y(new_n13273_));
  AND2X1   g13081(.A(new_n12699_), .B(new_n12692_), .Y(new_n13274_));
  NOR3X1   g13082(.A(new_n13274_), .B(new_n12722_), .C(new_n12681_), .Y(new_n13275_));
  NOR3X1   g13083(.A(new_n13000_), .B(new_n13274_), .C(new_n12681_), .Y(new_n13276_));
  NOR2X1   g13084(.A(new_n13276_), .B(new_n12697_), .Y(new_n13277_));
  AOI21X1  g13085(.A0(new_n13275_), .A1(\asqrt[19] ), .B0(new_n13277_), .Y(new_n13278_));
  INVX1    g13086(.A(new_n13278_), .Y(new_n13279_));
  AOI21X1  g13087(.A0(new_n13264_), .A1(new_n13255_), .B0(new_n13270_), .Y(new_n13280_));
  OAI21X1  g13088(.A0(new_n13280_), .A1(new_n4165_), .B0(new_n3863_), .Y(new_n13281_));
  OAI21X1  g13089(.A0(new_n13281_), .A1(new_n13272_), .B0(new_n13279_), .Y(new_n13282_));
  AOI21X1  g13090(.A0(new_n13282_), .A1(new_n13273_), .B0(new_n3564_), .Y(new_n13283_));
  AND2X1   g13091(.A(new_n12726_), .B(new_n12724_), .Y(new_n13284_));
  NOR3X1   g13092(.A(new_n13284_), .B(new_n12707_), .C(new_n12725_), .Y(new_n13285_));
  NOR3X1   g13093(.A(new_n13000_), .B(new_n13284_), .C(new_n12725_), .Y(new_n13286_));
  NOR2X1   g13094(.A(new_n13286_), .B(new_n12706_), .Y(new_n13287_));
  AOI21X1  g13095(.A0(new_n13285_), .A1(\asqrt[19] ), .B0(new_n13287_), .Y(new_n13288_));
  INVX1    g13096(.A(new_n13288_), .Y(new_n13289_));
  NAND3X1  g13097(.A(new_n13282_), .B(new_n13273_), .C(new_n3564_), .Y(new_n13290_));
  AOI21X1  g13098(.A0(new_n13290_), .A1(new_n13289_), .B0(new_n13283_), .Y(new_n13291_));
  OR2X1    g13099(.A(new_n13291_), .B(new_n3276_), .Y(new_n13292_));
  OR2X1    g13100(.A(new_n13280_), .B(new_n4165_), .Y(new_n13293_));
  AND2X1   g13101(.A(new_n13264_), .B(new_n13255_), .Y(new_n13294_));
  INVX1    g13102(.A(new_n13269_), .Y(new_n13295_));
  OR2X1    g13103(.A(new_n13270_), .B(\asqrt[39] ), .Y(new_n13296_));
  OAI21X1  g13104(.A0(new_n13296_), .A1(new_n13294_), .B0(new_n13295_), .Y(new_n13297_));
  AOI21X1  g13105(.A0(new_n13297_), .A1(new_n13293_), .B0(new_n3863_), .Y(new_n13298_));
  AOI21X1  g13106(.A0(new_n13253_), .A1(\asqrt[39] ), .B0(\asqrt[40] ), .Y(new_n13299_));
  AOI21X1  g13107(.A0(new_n13299_), .A1(new_n13297_), .B0(new_n13278_), .Y(new_n13300_));
  NOR3X1   g13108(.A(new_n13300_), .B(new_n13298_), .C(\asqrt[41] ), .Y(new_n13301_));
  NOR2X1   g13109(.A(new_n13301_), .B(new_n13288_), .Y(new_n13302_));
  OR4X1    g13110(.A(new_n13000_), .B(new_n12728_), .C(new_n12716_), .D(new_n12711_), .Y(new_n13303_));
  OR2X1    g13111(.A(new_n12728_), .B(new_n12711_), .Y(new_n13304_));
  OAI21X1  g13112(.A0(new_n13304_), .A1(new_n13000_), .B0(new_n12716_), .Y(new_n13305_));
  AND2X1   g13113(.A(new_n13305_), .B(new_n13303_), .Y(new_n13306_));
  INVX1    g13114(.A(new_n13306_), .Y(new_n13307_));
  OAI21X1  g13115(.A0(new_n13300_), .A1(new_n13298_), .B0(\asqrt[41] ), .Y(new_n13308_));
  NAND2X1  g13116(.A(new_n13308_), .B(new_n3276_), .Y(new_n13309_));
  OAI21X1  g13117(.A0(new_n13309_), .A1(new_n13302_), .B0(new_n13307_), .Y(new_n13310_));
  AOI21X1  g13118(.A0(new_n13310_), .A1(new_n13292_), .B0(new_n3008_), .Y(new_n13311_));
  AOI21X1  g13119(.A0(new_n12773_), .A1(new_n12772_), .B0(new_n12735_), .Y(new_n13312_));
  AND2X1   g13120(.A(new_n13312_), .B(new_n12719_), .Y(new_n13313_));
  AOI22X1  g13121(.A0(new_n12773_), .A1(new_n12772_), .B0(new_n12745_), .B1(\asqrt[42] ), .Y(new_n13314_));
  AOI21X1  g13122(.A0(new_n13314_), .A1(\asqrt[19] ), .B0(new_n12734_), .Y(new_n13315_));
  AOI21X1  g13123(.A0(new_n13313_), .A1(\asqrt[19] ), .B0(new_n13315_), .Y(new_n13316_));
  OAI21X1  g13124(.A0(new_n13301_), .A1(new_n13288_), .B0(new_n13308_), .Y(new_n13317_));
  AOI21X1  g13125(.A0(new_n13317_), .A1(\asqrt[42] ), .B0(\asqrt[43] ), .Y(new_n13318_));
  AOI21X1  g13126(.A0(new_n13318_), .A1(new_n13310_), .B0(new_n13316_), .Y(new_n13319_));
  OAI21X1  g13127(.A0(new_n13319_), .A1(new_n13311_), .B0(\asqrt[44] ), .Y(new_n13320_));
  AND2X1   g13128(.A(new_n12746_), .B(new_n12738_), .Y(new_n13321_));
  NOR3X1   g13129(.A(new_n13321_), .B(new_n12776_), .C(new_n12739_), .Y(new_n13322_));
  NOR3X1   g13130(.A(new_n13000_), .B(new_n13321_), .C(new_n12739_), .Y(new_n13323_));
  NOR2X1   g13131(.A(new_n13323_), .B(new_n12744_), .Y(new_n13324_));
  AOI21X1  g13132(.A0(new_n13322_), .A1(\asqrt[19] ), .B0(new_n13324_), .Y(new_n13325_));
  NOR3X1   g13133(.A(new_n13319_), .B(new_n13311_), .C(\asqrt[44] ), .Y(new_n13326_));
  OAI21X1  g13134(.A0(new_n13326_), .A1(new_n13325_), .B0(new_n13320_), .Y(new_n13327_));
  AND2X1   g13135(.A(new_n13327_), .B(\asqrt[45] ), .Y(new_n13328_));
  OR2X1    g13136(.A(new_n13326_), .B(new_n13325_), .Y(new_n13329_));
  OR4X1    g13137(.A(new_n13000_), .B(new_n12753_), .C(new_n12780_), .D(new_n12779_), .Y(new_n13330_));
  OR2X1    g13138(.A(new_n12753_), .B(new_n12779_), .Y(new_n13331_));
  OAI21X1  g13139(.A0(new_n13331_), .A1(new_n13000_), .B0(new_n12780_), .Y(new_n13332_));
  AND2X1   g13140(.A(new_n13332_), .B(new_n13330_), .Y(new_n13333_));
  AND2X1   g13141(.A(new_n13320_), .B(new_n2570_), .Y(new_n13334_));
  AOI21X1  g13142(.A0(new_n13334_), .A1(new_n13329_), .B0(new_n13333_), .Y(new_n13335_));
  OAI21X1  g13143(.A0(new_n13335_), .A1(new_n13328_), .B0(\asqrt[46] ), .Y(new_n13336_));
  AND2X1   g13144(.A(new_n13317_), .B(\asqrt[42] ), .Y(new_n13337_));
  OR2X1    g13145(.A(new_n13301_), .B(new_n13288_), .Y(new_n13338_));
  AND2X1   g13146(.A(new_n13308_), .B(new_n3276_), .Y(new_n13339_));
  AOI21X1  g13147(.A0(new_n13339_), .A1(new_n13338_), .B0(new_n13306_), .Y(new_n13340_));
  OAI21X1  g13148(.A0(new_n13340_), .A1(new_n13337_), .B0(\asqrt[43] ), .Y(new_n13341_));
  INVX1    g13149(.A(new_n13316_), .Y(new_n13342_));
  OAI21X1  g13150(.A0(new_n13291_), .A1(new_n3276_), .B0(new_n3008_), .Y(new_n13343_));
  OAI21X1  g13151(.A0(new_n13343_), .A1(new_n13340_), .B0(new_n13342_), .Y(new_n13344_));
  AOI21X1  g13152(.A0(new_n13344_), .A1(new_n13341_), .B0(new_n2769_), .Y(new_n13345_));
  INVX1    g13153(.A(new_n13325_), .Y(new_n13346_));
  NAND3X1  g13154(.A(new_n13344_), .B(new_n13341_), .C(new_n2769_), .Y(new_n13347_));
  AOI21X1  g13155(.A0(new_n13347_), .A1(new_n13346_), .B0(new_n13345_), .Y(new_n13348_));
  OAI21X1  g13156(.A0(new_n13348_), .A1(new_n2570_), .B0(new_n2263_), .Y(new_n13349_));
  AND2X1   g13157(.A(new_n12757_), .B(new_n12756_), .Y(new_n13350_));
  NOR3X1   g13158(.A(new_n12802_), .B(new_n13350_), .C(new_n12755_), .Y(new_n13351_));
  NOR3X1   g13159(.A(new_n13000_), .B(new_n13350_), .C(new_n12755_), .Y(new_n13352_));
  NOR2X1   g13160(.A(new_n13352_), .B(new_n12762_), .Y(new_n13353_));
  AOI21X1  g13161(.A0(new_n13351_), .A1(\asqrt[19] ), .B0(new_n13353_), .Y(new_n13354_));
  INVX1    g13162(.A(new_n13354_), .Y(new_n13355_));
  OAI21X1  g13163(.A0(new_n13349_), .A1(new_n13335_), .B0(new_n13355_), .Y(new_n13356_));
  AOI21X1  g13164(.A0(new_n13356_), .A1(new_n13336_), .B0(new_n2040_), .Y(new_n13357_));
  AND2X1   g13165(.A(new_n12805_), .B(new_n12803_), .Y(new_n13358_));
  NOR3X1   g13166(.A(new_n13358_), .B(new_n12770_), .C(new_n12804_), .Y(new_n13359_));
  NOR3X1   g13167(.A(new_n13000_), .B(new_n13358_), .C(new_n12804_), .Y(new_n13360_));
  NOR2X1   g13168(.A(new_n13360_), .B(new_n12769_), .Y(new_n13361_));
  AOI21X1  g13169(.A0(new_n13359_), .A1(\asqrt[19] ), .B0(new_n13361_), .Y(new_n13362_));
  INVX1    g13170(.A(new_n13362_), .Y(new_n13363_));
  NAND3X1  g13171(.A(new_n13356_), .B(new_n13336_), .C(new_n2040_), .Y(new_n13364_));
  AOI21X1  g13172(.A0(new_n13364_), .A1(new_n13363_), .B0(new_n13357_), .Y(new_n13365_));
  OR2X1    g13173(.A(new_n13365_), .B(new_n1834_), .Y(new_n13366_));
  OR2X1    g13174(.A(new_n13348_), .B(new_n2570_), .Y(new_n13367_));
  NOR2X1   g13175(.A(new_n13326_), .B(new_n13325_), .Y(new_n13368_));
  INVX1    g13176(.A(new_n13333_), .Y(new_n13369_));
  NAND2X1  g13177(.A(new_n13320_), .B(new_n2570_), .Y(new_n13370_));
  OAI21X1  g13178(.A0(new_n13370_), .A1(new_n13368_), .B0(new_n13369_), .Y(new_n13371_));
  AOI21X1  g13179(.A0(new_n13371_), .A1(new_n13367_), .B0(new_n2263_), .Y(new_n13372_));
  AOI21X1  g13180(.A0(new_n13327_), .A1(\asqrt[45] ), .B0(\asqrt[46] ), .Y(new_n13373_));
  AOI21X1  g13181(.A0(new_n13373_), .A1(new_n13371_), .B0(new_n13354_), .Y(new_n13374_));
  NOR3X1   g13182(.A(new_n13374_), .B(new_n13372_), .C(\asqrt[47] ), .Y(new_n13375_));
  NOR2X1   g13183(.A(new_n13375_), .B(new_n13362_), .Y(new_n13376_));
  OR4X1    g13184(.A(new_n13000_), .B(new_n12817_), .C(new_n12788_), .D(new_n12785_), .Y(new_n13377_));
  OR2X1    g13185(.A(new_n12817_), .B(new_n12785_), .Y(new_n13378_));
  OAI21X1  g13186(.A0(new_n13378_), .A1(new_n13000_), .B0(new_n12788_), .Y(new_n13379_));
  AND2X1   g13187(.A(new_n13379_), .B(new_n13377_), .Y(new_n13380_));
  INVX1    g13188(.A(new_n13380_), .Y(new_n13381_));
  OAI21X1  g13189(.A0(new_n13374_), .A1(new_n13372_), .B0(\asqrt[47] ), .Y(new_n13382_));
  NAND2X1  g13190(.A(new_n13382_), .B(new_n1834_), .Y(new_n13383_));
  OAI21X1  g13191(.A0(new_n13383_), .A1(new_n13376_), .B0(new_n13381_), .Y(new_n13384_));
  AOI21X1  g13192(.A0(new_n13384_), .A1(new_n13366_), .B0(new_n1632_), .Y(new_n13385_));
  AOI21X1  g13193(.A0(new_n12846_), .A1(new_n12845_), .B0(new_n12798_), .Y(new_n13386_));
  AND2X1   g13194(.A(new_n13386_), .B(new_n12791_), .Y(new_n13387_));
  AOI22X1  g13195(.A0(new_n12846_), .A1(new_n12845_), .B0(new_n12818_), .B1(\asqrt[48] ), .Y(new_n13388_));
  AOI21X1  g13196(.A0(new_n13388_), .A1(\asqrt[19] ), .B0(new_n12797_), .Y(new_n13389_));
  AOI21X1  g13197(.A0(new_n13387_), .A1(\asqrt[19] ), .B0(new_n13389_), .Y(new_n13390_));
  OAI21X1  g13198(.A0(new_n13375_), .A1(new_n13362_), .B0(new_n13382_), .Y(new_n13391_));
  AOI21X1  g13199(.A0(new_n13391_), .A1(\asqrt[48] ), .B0(\asqrt[49] ), .Y(new_n13392_));
  AOI21X1  g13200(.A0(new_n13392_), .A1(new_n13384_), .B0(new_n13390_), .Y(new_n13393_));
  OAI21X1  g13201(.A0(new_n13393_), .A1(new_n13385_), .B0(\asqrt[50] ), .Y(new_n13394_));
  AND2X1   g13202(.A(new_n12819_), .B(new_n12809_), .Y(new_n13395_));
  NOR3X1   g13203(.A(new_n13395_), .B(new_n12849_), .C(new_n12810_), .Y(new_n13396_));
  NOR3X1   g13204(.A(new_n13000_), .B(new_n13395_), .C(new_n12810_), .Y(new_n13397_));
  NOR2X1   g13205(.A(new_n13397_), .B(new_n12815_), .Y(new_n13398_));
  AOI21X1  g13206(.A0(new_n13396_), .A1(\asqrt[19] ), .B0(new_n13398_), .Y(new_n13399_));
  NOR3X1   g13207(.A(new_n13393_), .B(new_n13385_), .C(\asqrt[50] ), .Y(new_n13400_));
  OAI21X1  g13208(.A0(new_n13400_), .A1(new_n13399_), .B0(new_n13394_), .Y(new_n13401_));
  AND2X1   g13209(.A(new_n13401_), .B(\asqrt[51] ), .Y(new_n13402_));
  OR2X1    g13210(.A(new_n13400_), .B(new_n13399_), .Y(new_n13403_));
  OR4X1    g13211(.A(new_n13000_), .B(new_n12826_), .C(new_n12853_), .D(new_n12852_), .Y(new_n13404_));
  OR2X1    g13212(.A(new_n12826_), .B(new_n12852_), .Y(new_n13405_));
  OAI21X1  g13213(.A0(new_n13405_), .A1(new_n13000_), .B0(new_n12853_), .Y(new_n13406_));
  AND2X1   g13214(.A(new_n13406_), .B(new_n13404_), .Y(new_n13407_));
  AND2X1   g13215(.A(new_n13394_), .B(new_n1277_), .Y(new_n13408_));
  AOI21X1  g13216(.A0(new_n13408_), .A1(new_n13403_), .B0(new_n13407_), .Y(new_n13409_));
  OAI21X1  g13217(.A0(new_n13409_), .A1(new_n13402_), .B0(\asqrt[52] ), .Y(new_n13410_));
  AND2X1   g13218(.A(new_n12835_), .B(new_n12829_), .Y(new_n13411_));
  NOR3X1   g13219(.A(new_n13411_), .B(new_n12869_), .C(new_n12828_), .Y(new_n13412_));
  NOR3X1   g13220(.A(new_n13000_), .B(new_n13411_), .C(new_n12828_), .Y(new_n13413_));
  NOR2X1   g13221(.A(new_n13413_), .B(new_n12834_), .Y(new_n13414_));
  AOI21X1  g13222(.A0(new_n13412_), .A1(\asqrt[19] ), .B0(new_n13414_), .Y(new_n13415_));
  INVX1    g13223(.A(new_n13415_), .Y(new_n13416_));
  AND2X1   g13224(.A(new_n13391_), .B(\asqrt[48] ), .Y(new_n13417_));
  OR2X1    g13225(.A(new_n13375_), .B(new_n13362_), .Y(new_n13418_));
  AND2X1   g13226(.A(new_n13382_), .B(new_n1834_), .Y(new_n13419_));
  AOI21X1  g13227(.A0(new_n13419_), .A1(new_n13418_), .B0(new_n13380_), .Y(new_n13420_));
  OAI21X1  g13228(.A0(new_n13420_), .A1(new_n13417_), .B0(\asqrt[49] ), .Y(new_n13421_));
  INVX1    g13229(.A(new_n13390_), .Y(new_n13422_));
  OAI21X1  g13230(.A0(new_n13365_), .A1(new_n1834_), .B0(new_n1632_), .Y(new_n13423_));
  OAI21X1  g13231(.A0(new_n13423_), .A1(new_n13420_), .B0(new_n13422_), .Y(new_n13424_));
  AOI21X1  g13232(.A0(new_n13424_), .A1(new_n13421_), .B0(new_n1469_), .Y(new_n13425_));
  INVX1    g13233(.A(new_n13399_), .Y(new_n13426_));
  NAND3X1  g13234(.A(new_n13424_), .B(new_n13421_), .C(new_n1469_), .Y(new_n13427_));
  AOI21X1  g13235(.A0(new_n13427_), .A1(new_n13426_), .B0(new_n13425_), .Y(new_n13428_));
  OAI21X1  g13236(.A0(new_n13428_), .A1(new_n1277_), .B0(new_n1111_), .Y(new_n13429_));
  OAI21X1  g13237(.A0(new_n13429_), .A1(new_n13409_), .B0(new_n13416_), .Y(new_n13430_));
  AOI21X1  g13238(.A0(new_n13430_), .A1(new_n13410_), .B0(new_n968_), .Y(new_n13431_));
  AND2X1   g13239(.A(new_n12873_), .B(new_n12871_), .Y(new_n13432_));
  NOR3X1   g13240(.A(new_n13432_), .B(new_n12843_), .C(new_n12872_), .Y(new_n13433_));
  NOR3X1   g13241(.A(new_n13000_), .B(new_n13432_), .C(new_n12872_), .Y(new_n13434_));
  NOR2X1   g13242(.A(new_n13434_), .B(new_n12842_), .Y(new_n13435_));
  AOI21X1  g13243(.A0(new_n13433_), .A1(\asqrt[19] ), .B0(new_n13435_), .Y(new_n13436_));
  INVX1    g13244(.A(new_n13436_), .Y(new_n13437_));
  NAND3X1  g13245(.A(new_n13430_), .B(new_n13410_), .C(new_n968_), .Y(new_n13438_));
  AOI21X1  g13246(.A0(new_n13438_), .A1(new_n13437_), .B0(new_n13431_), .Y(new_n13439_));
  OR2X1    g13247(.A(new_n13439_), .B(new_n902_), .Y(new_n13440_));
  OR2X1    g13248(.A(new_n13428_), .B(new_n1277_), .Y(new_n13441_));
  NOR2X1   g13249(.A(new_n13400_), .B(new_n13399_), .Y(new_n13442_));
  INVX1    g13250(.A(new_n13407_), .Y(new_n13443_));
  NAND2X1  g13251(.A(new_n13394_), .B(new_n1277_), .Y(new_n13444_));
  OAI21X1  g13252(.A0(new_n13444_), .A1(new_n13442_), .B0(new_n13443_), .Y(new_n13445_));
  AOI21X1  g13253(.A0(new_n13445_), .A1(new_n13441_), .B0(new_n1111_), .Y(new_n13446_));
  AOI21X1  g13254(.A0(new_n13401_), .A1(\asqrt[51] ), .B0(\asqrt[52] ), .Y(new_n13447_));
  AOI21X1  g13255(.A0(new_n13447_), .A1(new_n13445_), .B0(new_n13415_), .Y(new_n13448_));
  NOR3X1   g13256(.A(new_n13448_), .B(new_n13446_), .C(\asqrt[53] ), .Y(new_n13449_));
  NOR2X1   g13257(.A(new_n13449_), .B(new_n13436_), .Y(new_n13450_));
  OR4X1    g13258(.A(new_n13000_), .B(new_n12875_), .C(new_n12863_), .D(new_n12858_), .Y(new_n13451_));
  OR2X1    g13259(.A(new_n12875_), .B(new_n12858_), .Y(new_n13452_));
  OAI21X1  g13260(.A0(new_n13452_), .A1(new_n13000_), .B0(new_n12863_), .Y(new_n13453_));
  AND2X1   g13261(.A(new_n13453_), .B(new_n13451_), .Y(new_n13454_));
  INVX1    g13262(.A(new_n13454_), .Y(new_n13455_));
  OAI21X1  g13263(.A0(new_n13448_), .A1(new_n13446_), .B0(\asqrt[53] ), .Y(new_n13456_));
  NAND2X1  g13264(.A(new_n13456_), .B(new_n902_), .Y(new_n13457_));
  OAI21X1  g13265(.A0(new_n13457_), .A1(new_n13450_), .B0(new_n13455_), .Y(new_n13458_));
  AOI21X1  g13266(.A0(new_n13458_), .A1(new_n13440_), .B0(new_n697_), .Y(new_n13459_));
  AOI21X1  g13267(.A0(new_n12905_), .A1(new_n12904_), .B0(new_n12882_), .Y(new_n13460_));
  AND2X1   g13268(.A(new_n13460_), .B(new_n12866_), .Y(new_n13461_));
  AOI22X1  g13269(.A0(new_n12905_), .A1(new_n12904_), .B0(new_n12892_), .B1(\asqrt[54] ), .Y(new_n13462_));
  AOI21X1  g13270(.A0(new_n13462_), .A1(\asqrt[19] ), .B0(new_n12881_), .Y(new_n13463_));
  AOI21X1  g13271(.A0(new_n13461_), .A1(\asqrt[19] ), .B0(new_n13463_), .Y(new_n13464_));
  OAI21X1  g13272(.A0(new_n13449_), .A1(new_n13436_), .B0(new_n13456_), .Y(new_n13465_));
  AOI21X1  g13273(.A0(new_n13465_), .A1(\asqrt[54] ), .B0(\asqrt[55] ), .Y(new_n13466_));
  AOI21X1  g13274(.A0(new_n13466_), .A1(new_n13458_), .B0(new_n13464_), .Y(new_n13467_));
  OAI21X1  g13275(.A0(new_n13467_), .A1(new_n13459_), .B0(\asqrt[56] ), .Y(new_n13468_));
  AND2X1   g13276(.A(new_n12893_), .B(new_n12885_), .Y(new_n13469_));
  NOR3X1   g13277(.A(new_n13469_), .B(new_n12908_), .C(new_n12886_), .Y(new_n13470_));
  NOR3X1   g13278(.A(new_n13000_), .B(new_n13469_), .C(new_n12886_), .Y(new_n13471_));
  NOR2X1   g13279(.A(new_n13471_), .B(new_n12891_), .Y(new_n13472_));
  AOI21X1  g13280(.A0(new_n13470_), .A1(\asqrt[19] ), .B0(new_n13472_), .Y(new_n13473_));
  NOR3X1   g13281(.A(new_n13467_), .B(new_n13459_), .C(\asqrt[56] ), .Y(new_n13474_));
  OAI21X1  g13282(.A0(new_n13474_), .A1(new_n13473_), .B0(new_n13468_), .Y(new_n13475_));
  AND2X1   g13283(.A(new_n13475_), .B(\asqrt[57] ), .Y(new_n13476_));
  OR2X1    g13284(.A(new_n13474_), .B(new_n13473_), .Y(new_n13477_));
  OR4X1    g13285(.A(new_n13000_), .B(new_n12900_), .C(new_n12898_), .D(new_n12927_), .Y(new_n13478_));
  OR2X1    g13286(.A(new_n12900_), .B(new_n12927_), .Y(new_n13479_));
  OAI21X1  g13287(.A0(new_n13479_), .A1(new_n13000_), .B0(new_n12898_), .Y(new_n13480_));
  AND2X1   g13288(.A(new_n13480_), .B(new_n13478_), .Y(new_n13481_));
  AND2X1   g13289(.A(new_n13468_), .B(new_n481_), .Y(new_n13482_));
  AOI21X1  g13290(.A0(new_n13482_), .A1(new_n13477_), .B0(new_n13481_), .Y(new_n13483_));
  OAI21X1  g13291(.A0(new_n13483_), .A1(new_n13476_), .B0(\asqrt[58] ), .Y(new_n13484_));
  AND2X1   g13292(.A(new_n12918_), .B(new_n12912_), .Y(new_n13485_));
  NOR3X1   g13293(.A(new_n13485_), .B(new_n12942_), .C(new_n12902_), .Y(new_n13486_));
  NOR3X1   g13294(.A(new_n13000_), .B(new_n13485_), .C(new_n12902_), .Y(new_n13487_));
  NOR2X1   g13295(.A(new_n13487_), .B(new_n12917_), .Y(new_n13488_));
  AOI21X1  g13296(.A0(new_n13486_), .A1(\asqrt[19] ), .B0(new_n13488_), .Y(new_n13489_));
  INVX1    g13297(.A(new_n13489_), .Y(new_n13490_));
  AND2X1   g13298(.A(new_n13465_), .B(\asqrt[54] ), .Y(new_n13491_));
  OR2X1    g13299(.A(new_n13449_), .B(new_n13436_), .Y(new_n13492_));
  AND2X1   g13300(.A(new_n13456_), .B(new_n902_), .Y(new_n13493_));
  AOI21X1  g13301(.A0(new_n13493_), .A1(new_n13492_), .B0(new_n13454_), .Y(new_n13494_));
  OAI21X1  g13302(.A0(new_n13494_), .A1(new_n13491_), .B0(\asqrt[55] ), .Y(new_n13495_));
  INVX1    g13303(.A(new_n13464_), .Y(new_n13496_));
  OAI21X1  g13304(.A0(new_n13439_), .A1(new_n902_), .B0(new_n697_), .Y(new_n13497_));
  OAI21X1  g13305(.A0(new_n13497_), .A1(new_n13494_), .B0(new_n13496_), .Y(new_n13498_));
  AOI21X1  g13306(.A0(new_n13498_), .A1(new_n13495_), .B0(new_n582_), .Y(new_n13499_));
  INVX1    g13307(.A(new_n13473_), .Y(new_n13500_));
  NAND3X1  g13308(.A(new_n13498_), .B(new_n13495_), .C(new_n582_), .Y(new_n13501_));
  AOI21X1  g13309(.A0(new_n13501_), .A1(new_n13500_), .B0(new_n13499_), .Y(new_n13502_));
  OAI21X1  g13310(.A0(new_n13502_), .A1(new_n481_), .B0(new_n399_), .Y(new_n13503_));
  OAI21X1  g13311(.A0(new_n13503_), .A1(new_n13483_), .B0(new_n13490_), .Y(new_n13504_));
  AOI21X1  g13312(.A0(new_n13504_), .A1(new_n13484_), .B0(new_n328_), .Y(new_n13505_));
  AND2X1   g13313(.A(new_n12946_), .B(new_n12944_), .Y(new_n13506_));
  NOR3X1   g13314(.A(new_n13506_), .B(new_n12926_), .C(new_n12945_), .Y(new_n13507_));
  NOR3X1   g13315(.A(new_n13000_), .B(new_n13506_), .C(new_n12945_), .Y(new_n13508_));
  NOR2X1   g13316(.A(new_n13508_), .B(new_n12925_), .Y(new_n13509_));
  AOI21X1  g13317(.A0(new_n13507_), .A1(\asqrt[19] ), .B0(new_n13509_), .Y(new_n13510_));
  INVX1    g13318(.A(new_n13510_), .Y(new_n13511_));
  NAND3X1  g13319(.A(new_n13504_), .B(new_n13484_), .C(new_n328_), .Y(new_n13512_));
  AOI21X1  g13320(.A0(new_n13512_), .A1(new_n13511_), .B0(new_n13505_), .Y(new_n13513_));
  OR2X1    g13321(.A(new_n13513_), .B(new_n292_), .Y(new_n13514_));
  OR2X1    g13322(.A(new_n13502_), .B(new_n481_), .Y(new_n13515_));
  NOR2X1   g13323(.A(new_n13474_), .B(new_n13473_), .Y(new_n13516_));
  INVX1    g13324(.A(new_n13481_), .Y(new_n13517_));
  NAND2X1  g13325(.A(new_n13468_), .B(new_n481_), .Y(new_n13518_));
  OAI21X1  g13326(.A0(new_n13518_), .A1(new_n13516_), .B0(new_n13517_), .Y(new_n13519_));
  AOI21X1  g13327(.A0(new_n13519_), .A1(new_n13515_), .B0(new_n399_), .Y(new_n13520_));
  AOI21X1  g13328(.A0(new_n13475_), .A1(\asqrt[57] ), .B0(\asqrt[58] ), .Y(new_n13521_));
  AOI21X1  g13329(.A0(new_n13521_), .A1(new_n13519_), .B0(new_n13489_), .Y(new_n13522_));
  NOR3X1   g13330(.A(new_n13522_), .B(new_n13520_), .C(\asqrt[59] ), .Y(new_n13523_));
  NOR2X1   g13331(.A(new_n13523_), .B(new_n13510_), .Y(new_n13524_));
  OR4X1    g13332(.A(new_n13000_), .B(new_n12948_), .C(new_n12936_), .D(new_n12931_), .Y(new_n13525_));
  OR2X1    g13333(.A(new_n12948_), .B(new_n12931_), .Y(new_n13526_));
  OAI21X1  g13334(.A0(new_n13526_), .A1(new_n13000_), .B0(new_n12936_), .Y(new_n13527_));
  AND2X1   g13335(.A(new_n13527_), .B(new_n13525_), .Y(new_n13528_));
  INVX1    g13336(.A(new_n13528_), .Y(new_n13529_));
  OAI21X1  g13337(.A0(new_n13522_), .A1(new_n13520_), .B0(\asqrt[59] ), .Y(new_n13530_));
  NAND2X1  g13338(.A(new_n13530_), .B(new_n292_), .Y(new_n13531_));
  OAI21X1  g13339(.A0(new_n13531_), .A1(new_n13524_), .B0(new_n13529_), .Y(new_n13532_));
  AOI21X1  g13340(.A0(new_n13532_), .A1(new_n13514_), .B0(new_n217_), .Y(new_n13533_));
  AOI21X1  g13341(.A0(new_n13009_), .A1(new_n13008_), .B0(new_n12955_), .Y(new_n13534_));
  AND2X1   g13342(.A(new_n13534_), .B(new_n12939_), .Y(new_n13535_));
  AOI22X1  g13343(.A0(new_n13009_), .A1(new_n13008_), .B0(new_n12965_), .B1(\asqrt[60] ), .Y(new_n13536_));
  AOI21X1  g13344(.A0(new_n13536_), .A1(\asqrt[19] ), .B0(new_n12954_), .Y(new_n13537_));
  AOI21X1  g13345(.A0(new_n13535_), .A1(\asqrt[19] ), .B0(new_n13537_), .Y(new_n13538_));
  OAI21X1  g13346(.A0(new_n13523_), .A1(new_n13510_), .B0(new_n13530_), .Y(new_n13539_));
  AOI21X1  g13347(.A0(new_n13539_), .A1(\asqrt[60] ), .B0(\asqrt[61] ), .Y(new_n13540_));
  AOI21X1  g13348(.A0(new_n13540_), .A1(new_n13532_), .B0(new_n13538_), .Y(new_n13541_));
  OAI21X1  g13349(.A0(new_n13541_), .A1(new_n13533_), .B0(\asqrt[62] ), .Y(new_n13542_));
  AND2X1   g13350(.A(new_n12966_), .B(new_n12958_), .Y(new_n13543_));
  NOR3X1   g13351(.A(new_n13543_), .B(new_n13012_), .C(new_n12959_), .Y(new_n13544_));
  NOR3X1   g13352(.A(new_n13000_), .B(new_n13543_), .C(new_n12959_), .Y(new_n13545_));
  NOR2X1   g13353(.A(new_n13545_), .B(new_n12964_), .Y(new_n13546_));
  AOI21X1  g13354(.A0(new_n13544_), .A1(\asqrt[19] ), .B0(new_n13546_), .Y(new_n13547_));
  NOR3X1   g13355(.A(new_n13541_), .B(new_n13533_), .C(\asqrt[62] ), .Y(new_n13548_));
  OAI21X1  g13356(.A0(new_n13548_), .A1(new_n13547_), .B0(new_n13542_), .Y(new_n13549_));
  NOR4X1   g13357(.A(new_n13000_), .B(new_n12973_), .C(new_n13016_), .D(new_n13015_), .Y(new_n13550_));
  NOR3X1   g13358(.A(new_n13000_), .B(new_n12973_), .C(new_n13015_), .Y(new_n13551_));
  NOR2X1   g13359(.A(new_n13551_), .B(new_n12972_), .Y(new_n13552_));
  NOR2X1   g13360(.A(new_n13552_), .B(new_n13550_), .Y(new_n13553_));
  INVX1    g13361(.A(new_n13553_), .Y(new_n13554_));
  AND2X1   g13362(.A(new_n12981_), .B(new_n12974_), .Y(new_n13555_));
  AOI21X1  g13363(.A0(new_n13555_), .A1(\asqrt[19] ), .B0(new_n13041_), .Y(new_n13556_));
  AND2X1   g13364(.A(new_n13556_), .B(new_n13554_), .Y(new_n13557_));
  AOI21X1  g13365(.A0(new_n13557_), .A1(new_n13549_), .B0(\asqrt[63] ), .Y(new_n13558_));
  NOR2X1   g13366(.A(new_n13548_), .B(new_n13547_), .Y(new_n13559_));
  NAND2X1  g13367(.A(new_n13553_), .B(new_n13542_), .Y(new_n13560_));
  AOI21X1  g13368(.A0(new_n13024_), .A1(new_n13020_), .B0(new_n12980_), .Y(new_n13561_));
  AOI21X1  g13369(.A0(new_n12981_), .A1(new_n12974_), .B0(new_n193_), .Y(new_n13562_));
  OAI21X1  g13370(.A0(new_n13561_), .A1(new_n12974_), .B0(new_n13562_), .Y(new_n13563_));
  INVX1    g13371(.A(new_n12979_), .Y(new_n13564_));
  NOR4X1   g13372(.A(new_n12997_), .B(new_n12991_), .C(new_n13564_), .D(new_n12976_), .Y(new_n13565_));
  OAI21X1  g13373(.A0(new_n12988_), .A1(new_n12987_), .B0(new_n13565_), .Y(new_n13566_));
  NOR2X1   g13374(.A(new_n13566_), .B(new_n12986_), .Y(new_n13567_));
  INVX1    g13375(.A(new_n13567_), .Y(new_n13568_));
  AND2X1   g13376(.A(new_n13568_), .B(new_n13563_), .Y(new_n13569_));
  OAI21X1  g13377(.A0(new_n13560_), .A1(new_n13559_), .B0(new_n13569_), .Y(new_n13570_));
  NOR2X1   g13378(.A(new_n13570_), .B(new_n13558_), .Y(new_n13571_));
  INVX1    g13379(.A(\a[36] ), .Y(new_n13572_));
  AND2X1   g13380(.A(new_n13539_), .B(\asqrt[60] ), .Y(new_n13573_));
  OR2X1    g13381(.A(new_n13523_), .B(new_n13510_), .Y(new_n13574_));
  AND2X1   g13382(.A(new_n13530_), .B(new_n292_), .Y(new_n13575_));
  AOI21X1  g13383(.A0(new_n13575_), .A1(new_n13574_), .B0(new_n13528_), .Y(new_n13576_));
  OAI21X1  g13384(.A0(new_n13576_), .A1(new_n13573_), .B0(\asqrt[61] ), .Y(new_n13577_));
  INVX1    g13385(.A(new_n13538_), .Y(new_n13578_));
  OAI21X1  g13386(.A0(new_n13513_), .A1(new_n292_), .B0(new_n217_), .Y(new_n13579_));
  OAI21X1  g13387(.A0(new_n13579_), .A1(new_n13576_), .B0(new_n13578_), .Y(new_n13580_));
  AOI21X1  g13388(.A0(new_n13580_), .A1(new_n13577_), .B0(new_n199_), .Y(new_n13581_));
  INVX1    g13389(.A(new_n13547_), .Y(new_n13582_));
  NAND3X1  g13390(.A(new_n13580_), .B(new_n13577_), .C(new_n199_), .Y(new_n13583_));
  AOI21X1  g13391(.A0(new_n13583_), .A1(new_n13582_), .B0(new_n13581_), .Y(new_n13584_));
  INVX1    g13392(.A(new_n13557_), .Y(new_n13585_));
  OAI21X1  g13393(.A0(new_n13585_), .A1(new_n13584_), .B0(new_n193_), .Y(new_n13586_));
  OR2X1    g13394(.A(new_n13548_), .B(new_n13547_), .Y(new_n13587_));
  AND2X1   g13395(.A(new_n13553_), .B(new_n13542_), .Y(new_n13588_));
  INVX1    g13396(.A(new_n13569_), .Y(new_n13589_));
  AOI21X1  g13397(.A0(new_n13588_), .A1(new_n13587_), .B0(new_n13589_), .Y(new_n13590_));
  AOI21X1  g13398(.A0(new_n13590_), .A1(new_n13586_), .B0(new_n13572_), .Y(new_n13591_));
  NOR3X1   g13399(.A(\a[36] ), .B(\a[35] ), .C(\a[34] ), .Y(new_n13592_));
  OAI21X1  g13400(.A0(new_n13592_), .A1(new_n13591_), .B0(\asqrt[19] ), .Y(new_n13593_));
  OAI21X1  g13401(.A0(new_n13570_), .A1(new_n13558_), .B0(\a[36] ), .Y(new_n13594_));
  OR2X1    g13402(.A(new_n13592_), .B(new_n12997_), .Y(new_n13595_));
  NOR4X1   g13403(.A(new_n13595_), .B(new_n12991_), .C(new_n13041_), .D(new_n12986_), .Y(new_n13596_));
  AND2X1   g13404(.A(new_n13596_), .B(new_n13594_), .Y(new_n13597_));
  INVX1    g13405(.A(\a[37] ), .Y(new_n13598_));
  AOI21X1  g13406(.A0(new_n13590_), .A1(new_n13586_), .B0(\a[36] ), .Y(new_n13599_));
  OAI21X1  g13407(.A0(new_n13570_), .A1(new_n13558_), .B0(new_n13004_), .Y(new_n13600_));
  OAI21X1  g13408(.A0(new_n13599_), .A1(new_n13598_), .B0(new_n13600_), .Y(new_n13601_));
  OAI21X1  g13409(.A0(new_n13601_), .A1(new_n13597_), .B0(new_n13593_), .Y(new_n13602_));
  AND2X1   g13410(.A(new_n13602_), .B(\asqrt[20] ), .Y(new_n13603_));
  NAND2X1  g13411(.A(new_n13596_), .B(new_n13594_), .Y(new_n13604_));
  OAI21X1  g13412(.A0(new_n13570_), .A1(new_n13558_), .B0(new_n13572_), .Y(new_n13605_));
  INVX1    g13413(.A(new_n13004_), .Y(new_n13606_));
  AOI21X1  g13414(.A0(new_n13590_), .A1(new_n13586_), .B0(new_n13606_), .Y(new_n13607_));
  AOI21X1  g13415(.A0(new_n13605_), .A1(\a[37] ), .B0(new_n13607_), .Y(new_n13608_));
  NAND2X1  g13416(.A(new_n13608_), .B(new_n13604_), .Y(new_n13609_));
  AND2X1   g13417(.A(new_n13593_), .B(new_n12447_), .Y(new_n13610_));
  INVX1    g13418(.A(new_n13563_), .Y(new_n13611_));
  NOR3X1   g13419(.A(new_n13567_), .B(new_n13611_), .C(new_n13000_), .Y(new_n13612_));
  OAI21X1  g13420(.A0(new_n13560_), .A1(new_n13559_), .B0(new_n13612_), .Y(new_n13613_));
  OR2X1    g13421(.A(new_n13613_), .B(new_n13558_), .Y(new_n13614_));
  AOI21X1  g13422(.A0(new_n13614_), .A1(new_n13600_), .B0(new_n13003_), .Y(new_n13615_));
  OAI21X1  g13423(.A0(new_n13613_), .A1(new_n13558_), .B0(new_n13003_), .Y(new_n13616_));
  NOR2X1   g13424(.A(new_n13616_), .B(new_n13607_), .Y(new_n13617_));
  NOR2X1   g13425(.A(new_n13617_), .B(new_n13615_), .Y(new_n13618_));
  AOI21X1  g13426(.A0(new_n13610_), .A1(new_n13609_), .B0(new_n13618_), .Y(new_n13619_));
  OAI21X1  g13427(.A0(new_n13619_), .A1(new_n13603_), .B0(\asqrt[21] ), .Y(new_n13620_));
  NOR3X1   g13428(.A(new_n13037_), .B(new_n13027_), .C(new_n13039_), .Y(new_n13621_));
  OAI21X1  g13429(.A0(new_n13570_), .A1(new_n13558_), .B0(new_n13621_), .Y(new_n13622_));
  NOR2X1   g13430(.A(new_n13027_), .B(new_n13039_), .Y(new_n13623_));
  OAI21X1  g13431(.A0(new_n13570_), .A1(new_n13558_), .B0(new_n13623_), .Y(new_n13624_));
  NAND2X1  g13432(.A(new_n13624_), .B(new_n13037_), .Y(new_n13625_));
  NAND2X1  g13433(.A(new_n13625_), .B(new_n13622_), .Y(new_n13626_));
  INVX1    g13434(.A(new_n13592_), .Y(new_n13627_));
  AOI21X1  g13435(.A0(new_n13627_), .A1(new_n13594_), .B0(new_n13000_), .Y(new_n13628_));
  AOI21X1  g13436(.A0(new_n13608_), .A1(new_n13604_), .B0(new_n13628_), .Y(new_n13629_));
  OAI21X1  g13437(.A0(new_n13629_), .A1(new_n12447_), .B0(new_n11896_), .Y(new_n13630_));
  OAI21X1  g13438(.A0(new_n13630_), .A1(new_n13619_), .B0(new_n13626_), .Y(new_n13631_));
  AOI21X1  g13439(.A0(new_n13631_), .A1(new_n13620_), .B0(new_n11362_), .Y(new_n13632_));
  AOI21X1  g13440(.A0(new_n13040_), .A1(new_n13038_), .B0(new_n13075_), .Y(new_n13633_));
  AND2X1   g13441(.A(new_n13633_), .B(new_n13072_), .Y(new_n13634_));
  OAI21X1  g13442(.A0(new_n13570_), .A1(new_n13558_), .B0(new_n13634_), .Y(new_n13635_));
  AOI22X1  g13443(.A0(new_n13040_), .A1(new_n13038_), .B0(new_n13032_), .B1(\asqrt[21] ), .Y(new_n13636_));
  OAI21X1  g13444(.A0(new_n13570_), .A1(new_n13558_), .B0(new_n13636_), .Y(new_n13637_));
  NAND2X1  g13445(.A(new_n13637_), .B(new_n13075_), .Y(new_n13638_));
  AND2X1   g13446(.A(new_n13638_), .B(new_n13635_), .Y(new_n13639_));
  INVX1    g13447(.A(new_n13639_), .Y(new_n13640_));
  NAND3X1  g13448(.A(new_n13631_), .B(new_n13620_), .C(new_n11362_), .Y(new_n13641_));
  AOI21X1  g13449(.A0(new_n13641_), .A1(new_n13640_), .B0(new_n13632_), .Y(new_n13642_));
  OR2X1    g13450(.A(new_n13642_), .B(new_n10849_), .Y(new_n13643_));
  OR2X1    g13451(.A(new_n13629_), .B(new_n12447_), .Y(new_n13644_));
  AND2X1   g13452(.A(new_n13608_), .B(new_n13604_), .Y(new_n13645_));
  OR2X1    g13453(.A(new_n13628_), .B(\asqrt[20] ), .Y(new_n13646_));
  OR2X1    g13454(.A(new_n13617_), .B(new_n13615_), .Y(new_n13647_));
  OAI21X1  g13455(.A0(new_n13646_), .A1(new_n13645_), .B0(new_n13647_), .Y(new_n13648_));
  AOI21X1  g13456(.A0(new_n13648_), .A1(new_n13644_), .B0(new_n11896_), .Y(new_n13649_));
  AND2X1   g13457(.A(new_n13625_), .B(new_n13622_), .Y(new_n13650_));
  AOI21X1  g13458(.A0(new_n13602_), .A1(\asqrt[20] ), .B0(\asqrt[21] ), .Y(new_n13651_));
  AOI21X1  g13459(.A0(new_n13651_), .A1(new_n13648_), .B0(new_n13650_), .Y(new_n13652_));
  NOR3X1   g13460(.A(new_n13652_), .B(new_n13649_), .C(\asqrt[22] ), .Y(new_n13653_));
  NOR2X1   g13461(.A(new_n13653_), .B(new_n13639_), .Y(new_n13654_));
  INVX1    g13462(.A(new_n13571_), .Y(\asqrt[18] ));
  AND2X1   g13463(.A(new_n13078_), .B(new_n13076_), .Y(new_n13656_));
  NOR3X1   g13464(.A(new_n13656_), .B(new_n13056_), .C(new_n13077_), .Y(new_n13657_));
  NOR2X1   g13465(.A(new_n13656_), .B(new_n13077_), .Y(new_n13658_));
  OAI21X1  g13466(.A0(new_n13570_), .A1(new_n13558_), .B0(new_n13658_), .Y(new_n13659_));
  AOI22X1  g13467(.A0(new_n13659_), .A1(new_n13056_), .B0(new_n13657_), .B1(\asqrt[18] ), .Y(new_n13660_));
  INVX1    g13468(.A(new_n13660_), .Y(new_n13661_));
  OAI21X1  g13469(.A0(new_n13652_), .A1(new_n13649_), .B0(\asqrt[22] ), .Y(new_n13662_));
  NAND2X1  g13470(.A(new_n13662_), .B(new_n10849_), .Y(new_n13663_));
  OAI21X1  g13471(.A0(new_n13663_), .A1(new_n13654_), .B0(new_n13661_), .Y(new_n13664_));
  AOI21X1  g13472(.A0(new_n13664_), .A1(new_n13643_), .B0(new_n10332_), .Y(new_n13665_));
  NAND4X1  g13473(.A(\asqrt[18] ), .B(new_n13069_), .C(new_n13067_), .D(new_n13094_), .Y(new_n13666_));
  NOR3X1   g13474(.A(new_n13571_), .B(new_n13080_), .C(new_n13060_), .Y(new_n13667_));
  OAI21X1  g13475(.A0(new_n13667_), .A1(new_n13067_), .B0(new_n13666_), .Y(new_n13668_));
  INVX1    g13476(.A(new_n13668_), .Y(new_n13669_));
  OAI21X1  g13477(.A0(new_n13653_), .A1(new_n13639_), .B0(new_n13662_), .Y(new_n13670_));
  AOI21X1  g13478(.A0(new_n13670_), .A1(\asqrt[23] ), .B0(\asqrt[24] ), .Y(new_n13671_));
  AOI21X1  g13479(.A0(new_n13671_), .A1(new_n13664_), .B0(new_n13669_), .Y(new_n13672_));
  OAI21X1  g13480(.A0(new_n13672_), .A1(new_n13665_), .B0(\asqrt[25] ), .Y(new_n13673_));
  AND2X1   g13481(.A(new_n13123_), .B(new_n13122_), .Y(new_n13674_));
  NOR3X1   g13482(.A(new_n13674_), .B(new_n13085_), .C(new_n13121_), .Y(new_n13675_));
  NOR3X1   g13483(.A(new_n13571_), .B(new_n13674_), .C(new_n13121_), .Y(new_n13676_));
  NOR2X1   g13484(.A(new_n13676_), .B(new_n13084_), .Y(new_n13677_));
  AOI21X1  g13485(.A0(new_n13675_), .A1(\asqrt[18] ), .B0(new_n13677_), .Y(new_n13678_));
  NOR3X1   g13486(.A(new_n13672_), .B(new_n13665_), .C(\asqrt[25] ), .Y(new_n13679_));
  OAI21X1  g13487(.A0(new_n13679_), .A1(new_n13678_), .B0(new_n13673_), .Y(new_n13680_));
  AND2X1   g13488(.A(new_n13680_), .B(\asqrt[26] ), .Y(new_n13681_));
  INVX1    g13489(.A(new_n13678_), .Y(new_n13682_));
  AND2X1   g13490(.A(new_n13670_), .B(\asqrt[23] ), .Y(new_n13683_));
  OR2X1    g13491(.A(new_n13653_), .B(new_n13639_), .Y(new_n13684_));
  AND2X1   g13492(.A(new_n13662_), .B(new_n10849_), .Y(new_n13685_));
  AOI21X1  g13493(.A0(new_n13685_), .A1(new_n13684_), .B0(new_n13660_), .Y(new_n13686_));
  OAI21X1  g13494(.A0(new_n13686_), .A1(new_n13683_), .B0(\asqrt[24] ), .Y(new_n13687_));
  OAI21X1  g13495(.A0(new_n13642_), .A1(new_n10849_), .B0(new_n10332_), .Y(new_n13688_));
  OAI21X1  g13496(.A0(new_n13688_), .A1(new_n13686_), .B0(new_n13668_), .Y(new_n13689_));
  NAND3X1  g13497(.A(new_n13689_), .B(new_n13687_), .C(new_n9833_), .Y(new_n13690_));
  NAND2X1  g13498(.A(new_n13690_), .B(new_n13682_), .Y(new_n13691_));
  AND2X1   g13499(.A(new_n13096_), .B(new_n13087_), .Y(new_n13692_));
  NOR3X1   g13500(.A(new_n13692_), .B(new_n13126_), .C(new_n13088_), .Y(new_n13693_));
  NOR3X1   g13501(.A(new_n13571_), .B(new_n13692_), .C(new_n13088_), .Y(new_n13694_));
  NOR2X1   g13502(.A(new_n13694_), .B(new_n13093_), .Y(new_n13695_));
  AOI21X1  g13503(.A0(new_n13693_), .A1(\asqrt[18] ), .B0(new_n13695_), .Y(new_n13696_));
  AND2X1   g13504(.A(new_n13673_), .B(new_n9353_), .Y(new_n13697_));
  AOI21X1  g13505(.A0(new_n13697_), .A1(new_n13691_), .B0(new_n13696_), .Y(new_n13698_));
  OAI21X1  g13506(.A0(new_n13698_), .A1(new_n13681_), .B0(\asqrt[27] ), .Y(new_n13699_));
  OR4X1    g13507(.A(new_n13571_), .B(new_n13104_), .C(new_n13130_), .D(new_n13129_), .Y(new_n13700_));
  OR2X1    g13508(.A(new_n13104_), .B(new_n13129_), .Y(new_n13701_));
  OAI21X1  g13509(.A0(new_n13701_), .A1(new_n13571_), .B0(new_n13130_), .Y(new_n13702_));
  AND2X1   g13510(.A(new_n13702_), .B(new_n13700_), .Y(new_n13703_));
  INVX1    g13511(.A(new_n13703_), .Y(new_n13704_));
  AOI21X1  g13512(.A0(new_n13689_), .A1(new_n13687_), .B0(new_n9833_), .Y(new_n13705_));
  AOI21X1  g13513(.A0(new_n13690_), .A1(new_n13682_), .B0(new_n13705_), .Y(new_n13706_));
  OAI21X1  g13514(.A0(new_n13706_), .A1(new_n9353_), .B0(new_n8874_), .Y(new_n13707_));
  OAI21X1  g13515(.A0(new_n13707_), .A1(new_n13698_), .B0(new_n13704_), .Y(new_n13708_));
  AOI21X1  g13516(.A0(new_n13708_), .A1(new_n13699_), .B0(new_n8412_), .Y(new_n13709_));
  AOI21X1  g13517(.A0(new_n13112_), .A1(new_n13107_), .B0(new_n13147_), .Y(new_n13710_));
  AND2X1   g13518(.A(new_n13710_), .B(new_n13145_), .Y(new_n13711_));
  AOI22X1  g13519(.A0(new_n13112_), .A1(new_n13107_), .B0(new_n13105_), .B1(\asqrt[27] ), .Y(new_n13712_));
  AOI21X1  g13520(.A0(new_n13712_), .A1(\asqrt[18] ), .B0(new_n13111_), .Y(new_n13713_));
  AOI21X1  g13521(.A0(new_n13711_), .A1(\asqrt[18] ), .B0(new_n13713_), .Y(new_n13714_));
  INVX1    g13522(.A(new_n13714_), .Y(new_n13715_));
  NAND3X1  g13523(.A(new_n13708_), .B(new_n13699_), .C(new_n8412_), .Y(new_n13716_));
  AOI21X1  g13524(.A0(new_n13716_), .A1(new_n13715_), .B0(new_n13709_), .Y(new_n13717_));
  OR2X1    g13525(.A(new_n13717_), .B(new_n7970_), .Y(new_n13718_));
  AND2X1   g13526(.A(new_n13716_), .B(new_n13715_), .Y(new_n13719_));
  AND2X1   g13527(.A(new_n13151_), .B(new_n13149_), .Y(new_n13720_));
  NOR3X1   g13528(.A(new_n13720_), .B(new_n13120_), .C(new_n13150_), .Y(new_n13721_));
  NOR3X1   g13529(.A(new_n13571_), .B(new_n13720_), .C(new_n13150_), .Y(new_n13722_));
  NOR2X1   g13530(.A(new_n13722_), .B(new_n13119_), .Y(new_n13723_));
  AOI21X1  g13531(.A0(new_n13721_), .A1(\asqrt[18] ), .B0(new_n13723_), .Y(new_n13724_));
  INVX1    g13532(.A(new_n13724_), .Y(new_n13725_));
  OR2X1    g13533(.A(new_n13706_), .B(new_n9353_), .Y(new_n13726_));
  AND2X1   g13534(.A(new_n13690_), .B(new_n13682_), .Y(new_n13727_));
  INVX1    g13535(.A(new_n13696_), .Y(new_n13728_));
  NAND2X1  g13536(.A(new_n13673_), .B(new_n9353_), .Y(new_n13729_));
  OAI21X1  g13537(.A0(new_n13729_), .A1(new_n13727_), .B0(new_n13728_), .Y(new_n13730_));
  AOI21X1  g13538(.A0(new_n13730_), .A1(new_n13726_), .B0(new_n8874_), .Y(new_n13731_));
  AOI21X1  g13539(.A0(new_n13680_), .A1(\asqrt[26] ), .B0(\asqrt[27] ), .Y(new_n13732_));
  AOI21X1  g13540(.A0(new_n13732_), .A1(new_n13730_), .B0(new_n13703_), .Y(new_n13733_));
  OAI21X1  g13541(.A0(new_n13733_), .A1(new_n13731_), .B0(\asqrt[28] ), .Y(new_n13734_));
  NAND2X1  g13542(.A(new_n13734_), .B(new_n7970_), .Y(new_n13735_));
  OAI21X1  g13543(.A0(new_n13735_), .A1(new_n13719_), .B0(new_n13725_), .Y(new_n13736_));
  AOI21X1  g13544(.A0(new_n13736_), .A1(new_n13718_), .B0(new_n7527_), .Y(new_n13737_));
  OR4X1    g13545(.A(new_n13571_), .B(new_n13153_), .C(new_n13141_), .D(new_n13135_), .Y(new_n13738_));
  OR2X1    g13546(.A(new_n13153_), .B(new_n13135_), .Y(new_n13739_));
  OAI21X1  g13547(.A0(new_n13739_), .A1(new_n13571_), .B0(new_n13141_), .Y(new_n13740_));
  AND2X1   g13548(.A(new_n13740_), .B(new_n13738_), .Y(new_n13741_));
  NOR3X1   g13549(.A(new_n13733_), .B(new_n13731_), .C(\asqrt[28] ), .Y(new_n13742_));
  OAI21X1  g13550(.A0(new_n13742_), .A1(new_n13714_), .B0(new_n13734_), .Y(new_n13743_));
  AOI21X1  g13551(.A0(new_n13743_), .A1(\asqrt[29] ), .B0(\asqrt[30] ), .Y(new_n13744_));
  AOI21X1  g13552(.A0(new_n13744_), .A1(new_n13736_), .B0(new_n13741_), .Y(new_n13745_));
  OAI21X1  g13553(.A0(new_n13745_), .A1(new_n13737_), .B0(\asqrt[31] ), .Y(new_n13746_));
  AND2X1   g13554(.A(new_n13184_), .B(new_n13183_), .Y(new_n13747_));
  NOR3X1   g13555(.A(new_n13747_), .B(new_n13159_), .C(new_n13182_), .Y(new_n13748_));
  NOR3X1   g13556(.A(new_n13571_), .B(new_n13747_), .C(new_n13182_), .Y(new_n13749_));
  NOR2X1   g13557(.A(new_n13749_), .B(new_n13158_), .Y(new_n13750_));
  AOI21X1  g13558(.A0(new_n13748_), .A1(\asqrt[18] ), .B0(new_n13750_), .Y(new_n13751_));
  NOR3X1   g13559(.A(new_n13745_), .B(new_n13737_), .C(\asqrt[31] ), .Y(new_n13752_));
  OAI21X1  g13560(.A0(new_n13752_), .A1(new_n13751_), .B0(new_n13746_), .Y(new_n13753_));
  AND2X1   g13561(.A(new_n13753_), .B(\asqrt[32] ), .Y(new_n13754_));
  INVX1    g13562(.A(new_n13751_), .Y(new_n13755_));
  AND2X1   g13563(.A(new_n13743_), .B(\asqrt[29] ), .Y(new_n13756_));
  NAND2X1  g13564(.A(new_n13716_), .B(new_n13715_), .Y(new_n13757_));
  AND2X1   g13565(.A(new_n13734_), .B(new_n7970_), .Y(new_n13758_));
  AOI21X1  g13566(.A0(new_n13758_), .A1(new_n13757_), .B0(new_n13724_), .Y(new_n13759_));
  OAI21X1  g13567(.A0(new_n13759_), .A1(new_n13756_), .B0(\asqrt[30] ), .Y(new_n13760_));
  INVX1    g13568(.A(new_n13741_), .Y(new_n13761_));
  OAI21X1  g13569(.A0(new_n13717_), .A1(new_n7970_), .B0(new_n7527_), .Y(new_n13762_));
  OAI21X1  g13570(.A0(new_n13762_), .A1(new_n13759_), .B0(new_n13761_), .Y(new_n13763_));
  NAND3X1  g13571(.A(new_n13763_), .B(new_n13760_), .C(new_n7103_), .Y(new_n13764_));
  NAND2X1  g13572(.A(new_n13764_), .B(new_n13755_), .Y(new_n13765_));
  AND2X1   g13573(.A(new_n13170_), .B(new_n13162_), .Y(new_n13766_));
  NOR3X1   g13574(.A(new_n13766_), .B(new_n13187_), .C(new_n13163_), .Y(new_n13767_));
  NOR3X1   g13575(.A(new_n13571_), .B(new_n13766_), .C(new_n13163_), .Y(new_n13768_));
  NOR2X1   g13576(.A(new_n13768_), .B(new_n13168_), .Y(new_n13769_));
  AOI21X1  g13577(.A0(new_n13767_), .A1(\asqrt[18] ), .B0(new_n13769_), .Y(new_n13770_));
  AND2X1   g13578(.A(new_n13746_), .B(new_n6699_), .Y(new_n13771_));
  AOI21X1  g13579(.A0(new_n13771_), .A1(new_n13765_), .B0(new_n13770_), .Y(new_n13772_));
  OAI21X1  g13580(.A0(new_n13772_), .A1(new_n13754_), .B0(\asqrt[33] ), .Y(new_n13773_));
  NAND4X1  g13581(.A(\asqrt[18] ), .B(new_n13190_), .C(new_n13177_), .D(new_n13172_), .Y(new_n13774_));
  NAND2X1  g13582(.A(new_n13190_), .B(new_n13172_), .Y(new_n13775_));
  OAI21X1  g13583(.A0(new_n13775_), .A1(new_n13571_), .B0(new_n13181_), .Y(new_n13776_));
  AND2X1   g13584(.A(new_n13776_), .B(new_n13774_), .Y(new_n13777_));
  INVX1    g13585(.A(new_n13777_), .Y(new_n13778_));
  AOI21X1  g13586(.A0(new_n13763_), .A1(new_n13760_), .B0(new_n7103_), .Y(new_n13779_));
  AOI21X1  g13587(.A0(new_n13764_), .A1(new_n13755_), .B0(new_n13779_), .Y(new_n13780_));
  OAI21X1  g13588(.A0(new_n13780_), .A1(new_n6699_), .B0(new_n6294_), .Y(new_n13781_));
  OAI21X1  g13589(.A0(new_n13781_), .A1(new_n13772_), .B0(new_n13778_), .Y(new_n13782_));
  AOI21X1  g13590(.A0(new_n13782_), .A1(new_n13773_), .B0(new_n5941_), .Y(new_n13783_));
  AOI21X1  g13591(.A0(new_n13197_), .A1(new_n13191_), .B0(new_n13221_), .Y(new_n13784_));
  AND2X1   g13592(.A(new_n13784_), .B(new_n13219_), .Y(new_n13785_));
  AOI22X1  g13593(.A0(new_n13197_), .A1(new_n13191_), .B0(new_n13179_), .B1(\asqrt[33] ), .Y(new_n13786_));
  AOI21X1  g13594(.A0(new_n13786_), .A1(\asqrt[18] ), .B0(new_n13195_), .Y(new_n13787_));
  AOI21X1  g13595(.A0(new_n13785_), .A1(\asqrt[18] ), .B0(new_n13787_), .Y(new_n13788_));
  INVX1    g13596(.A(new_n13788_), .Y(new_n13789_));
  NAND3X1  g13597(.A(new_n13782_), .B(new_n13773_), .C(new_n5941_), .Y(new_n13790_));
  AOI21X1  g13598(.A0(new_n13790_), .A1(new_n13789_), .B0(new_n13783_), .Y(new_n13791_));
  OR2X1    g13599(.A(new_n13791_), .B(new_n5541_), .Y(new_n13792_));
  AND2X1   g13600(.A(new_n13790_), .B(new_n13789_), .Y(new_n13793_));
  AND2X1   g13601(.A(new_n13225_), .B(new_n13223_), .Y(new_n13794_));
  NOR3X1   g13602(.A(new_n13794_), .B(new_n13205_), .C(new_n13224_), .Y(new_n13795_));
  NOR3X1   g13603(.A(new_n13571_), .B(new_n13794_), .C(new_n13224_), .Y(new_n13796_));
  NOR2X1   g13604(.A(new_n13796_), .B(new_n13204_), .Y(new_n13797_));
  AOI21X1  g13605(.A0(new_n13795_), .A1(\asqrt[18] ), .B0(new_n13797_), .Y(new_n13798_));
  INVX1    g13606(.A(new_n13798_), .Y(new_n13799_));
  OR2X1    g13607(.A(new_n13780_), .B(new_n6699_), .Y(new_n13800_));
  AND2X1   g13608(.A(new_n13764_), .B(new_n13755_), .Y(new_n13801_));
  INVX1    g13609(.A(new_n13770_), .Y(new_n13802_));
  NAND2X1  g13610(.A(new_n13746_), .B(new_n6699_), .Y(new_n13803_));
  OAI21X1  g13611(.A0(new_n13803_), .A1(new_n13801_), .B0(new_n13802_), .Y(new_n13804_));
  AOI21X1  g13612(.A0(new_n13804_), .A1(new_n13800_), .B0(new_n6294_), .Y(new_n13805_));
  AOI21X1  g13613(.A0(new_n13753_), .A1(\asqrt[32] ), .B0(\asqrt[33] ), .Y(new_n13806_));
  AOI21X1  g13614(.A0(new_n13806_), .A1(new_n13804_), .B0(new_n13777_), .Y(new_n13807_));
  OAI21X1  g13615(.A0(new_n13807_), .A1(new_n13805_), .B0(\asqrt[34] ), .Y(new_n13808_));
  NAND2X1  g13616(.A(new_n13808_), .B(new_n5541_), .Y(new_n13809_));
  OAI21X1  g13617(.A0(new_n13809_), .A1(new_n13793_), .B0(new_n13799_), .Y(new_n13810_));
  AOI21X1  g13618(.A0(new_n13810_), .A1(new_n13792_), .B0(new_n5176_), .Y(new_n13811_));
  NAND4X1  g13619(.A(\asqrt[18] ), .B(new_n13216_), .C(new_n13214_), .D(new_n13242_), .Y(new_n13812_));
  NAND2X1  g13620(.A(new_n13216_), .B(new_n13242_), .Y(new_n13813_));
  OAI21X1  g13621(.A0(new_n13813_), .A1(new_n13571_), .B0(new_n13215_), .Y(new_n13814_));
  AND2X1   g13622(.A(new_n13814_), .B(new_n13812_), .Y(new_n13815_));
  NOR3X1   g13623(.A(new_n13807_), .B(new_n13805_), .C(\asqrt[34] ), .Y(new_n13816_));
  OAI21X1  g13624(.A0(new_n13816_), .A1(new_n13788_), .B0(new_n13808_), .Y(new_n13817_));
  AOI21X1  g13625(.A0(new_n13817_), .A1(\asqrt[35] ), .B0(\asqrt[36] ), .Y(new_n13818_));
  AOI21X1  g13626(.A0(new_n13818_), .A1(new_n13810_), .B0(new_n13815_), .Y(new_n13819_));
  OAI21X1  g13627(.A0(new_n13819_), .A1(new_n13811_), .B0(\asqrt[37] ), .Y(new_n13820_));
  AND2X1   g13628(.A(new_n13258_), .B(new_n13257_), .Y(new_n13821_));
  NOR3X1   g13629(.A(new_n13821_), .B(new_n13233_), .C(new_n13256_), .Y(new_n13822_));
  NOR3X1   g13630(.A(new_n13571_), .B(new_n13821_), .C(new_n13256_), .Y(new_n13823_));
  NOR2X1   g13631(.A(new_n13823_), .B(new_n13232_), .Y(new_n13824_));
  AOI21X1  g13632(.A0(new_n13822_), .A1(\asqrt[18] ), .B0(new_n13824_), .Y(new_n13825_));
  NOR3X1   g13633(.A(new_n13819_), .B(new_n13811_), .C(\asqrt[37] ), .Y(new_n13826_));
  OAI21X1  g13634(.A0(new_n13826_), .A1(new_n13825_), .B0(new_n13820_), .Y(new_n13827_));
  AND2X1   g13635(.A(new_n13827_), .B(\asqrt[38] ), .Y(new_n13828_));
  INVX1    g13636(.A(new_n13825_), .Y(new_n13829_));
  AND2X1   g13637(.A(new_n13817_), .B(\asqrt[35] ), .Y(new_n13830_));
  NAND2X1  g13638(.A(new_n13790_), .B(new_n13789_), .Y(new_n13831_));
  AND2X1   g13639(.A(new_n13808_), .B(new_n5541_), .Y(new_n13832_));
  AOI21X1  g13640(.A0(new_n13832_), .A1(new_n13831_), .B0(new_n13798_), .Y(new_n13833_));
  OAI21X1  g13641(.A0(new_n13833_), .A1(new_n13830_), .B0(\asqrt[36] ), .Y(new_n13834_));
  INVX1    g13642(.A(new_n13815_), .Y(new_n13835_));
  OAI21X1  g13643(.A0(new_n13791_), .A1(new_n5541_), .B0(new_n5176_), .Y(new_n13836_));
  OAI21X1  g13644(.A0(new_n13836_), .A1(new_n13833_), .B0(new_n13835_), .Y(new_n13837_));
  NAND3X1  g13645(.A(new_n13837_), .B(new_n13834_), .C(new_n4826_), .Y(new_n13838_));
  NAND2X1  g13646(.A(new_n13838_), .B(new_n13829_), .Y(new_n13839_));
  AND2X1   g13647(.A(new_n13244_), .B(new_n13235_), .Y(new_n13840_));
  NOR3X1   g13648(.A(new_n13840_), .B(new_n13261_), .C(new_n13236_), .Y(new_n13841_));
  NOR3X1   g13649(.A(new_n13571_), .B(new_n13840_), .C(new_n13236_), .Y(new_n13842_));
  NOR2X1   g13650(.A(new_n13842_), .B(new_n13241_), .Y(new_n13843_));
  AOI21X1  g13651(.A0(new_n13841_), .A1(\asqrt[18] ), .B0(new_n13843_), .Y(new_n13844_));
  AND2X1   g13652(.A(new_n13820_), .B(new_n4493_), .Y(new_n13845_));
  AOI21X1  g13653(.A0(new_n13845_), .A1(new_n13839_), .B0(new_n13844_), .Y(new_n13846_));
  OAI21X1  g13654(.A0(new_n13846_), .A1(new_n13828_), .B0(\asqrt[39] ), .Y(new_n13847_));
  NAND4X1  g13655(.A(\asqrt[18] ), .B(new_n13264_), .C(new_n13251_), .D(new_n13246_), .Y(new_n13848_));
  NAND2X1  g13656(.A(new_n13264_), .B(new_n13246_), .Y(new_n13849_));
  OAI21X1  g13657(.A0(new_n13849_), .A1(new_n13571_), .B0(new_n13255_), .Y(new_n13850_));
  AND2X1   g13658(.A(new_n13850_), .B(new_n13848_), .Y(new_n13851_));
  INVX1    g13659(.A(new_n13851_), .Y(new_n13852_));
  AOI21X1  g13660(.A0(new_n13837_), .A1(new_n13834_), .B0(new_n4826_), .Y(new_n13853_));
  AOI21X1  g13661(.A0(new_n13838_), .A1(new_n13829_), .B0(new_n13853_), .Y(new_n13854_));
  OAI21X1  g13662(.A0(new_n13854_), .A1(new_n4493_), .B0(new_n4165_), .Y(new_n13855_));
  OAI21X1  g13663(.A0(new_n13855_), .A1(new_n13846_), .B0(new_n13852_), .Y(new_n13856_));
  AOI21X1  g13664(.A0(new_n13856_), .A1(new_n13847_), .B0(new_n3863_), .Y(new_n13857_));
  AOI21X1  g13665(.A0(new_n13271_), .A1(new_n13265_), .B0(new_n13295_), .Y(new_n13858_));
  AND2X1   g13666(.A(new_n13858_), .B(new_n13293_), .Y(new_n13859_));
  AOI22X1  g13667(.A0(new_n13271_), .A1(new_n13265_), .B0(new_n13253_), .B1(\asqrt[39] ), .Y(new_n13860_));
  AOI21X1  g13668(.A0(new_n13860_), .A1(\asqrt[18] ), .B0(new_n13269_), .Y(new_n13861_));
  AOI21X1  g13669(.A0(new_n13859_), .A1(\asqrt[18] ), .B0(new_n13861_), .Y(new_n13862_));
  INVX1    g13670(.A(new_n13862_), .Y(new_n13863_));
  NAND3X1  g13671(.A(new_n13856_), .B(new_n13847_), .C(new_n3863_), .Y(new_n13864_));
  AOI21X1  g13672(.A0(new_n13864_), .A1(new_n13863_), .B0(new_n13857_), .Y(new_n13865_));
  OR2X1    g13673(.A(new_n13865_), .B(new_n3564_), .Y(new_n13866_));
  AND2X1   g13674(.A(new_n13864_), .B(new_n13863_), .Y(new_n13867_));
  AND2X1   g13675(.A(new_n13299_), .B(new_n13297_), .Y(new_n13868_));
  NOR3X1   g13676(.A(new_n13868_), .B(new_n13279_), .C(new_n13298_), .Y(new_n13869_));
  NOR3X1   g13677(.A(new_n13571_), .B(new_n13868_), .C(new_n13298_), .Y(new_n13870_));
  NOR2X1   g13678(.A(new_n13870_), .B(new_n13278_), .Y(new_n13871_));
  AOI21X1  g13679(.A0(new_n13869_), .A1(\asqrt[18] ), .B0(new_n13871_), .Y(new_n13872_));
  INVX1    g13680(.A(new_n13872_), .Y(new_n13873_));
  OR2X1    g13681(.A(new_n13854_), .B(new_n4493_), .Y(new_n13874_));
  AND2X1   g13682(.A(new_n13838_), .B(new_n13829_), .Y(new_n13875_));
  INVX1    g13683(.A(new_n13844_), .Y(new_n13876_));
  NAND2X1  g13684(.A(new_n13820_), .B(new_n4493_), .Y(new_n13877_));
  OAI21X1  g13685(.A0(new_n13877_), .A1(new_n13875_), .B0(new_n13876_), .Y(new_n13878_));
  AOI21X1  g13686(.A0(new_n13878_), .A1(new_n13874_), .B0(new_n4165_), .Y(new_n13879_));
  AOI21X1  g13687(.A0(new_n13827_), .A1(\asqrt[38] ), .B0(\asqrt[39] ), .Y(new_n13880_));
  AOI21X1  g13688(.A0(new_n13880_), .A1(new_n13878_), .B0(new_n13851_), .Y(new_n13881_));
  OAI21X1  g13689(.A0(new_n13881_), .A1(new_n13879_), .B0(\asqrt[40] ), .Y(new_n13882_));
  NAND2X1  g13690(.A(new_n13882_), .B(new_n3564_), .Y(new_n13883_));
  OAI21X1  g13691(.A0(new_n13883_), .A1(new_n13867_), .B0(new_n13873_), .Y(new_n13884_));
  AOI21X1  g13692(.A0(new_n13884_), .A1(new_n13866_), .B0(new_n3276_), .Y(new_n13885_));
  OR4X1    g13693(.A(new_n13571_), .B(new_n13301_), .C(new_n13289_), .D(new_n13283_), .Y(new_n13886_));
  OR2X1    g13694(.A(new_n13301_), .B(new_n13283_), .Y(new_n13887_));
  OAI21X1  g13695(.A0(new_n13887_), .A1(new_n13571_), .B0(new_n13289_), .Y(new_n13888_));
  AND2X1   g13696(.A(new_n13888_), .B(new_n13886_), .Y(new_n13889_));
  NOR3X1   g13697(.A(new_n13881_), .B(new_n13879_), .C(\asqrt[40] ), .Y(new_n13890_));
  OAI21X1  g13698(.A0(new_n13890_), .A1(new_n13862_), .B0(new_n13882_), .Y(new_n13891_));
  AOI21X1  g13699(.A0(new_n13891_), .A1(\asqrt[41] ), .B0(\asqrt[42] ), .Y(new_n13892_));
  AOI21X1  g13700(.A0(new_n13892_), .A1(new_n13884_), .B0(new_n13889_), .Y(new_n13893_));
  OAI21X1  g13701(.A0(new_n13893_), .A1(new_n13885_), .B0(\asqrt[43] ), .Y(new_n13894_));
  AND2X1   g13702(.A(new_n13339_), .B(new_n13338_), .Y(new_n13895_));
  NOR3X1   g13703(.A(new_n13895_), .B(new_n13307_), .C(new_n13337_), .Y(new_n13896_));
  NOR3X1   g13704(.A(new_n13571_), .B(new_n13895_), .C(new_n13337_), .Y(new_n13897_));
  NOR2X1   g13705(.A(new_n13897_), .B(new_n13306_), .Y(new_n13898_));
  AOI21X1  g13706(.A0(new_n13896_), .A1(\asqrt[18] ), .B0(new_n13898_), .Y(new_n13899_));
  NOR3X1   g13707(.A(new_n13893_), .B(new_n13885_), .C(\asqrt[43] ), .Y(new_n13900_));
  OAI21X1  g13708(.A0(new_n13900_), .A1(new_n13899_), .B0(new_n13894_), .Y(new_n13901_));
  AND2X1   g13709(.A(new_n13901_), .B(\asqrt[44] ), .Y(new_n13902_));
  OR2X1    g13710(.A(new_n13900_), .B(new_n13899_), .Y(new_n13903_));
  AND2X1   g13711(.A(new_n13318_), .B(new_n13310_), .Y(new_n13904_));
  NOR3X1   g13712(.A(new_n13904_), .B(new_n13342_), .C(new_n13311_), .Y(new_n13905_));
  NOR3X1   g13713(.A(new_n13571_), .B(new_n13904_), .C(new_n13311_), .Y(new_n13906_));
  NOR2X1   g13714(.A(new_n13906_), .B(new_n13316_), .Y(new_n13907_));
  AOI21X1  g13715(.A0(new_n13905_), .A1(\asqrt[18] ), .B0(new_n13907_), .Y(new_n13908_));
  AND2X1   g13716(.A(new_n13894_), .B(new_n2769_), .Y(new_n13909_));
  AOI21X1  g13717(.A0(new_n13909_), .A1(new_n13903_), .B0(new_n13908_), .Y(new_n13910_));
  OAI21X1  g13718(.A0(new_n13910_), .A1(new_n13902_), .B0(\asqrt[45] ), .Y(new_n13911_));
  OR4X1    g13719(.A(new_n13571_), .B(new_n13326_), .C(new_n13346_), .D(new_n13345_), .Y(new_n13912_));
  OR2X1    g13720(.A(new_n13326_), .B(new_n13345_), .Y(new_n13913_));
  OAI21X1  g13721(.A0(new_n13913_), .A1(new_n13571_), .B0(new_n13346_), .Y(new_n13914_));
  AND2X1   g13722(.A(new_n13914_), .B(new_n13912_), .Y(new_n13915_));
  INVX1    g13723(.A(new_n13915_), .Y(new_n13916_));
  AND2X1   g13724(.A(new_n13891_), .B(\asqrt[41] ), .Y(new_n13917_));
  NAND2X1  g13725(.A(new_n13864_), .B(new_n13863_), .Y(new_n13918_));
  AND2X1   g13726(.A(new_n13882_), .B(new_n3564_), .Y(new_n13919_));
  AOI21X1  g13727(.A0(new_n13919_), .A1(new_n13918_), .B0(new_n13872_), .Y(new_n13920_));
  OAI21X1  g13728(.A0(new_n13920_), .A1(new_n13917_), .B0(\asqrt[42] ), .Y(new_n13921_));
  INVX1    g13729(.A(new_n13889_), .Y(new_n13922_));
  OAI21X1  g13730(.A0(new_n13865_), .A1(new_n3564_), .B0(new_n3276_), .Y(new_n13923_));
  OAI21X1  g13731(.A0(new_n13923_), .A1(new_n13920_), .B0(new_n13922_), .Y(new_n13924_));
  AOI21X1  g13732(.A0(new_n13924_), .A1(new_n13921_), .B0(new_n3008_), .Y(new_n13925_));
  INVX1    g13733(.A(new_n13899_), .Y(new_n13926_));
  NAND3X1  g13734(.A(new_n13924_), .B(new_n13921_), .C(new_n3008_), .Y(new_n13927_));
  AOI21X1  g13735(.A0(new_n13927_), .A1(new_n13926_), .B0(new_n13925_), .Y(new_n13928_));
  OAI21X1  g13736(.A0(new_n13928_), .A1(new_n2769_), .B0(new_n2570_), .Y(new_n13929_));
  OAI21X1  g13737(.A0(new_n13929_), .A1(new_n13910_), .B0(new_n13916_), .Y(new_n13930_));
  AOI21X1  g13738(.A0(new_n13930_), .A1(new_n13911_), .B0(new_n2263_), .Y(new_n13931_));
  AOI21X1  g13739(.A0(new_n13334_), .A1(new_n13329_), .B0(new_n13369_), .Y(new_n13932_));
  AND2X1   g13740(.A(new_n13932_), .B(new_n13367_), .Y(new_n13933_));
  AOI22X1  g13741(.A0(new_n13334_), .A1(new_n13329_), .B0(new_n13327_), .B1(\asqrt[45] ), .Y(new_n13934_));
  AOI21X1  g13742(.A0(new_n13934_), .A1(\asqrt[18] ), .B0(new_n13333_), .Y(new_n13935_));
  AOI21X1  g13743(.A0(new_n13933_), .A1(\asqrt[18] ), .B0(new_n13935_), .Y(new_n13936_));
  INVX1    g13744(.A(new_n13936_), .Y(new_n13937_));
  NAND3X1  g13745(.A(new_n13930_), .B(new_n13911_), .C(new_n2263_), .Y(new_n13938_));
  AOI21X1  g13746(.A0(new_n13938_), .A1(new_n13937_), .B0(new_n13931_), .Y(new_n13939_));
  OR2X1    g13747(.A(new_n13939_), .B(new_n2040_), .Y(new_n13940_));
  OR2X1    g13748(.A(new_n13928_), .B(new_n2769_), .Y(new_n13941_));
  AND2X1   g13749(.A(new_n13927_), .B(new_n13926_), .Y(new_n13942_));
  INVX1    g13750(.A(new_n13908_), .Y(new_n13943_));
  NAND2X1  g13751(.A(new_n13894_), .B(new_n2769_), .Y(new_n13944_));
  OAI21X1  g13752(.A0(new_n13944_), .A1(new_n13942_), .B0(new_n13943_), .Y(new_n13945_));
  AOI21X1  g13753(.A0(new_n13945_), .A1(new_n13941_), .B0(new_n2570_), .Y(new_n13946_));
  AOI21X1  g13754(.A0(new_n13901_), .A1(\asqrt[44] ), .B0(\asqrt[45] ), .Y(new_n13947_));
  AOI21X1  g13755(.A0(new_n13947_), .A1(new_n13945_), .B0(new_n13915_), .Y(new_n13948_));
  NOR3X1   g13756(.A(new_n13948_), .B(new_n13946_), .C(\asqrt[46] ), .Y(new_n13949_));
  NOR2X1   g13757(.A(new_n13949_), .B(new_n13936_), .Y(new_n13950_));
  OAI21X1  g13758(.A0(new_n13948_), .A1(new_n13946_), .B0(\asqrt[46] ), .Y(new_n13951_));
  NAND2X1  g13759(.A(new_n13951_), .B(new_n2040_), .Y(new_n13952_));
  AND2X1   g13760(.A(new_n13373_), .B(new_n13371_), .Y(new_n13953_));
  NOR3X1   g13761(.A(new_n13355_), .B(new_n13953_), .C(new_n13372_), .Y(new_n13954_));
  NOR3X1   g13762(.A(new_n13571_), .B(new_n13953_), .C(new_n13372_), .Y(new_n13955_));
  NOR2X1   g13763(.A(new_n13955_), .B(new_n13354_), .Y(new_n13956_));
  AOI21X1  g13764(.A0(new_n13954_), .A1(\asqrt[18] ), .B0(new_n13956_), .Y(new_n13957_));
  INVX1    g13765(.A(new_n13957_), .Y(new_n13958_));
  OAI21X1  g13766(.A0(new_n13952_), .A1(new_n13950_), .B0(new_n13958_), .Y(new_n13959_));
  AOI21X1  g13767(.A0(new_n13959_), .A1(new_n13940_), .B0(new_n1834_), .Y(new_n13960_));
  OR4X1    g13768(.A(new_n13571_), .B(new_n13375_), .C(new_n13363_), .D(new_n13357_), .Y(new_n13961_));
  OR2X1    g13769(.A(new_n13375_), .B(new_n13357_), .Y(new_n13962_));
  OAI21X1  g13770(.A0(new_n13962_), .A1(new_n13571_), .B0(new_n13363_), .Y(new_n13963_));
  AND2X1   g13771(.A(new_n13963_), .B(new_n13961_), .Y(new_n13964_));
  OAI21X1  g13772(.A0(new_n13949_), .A1(new_n13936_), .B0(new_n13951_), .Y(new_n13965_));
  AOI21X1  g13773(.A0(new_n13965_), .A1(\asqrt[47] ), .B0(\asqrt[48] ), .Y(new_n13966_));
  AOI21X1  g13774(.A0(new_n13966_), .A1(new_n13959_), .B0(new_n13964_), .Y(new_n13967_));
  OAI21X1  g13775(.A0(new_n13967_), .A1(new_n13960_), .B0(\asqrt[49] ), .Y(new_n13968_));
  AND2X1   g13776(.A(new_n13419_), .B(new_n13418_), .Y(new_n13969_));
  NOR3X1   g13777(.A(new_n13969_), .B(new_n13381_), .C(new_n13417_), .Y(new_n13970_));
  NOR3X1   g13778(.A(new_n13571_), .B(new_n13969_), .C(new_n13417_), .Y(new_n13971_));
  NOR2X1   g13779(.A(new_n13971_), .B(new_n13380_), .Y(new_n13972_));
  AOI21X1  g13780(.A0(new_n13970_), .A1(\asqrt[18] ), .B0(new_n13972_), .Y(new_n13973_));
  NOR3X1   g13781(.A(new_n13967_), .B(new_n13960_), .C(\asqrt[49] ), .Y(new_n13974_));
  OAI21X1  g13782(.A0(new_n13974_), .A1(new_n13973_), .B0(new_n13968_), .Y(new_n13975_));
  AND2X1   g13783(.A(new_n13975_), .B(\asqrt[50] ), .Y(new_n13976_));
  INVX1    g13784(.A(new_n13973_), .Y(new_n13977_));
  AND2X1   g13785(.A(new_n13965_), .B(\asqrt[47] ), .Y(new_n13978_));
  OR2X1    g13786(.A(new_n13949_), .B(new_n13936_), .Y(new_n13979_));
  AND2X1   g13787(.A(new_n13951_), .B(new_n2040_), .Y(new_n13980_));
  AOI21X1  g13788(.A0(new_n13980_), .A1(new_n13979_), .B0(new_n13957_), .Y(new_n13981_));
  OAI21X1  g13789(.A0(new_n13981_), .A1(new_n13978_), .B0(\asqrt[48] ), .Y(new_n13982_));
  INVX1    g13790(.A(new_n13964_), .Y(new_n13983_));
  OAI21X1  g13791(.A0(new_n13939_), .A1(new_n2040_), .B0(new_n1834_), .Y(new_n13984_));
  OAI21X1  g13792(.A0(new_n13984_), .A1(new_n13981_), .B0(new_n13983_), .Y(new_n13985_));
  NAND3X1  g13793(.A(new_n13985_), .B(new_n13982_), .C(new_n1632_), .Y(new_n13986_));
  NAND2X1  g13794(.A(new_n13986_), .B(new_n13977_), .Y(new_n13987_));
  AND2X1   g13795(.A(new_n13392_), .B(new_n13384_), .Y(new_n13988_));
  NOR3X1   g13796(.A(new_n13988_), .B(new_n13422_), .C(new_n13385_), .Y(new_n13989_));
  NOR3X1   g13797(.A(new_n13571_), .B(new_n13988_), .C(new_n13385_), .Y(new_n13990_));
  NOR2X1   g13798(.A(new_n13990_), .B(new_n13390_), .Y(new_n13991_));
  AOI21X1  g13799(.A0(new_n13989_), .A1(\asqrt[18] ), .B0(new_n13991_), .Y(new_n13992_));
  AND2X1   g13800(.A(new_n13968_), .B(new_n1469_), .Y(new_n13993_));
  AOI21X1  g13801(.A0(new_n13993_), .A1(new_n13987_), .B0(new_n13992_), .Y(new_n13994_));
  OAI21X1  g13802(.A0(new_n13994_), .A1(new_n13976_), .B0(\asqrt[51] ), .Y(new_n13995_));
  OR4X1    g13803(.A(new_n13571_), .B(new_n13400_), .C(new_n13426_), .D(new_n13425_), .Y(new_n13996_));
  OR2X1    g13804(.A(new_n13400_), .B(new_n13425_), .Y(new_n13997_));
  OAI21X1  g13805(.A0(new_n13997_), .A1(new_n13571_), .B0(new_n13426_), .Y(new_n13998_));
  AND2X1   g13806(.A(new_n13998_), .B(new_n13996_), .Y(new_n13999_));
  INVX1    g13807(.A(new_n13999_), .Y(new_n14000_));
  AOI21X1  g13808(.A0(new_n13985_), .A1(new_n13982_), .B0(new_n1632_), .Y(new_n14001_));
  AOI21X1  g13809(.A0(new_n13986_), .A1(new_n13977_), .B0(new_n14001_), .Y(new_n14002_));
  OAI21X1  g13810(.A0(new_n14002_), .A1(new_n1469_), .B0(new_n1277_), .Y(new_n14003_));
  OAI21X1  g13811(.A0(new_n14003_), .A1(new_n13994_), .B0(new_n14000_), .Y(new_n14004_));
  AOI21X1  g13812(.A0(new_n14004_), .A1(new_n13995_), .B0(new_n1111_), .Y(new_n14005_));
  AOI21X1  g13813(.A0(new_n13408_), .A1(new_n13403_), .B0(new_n13443_), .Y(new_n14006_));
  AND2X1   g13814(.A(new_n14006_), .B(new_n13441_), .Y(new_n14007_));
  AOI22X1  g13815(.A0(new_n13408_), .A1(new_n13403_), .B0(new_n13401_), .B1(\asqrt[51] ), .Y(new_n14008_));
  AOI21X1  g13816(.A0(new_n14008_), .A1(\asqrt[18] ), .B0(new_n13407_), .Y(new_n14009_));
  AOI21X1  g13817(.A0(new_n14007_), .A1(\asqrt[18] ), .B0(new_n14009_), .Y(new_n14010_));
  INVX1    g13818(.A(new_n14010_), .Y(new_n14011_));
  NAND3X1  g13819(.A(new_n14004_), .B(new_n13995_), .C(new_n1111_), .Y(new_n14012_));
  AOI21X1  g13820(.A0(new_n14012_), .A1(new_n14011_), .B0(new_n14005_), .Y(new_n14013_));
  OR2X1    g13821(.A(new_n14013_), .B(new_n968_), .Y(new_n14014_));
  OR2X1    g13822(.A(new_n14002_), .B(new_n1469_), .Y(new_n14015_));
  AND2X1   g13823(.A(new_n13986_), .B(new_n13977_), .Y(new_n14016_));
  INVX1    g13824(.A(new_n13992_), .Y(new_n14017_));
  NAND2X1  g13825(.A(new_n13968_), .B(new_n1469_), .Y(new_n14018_));
  OAI21X1  g13826(.A0(new_n14018_), .A1(new_n14016_), .B0(new_n14017_), .Y(new_n14019_));
  AOI21X1  g13827(.A0(new_n14019_), .A1(new_n14015_), .B0(new_n1277_), .Y(new_n14020_));
  AOI21X1  g13828(.A0(new_n13975_), .A1(\asqrt[50] ), .B0(\asqrt[51] ), .Y(new_n14021_));
  AOI21X1  g13829(.A0(new_n14021_), .A1(new_n14019_), .B0(new_n13999_), .Y(new_n14022_));
  NOR3X1   g13830(.A(new_n14022_), .B(new_n14020_), .C(\asqrt[52] ), .Y(new_n14023_));
  NOR2X1   g13831(.A(new_n14023_), .B(new_n14010_), .Y(new_n14024_));
  AND2X1   g13832(.A(new_n13447_), .B(new_n13445_), .Y(new_n14025_));
  NOR3X1   g13833(.A(new_n14025_), .B(new_n13416_), .C(new_n13446_), .Y(new_n14026_));
  NOR3X1   g13834(.A(new_n13571_), .B(new_n14025_), .C(new_n13446_), .Y(new_n14027_));
  NOR2X1   g13835(.A(new_n14027_), .B(new_n13415_), .Y(new_n14028_));
  AOI21X1  g13836(.A0(new_n14026_), .A1(\asqrt[18] ), .B0(new_n14028_), .Y(new_n14029_));
  INVX1    g13837(.A(new_n14029_), .Y(new_n14030_));
  OAI21X1  g13838(.A0(new_n14022_), .A1(new_n14020_), .B0(\asqrt[52] ), .Y(new_n14031_));
  NAND2X1  g13839(.A(new_n14031_), .B(new_n968_), .Y(new_n14032_));
  OAI21X1  g13840(.A0(new_n14032_), .A1(new_n14024_), .B0(new_n14030_), .Y(new_n14033_));
  AOI21X1  g13841(.A0(new_n14033_), .A1(new_n14014_), .B0(new_n902_), .Y(new_n14034_));
  OR4X1    g13842(.A(new_n13571_), .B(new_n13449_), .C(new_n13437_), .D(new_n13431_), .Y(new_n14035_));
  OR2X1    g13843(.A(new_n13449_), .B(new_n13431_), .Y(new_n14036_));
  OAI21X1  g13844(.A0(new_n14036_), .A1(new_n13571_), .B0(new_n13437_), .Y(new_n14037_));
  AND2X1   g13845(.A(new_n14037_), .B(new_n14035_), .Y(new_n14038_));
  OAI21X1  g13846(.A0(new_n14023_), .A1(new_n14010_), .B0(new_n14031_), .Y(new_n14039_));
  AOI21X1  g13847(.A0(new_n14039_), .A1(\asqrt[53] ), .B0(\asqrt[54] ), .Y(new_n14040_));
  AOI21X1  g13848(.A0(new_n14040_), .A1(new_n14033_), .B0(new_n14038_), .Y(new_n14041_));
  OAI21X1  g13849(.A0(new_n14041_), .A1(new_n14034_), .B0(\asqrt[55] ), .Y(new_n14042_));
  AND2X1   g13850(.A(new_n13493_), .B(new_n13492_), .Y(new_n14043_));
  NOR3X1   g13851(.A(new_n14043_), .B(new_n13455_), .C(new_n13491_), .Y(new_n14044_));
  NOR3X1   g13852(.A(new_n13571_), .B(new_n14043_), .C(new_n13491_), .Y(new_n14045_));
  NOR2X1   g13853(.A(new_n14045_), .B(new_n13454_), .Y(new_n14046_));
  AOI21X1  g13854(.A0(new_n14044_), .A1(\asqrt[18] ), .B0(new_n14046_), .Y(new_n14047_));
  NOR3X1   g13855(.A(new_n14041_), .B(new_n14034_), .C(\asqrt[55] ), .Y(new_n14048_));
  OAI21X1  g13856(.A0(new_n14048_), .A1(new_n14047_), .B0(new_n14042_), .Y(new_n14049_));
  AND2X1   g13857(.A(new_n14049_), .B(\asqrt[56] ), .Y(new_n14050_));
  OR2X1    g13858(.A(new_n14048_), .B(new_n14047_), .Y(new_n14051_));
  AND2X1   g13859(.A(new_n13466_), .B(new_n13458_), .Y(new_n14052_));
  NOR3X1   g13860(.A(new_n14052_), .B(new_n13496_), .C(new_n13459_), .Y(new_n14053_));
  NOR3X1   g13861(.A(new_n13571_), .B(new_n14052_), .C(new_n13459_), .Y(new_n14054_));
  NOR2X1   g13862(.A(new_n14054_), .B(new_n13464_), .Y(new_n14055_));
  AOI21X1  g13863(.A0(new_n14053_), .A1(\asqrt[18] ), .B0(new_n14055_), .Y(new_n14056_));
  AND2X1   g13864(.A(new_n14042_), .B(new_n582_), .Y(new_n14057_));
  AOI21X1  g13865(.A0(new_n14057_), .A1(new_n14051_), .B0(new_n14056_), .Y(new_n14058_));
  OAI21X1  g13866(.A0(new_n14058_), .A1(new_n14050_), .B0(\asqrt[57] ), .Y(new_n14059_));
  OR4X1    g13867(.A(new_n13571_), .B(new_n13474_), .C(new_n13500_), .D(new_n13499_), .Y(new_n14060_));
  OR2X1    g13868(.A(new_n13474_), .B(new_n13499_), .Y(new_n14061_));
  OAI21X1  g13869(.A0(new_n14061_), .A1(new_n13571_), .B0(new_n13500_), .Y(new_n14062_));
  AND2X1   g13870(.A(new_n14062_), .B(new_n14060_), .Y(new_n14063_));
  INVX1    g13871(.A(new_n14063_), .Y(new_n14064_));
  AND2X1   g13872(.A(new_n14039_), .B(\asqrt[53] ), .Y(new_n14065_));
  OR2X1    g13873(.A(new_n14023_), .B(new_n14010_), .Y(new_n14066_));
  AND2X1   g13874(.A(new_n14031_), .B(new_n968_), .Y(new_n14067_));
  AOI21X1  g13875(.A0(new_n14067_), .A1(new_n14066_), .B0(new_n14029_), .Y(new_n14068_));
  OAI21X1  g13876(.A0(new_n14068_), .A1(new_n14065_), .B0(\asqrt[54] ), .Y(new_n14069_));
  INVX1    g13877(.A(new_n14038_), .Y(new_n14070_));
  OAI21X1  g13878(.A0(new_n14013_), .A1(new_n968_), .B0(new_n902_), .Y(new_n14071_));
  OAI21X1  g13879(.A0(new_n14071_), .A1(new_n14068_), .B0(new_n14070_), .Y(new_n14072_));
  AOI21X1  g13880(.A0(new_n14072_), .A1(new_n14069_), .B0(new_n697_), .Y(new_n14073_));
  INVX1    g13881(.A(new_n14047_), .Y(new_n14074_));
  NAND3X1  g13882(.A(new_n14072_), .B(new_n14069_), .C(new_n697_), .Y(new_n14075_));
  AOI21X1  g13883(.A0(new_n14075_), .A1(new_n14074_), .B0(new_n14073_), .Y(new_n14076_));
  OAI21X1  g13884(.A0(new_n14076_), .A1(new_n582_), .B0(new_n481_), .Y(new_n14077_));
  OAI21X1  g13885(.A0(new_n14077_), .A1(new_n14058_), .B0(new_n14064_), .Y(new_n14078_));
  AOI21X1  g13886(.A0(new_n14078_), .A1(new_n14059_), .B0(new_n399_), .Y(new_n14079_));
  AOI21X1  g13887(.A0(new_n13482_), .A1(new_n13477_), .B0(new_n13517_), .Y(new_n14080_));
  AND2X1   g13888(.A(new_n14080_), .B(new_n13515_), .Y(new_n14081_));
  AOI22X1  g13889(.A0(new_n13482_), .A1(new_n13477_), .B0(new_n13475_), .B1(\asqrt[57] ), .Y(new_n14082_));
  AOI21X1  g13890(.A0(new_n14082_), .A1(\asqrt[18] ), .B0(new_n13481_), .Y(new_n14083_));
  AOI21X1  g13891(.A0(new_n14081_), .A1(\asqrt[18] ), .B0(new_n14083_), .Y(new_n14084_));
  INVX1    g13892(.A(new_n14084_), .Y(new_n14085_));
  NAND3X1  g13893(.A(new_n14078_), .B(new_n14059_), .C(new_n399_), .Y(new_n14086_));
  AOI21X1  g13894(.A0(new_n14086_), .A1(new_n14085_), .B0(new_n14079_), .Y(new_n14087_));
  OR2X1    g13895(.A(new_n14087_), .B(new_n328_), .Y(new_n14088_));
  AND2X1   g13896(.A(new_n14086_), .B(new_n14085_), .Y(new_n14089_));
  AND2X1   g13897(.A(new_n13521_), .B(new_n13519_), .Y(new_n14090_));
  NOR3X1   g13898(.A(new_n14090_), .B(new_n13490_), .C(new_n13520_), .Y(new_n14091_));
  NOR3X1   g13899(.A(new_n13571_), .B(new_n14090_), .C(new_n13520_), .Y(new_n14092_));
  NOR2X1   g13900(.A(new_n14092_), .B(new_n13489_), .Y(new_n14093_));
  AOI21X1  g13901(.A0(new_n14091_), .A1(\asqrt[18] ), .B0(new_n14093_), .Y(new_n14094_));
  INVX1    g13902(.A(new_n14094_), .Y(new_n14095_));
  OR2X1    g13903(.A(new_n14076_), .B(new_n582_), .Y(new_n14096_));
  NOR2X1   g13904(.A(new_n14048_), .B(new_n14047_), .Y(new_n14097_));
  INVX1    g13905(.A(new_n14056_), .Y(new_n14098_));
  NAND2X1  g13906(.A(new_n14042_), .B(new_n582_), .Y(new_n14099_));
  OAI21X1  g13907(.A0(new_n14099_), .A1(new_n14097_), .B0(new_n14098_), .Y(new_n14100_));
  AOI21X1  g13908(.A0(new_n14100_), .A1(new_n14096_), .B0(new_n481_), .Y(new_n14101_));
  AOI21X1  g13909(.A0(new_n14049_), .A1(\asqrt[56] ), .B0(\asqrt[57] ), .Y(new_n14102_));
  AOI21X1  g13910(.A0(new_n14102_), .A1(new_n14100_), .B0(new_n14063_), .Y(new_n14103_));
  OAI21X1  g13911(.A0(new_n14103_), .A1(new_n14101_), .B0(\asqrt[58] ), .Y(new_n14104_));
  NAND2X1  g13912(.A(new_n14104_), .B(new_n328_), .Y(new_n14105_));
  OAI21X1  g13913(.A0(new_n14105_), .A1(new_n14089_), .B0(new_n14095_), .Y(new_n14106_));
  AOI21X1  g13914(.A0(new_n14106_), .A1(new_n14088_), .B0(new_n292_), .Y(new_n14107_));
  OR4X1    g13915(.A(new_n13571_), .B(new_n13523_), .C(new_n13511_), .D(new_n13505_), .Y(new_n14108_));
  OR2X1    g13916(.A(new_n13523_), .B(new_n13505_), .Y(new_n14109_));
  OAI21X1  g13917(.A0(new_n14109_), .A1(new_n13571_), .B0(new_n13511_), .Y(new_n14110_));
  AND2X1   g13918(.A(new_n14110_), .B(new_n14108_), .Y(new_n14111_));
  NOR3X1   g13919(.A(new_n14103_), .B(new_n14101_), .C(\asqrt[58] ), .Y(new_n14112_));
  OAI21X1  g13920(.A0(new_n14112_), .A1(new_n14084_), .B0(new_n14104_), .Y(new_n14113_));
  AOI21X1  g13921(.A0(new_n14113_), .A1(\asqrt[59] ), .B0(\asqrt[60] ), .Y(new_n14114_));
  AOI21X1  g13922(.A0(new_n14114_), .A1(new_n14106_), .B0(new_n14111_), .Y(new_n14115_));
  OAI21X1  g13923(.A0(new_n14115_), .A1(new_n14107_), .B0(\asqrt[61] ), .Y(new_n14116_));
  AND2X1   g13924(.A(new_n13575_), .B(new_n13574_), .Y(new_n14117_));
  NOR3X1   g13925(.A(new_n14117_), .B(new_n13529_), .C(new_n13573_), .Y(new_n14118_));
  NOR3X1   g13926(.A(new_n13571_), .B(new_n14117_), .C(new_n13573_), .Y(new_n14119_));
  NOR2X1   g13927(.A(new_n14119_), .B(new_n13528_), .Y(new_n14120_));
  AOI21X1  g13928(.A0(new_n14118_), .A1(\asqrt[18] ), .B0(new_n14120_), .Y(new_n14121_));
  NOR3X1   g13929(.A(new_n14115_), .B(new_n14107_), .C(\asqrt[61] ), .Y(new_n14122_));
  OAI21X1  g13930(.A0(new_n14122_), .A1(new_n14121_), .B0(new_n14116_), .Y(new_n14123_));
  AND2X1   g13931(.A(new_n14123_), .B(\asqrt[62] ), .Y(new_n14124_));
  OR2X1    g13932(.A(new_n14122_), .B(new_n14121_), .Y(new_n14125_));
  AND2X1   g13933(.A(new_n13540_), .B(new_n13532_), .Y(new_n14126_));
  NOR3X1   g13934(.A(new_n14126_), .B(new_n13578_), .C(new_n13533_), .Y(new_n14127_));
  NOR3X1   g13935(.A(new_n13571_), .B(new_n14126_), .C(new_n13533_), .Y(new_n14128_));
  NOR2X1   g13936(.A(new_n14128_), .B(new_n13538_), .Y(new_n14129_));
  AOI21X1  g13937(.A0(new_n14127_), .A1(\asqrt[18] ), .B0(new_n14129_), .Y(new_n14130_));
  AND2X1   g13938(.A(new_n14116_), .B(new_n199_), .Y(new_n14131_));
  AOI21X1  g13939(.A0(new_n14131_), .A1(new_n14125_), .B0(new_n14130_), .Y(new_n14132_));
  NOR4X1   g13940(.A(new_n13571_), .B(new_n13548_), .C(new_n13582_), .D(new_n13581_), .Y(new_n14133_));
  NAND3X1  g13941(.A(\asqrt[18] ), .B(new_n13583_), .C(new_n13542_), .Y(new_n14134_));
  AOI21X1  g13942(.A0(new_n14134_), .A1(new_n13582_), .B0(new_n14133_), .Y(new_n14135_));
  INVX1    g13943(.A(new_n14135_), .Y(new_n14136_));
  OR2X1    g13944(.A(new_n13560_), .B(new_n13559_), .Y(new_n14137_));
  INVX1    g13945(.A(new_n14137_), .Y(new_n14138_));
  AND2X1   g13946(.A(new_n13554_), .B(new_n13549_), .Y(new_n14139_));
  AOI21X1  g13947(.A0(new_n14139_), .A1(\asqrt[18] ), .B0(new_n14138_), .Y(new_n14140_));
  AND2X1   g13948(.A(new_n14140_), .B(new_n14136_), .Y(new_n14141_));
  OAI21X1  g13949(.A0(new_n14132_), .A1(new_n14124_), .B0(new_n14141_), .Y(new_n14142_));
  AND2X1   g13950(.A(new_n14113_), .B(\asqrt[59] ), .Y(new_n14143_));
  NAND2X1  g13951(.A(new_n14086_), .B(new_n14085_), .Y(new_n14144_));
  AND2X1   g13952(.A(new_n14104_), .B(new_n328_), .Y(new_n14145_));
  AOI21X1  g13953(.A0(new_n14145_), .A1(new_n14144_), .B0(new_n14094_), .Y(new_n14146_));
  OAI21X1  g13954(.A0(new_n14146_), .A1(new_n14143_), .B0(\asqrt[60] ), .Y(new_n14147_));
  INVX1    g13955(.A(new_n14111_), .Y(new_n14148_));
  OAI21X1  g13956(.A0(new_n14087_), .A1(new_n328_), .B0(new_n292_), .Y(new_n14149_));
  OAI21X1  g13957(.A0(new_n14149_), .A1(new_n14146_), .B0(new_n14148_), .Y(new_n14150_));
  AOI21X1  g13958(.A0(new_n14150_), .A1(new_n14147_), .B0(new_n217_), .Y(new_n14151_));
  INVX1    g13959(.A(new_n14121_), .Y(new_n14152_));
  NAND3X1  g13960(.A(new_n14150_), .B(new_n14147_), .C(new_n217_), .Y(new_n14153_));
  AOI21X1  g13961(.A0(new_n14153_), .A1(new_n14152_), .B0(new_n14151_), .Y(new_n14154_));
  OAI21X1  g13962(.A0(new_n14154_), .A1(new_n199_), .B0(new_n14135_), .Y(new_n14155_));
  AOI21X1  g13963(.A0(new_n13590_), .A1(new_n13586_), .B0(new_n13553_), .Y(new_n14156_));
  AOI21X1  g13964(.A0(new_n13554_), .A1(new_n13549_), .B0(new_n193_), .Y(new_n14157_));
  OAI21X1  g13965(.A0(new_n14156_), .A1(new_n13549_), .B0(new_n14157_), .Y(new_n14158_));
  OR2X1    g13966(.A(new_n13567_), .B(new_n13550_), .Y(new_n14159_));
  OR2X1    g13967(.A(new_n14159_), .B(new_n13552_), .Y(new_n14160_));
  NOR4X1   g13968(.A(new_n14160_), .B(new_n13611_), .C(new_n14138_), .D(new_n13558_), .Y(new_n14161_));
  INVX1    g13969(.A(new_n14161_), .Y(new_n14162_));
  AND2X1   g13970(.A(new_n14162_), .B(new_n14158_), .Y(new_n14163_));
  OAI21X1  g13971(.A0(new_n14155_), .A1(new_n14132_), .B0(new_n14163_), .Y(new_n14164_));
  AOI21X1  g13972(.A0(new_n14142_), .A1(new_n193_), .B0(new_n14164_), .Y(new_n14165_));
  NOR2X1   g13973(.A(\a[33] ), .B(\a[32] ), .Y(new_n14166_));
  INVX1    g13974(.A(new_n14166_), .Y(new_n14167_));
  MX2X1    g13975(.A(new_n14167_), .B(new_n14165_), .S0(\a[34] ), .Y(new_n14168_));
  OR2X1    g13976(.A(new_n14168_), .B(new_n13571_), .Y(new_n14169_));
  INVX1    g13977(.A(\a[34] ), .Y(new_n14170_));
  NOR3X1   g13978(.A(\a[34] ), .B(\a[33] ), .C(\a[32] ), .Y(new_n14171_));
  NOR3X1   g13979(.A(new_n14171_), .B(new_n13567_), .C(new_n13611_), .Y(new_n14172_));
  NAND3X1  g13980(.A(new_n14172_), .B(new_n14137_), .C(new_n13586_), .Y(new_n14173_));
  INVX1    g13981(.A(new_n14173_), .Y(new_n14174_));
  OAI21X1  g13982(.A0(new_n14165_), .A1(new_n14170_), .B0(new_n14174_), .Y(new_n14175_));
  OAI21X1  g13983(.A0(new_n14165_), .A1(\a[34] ), .B0(\a[35] ), .Y(new_n14176_));
  NOR2X1   g13984(.A(\a[35] ), .B(\a[34] ), .Y(new_n14177_));
  INVX1    g13985(.A(new_n14177_), .Y(new_n14178_));
  OR2X1    g13986(.A(new_n14165_), .B(new_n14178_), .Y(new_n14179_));
  NAND3X1  g13987(.A(new_n14179_), .B(new_n14176_), .C(new_n14175_), .Y(new_n14180_));
  AOI21X1  g13988(.A0(new_n14180_), .A1(new_n14169_), .B0(new_n13000_), .Y(new_n14181_));
  OR2X1    g13989(.A(new_n14154_), .B(new_n199_), .Y(new_n14182_));
  NOR2X1   g13990(.A(new_n14122_), .B(new_n14121_), .Y(new_n14183_));
  INVX1    g13991(.A(new_n14130_), .Y(new_n14184_));
  NAND2X1  g13992(.A(new_n14116_), .B(new_n199_), .Y(new_n14185_));
  OAI21X1  g13993(.A0(new_n14185_), .A1(new_n14183_), .B0(new_n14184_), .Y(new_n14186_));
  INVX1    g13994(.A(new_n14141_), .Y(new_n14187_));
  AOI21X1  g13995(.A0(new_n14186_), .A1(new_n14182_), .B0(new_n14187_), .Y(new_n14188_));
  AOI21X1  g13996(.A0(new_n14123_), .A1(\asqrt[62] ), .B0(new_n14136_), .Y(new_n14189_));
  INVX1    g13997(.A(new_n14163_), .Y(new_n14190_));
  AOI21X1  g13998(.A0(new_n14189_), .A1(new_n14186_), .B0(new_n14190_), .Y(new_n14191_));
  OAI21X1  g13999(.A0(new_n14188_), .A1(\asqrt[63] ), .B0(new_n14191_), .Y(\asqrt[17] ));
  MX2X1    g14000(.A(new_n14166_), .B(\asqrt[17] ), .S0(\a[34] ), .Y(new_n14193_));
  AOI21X1  g14001(.A0(new_n14193_), .A1(\asqrt[18] ), .B0(\asqrt[19] ), .Y(new_n14194_));
  NAND3X1  g14002(.A(new_n14162_), .B(new_n14158_), .C(\asqrt[18] ), .Y(new_n14195_));
  INVX1    g14003(.A(new_n14195_), .Y(new_n14196_));
  OAI21X1  g14004(.A0(new_n14155_), .A1(new_n14132_), .B0(new_n14196_), .Y(new_n14197_));
  AOI21X1  g14005(.A0(new_n14142_), .A1(new_n193_), .B0(new_n14197_), .Y(new_n14198_));
  AOI21X1  g14006(.A0(\asqrt[17] ), .A1(new_n14177_), .B0(new_n14198_), .Y(new_n14199_));
  OR2X1    g14007(.A(new_n14199_), .B(new_n13572_), .Y(new_n14200_));
  AND2X1   g14008(.A(\asqrt[17] ), .B(new_n14177_), .Y(new_n14201_));
  OR2X1    g14009(.A(new_n14198_), .B(\a[36] ), .Y(new_n14202_));
  OR2X1    g14010(.A(new_n14202_), .B(new_n14201_), .Y(new_n14203_));
  AOI22X1  g14011(.A0(new_n14203_), .A1(new_n14200_), .B0(new_n14194_), .B1(new_n14180_), .Y(new_n14204_));
  OAI21X1  g14012(.A0(new_n14204_), .A1(new_n14181_), .B0(\asqrt[20] ), .Y(new_n14205_));
  AND2X1   g14013(.A(new_n13604_), .B(new_n13593_), .Y(new_n14206_));
  NAND3X1  g14014(.A(new_n14206_), .B(\asqrt[17] ), .C(new_n13601_), .Y(new_n14207_));
  INVX1    g14015(.A(new_n14206_), .Y(new_n14208_));
  OAI21X1  g14016(.A0(new_n14208_), .A1(new_n14165_), .B0(new_n13608_), .Y(new_n14209_));
  AND2X1   g14017(.A(new_n14209_), .B(new_n14207_), .Y(new_n14210_));
  NOR3X1   g14018(.A(new_n14204_), .B(new_n14181_), .C(\asqrt[20] ), .Y(new_n14211_));
  OAI21X1  g14019(.A0(new_n14211_), .A1(new_n14210_), .B0(new_n14205_), .Y(new_n14212_));
  AND2X1   g14020(.A(new_n14212_), .B(\asqrt[21] ), .Y(new_n14213_));
  INVX1    g14021(.A(new_n14210_), .Y(new_n14214_));
  AND2X1   g14022(.A(new_n14193_), .B(\asqrt[18] ), .Y(new_n14215_));
  AOI21X1  g14023(.A0(\asqrt[17] ), .A1(\a[34] ), .B0(new_n14173_), .Y(new_n14216_));
  INVX1    g14024(.A(\a[35] ), .Y(new_n14217_));
  AOI21X1  g14025(.A0(\asqrt[17] ), .A1(new_n14170_), .B0(new_n14217_), .Y(new_n14218_));
  NOR3X1   g14026(.A(new_n14201_), .B(new_n14218_), .C(new_n14216_), .Y(new_n14219_));
  OAI21X1  g14027(.A0(new_n14219_), .A1(new_n14215_), .B0(\asqrt[19] ), .Y(new_n14220_));
  OAI21X1  g14028(.A0(new_n14168_), .A1(new_n13571_), .B0(new_n13000_), .Y(new_n14221_));
  OAI22X1  g14029(.A0(new_n14202_), .A1(new_n14201_), .B0(new_n14199_), .B1(new_n13572_), .Y(new_n14222_));
  OAI21X1  g14030(.A0(new_n14221_), .A1(new_n14219_), .B0(new_n14222_), .Y(new_n14223_));
  NAND3X1  g14031(.A(new_n14223_), .B(new_n14220_), .C(new_n12447_), .Y(new_n14224_));
  NAND2X1  g14032(.A(new_n14224_), .B(new_n14214_), .Y(new_n14225_));
  AOI21X1  g14033(.A0(new_n13610_), .A1(new_n13609_), .B0(new_n13647_), .Y(new_n14226_));
  NAND3X1  g14034(.A(new_n14226_), .B(\asqrt[17] ), .C(new_n13644_), .Y(new_n14227_));
  OAI22X1  g14035(.A0(new_n13646_), .A1(new_n13645_), .B0(new_n13629_), .B1(new_n12447_), .Y(new_n14228_));
  OAI21X1  g14036(.A0(new_n14228_), .A1(new_n14165_), .B0(new_n13647_), .Y(new_n14229_));
  AND2X1   g14037(.A(new_n14229_), .B(new_n14227_), .Y(new_n14230_));
  AOI21X1  g14038(.A0(new_n14223_), .A1(new_n14220_), .B0(new_n12447_), .Y(new_n14231_));
  NOR2X1   g14039(.A(new_n14231_), .B(\asqrt[21] ), .Y(new_n14232_));
  AOI21X1  g14040(.A0(new_n14232_), .A1(new_n14225_), .B0(new_n14230_), .Y(new_n14233_));
  OAI21X1  g14041(.A0(new_n14233_), .A1(new_n14213_), .B0(\asqrt[22] ), .Y(new_n14234_));
  OR2X1    g14042(.A(new_n13630_), .B(new_n13619_), .Y(new_n14235_));
  NAND4X1  g14043(.A(\asqrt[17] ), .B(new_n14235_), .C(new_n13650_), .D(new_n13620_), .Y(new_n14236_));
  NAND2X1  g14044(.A(new_n14235_), .B(new_n13620_), .Y(new_n14237_));
  OAI21X1  g14045(.A0(new_n14237_), .A1(new_n14165_), .B0(new_n13626_), .Y(new_n14238_));
  AND2X1   g14046(.A(new_n14238_), .B(new_n14236_), .Y(new_n14239_));
  INVX1    g14047(.A(new_n14239_), .Y(new_n14240_));
  AOI21X1  g14048(.A0(new_n14224_), .A1(new_n14214_), .B0(new_n14231_), .Y(new_n14241_));
  OAI21X1  g14049(.A0(new_n14241_), .A1(new_n11896_), .B0(new_n11362_), .Y(new_n14242_));
  OAI21X1  g14050(.A0(new_n14242_), .A1(new_n14233_), .B0(new_n14240_), .Y(new_n14243_));
  AOI21X1  g14051(.A0(new_n14243_), .A1(new_n14234_), .B0(new_n10849_), .Y(new_n14244_));
  OR4X1    g14052(.A(new_n14165_), .B(new_n13653_), .C(new_n13640_), .D(new_n13632_), .Y(new_n14245_));
  NAND2X1  g14053(.A(new_n13641_), .B(new_n13662_), .Y(new_n14246_));
  OAI21X1  g14054(.A0(new_n14246_), .A1(new_n14165_), .B0(new_n13640_), .Y(new_n14247_));
  AND2X1   g14055(.A(new_n14247_), .B(new_n14245_), .Y(new_n14248_));
  INVX1    g14056(.A(new_n14248_), .Y(new_n14249_));
  NAND3X1  g14057(.A(new_n14243_), .B(new_n14234_), .C(new_n10849_), .Y(new_n14250_));
  AOI21X1  g14058(.A0(new_n14250_), .A1(new_n14249_), .B0(new_n14244_), .Y(new_n14251_));
  OR2X1    g14059(.A(new_n14251_), .B(new_n10332_), .Y(new_n14252_));
  AND2X1   g14060(.A(new_n14250_), .B(new_n14249_), .Y(new_n14253_));
  AND2X1   g14061(.A(new_n13685_), .B(new_n13684_), .Y(new_n14254_));
  NOR4X1   g14062(.A(new_n14165_), .B(new_n14254_), .C(new_n13661_), .D(new_n13683_), .Y(new_n14255_));
  AOI22X1  g14063(.A0(new_n13685_), .A1(new_n13684_), .B0(new_n13670_), .B1(\asqrt[23] ), .Y(new_n14256_));
  AOI21X1  g14064(.A0(new_n14256_), .A1(\asqrt[17] ), .B0(new_n13660_), .Y(new_n14257_));
  NOR2X1   g14065(.A(new_n14257_), .B(new_n14255_), .Y(new_n14258_));
  INVX1    g14066(.A(new_n14258_), .Y(new_n14259_));
  OR2X1    g14067(.A(new_n14244_), .B(\asqrt[24] ), .Y(new_n14260_));
  OAI21X1  g14068(.A0(new_n14260_), .A1(new_n14253_), .B0(new_n14259_), .Y(new_n14261_));
  AOI21X1  g14069(.A0(new_n14261_), .A1(new_n14252_), .B0(new_n9833_), .Y(new_n14262_));
  AND2X1   g14070(.A(new_n13671_), .B(new_n13664_), .Y(new_n14263_));
  OR4X1    g14071(.A(new_n14165_), .B(new_n14263_), .C(new_n13668_), .D(new_n13665_), .Y(new_n14264_));
  OR2X1    g14072(.A(new_n14263_), .B(new_n13665_), .Y(new_n14265_));
  OAI21X1  g14073(.A0(new_n14265_), .A1(new_n14165_), .B0(new_n13668_), .Y(new_n14266_));
  AND2X1   g14074(.A(new_n14266_), .B(new_n14264_), .Y(new_n14267_));
  OR2X1    g14075(.A(new_n14241_), .B(new_n11896_), .Y(new_n14268_));
  AND2X1   g14076(.A(new_n14224_), .B(new_n14214_), .Y(new_n14269_));
  INVX1    g14077(.A(new_n14230_), .Y(new_n14270_));
  OR2X1    g14078(.A(new_n14231_), .B(\asqrt[21] ), .Y(new_n14271_));
  OAI21X1  g14079(.A0(new_n14271_), .A1(new_n14269_), .B0(new_n14270_), .Y(new_n14272_));
  AOI21X1  g14080(.A0(new_n14272_), .A1(new_n14268_), .B0(new_n11362_), .Y(new_n14273_));
  AOI21X1  g14081(.A0(new_n14212_), .A1(\asqrt[21] ), .B0(\asqrt[22] ), .Y(new_n14274_));
  AOI21X1  g14082(.A0(new_n14274_), .A1(new_n14272_), .B0(new_n14239_), .Y(new_n14275_));
  OAI21X1  g14083(.A0(new_n14275_), .A1(new_n14273_), .B0(\asqrt[23] ), .Y(new_n14276_));
  NOR3X1   g14084(.A(new_n14275_), .B(new_n14273_), .C(\asqrt[23] ), .Y(new_n14277_));
  OAI21X1  g14085(.A0(new_n14277_), .A1(new_n14248_), .B0(new_n14276_), .Y(new_n14278_));
  AOI21X1  g14086(.A0(new_n14278_), .A1(\asqrt[24] ), .B0(\asqrt[25] ), .Y(new_n14279_));
  AOI21X1  g14087(.A0(new_n14279_), .A1(new_n14261_), .B0(new_n14267_), .Y(new_n14280_));
  OAI21X1  g14088(.A0(new_n14280_), .A1(new_n14262_), .B0(\asqrt[26] ), .Y(new_n14281_));
  OR4X1    g14089(.A(new_n14165_), .B(new_n13679_), .C(new_n13682_), .D(new_n13705_), .Y(new_n14282_));
  NAND2X1  g14090(.A(new_n13690_), .B(new_n13673_), .Y(new_n14283_));
  OAI21X1  g14091(.A0(new_n14283_), .A1(new_n14165_), .B0(new_n13682_), .Y(new_n14284_));
  AND2X1   g14092(.A(new_n14284_), .B(new_n14282_), .Y(new_n14285_));
  NOR3X1   g14093(.A(new_n14280_), .B(new_n14262_), .C(\asqrt[26] ), .Y(new_n14286_));
  OAI21X1  g14094(.A0(new_n14286_), .A1(new_n14285_), .B0(new_n14281_), .Y(new_n14287_));
  AND2X1   g14095(.A(new_n14287_), .B(\asqrt[27] ), .Y(new_n14288_));
  INVX1    g14096(.A(new_n14285_), .Y(new_n14289_));
  AND2X1   g14097(.A(new_n14278_), .B(\asqrt[24] ), .Y(new_n14290_));
  NAND2X1  g14098(.A(new_n14250_), .B(new_n14249_), .Y(new_n14291_));
  NOR2X1   g14099(.A(new_n14244_), .B(\asqrt[24] ), .Y(new_n14292_));
  AOI21X1  g14100(.A0(new_n14292_), .A1(new_n14291_), .B0(new_n14258_), .Y(new_n14293_));
  OAI21X1  g14101(.A0(new_n14293_), .A1(new_n14290_), .B0(\asqrt[25] ), .Y(new_n14294_));
  INVX1    g14102(.A(new_n14267_), .Y(new_n14295_));
  OAI21X1  g14103(.A0(new_n14251_), .A1(new_n10332_), .B0(new_n9833_), .Y(new_n14296_));
  OAI21X1  g14104(.A0(new_n14296_), .A1(new_n14293_), .B0(new_n14295_), .Y(new_n14297_));
  NAND3X1  g14105(.A(new_n14297_), .B(new_n14294_), .C(new_n9353_), .Y(new_n14298_));
  NAND2X1  g14106(.A(new_n14298_), .B(new_n14289_), .Y(new_n14299_));
  OAI21X1  g14107(.A0(new_n13729_), .A1(new_n13727_), .B0(new_n13696_), .Y(new_n14300_));
  NOR3X1   g14108(.A(new_n14300_), .B(new_n14165_), .C(new_n13681_), .Y(new_n14301_));
  AOI22X1  g14109(.A0(new_n13697_), .A1(new_n13691_), .B0(new_n13680_), .B1(\asqrt[26] ), .Y(new_n14302_));
  AOI21X1  g14110(.A0(new_n14302_), .A1(\asqrt[17] ), .B0(new_n13696_), .Y(new_n14303_));
  NOR2X1   g14111(.A(new_n14303_), .B(new_n14301_), .Y(new_n14304_));
  AOI21X1  g14112(.A0(new_n14297_), .A1(new_n14294_), .B0(new_n9353_), .Y(new_n14305_));
  NOR2X1   g14113(.A(new_n14305_), .B(\asqrt[27] ), .Y(new_n14306_));
  AOI21X1  g14114(.A0(new_n14306_), .A1(new_n14299_), .B0(new_n14304_), .Y(new_n14307_));
  OAI21X1  g14115(.A0(new_n14307_), .A1(new_n14288_), .B0(\asqrt[28] ), .Y(new_n14308_));
  AND2X1   g14116(.A(new_n13732_), .B(new_n13730_), .Y(new_n14309_));
  OR4X1    g14117(.A(new_n14165_), .B(new_n14309_), .C(new_n13704_), .D(new_n13731_), .Y(new_n14310_));
  OR2X1    g14118(.A(new_n14309_), .B(new_n13731_), .Y(new_n14311_));
  OAI21X1  g14119(.A0(new_n14311_), .A1(new_n14165_), .B0(new_n13704_), .Y(new_n14312_));
  AND2X1   g14120(.A(new_n14312_), .B(new_n14310_), .Y(new_n14313_));
  INVX1    g14121(.A(new_n14313_), .Y(new_n14314_));
  AOI21X1  g14122(.A0(new_n14298_), .A1(new_n14289_), .B0(new_n14305_), .Y(new_n14315_));
  OAI21X1  g14123(.A0(new_n14315_), .A1(new_n8874_), .B0(new_n8412_), .Y(new_n14316_));
  OAI21X1  g14124(.A0(new_n14316_), .A1(new_n14307_), .B0(new_n14314_), .Y(new_n14317_));
  AOI21X1  g14125(.A0(new_n14317_), .A1(new_n14308_), .B0(new_n7970_), .Y(new_n14318_));
  OR4X1    g14126(.A(new_n14165_), .B(new_n13742_), .C(new_n13715_), .D(new_n13709_), .Y(new_n14319_));
  NAND2X1  g14127(.A(new_n13716_), .B(new_n13734_), .Y(new_n14320_));
  OAI21X1  g14128(.A0(new_n14320_), .A1(new_n14165_), .B0(new_n13715_), .Y(new_n14321_));
  AND2X1   g14129(.A(new_n14321_), .B(new_n14319_), .Y(new_n14322_));
  INVX1    g14130(.A(new_n14322_), .Y(new_n14323_));
  NAND3X1  g14131(.A(new_n14317_), .B(new_n14308_), .C(new_n7970_), .Y(new_n14324_));
  AOI21X1  g14132(.A0(new_n14324_), .A1(new_n14323_), .B0(new_n14318_), .Y(new_n14325_));
  OR2X1    g14133(.A(new_n14325_), .B(new_n7527_), .Y(new_n14326_));
  AND2X1   g14134(.A(new_n14324_), .B(new_n14323_), .Y(new_n14327_));
  AND2X1   g14135(.A(new_n13758_), .B(new_n13757_), .Y(new_n14328_));
  NOR4X1   g14136(.A(new_n14165_), .B(new_n14328_), .C(new_n13725_), .D(new_n13756_), .Y(new_n14329_));
  AOI22X1  g14137(.A0(new_n13758_), .A1(new_n13757_), .B0(new_n13743_), .B1(\asqrt[29] ), .Y(new_n14330_));
  AOI21X1  g14138(.A0(new_n14330_), .A1(\asqrt[17] ), .B0(new_n13724_), .Y(new_n14331_));
  NOR2X1   g14139(.A(new_n14331_), .B(new_n14329_), .Y(new_n14332_));
  INVX1    g14140(.A(new_n14332_), .Y(new_n14333_));
  OR2X1    g14141(.A(new_n14318_), .B(\asqrt[30] ), .Y(new_n14334_));
  OAI21X1  g14142(.A0(new_n14334_), .A1(new_n14327_), .B0(new_n14333_), .Y(new_n14335_));
  AOI21X1  g14143(.A0(new_n14335_), .A1(new_n14326_), .B0(new_n7103_), .Y(new_n14336_));
  OAI21X1  g14144(.A0(new_n13762_), .A1(new_n13759_), .B0(new_n13741_), .Y(new_n14337_));
  OR2X1    g14145(.A(new_n14337_), .B(new_n13737_), .Y(new_n14338_));
  AND2X1   g14146(.A(new_n13744_), .B(new_n13736_), .Y(new_n14339_));
  NOR3X1   g14147(.A(new_n14165_), .B(new_n14339_), .C(new_n13737_), .Y(new_n14340_));
  OAI22X1  g14148(.A0(new_n14340_), .A1(new_n13741_), .B0(new_n14338_), .B1(new_n14165_), .Y(new_n14341_));
  INVX1    g14149(.A(new_n14341_), .Y(new_n14342_));
  OR2X1    g14150(.A(new_n14315_), .B(new_n8874_), .Y(new_n14343_));
  AND2X1   g14151(.A(new_n14298_), .B(new_n14289_), .Y(new_n14344_));
  INVX1    g14152(.A(new_n14304_), .Y(new_n14345_));
  OR2X1    g14153(.A(new_n14305_), .B(\asqrt[27] ), .Y(new_n14346_));
  OAI21X1  g14154(.A0(new_n14346_), .A1(new_n14344_), .B0(new_n14345_), .Y(new_n14347_));
  AOI21X1  g14155(.A0(new_n14347_), .A1(new_n14343_), .B0(new_n8412_), .Y(new_n14348_));
  AOI21X1  g14156(.A0(new_n14287_), .A1(\asqrt[27] ), .B0(\asqrt[28] ), .Y(new_n14349_));
  AOI21X1  g14157(.A0(new_n14349_), .A1(new_n14347_), .B0(new_n14313_), .Y(new_n14350_));
  OAI21X1  g14158(.A0(new_n14350_), .A1(new_n14348_), .B0(\asqrt[29] ), .Y(new_n14351_));
  NOR3X1   g14159(.A(new_n14350_), .B(new_n14348_), .C(\asqrt[29] ), .Y(new_n14352_));
  OAI21X1  g14160(.A0(new_n14352_), .A1(new_n14322_), .B0(new_n14351_), .Y(new_n14353_));
  AOI21X1  g14161(.A0(new_n14353_), .A1(\asqrt[30] ), .B0(\asqrt[31] ), .Y(new_n14354_));
  AOI21X1  g14162(.A0(new_n14354_), .A1(new_n14335_), .B0(new_n14342_), .Y(new_n14355_));
  OAI21X1  g14163(.A0(new_n14355_), .A1(new_n14336_), .B0(\asqrt[32] ), .Y(new_n14356_));
  OR4X1    g14164(.A(new_n14165_), .B(new_n13752_), .C(new_n13755_), .D(new_n13779_), .Y(new_n14357_));
  NAND2X1  g14165(.A(new_n13764_), .B(new_n13746_), .Y(new_n14358_));
  OAI21X1  g14166(.A0(new_n14358_), .A1(new_n14165_), .B0(new_n13755_), .Y(new_n14359_));
  AND2X1   g14167(.A(new_n14359_), .B(new_n14357_), .Y(new_n14360_));
  NOR3X1   g14168(.A(new_n14355_), .B(new_n14336_), .C(\asqrt[32] ), .Y(new_n14361_));
  OAI21X1  g14169(.A0(new_n14361_), .A1(new_n14360_), .B0(new_n14356_), .Y(new_n14362_));
  AND2X1   g14170(.A(new_n14362_), .B(\asqrt[33] ), .Y(new_n14363_));
  INVX1    g14171(.A(new_n14360_), .Y(new_n14364_));
  AND2X1   g14172(.A(new_n14353_), .B(\asqrt[30] ), .Y(new_n14365_));
  NAND2X1  g14173(.A(new_n14324_), .B(new_n14323_), .Y(new_n14366_));
  NOR2X1   g14174(.A(new_n14318_), .B(\asqrt[30] ), .Y(new_n14367_));
  AOI21X1  g14175(.A0(new_n14367_), .A1(new_n14366_), .B0(new_n14332_), .Y(new_n14368_));
  OAI21X1  g14176(.A0(new_n14368_), .A1(new_n14365_), .B0(\asqrt[31] ), .Y(new_n14369_));
  OAI21X1  g14177(.A0(new_n14325_), .A1(new_n7527_), .B0(new_n7103_), .Y(new_n14370_));
  OAI21X1  g14178(.A0(new_n14370_), .A1(new_n14368_), .B0(new_n14341_), .Y(new_n14371_));
  NAND3X1  g14179(.A(new_n14371_), .B(new_n14369_), .C(new_n6699_), .Y(new_n14372_));
  NAND2X1  g14180(.A(new_n14372_), .B(new_n14364_), .Y(new_n14373_));
  OAI21X1  g14181(.A0(new_n13803_), .A1(new_n13801_), .B0(new_n13770_), .Y(new_n14374_));
  NOR3X1   g14182(.A(new_n14374_), .B(new_n14165_), .C(new_n13754_), .Y(new_n14375_));
  AOI22X1  g14183(.A0(new_n13771_), .A1(new_n13765_), .B0(new_n13753_), .B1(\asqrt[32] ), .Y(new_n14376_));
  AOI21X1  g14184(.A0(new_n14376_), .A1(\asqrt[17] ), .B0(new_n13770_), .Y(new_n14377_));
  NOR2X1   g14185(.A(new_n14377_), .B(new_n14375_), .Y(new_n14378_));
  AOI21X1  g14186(.A0(new_n14371_), .A1(new_n14369_), .B0(new_n6699_), .Y(new_n14379_));
  NOR2X1   g14187(.A(new_n14379_), .B(\asqrt[33] ), .Y(new_n14380_));
  AOI21X1  g14188(.A0(new_n14380_), .A1(new_n14373_), .B0(new_n14378_), .Y(new_n14381_));
  OAI21X1  g14189(.A0(new_n14381_), .A1(new_n14363_), .B0(\asqrt[34] ), .Y(new_n14382_));
  AND2X1   g14190(.A(new_n13806_), .B(new_n13804_), .Y(new_n14383_));
  OR4X1    g14191(.A(new_n14165_), .B(new_n14383_), .C(new_n13778_), .D(new_n13805_), .Y(new_n14384_));
  OR2X1    g14192(.A(new_n14383_), .B(new_n13805_), .Y(new_n14385_));
  OAI21X1  g14193(.A0(new_n14385_), .A1(new_n14165_), .B0(new_n13778_), .Y(new_n14386_));
  AND2X1   g14194(.A(new_n14386_), .B(new_n14384_), .Y(new_n14387_));
  INVX1    g14195(.A(new_n14387_), .Y(new_n14388_));
  AOI21X1  g14196(.A0(new_n14372_), .A1(new_n14364_), .B0(new_n14379_), .Y(new_n14389_));
  OAI21X1  g14197(.A0(new_n14389_), .A1(new_n6294_), .B0(new_n5941_), .Y(new_n14390_));
  OAI21X1  g14198(.A0(new_n14390_), .A1(new_n14381_), .B0(new_n14388_), .Y(new_n14391_));
  AOI21X1  g14199(.A0(new_n14391_), .A1(new_n14382_), .B0(new_n5541_), .Y(new_n14392_));
  NAND3X1  g14200(.A(new_n13790_), .B(new_n13788_), .C(new_n13808_), .Y(new_n14393_));
  NOR3X1   g14201(.A(new_n14165_), .B(new_n13816_), .C(new_n13783_), .Y(new_n14394_));
  OAI22X1  g14202(.A0(new_n14394_), .A1(new_n13788_), .B0(new_n14393_), .B1(new_n14165_), .Y(new_n14395_));
  NAND3X1  g14203(.A(new_n14391_), .B(new_n14382_), .C(new_n5541_), .Y(new_n14396_));
  AOI21X1  g14204(.A0(new_n14396_), .A1(new_n14395_), .B0(new_n14392_), .Y(new_n14397_));
  OR2X1    g14205(.A(new_n14397_), .B(new_n5176_), .Y(new_n14398_));
  AND2X1   g14206(.A(new_n14396_), .B(new_n14395_), .Y(new_n14399_));
  AND2X1   g14207(.A(new_n13832_), .B(new_n13831_), .Y(new_n14400_));
  NOR4X1   g14208(.A(new_n14165_), .B(new_n14400_), .C(new_n13799_), .D(new_n13830_), .Y(new_n14401_));
  AOI22X1  g14209(.A0(new_n13832_), .A1(new_n13831_), .B0(new_n13817_), .B1(\asqrt[35] ), .Y(new_n14402_));
  AOI21X1  g14210(.A0(new_n14402_), .A1(\asqrt[17] ), .B0(new_n13798_), .Y(new_n14403_));
  NOR2X1   g14211(.A(new_n14403_), .B(new_n14401_), .Y(new_n14404_));
  INVX1    g14212(.A(new_n14404_), .Y(new_n14405_));
  OR2X1    g14213(.A(new_n14392_), .B(\asqrt[36] ), .Y(new_n14406_));
  OAI21X1  g14214(.A0(new_n14406_), .A1(new_n14399_), .B0(new_n14405_), .Y(new_n14407_));
  AOI21X1  g14215(.A0(new_n14407_), .A1(new_n14398_), .B0(new_n4826_), .Y(new_n14408_));
  AND2X1   g14216(.A(new_n13818_), .B(new_n13810_), .Y(new_n14409_));
  NOR4X1   g14217(.A(new_n14165_), .B(new_n14409_), .C(new_n13835_), .D(new_n13811_), .Y(new_n14410_));
  NOR2X1   g14218(.A(new_n14409_), .B(new_n13811_), .Y(new_n14411_));
  AOI21X1  g14219(.A0(new_n14411_), .A1(\asqrt[17] ), .B0(new_n13815_), .Y(new_n14412_));
  NOR2X1   g14220(.A(new_n14412_), .B(new_n14410_), .Y(new_n14413_));
  OR2X1    g14221(.A(new_n14389_), .B(new_n6294_), .Y(new_n14414_));
  AND2X1   g14222(.A(new_n14372_), .B(new_n14364_), .Y(new_n14415_));
  INVX1    g14223(.A(new_n14378_), .Y(new_n14416_));
  OR2X1    g14224(.A(new_n14379_), .B(\asqrt[33] ), .Y(new_n14417_));
  OAI21X1  g14225(.A0(new_n14417_), .A1(new_n14415_), .B0(new_n14416_), .Y(new_n14418_));
  AOI21X1  g14226(.A0(new_n14418_), .A1(new_n14414_), .B0(new_n5941_), .Y(new_n14419_));
  AOI21X1  g14227(.A0(new_n14362_), .A1(\asqrt[33] ), .B0(\asqrt[34] ), .Y(new_n14420_));
  AOI21X1  g14228(.A0(new_n14420_), .A1(new_n14418_), .B0(new_n14387_), .Y(new_n14421_));
  OAI21X1  g14229(.A0(new_n14421_), .A1(new_n14419_), .B0(\asqrt[35] ), .Y(new_n14422_));
  INVX1    g14230(.A(new_n14395_), .Y(new_n14423_));
  NOR3X1   g14231(.A(new_n14421_), .B(new_n14419_), .C(\asqrt[35] ), .Y(new_n14424_));
  OAI21X1  g14232(.A0(new_n14424_), .A1(new_n14423_), .B0(new_n14422_), .Y(new_n14425_));
  AOI21X1  g14233(.A0(new_n14425_), .A1(\asqrt[36] ), .B0(\asqrt[37] ), .Y(new_n14426_));
  AOI21X1  g14234(.A0(new_n14426_), .A1(new_n14407_), .B0(new_n14413_), .Y(new_n14427_));
  OAI21X1  g14235(.A0(new_n14427_), .A1(new_n14408_), .B0(\asqrt[38] ), .Y(new_n14428_));
  OR4X1    g14236(.A(new_n14165_), .B(new_n13826_), .C(new_n13829_), .D(new_n13853_), .Y(new_n14429_));
  NAND2X1  g14237(.A(new_n13838_), .B(new_n13820_), .Y(new_n14430_));
  OAI21X1  g14238(.A0(new_n14430_), .A1(new_n14165_), .B0(new_n13829_), .Y(new_n14431_));
  AND2X1   g14239(.A(new_n14431_), .B(new_n14429_), .Y(new_n14432_));
  NOR3X1   g14240(.A(new_n14427_), .B(new_n14408_), .C(\asqrt[38] ), .Y(new_n14433_));
  OAI21X1  g14241(.A0(new_n14433_), .A1(new_n14432_), .B0(new_n14428_), .Y(new_n14434_));
  AND2X1   g14242(.A(new_n14434_), .B(\asqrt[39] ), .Y(new_n14435_));
  OR2X1    g14243(.A(new_n14433_), .B(new_n14432_), .Y(new_n14436_));
  OAI21X1  g14244(.A0(new_n13877_), .A1(new_n13875_), .B0(new_n13844_), .Y(new_n14437_));
  NOR3X1   g14245(.A(new_n14437_), .B(new_n14165_), .C(new_n13828_), .Y(new_n14438_));
  AOI22X1  g14246(.A0(new_n13845_), .A1(new_n13839_), .B0(new_n13827_), .B1(\asqrt[38] ), .Y(new_n14439_));
  AOI21X1  g14247(.A0(new_n14439_), .A1(\asqrt[17] ), .B0(new_n13844_), .Y(new_n14440_));
  NOR2X1   g14248(.A(new_n14440_), .B(new_n14438_), .Y(new_n14441_));
  AND2X1   g14249(.A(new_n14428_), .B(new_n4165_), .Y(new_n14442_));
  AOI21X1  g14250(.A0(new_n14442_), .A1(new_n14436_), .B0(new_n14441_), .Y(new_n14443_));
  OAI21X1  g14251(.A0(new_n14443_), .A1(new_n14435_), .B0(\asqrt[40] ), .Y(new_n14444_));
  AND2X1   g14252(.A(new_n13880_), .B(new_n13878_), .Y(new_n14445_));
  OR2X1    g14253(.A(new_n13852_), .B(new_n13879_), .Y(new_n14446_));
  OR2X1    g14254(.A(new_n14446_), .B(new_n14445_), .Y(new_n14447_));
  NOR3X1   g14255(.A(new_n14165_), .B(new_n14445_), .C(new_n13879_), .Y(new_n14448_));
  OAI22X1  g14256(.A0(new_n14448_), .A1(new_n13851_), .B0(new_n14447_), .B1(new_n14165_), .Y(new_n14449_));
  AND2X1   g14257(.A(new_n14425_), .B(\asqrt[36] ), .Y(new_n14450_));
  NAND2X1  g14258(.A(new_n14396_), .B(new_n14395_), .Y(new_n14451_));
  NOR2X1   g14259(.A(new_n14392_), .B(\asqrt[36] ), .Y(new_n14452_));
  AOI21X1  g14260(.A0(new_n14452_), .A1(new_n14451_), .B0(new_n14404_), .Y(new_n14453_));
  OAI21X1  g14261(.A0(new_n14453_), .A1(new_n14450_), .B0(\asqrt[37] ), .Y(new_n14454_));
  INVX1    g14262(.A(new_n14413_), .Y(new_n14455_));
  OAI21X1  g14263(.A0(new_n14397_), .A1(new_n5176_), .B0(new_n4826_), .Y(new_n14456_));
  OAI21X1  g14264(.A0(new_n14456_), .A1(new_n14453_), .B0(new_n14455_), .Y(new_n14457_));
  AOI21X1  g14265(.A0(new_n14457_), .A1(new_n14454_), .B0(new_n4493_), .Y(new_n14458_));
  INVX1    g14266(.A(new_n14432_), .Y(new_n14459_));
  NAND3X1  g14267(.A(new_n14457_), .B(new_n14454_), .C(new_n4493_), .Y(new_n14460_));
  AOI21X1  g14268(.A0(new_n14460_), .A1(new_n14459_), .B0(new_n14458_), .Y(new_n14461_));
  OAI21X1  g14269(.A0(new_n14461_), .A1(new_n4165_), .B0(new_n3863_), .Y(new_n14462_));
  OAI21X1  g14270(.A0(new_n14462_), .A1(new_n14443_), .B0(new_n14449_), .Y(new_n14463_));
  AOI21X1  g14271(.A0(new_n14463_), .A1(new_n14444_), .B0(new_n3564_), .Y(new_n14464_));
  OR4X1    g14272(.A(new_n14165_), .B(new_n13890_), .C(new_n13863_), .D(new_n13857_), .Y(new_n14465_));
  NAND2X1  g14273(.A(new_n13864_), .B(new_n13882_), .Y(new_n14466_));
  OAI21X1  g14274(.A0(new_n14466_), .A1(new_n14165_), .B0(new_n13863_), .Y(new_n14467_));
  AND2X1   g14275(.A(new_n14467_), .B(new_n14465_), .Y(new_n14468_));
  INVX1    g14276(.A(new_n14468_), .Y(new_n14469_));
  NAND3X1  g14277(.A(new_n14463_), .B(new_n14444_), .C(new_n3564_), .Y(new_n14470_));
  AOI21X1  g14278(.A0(new_n14470_), .A1(new_n14469_), .B0(new_n14464_), .Y(new_n14471_));
  OR2X1    g14279(.A(new_n14471_), .B(new_n3276_), .Y(new_n14472_));
  OR2X1    g14280(.A(new_n14461_), .B(new_n4165_), .Y(new_n14473_));
  NOR2X1   g14281(.A(new_n14433_), .B(new_n14432_), .Y(new_n14474_));
  INVX1    g14282(.A(new_n14441_), .Y(new_n14475_));
  NAND2X1  g14283(.A(new_n14428_), .B(new_n4165_), .Y(new_n14476_));
  OAI21X1  g14284(.A0(new_n14476_), .A1(new_n14474_), .B0(new_n14475_), .Y(new_n14477_));
  AOI21X1  g14285(.A0(new_n14477_), .A1(new_n14473_), .B0(new_n3863_), .Y(new_n14478_));
  INVX1    g14286(.A(new_n14449_), .Y(new_n14479_));
  AOI21X1  g14287(.A0(new_n14434_), .A1(\asqrt[39] ), .B0(\asqrt[40] ), .Y(new_n14480_));
  AOI21X1  g14288(.A0(new_n14480_), .A1(new_n14477_), .B0(new_n14479_), .Y(new_n14481_));
  NOR3X1   g14289(.A(new_n14481_), .B(new_n14478_), .C(\asqrt[41] ), .Y(new_n14482_));
  NOR2X1   g14290(.A(new_n14482_), .B(new_n14468_), .Y(new_n14483_));
  AND2X1   g14291(.A(new_n13919_), .B(new_n13918_), .Y(new_n14484_));
  NOR4X1   g14292(.A(new_n14165_), .B(new_n14484_), .C(new_n13873_), .D(new_n13917_), .Y(new_n14485_));
  AOI22X1  g14293(.A0(new_n13919_), .A1(new_n13918_), .B0(new_n13891_), .B1(\asqrt[41] ), .Y(new_n14486_));
  AOI21X1  g14294(.A0(new_n14486_), .A1(\asqrt[17] ), .B0(new_n13872_), .Y(new_n14487_));
  NOR2X1   g14295(.A(new_n14487_), .B(new_n14485_), .Y(new_n14488_));
  INVX1    g14296(.A(new_n14488_), .Y(new_n14489_));
  OAI21X1  g14297(.A0(new_n14481_), .A1(new_n14478_), .B0(\asqrt[41] ), .Y(new_n14490_));
  NAND2X1  g14298(.A(new_n14490_), .B(new_n3276_), .Y(new_n14491_));
  OAI21X1  g14299(.A0(new_n14491_), .A1(new_n14483_), .B0(new_n14489_), .Y(new_n14492_));
  AOI21X1  g14300(.A0(new_n14492_), .A1(new_n14472_), .B0(new_n3008_), .Y(new_n14493_));
  AND2X1   g14301(.A(new_n13892_), .B(new_n13884_), .Y(new_n14494_));
  OR4X1    g14302(.A(new_n14165_), .B(new_n14494_), .C(new_n13922_), .D(new_n13885_), .Y(new_n14495_));
  OR2X1    g14303(.A(new_n14494_), .B(new_n13885_), .Y(new_n14496_));
  OAI21X1  g14304(.A0(new_n14496_), .A1(new_n14165_), .B0(new_n13922_), .Y(new_n14497_));
  AND2X1   g14305(.A(new_n14497_), .B(new_n14495_), .Y(new_n14498_));
  OAI21X1  g14306(.A0(new_n14482_), .A1(new_n14468_), .B0(new_n14490_), .Y(new_n14499_));
  AOI21X1  g14307(.A0(new_n14499_), .A1(\asqrt[42] ), .B0(\asqrt[43] ), .Y(new_n14500_));
  AOI21X1  g14308(.A0(new_n14500_), .A1(new_n14492_), .B0(new_n14498_), .Y(new_n14501_));
  OAI21X1  g14309(.A0(new_n14501_), .A1(new_n14493_), .B0(\asqrt[44] ), .Y(new_n14502_));
  NAND3X1  g14310(.A(new_n13927_), .B(new_n13899_), .C(new_n13894_), .Y(new_n14503_));
  NOR3X1   g14311(.A(new_n14165_), .B(new_n13900_), .C(new_n13925_), .Y(new_n14504_));
  OAI22X1  g14312(.A0(new_n14504_), .A1(new_n13899_), .B0(new_n14503_), .B1(new_n14165_), .Y(new_n14505_));
  INVX1    g14313(.A(new_n14505_), .Y(new_n14506_));
  NOR3X1   g14314(.A(new_n14501_), .B(new_n14493_), .C(\asqrt[44] ), .Y(new_n14507_));
  OAI21X1  g14315(.A0(new_n14507_), .A1(new_n14506_), .B0(new_n14502_), .Y(new_n14508_));
  AND2X1   g14316(.A(new_n14508_), .B(\asqrt[45] ), .Y(new_n14509_));
  AND2X1   g14317(.A(new_n14499_), .B(\asqrt[42] ), .Y(new_n14510_));
  OR2X1    g14318(.A(new_n14482_), .B(new_n14468_), .Y(new_n14511_));
  AND2X1   g14319(.A(new_n14490_), .B(new_n3276_), .Y(new_n14512_));
  AOI21X1  g14320(.A0(new_n14512_), .A1(new_n14511_), .B0(new_n14488_), .Y(new_n14513_));
  OAI21X1  g14321(.A0(new_n14513_), .A1(new_n14510_), .B0(\asqrt[43] ), .Y(new_n14514_));
  INVX1    g14322(.A(new_n14498_), .Y(new_n14515_));
  OAI21X1  g14323(.A0(new_n14471_), .A1(new_n3276_), .B0(new_n3008_), .Y(new_n14516_));
  OAI21X1  g14324(.A0(new_n14516_), .A1(new_n14513_), .B0(new_n14515_), .Y(new_n14517_));
  NAND3X1  g14325(.A(new_n14517_), .B(new_n14514_), .C(new_n2769_), .Y(new_n14518_));
  NAND2X1  g14326(.A(new_n14518_), .B(new_n14505_), .Y(new_n14519_));
  OAI21X1  g14327(.A0(new_n13944_), .A1(new_n13942_), .B0(new_n13908_), .Y(new_n14520_));
  NOR3X1   g14328(.A(new_n14520_), .B(new_n14165_), .C(new_n13902_), .Y(new_n14521_));
  AOI22X1  g14329(.A0(new_n13909_), .A1(new_n13903_), .B0(new_n13901_), .B1(\asqrt[44] ), .Y(new_n14522_));
  AOI21X1  g14330(.A0(new_n14522_), .A1(\asqrt[17] ), .B0(new_n13908_), .Y(new_n14523_));
  NOR2X1   g14331(.A(new_n14523_), .B(new_n14521_), .Y(new_n14524_));
  AND2X1   g14332(.A(new_n14502_), .B(new_n2570_), .Y(new_n14525_));
  AOI21X1  g14333(.A0(new_n14525_), .A1(new_n14519_), .B0(new_n14524_), .Y(new_n14526_));
  OAI21X1  g14334(.A0(new_n14526_), .A1(new_n14509_), .B0(\asqrt[46] ), .Y(new_n14527_));
  AND2X1   g14335(.A(new_n13947_), .B(new_n13945_), .Y(new_n14528_));
  OR2X1    g14336(.A(new_n13916_), .B(new_n13946_), .Y(new_n14529_));
  OR2X1    g14337(.A(new_n14529_), .B(new_n14528_), .Y(new_n14530_));
  NOR3X1   g14338(.A(new_n14165_), .B(new_n14528_), .C(new_n13946_), .Y(new_n14531_));
  OAI22X1  g14339(.A0(new_n14531_), .A1(new_n13915_), .B0(new_n14530_), .B1(new_n14165_), .Y(new_n14532_));
  AOI21X1  g14340(.A0(new_n14517_), .A1(new_n14514_), .B0(new_n2769_), .Y(new_n14533_));
  AOI21X1  g14341(.A0(new_n14518_), .A1(new_n14505_), .B0(new_n14533_), .Y(new_n14534_));
  OAI21X1  g14342(.A0(new_n14534_), .A1(new_n2570_), .B0(new_n2263_), .Y(new_n14535_));
  OAI21X1  g14343(.A0(new_n14535_), .A1(new_n14526_), .B0(new_n14532_), .Y(new_n14536_));
  AOI21X1  g14344(.A0(new_n14536_), .A1(new_n14527_), .B0(new_n2040_), .Y(new_n14537_));
  OR4X1    g14345(.A(new_n14165_), .B(new_n13949_), .C(new_n13937_), .D(new_n13931_), .Y(new_n14538_));
  OR2X1    g14346(.A(new_n13949_), .B(new_n13931_), .Y(new_n14539_));
  OAI21X1  g14347(.A0(new_n14539_), .A1(new_n14165_), .B0(new_n13937_), .Y(new_n14540_));
  AND2X1   g14348(.A(new_n14540_), .B(new_n14538_), .Y(new_n14541_));
  INVX1    g14349(.A(new_n14541_), .Y(new_n14542_));
  NAND3X1  g14350(.A(new_n14536_), .B(new_n14527_), .C(new_n2040_), .Y(new_n14543_));
  AOI21X1  g14351(.A0(new_n14543_), .A1(new_n14542_), .B0(new_n14537_), .Y(new_n14544_));
  OR2X1    g14352(.A(new_n14544_), .B(new_n1834_), .Y(new_n14545_));
  OR2X1    g14353(.A(new_n14534_), .B(new_n2570_), .Y(new_n14546_));
  AND2X1   g14354(.A(new_n14518_), .B(new_n14505_), .Y(new_n14547_));
  INVX1    g14355(.A(new_n14524_), .Y(new_n14548_));
  NAND2X1  g14356(.A(new_n14502_), .B(new_n2570_), .Y(new_n14549_));
  OAI21X1  g14357(.A0(new_n14549_), .A1(new_n14547_), .B0(new_n14548_), .Y(new_n14550_));
  AOI21X1  g14358(.A0(new_n14550_), .A1(new_n14546_), .B0(new_n2263_), .Y(new_n14551_));
  INVX1    g14359(.A(new_n14532_), .Y(new_n14552_));
  AOI21X1  g14360(.A0(new_n14508_), .A1(\asqrt[45] ), .B0(\asqrt[46] ), .Y(new_n14553_));
  AOI21X1  g14361(.A0(new_n14553_), .A1(new_n14550_), .B0(new_n14552_), .Y(new_n14554_));
  NOR3X1   g14362(.A(new_n14554_), .B(new_n14551_), .C(\asqrt[47] ), .Y(new_n14555_));
  NOR2X1   g14363(.A(new_n14555_), .B(new_n14541_), .Y(new_n14556_));
  OAI21X1  g14364(.A0(new_n14554_), .A1(new_n14551_), .B0(\asqrt[47] ), .Y(new_n14557_));
  NAND2X1  g14365(.A(new_n14557_), .B(new_n1834_), .Y(new_n14558_));
  AND2X1   g14366(.A(new_n13980_), .B(new_n13979_), .Y(new_n14559_));
  NOR4X1   g14367(.A(new_n14165_), .B(new_n13958_), .C(new_n14559_), .D(new_n13978_), .Y(new_n14560_));
  AOI22X1  g14368(.A0(new_n13980_), .A1(new_n13979_), .B0(new_n13965_), .B1(\asqrt[47] ), .Y(new_n14561_));
  AOI21X1  g14369(.A0(new_n14561_), .A1(\asqrt[17] ), .B0(new_n13957_), .Y(new_n14562_));
  NOR2X1   g14370(.A(new_n14562_), .B(new_n14560_), .Y(new_n14563_));
  INVX1    g14371(.A(new_n14563_), .Y(new_n14564_));
  OAI21X1  g14372(.A0(new_n14558_), .A1(new_n14556_), .B0(new_n14564_), .Y(new_n14565_));
  AOI21X1  g14373(.A0(new_n14565_), .A1(new_n14545_), .B0(new_n1632_), .Y(new_n14566_));
  AND2X1   g14374(.A(new_n13966_), .B(new_n13959_), .Y(new_n14567_));
  OR4X1    g14375(.A(new_n14165_), .B(new_n14567_), .C(new_n13983_), .D(new_n13960_), .Y(new_n14568_));
  OR2X1    g14376(.A(new_n14567_), .B(new_n13960_), .Y(new_n14569_));
  OAI21X1  g14377(.A0(new_n14569_), .A1(new_n14165_), .B0(new_n13983_), .Y(new_n14570_));
  AND2X1   g14378(.A(new_n14570_), .B(new_n14568_), .Y(new_n14571_));
  OAI21X1  g14379(.A0(new_n14555_), .A1(new_n14541_), .B0(new_n14557_), .Y(new_n14572_));
  AOI21X1  g14380(.A0(new_n14572_), .A1(\asqrt[48] ), .B0(\asqrt[49] ), .Y(new_n14573_));
  AOI21X1  g14381(.A0(new_n14573_), .A1(new_n14565_), .B0(new_n14571_), .Y(new_n14574_));
  OAI21X1  g14382(.A0(new_n14574_), .A1(new_n14566_), .B0(\asqrt[50] ), .Y(new_n14575_));
  OR4X1    g14383(.A(new_n14165_), .B(new_n13974_), .C(new_n13977_), .D(new_n14001_), .Y(new_n14576_));
  OR2X1    g14384(.A(new_n13974_), .B(new_n14001_), .Y(new_n14577_));
  OAI21X1  g14385(.A0(new_n14577_), .A1(new_n14165_), .B0(new_n13977_), .Y(new_n14578_));
  AND2X1   g14386(.A(new_n14578_), .B(new_n14576_), .Y(new_n14579_));
  NOR3X1   g14387(.A(new_n14574_), .B(new_n14566_), .C(\asqrt[50] ), .Y(new_n14580_));
  OAI21X1  g14388(.A0(new_n14580_), .A1(new_n14579_), .B0(new_n14575_), .Y(new_n14581_));
  AND2X1   g14389(.A(new_n14581_), .B(\asqrt[51] ), .Y(new_n14582_));
  OR2X1    g14390(.A(new_n14580_), .B(new_n14579_), .Y(new_n14583_));
  OAI21X1  g14391(.A0(new_n14018_), .A1(new_n14016_), .B0(new_n13992_), .Y(new_n14584_));
  NOR3X1   g14392(.A(new_n14584_), .B(new_n14165_), .C(new_n13976_), .Y(new_n14585_));
  AOI22X1  g14393(.A0(new_n13993_), .A1(new_n13987_), .B0(new_n13975_), .B1(\asqrt[50] ), .Y(new_n14586_));
  AOI21X1  g14394(.A0(new_n14586_), .A1(\asqrt[17] ), .B0(new_n13992_), .Y(new_n14587_));
  NOR2X1   g14395(.A(new_n14587_), .B(new_n14585_), .Y(new_n14588_));
  AND2X1   g14396(.A(new_n14575_), .B(new_n1277_), .Y(new_n14589_));
  AOI21X1  g14397(.A0(new_n14589_), .A1(new_n14583_), .B0(new_n14588_), .Y(new_n14590_));
  OAI21X1  g14398(.A0(new_n14590_), .A1(new_n14582_), .B0(\asqrt[52] ), .Y(new_n14591_));
  AND2X1   g14399(.A(new_n14021_), .B(new_n14019_), .Y(new_n14592_));
  OR2X1    g14400(.A(new_n14000_), .B(new_n14020_), .Y(new_n14593_));
  OR2X1    g14401(.A(new_n14593_), .B(new_n14592_), .Y(new_n14594_));
  NOR3X1   g14402(.A(new_n14165_), .B(new_n14592_), .C(new_n14020_), .Y(new_n14595_));
  OAI22X1  g14403(.A0(new_n14595_), .A1(new_n13999_), .B0(new_n14594_), .B1(new_n14165_), .Y(new_n14596_));
  AND2X1   g14404(.A(new_n14572_), .B(\asqrt[48] ), .Y(new_n14597_));
  OR2X1    g14405(.A(new_n14555_), .B(new_n14541_), .Y(new_n14598_));
  AND2X1   g14406(.A(new_n14557_), .B(new_n1834_), .Y(new_n14599_));
  AOI21X1  g14407(.A0(new_n14599_), .A1(new_n14598_), .B0(new_n14563_), .Y(new_n14600_));
  OAI21X1  g14408(.A0(new_n14600_), .A1(new_n14597_), .B0(\asqrt[49] ), .Y(new_n14601_));
  INVX1    g14409(.A(new_n14571_), .Y(new_n14602_));
  OAI21X1  g14410(.A0(new_n14544_), .A1(new_n1834_), .B0(new_n1632_), .Y(new_n14603_));
  OAI21X1  g14411(.A0(new_n14603_), .A1(new_n14600_), .B0(new_n14602_), .Y(new_n14604_));
  AOI21X1  g14412(.A0(new_n14604_), .A1(new_n14601_), .B0(new_n1469_), .Y(new_n14605_));
  INVX1    g14413(.A(new_n14579_), .Y(new_n14606_));
  NAND3X1  g14414(.A(new_n14604_), .B(new_n14601_), .C(new_n1469_), .Y(new_n14607_));
  AOI21X1  g14415(.A0(new_n14607_), .A1(new_n14606_), .B0(new_n14605_), .Y(new_n14608_));
  OAI21X1  g14416(.A0(new_n14608_), .A1(new_n1277_), .B0(new_n1111_), .Y(new_n14609_));
  OAI21X1  g14417(.A0(new_n14609_), .A1(new_n14590_), .B0(new_n14596_), .Y(new_n14610_));
  AOI21X1  g14418(.A0(new_n14610_), .A1(new_n14591_), .B0(new_n968_), .Y(new_n14611_));
  OR4X1    g14419(.A(new_n14165_), .B(new_n14023_), .C(new_n14011_), .D(new_n14005_), .Y(new_n14612_));
  OR2X1    g14420(.A(new_n14023_), .B(new_n14005_), .Y(new_n14613_));
  OAI21X1  g14421(.A0(new_n14613_), .A1(new_n14165_), .B0(new_n14011_), .Y(new_n14614_));
  AND2X1   g14422(.A(new_n14614_), .B(new_n14612_), .Y(new_n14615_));
  INVX1    g14423(.A(new_n14615_), .Y(new_n14616_));
  NAND3X1  g14424(.A(new_n14610_), .B(new_n14591_), .C(new_n968_), .Y(new_n14617_));
  AOI21X1  g14425(.A0(new_n14617_), .A1(new_n14616_), .B0(new_n14611_), .Y(new_n14618_));
  OR2X1    g14426(.A(new_n14618_), .B(new_n902_), .Y(new_n14619_));
  OR2X1    g14427(.A(new_n14608_), .B(new_n1277_), .Y(new_n14620_));
  NOR2X1   g14428(.A(new_n14580_), .B(new_n14579_), .Y(new_n14621_));
  INVX1    g14429(.A(new_n14588_), .Y(new_n14622_));
  NAND2X1  g14430(.A(new_n14575_), .B(new_n1277_), .Y(new_n14623_));
  OAI21X1  g14431(.A0(new_n14623_), .A1(new_n14621_), .B0(new_n14622_), .Y(new_n14624_));
  AOI21X1  g14432(.A0(new_n14624_), .A1(new_n14620_), .B0(new_n1111_), .Y(new_n14625_));
  INVX1    g14433(.A(new_n14596_), .Y(new_n14626_));
  AOI21X1  g14434(.A0(new_n14581_), .A1(\asqrt[51] ), .B0(\asqrt[52] ), .Y(new_n14627_));
  AOI21X1  g14435(.A0(new_n14627_), .A1(new_n14624_), .B0(new_n14626_), .Y(new_n14628_));
  NOR3X1   g14436(.A(new_n14628_), .B(new_n14625_), .C(\asqrt[53] ), .Y(new_n14629_));
  NOR2X1   g14437(.A(new_n14629_), .B(new_n14615_), .Y(new_n14630_));
  AND2X1   g14438(.A(new_n14067_), .B(new_n14066_), .Y(new_n14631_));
  NOR4X1   g14439(.A(new_n14165_), .B(new_n14631_), .C(new_n14030_), .D(new_n14065_), .Y(new_n14632_));
  AOI22X1  g14440(.A0(new_n14067_), .A1(new_n14066_), .B0(new_n14039_), .B1(\asqrt[53] ), .Y(new_n14633_));
  AOI21X1  g14441(.A0(new_n14633_), .A1(\asqrt[17] ), .B0(new_n14029_), .Y(new_n14634_));
  NOR2X1   g14442(.A(new_n14634_), .B(new_n14632_), .Y(new_n14635_));
  INVX1    g14443(.A(new_n14635_), .Y(new_n14636_));
  OAI21X1  g14444(.A0(new_n14628_), .A1(new_n14625_), .B0(\asqrt[53] ), .Y(new_n14637_));
  NAND2X1  g14445(.A(new_n14637_), .B(new_n902_), .Y(new_n14638_));
  OAI21X1  g14446(.A0(new_n14638_), .A1(new_n14630_), .B0(new_n14636_), .Y(new_n14639_));
  AOI21X1  g14447(.A0(new_n14639_), .A1(new_n14619_), .B0(new_n697_), .Y(new_n14640_));
  AND2X1   g14448(.A(new_n14040_), .B(new_n14033_), .Y(new_n14641_));
  OR4X1    g14449(.A(new_n14165_), .B(new_n14641_), .C(new_n14070_), .D(new_n14034_), .Y(new_n14642_));
  OR2X1    g14450(.A(new_n14641_), .B(new_n14034_), .Y(new_n14643_));
  OAI21X1  g14451(.A0(new_n14643_), .A1(new_n14165_), .B0(new_n14070_), .Y(new_n14644_));
  AND2X1   g14452(.A(new_n14644_), .B(new_n14642_), .Y(new_n14645_));
  OAI21X1  g14453(.A0(new_n14629_), .A1(new_n14615_), .B0(new_n14637_), .Y(new_n14646_));
  AOI21X1  g14454(.A0(new_n14646_), .A1(\asqrt[54] ), .B0(\asqrt[55] ), .Y(new_n14647_));
  AOI21X1  g14455(.A0(new_n14647_), .A1(new_n14639_), .B0(new_n14645_), .Y(new_n14648_));
  OAI21X1  g14456(.A0(new_n14648_), .A1(new_n14640_), .B0(\asqrt[56] ), .Y(new_n14649_));
  OR4X1    g14457(.A(new_n14165_), .B(new_n14048_), .C(new_n14074_), .D(new_n14073_), .Y(new_n14650_));
  OR2X1    g14458(.A(new_n14048_), .B(new_n14073_), .Y(new_n14651_));
  OAI21X1  g14459(.A0(new_n14651_), .A1(new_n14165_), .B0(new_n14074_), .Y(new_n14652_));
  AND2X1   g14460(.A(new_n14652_), .B(new_n14650_), .Y(new_n14653_));
  NOR3X1   g14461(.A(new_n14648_), .B(new_n14640_), .C(\asqrt[56] ), .Y(new_n14654_));
  OAI21X1  g14462(.A0(new_n14654_), .A1(new_n14653_), .B0(new_n14649_), .Y(new_n14655_));
  AND2X1   g14463(.A(new_n14655_), .B(\asqrt[57] ), .Y(new_n14656_));
  OR2X1    g14464(.A(new_n14654_), .B(new_n14653_), .Y(new_n14657_));
  OAI21X1  g14465(.A0(new_n14099_), .A1(new_n14097_), .B0(new_n14056_), .Y(new_n14658_));
  NOR3X1   g14466(.A(new_n14658_), .B(new_n14165_), .C(new_n14050_), .Y(new_n14659_));
  AOI22X1  g14467(.A0(new_n14057_), .A1(new_n14051_), .B0(new_n14049_), .B1(\asqrt[56] ), .Y(new_n14660_));
  AOI21X1  g14468(.A0(new_n14660_), .A1(\asqrt[17] ), .B0(new_n14056_), .Y(new_n14661_));
  NOR2X1   g14469(.A(new_n14661_), .B(new_n14659_), .Y(new_n14662_));
  AND2X1   g14470(.A(new_n14649_), .B(new_n481_), .Y(new_n14663_));
  AOI21X1  g14471(.A0(new_n14663_), .A1(new_n14657_), .B0(new_n14662_), .Y(new_n14664_));
  OAI21X1  g14472(.A0(new_n14664_), .A1(new_n14656_), .B0(\asqrt[58] ), .Y(new_n14665_));
  AND2X1   g14473(.A(new_n14102_), .B(new_n14100_), .Y(new_n14666_));
  OR4X1    g14474(.A(new_n14165_), .B(new_n14666_), .C(new_n14064_), .D(new_n14101_), .Y(new_n14667_));
  OR2X1    g14475(.A(new_n14666_), .B(new_n14101_), .Y(new_n14668_));
  OAI21X1  g14476(.A0(new_n14668_), .A1(new_n14165_), .B0(new_n14064_), .Y(new_n14669_));
  AND2X1   g14477(.A(new_n14669_), .B(new_n14667_), .Y(new_n14670_));
  INVX1    g14478(.A(new_n14670_), .Y(new_n14671_));
  AND2X1   g14479(.A(new_n14646_), .B(\asqrt[54] ), .Y(new_n14672_));
  OR2X1    g14480(.A(new_n14629_), .B(new_n14615_), .Y(new_n14673_));
  AND2X1   g14481(.A(new_n14637_), .B(new_n902_), .Y(new_n14674_));
  AOI21X1  g14482(.A0(new_n14674_), .A1(new_n14673_), .B0(new_n14635_), .Y(new_n14675_));
  OAI21X1  g14483(.A0(new_n14675_), .A1(new_n14672_), .B0(\asqrt[55] ), .Y(new_n14676_));
  INVX1    g14484(.A(new_n14645_), .Y(new_n14677_));
  OAI21X1  g14485(.A0(new_n14618_), .A1(new_n902_), .B0(new_n697_), .Y(new_n14678_));
  OAI21X1  g14486(.A0(new_n14678_), .A1(new_n14675_), .B0(new_n14677_), .Y(new_n14679_));
  AOI21X1  g14487(.A0(new_n14679_), .A1(new_n14676_), .B0(new_n582_), .Y(new_n14680_));
  INVX1    g14488(.A(new_n14653_), .Y(new_n14681_));
  NAND3X1  g14489(.A(new_n14679_), .B(new_n14676_), .C(new_n582_), .Y(new_n14682_));
  AOI21X1  g14490(.A0(new_n14682_), .A1(new_n14681_), .B0(new_n14680_), .Y(new_n14683_));
  OAI21X1  g14491(.A0(new_n14683_), .A1(new_n481_), .B0(new_n399_), .Y(new_n14684_));
  OAI21X1  g14492(.A0(new_n14684_), .A1(new_n14664_), .B0(new_n14671_), .Y(new_n14685_));
  AOI21X1  g14493(.A0(new_n14685_), .A1(new_n14665_), .B0(new_n328_), .Y(new_n14686_));
  OR4X1    g14494(.A(new_n14165_), .B(new_n14112_), .C(new_n14085_), .D(new_n14079_), .Y(new_n14687_));
  OR2X1    g14495(.A(new_n14112_), .B(new_n14079_), .Y(new_n14688_));
  OAI21X1  g14496(.A0(new_n14688_), .A1(new_n14165_), .B0(new_n14085_), .Y(new_n14689_));
  AND2X1   g14497(.A(new_n14689_), .B(new_n14687_), .Y(new_n14690_));
  INVX1    g14498(.A(new_n14690_), .Y(new_n14691_));
  NAND3X1  g14499(.A(new_n14685_), .B(new_n14665_), .C(new_n328_), .Y(new_n14692_));
  AOI21X1  g14500(.A0(new_n14692_), .A1(new_n14691_), .B0(new_n14686_), .Y(new_n14693_));
  OR2X1    g14501(.A(new_n14693_), .B(new_n292_), .Y(new_n14694_));
  OR2X1    g14502(.A(new_n14683_), .B(new_n481_), .Y(new_n14695_));
  NOR2X1   g14503(.A(new_n14654_), .B(new_n14653_), .Y(new_n14696_));
  INVX1    g14504(.A(new_n14662_), .Y(new_n14697_));
  NAND2X1  g14505(.A(new_n14649_), .B(new_n481_), .Y(new_n14698_));
  OAI21X1  g14506(.A0(new_n14698_), .A1(new_n14696_), .B0(new_n14697_), .Y(new_n14699_));
  AOI21X1  g14507(.A0(new_n14699_), .A1(new_n14695_), .B0(new_n399_), .Y(new_n14700_));
  AOI21X1  g14508(.A0(new_n14655_), .A1(\asqrt[57] ), .B0(\asqrt[58] ), .Y(new_n14701_));
  AOI21X1  g14509(.A0(new_n14701_), .A1(new_n14699_), .B0(new_n14670_), .Y(new_n14702_));
  NOR3X1   g14510(.A(new_n14702_), .B(new_n14700_), .C(\asqrt[59] ), .Y(new_n14703_));
  NOR2X1   g14511(.A(new_n14703_), .B(new_n14690_), .Y(new_n14704_));
  AND2X1   g14512(.A(new_n14145_), .B(new_n14144_), .Y(new_n14705_));
  NOR4X1   g14513(.A(new_n14165_), .B(new_n14705_), .C(new_n14095_), .D(new_n14143_), .Y(new_n14706_));
  AOI22X1  g14514(.A0(new_n14145_), .A1(new_n14144_), .B0(new_n14113_), .B1(\asqrt[59] ), .Y(new_n14707_));
  AOI21X1  g14515(.A0(new_n14707_), .A1(\asqrt[17] ), .B0(new_n14094_), .Y(new_n14708_));
  NOR2X1   g14516(.A(new_n14708_), .B(new_n14706_), .Y(new_n14709_));
  INVX1    g14517(.A(new_n14709_), .Y(new_n14710_));
  OAI21X1  g14518(.A0(new_n14702_), .A1(new_n14700_), .B0(\asqrt[59] ), .Y(new_n14711_));
  NAND2X1  g14519(.A(new_n14711_), .B(new_n292_), .Y(new_n14712_));
  OAI21X1  g14520(.A0(new_n14712_), .A1(new_n14704_), .B0(new_n14710_), .Y(new_n14713_));
  AOI21X1  g14521(.A0(new_n14713_), .A1(new_n14694_), .B0(new_n217_), .Y(new_n14714_));
  AND2X1   g14522(.A(new_n14114_), .B(new_n14106_), .Y(new_n14715_));
  OR4X1    g14523(.A(new_n14165_), .B(new_n14715_), .C(new_n14148_), .D(new_n14107_), .Y(new_n14716_));
  OR2X1    g14524(.A(new_n14715_), .B(new_n14107_), .Y(new_n14717_));
  OAI21X1  g14525(.A0(new_n14717_), .A1(new_n14165_), .B0(new_n14148_), .Y(new_n14718_));
  AND2X1   g14526(.A(new_n14718_), .B(new_n14716_), .Y(new_n14719_));
  OAI21X1  g14527(.A0(new_n14703_), .A1(new_n14690_), .B0(new_n14711_), .Y(new_n14720_));
  AOI21X1  g14528(.A0(new_n14720_), .A1(\asqrt[60] ), .B0(\asqrt[61] ), .Y(new_n14721_));
  AOI21X1  g14529(.A0(new_n14721_), .A1(new_n14713_), .B0(new_n14719_), .Y(new_n14722_));
  OAI21X1  g14530(.A0(new_n14722_), .A1(new_n14714_), .B0(\asqrt[62] ), .Y(new_n14723_));
  OR4X1    g14531(.A(new_n14165_), .B(new_n14122_), .C(new_n14152_), .D(new_n14151_), .Y(new_n14724_));
  OR2X1    g14532(.A(new_n14122_), .B(new_n14151_), .Y(new_n14725_));
  OAI21X1  g14533(.A0(new_n14725_), .A1(new_n14165_), .B0(new_n14152_), .Y(new_n14726_));
  AND2X1   g14534(.A(new_n14726_), .B(new_n14724_), .Y(new_n14727_));
  NOR3X1   g14535(.A(new_n14722_), .B(new_n14714_), .C(\asqrt[62] ), .Y(new_n14728_));
  OAI21X1  g14536(.A0(new_n14728_), .A1(new_n14727_), .B0(new_n14723_), .Y(new_n14729_));
  AND2X1   g14537(.A(new_n14131_), .B(new_n14125_), .Y(new_n14730_));
  NOR4X1   g14538(.A(new_n14165_), .B(new_n14730_), .C(new_n14184_), .D(new_n14124_), .Y(new_n14731_));
  INVX1    g14539(.A(new_n14731_), .Y(new_n14732_));
  OAI22X1  g14540(.A0(new_n14185_), .A1(new_n14183_), .B0(new_n14154_), .B1(new_n199_), .Y(new_n14733_));
  OAI21X1  g14541(.A0(new_n14733_), .A1(new_n14165_), .B0(new_n14184_), .Y(new_n14734_));
  AND2X1   g14542(.A(new_n14734_), .B(new_n14732_), .Y(new_n14735_));
  INVX1    g14543(.A(new_n14735_), .Y(new_n14736_));
  AND2X1   g14544(.A(new_n14189_), .B(new_n14186_), .Y(new_n14737_));
  AOI21X1  g14545(.A0(new_n14186_), .A1(new_n14182_), .B0(new_n14135_), .Y(new_n14738_));
  AOI21X1  g14546(.A0(new_n14738_), .A1(\asqrt[17] ), .B0(new_n14737_), .Y(new_n14739_));
  AND2X1   g14547(.A(new_n14739_), .B(new_n14736_), .Y(new_n14740_));
  AOI21X1  g14548(.A0(new_n14740_), .A1(new_n14729_), .B0(\asqrt[63] ), .Y(new_n14741_));
  NOR2X1   g14549(.A(new_n14728_), .B(new_n14727_), .Y(new_n14742_));
  NAND2X1  g14550(.A(new_n14735_), .B(new_n14723_), .Y(new_n14743_));
  NAND2X1  g14551(.A(new_n14186_), .B(new_n14182_), .Y(new_n14744_));
  AOI21X1  g14552(.A0(\asqrt[17] ), .A1(new_n14136_), .B0(new_n14744_), .Y(new_n14745_));
  NOR3X1   g14553(.A(new_n14745_), .B(new_n14738_), .C(new_n193_), .Y(new_n14746_));
  AND2X1   g14554(.A(new_n14142_), .B(new_n193_), .Y(new_n14747_));
  OR2X1    g14555(.A(new_n14161_), .B(new_n14133_), .Y(new_n14748_));
  AOI21X1  g14556(.A0(new_n14134_), .A1(new_n13582_), .B0(new_n14748_), .Y(new_n14749_));
  NAND2X1  g14557(.A(new_n14749_), .B(new_n14158_), .Y(new_n14750_));
  NOR3X1   g14558(.A(new_n14750_), .B(new_n14737_), .C(new_n14747_), .Y(new_n14751_));
  NOR2X1   g14559(.A(new_n14751_), .B(new_n14746_), .Y(new_n14752_));
  OAI21X1  g14560(.A0(new_n14743_), .A1(new_n14742_), .B0(new_n14752_), .Y(new_n14753_));
  NOR2X1   g14561(.A(new_n14753_), .B(new_n14741_), .Y(new_n14754_));
  INVX1    g14562(.A(new_n14754_), .Y(\asqrt[16] ));
  OAI21X1  g14563(.A0(new_n14753_), .A1(new_n14741_), .B0(\a[32] ), .Y(new_n14756_));
  INVX1    g14564(.A(\a[32] ), .Y(new_n14757_));
  NOR2X1   g14565(.A(\a[31] ), .B(\a[30] ), .Y(new_n14758_));
  NAND2X1  g14566(.A(new_n14758_), .B(new_n14757_), .Y(new_n14759_));
  AOI21X1  g14567(.A0(new_n14759_), .A1(new_n14756_), .B0(new_n14165_), .Y(new_n14760_));
  AND2X1   g14568(.A(new_n14720_), .B(\asqrt[60] ), .Y(new_n14761_));
  OR2X1    g14569(.A(new_n14703_), .B(new_n14690_), .Y(new_n14762_));
  AND2X1   g14570(.A(new_n14711_), .B(new_n292_), .Y(new_n14763_));
  AOI21X1  g14571(.A0(new_n14763_), .A1(new_n14762_), .B0(new_n14709_), .Y(new_n14764_));
  OAI21X1  g14572(.A0(new_n14764_), .A1(new_n14761_), .B0(\asqrt[61] ), .Y(new_n14765_));
  INVX1    g14573(.A(new_n14719_), .Y(new_n14766_));
  OAI21X1  g14574(.A0(new_n14693_), .A1(new_n292_), .B0(new_n217_), .Y(new_n14767_));
  OAI21X1  g14575(.A0(new_n14767_), .A1(new_n14764_), .B0(new_n14766_), .Y(new_n14768_));
  AOI21X1  g14576(.A0(new_n14768_), .A1(new_n14765_), .B0(new_n199_), .Y(new_n14769_));
  INVX1    g14577(.A(new_n14727_), .Y(new_n14770_));
  NAND3X1  g14578(.A(new_n14768_), .B(new_n14765_), .C(new_n199_), .Y(new_n14771_));
  AOI21X1  g14579(.A0(new_n14771_), .A1(new_n14770_), .B0(new_n14769_), .Y(new_n14772_));
  INVX1    g14580(.A(new_n14740_), .Y(new_n14773_));
  OAI21X1  g14581(.A0(new_n14773_), .A1(new_n14772_), .B0(new_n193_), .Y(new_n14774_));
  OR2X1    g14582(.A(new_n14728_), .B(new_n14727_), .Y(new_n14775_));
  AND2X1   g14583(.A(new_n14735_), .B(new_n14723_), .Y(new_n14776_));
  INVX1    g14584(.A(new_n14752_), .Y(new_n14777_));
  AOI21X1  g14585(.A0(new_n14776_), .A1(new_n14775_), .B0(new_n14777_), .Y(new_n14778_));
  AOI21X1  g14586(.A0(new_n14778_), .A1(new_n14774_), .B0(new_n14757_), .Y(new_n14779_));
  NAND3X1  g14587(.A(new_n14759_), .B(new_n14162_), .C(new_n14158_), .Y(new_n14780_));
  OR4X1    g14588(.A(new_n14780_), .B(new_n14779_), .C(new_n14737_), .D(new_n14747_), .Y(new_n14781_));
  OAI21X1  g14589(.A0(new_n14753_), .A1(new_n14741_), .B0(new_n14757_), .Y(new_n14782_));
  AOI21X1  g14590(.A0(new_n14778_), .A1(new_n14774_), .B0(new_n14167_), .Y(new_n14783_));
  AOI21X1  g14591(.A0(new_n14782_), .A1(\a[33] ), .B0(new_n14783_), .Y(new_n14784_));
  AOI21X1  g14592(.A0(new_n14784_), .A1(new_n14781_), .B0(new_n14760_), .Y(new_n14785_));
  OR2X1    g14593(.A(new_n14785_), .B(new_n13571_), .Y(new_n14786_));
  AND2X1   g14594(.A(new_n14784_), .B(new_n14781_), .Y(new_n14787_));
  OR2X1    g14595(.A(new_n14760_), .B(\asqrt[18] ), .Y(new_n14788_));
  OAI21X1  g14596(.A0(new_n14753_), .A1(new_n14741_), .B0(new_n14166_), .Y(new_n14789_));
  AND2X1   g14597(.A(new_n14776_), .B(new_n14775_), .Y(new_n14790_));
  OR2X1    g14598(.A(new_n14751_), .B(new_n14165_), .Y(new_n14791_));
  OR4X1    g14599(.A(new_n14791_), .B(new_n14746_), .C(new_n14790_), .D(new_n14741_), .Y(new_n14792_));
  AOI21X1  g14600(.A0(new_n14792_), .A1(new_n14789_), .B0(new_n14170_), .Y(new_n14793_));
  NOR4X1   g14601(.A(new_n14791_), .B(new_n14746_), .C(new_n14790_), .D(new_n14741_), .Y(new_n14794_));
  NOR3X1   g14602(.A(new_n14794_), .B(new_n14783_), .C(\a[34] ), .Y(new_n14795_));
  OR2X1    g14603(.A(new_n14795_), .B(new_n14793_), .Y(new_n14796_));
  OAI21X1  g14604(.A0(new_n14788_), .A1(new_n14787_), .B0(new_n14796_), .Y(new_n14797_));
  AOI21X1  g14605(.A0(new_n14797_), .A1(new_n14786_), .B0(new_n13000_), .Y(new_n14798_));
  AND2X1   g14606(.A(new_n14179_), .B(new_n14176_), .Y(new_n14799_));
  NOR3X1   g14607(.A(new_n14799_), .B(new_n14216_), .C(new_n14215_), .Y(new_n14800_));
  OAI21X1  g14608(.A0(new_n14753_), .A1(new_n14741_), .B0(new_n14800_), .Y(new_n14801_));
  AOI21X1  g14609(.A0(new_n14193_), .A1(\asqrt[18] ), .B0(new_n14216_), .Y(new_n14802_));
  OAI21X1  g14610(.A0(new_n14753_), .A1(new_n14741_), .B0(new_n14802_), .Y(new_n14803_));
  NAND2X1  g14611(.A(new_n14803_), .B(new_n14799_), .Y(new_n14804_));
  AND2X1   g14612(.A(new_n14759_), .B(new_n14756_), .Y(new_n14805_));
  NOR4X1   g14613(.A(new_n14780_), .B(new_n14779_), .C(new_n14737_), .D(new_n14747_), .Y(new_n14806_));
  INVX1    g14614(.A(\a[33] ), .Y(new_n14807_));
  AOI21X1  g14615(.A0(new_n14778_), .A1(new_n14774_), .B0(\a[32] ), .Y(new_n14808_));
  OAI21X1  g14616(.A0(new_n14808_), .A1(new_n14807_), .B0(new_n14789_), .Y(new_n14809_));
  OAI22X1  g14617(.A0(new_n14809_), .A1(new_n14806_), .B0(new_n14805_), .B1(new_n14165_), .Y(new_n14810_));
  AOI21X1  g14618(.A0(new_n14810_), .A1(\asqrt[18] ), .B0(\asqrt[19] ), .Y(new_n14811_));
  AOI22X1  g14619(.A0(new_n14811_), .A1(new_n14797_), .B0(new_n14804_), .B1(new_n14801_), .Y(new_n14812_));
  OAI21X1  g14620(.A0(new_n14812_), .A1(new_n14798_), .B0(\asqrt[20] ), .Y(new_n14813_));
  AND2X1   g14621(.A(new_n14194_), .B(new_n14180_), .Y(new_n14814_));
  NOR3X1   g14622(.A(new_n14222_), .B(new_n14814_), .C(new_n14181_), .Y(new_n14815_));
  OAI21X1  g14623(.A0(new_n14753_), .A1(new_n14741_), .B0(new_n14815_), .Y(new_n14816_));
  NOR2X1   g14624(.A(new_n14814_), .B(new_n14181_), .Y(new_n14817_));
  OAI21X1  g14625(.A0(new_n14753_), .A1(new_n14741_), .B0(new_n14817_), .Y(new_n14818_));
  NAND2X1  g14626(.A(new_n14818_), .B(new_n14222_), .Y(new_n14819_));
  AND2X1   g14627(.A(new_n14819_), .B(new_n14816_), .Y(new_n14820_));
  NOR3X1   g14628(.A(new_n14812_), .B(new_n14798_), .C(\asqrt[20] ), .Y(new_n14821_));
  OAI21X1  g14629(.A0(new_n14821_), .A1(new_n14820_), .B0(new_n14813_), .Y(new_n14822_));
  AND2X1   g14630(.A(new_n14822_), .B(\asqrt[21] ), .Y(new_n14823_));
  OR2X1    g14631(.A(new_n14821_), .B(new_n14820_), .Y(new_n14824_));
  NOR3X1   g14632(.A(new_n14211_), .B(new_n14214_), .C(new_n14231_), .Y(new_n14825_));
  NAND3X1  g14633(.A(\asqrt[16] ), .B(new_n14224_), .C(new_n14205_), .Y(new_n14826_));
  AOI22X1  g14634(.A0(new_n14826_), .A1(new_n14214_), .B0(new_n14825_), .B1(\asqrt[16] ), .Y(new_n14827_));
  AND2X1   g14635(.A(new_n14810_), .B(\asqrt[18] ), .Y(new_n14828_));
  NAND2X1  g14636(.A(new_n14784_), .B(new_n14781_), .Y(new_n14829_));
  NOR2X1   g14637(.A(new_n14760_), .B(\asqrt[18] ), .Y(new_n14830_));
  NOR2X1   g14638(.A(new_n14795_), .B(new_n14793_), .Y(new_n14831_));
  AOI21X1  g14639(.A0(new_n14830_), .A1(new_n14829_), .B0(new_n14831_), .Y(new_n14832_));
  OAI21X1  g14640(.A0(new_n14832_), .A1(new_n14828_), .B0(\asqrt[19] ), .Y(new_n14833_));
  NAND2X1  g14641(.A(new_n14804_), .B(new_n14801_), .Y(new_n14834_));
  OAI21X1  g14642(.A0(new_n14785_), .A1(new_n13571_), .B0(new_n13000_), .Y(new_n14835_));
  OAI21X1  g14643(.A0(new_n14835_), .A1(new_n14832_), .B0(new_n14834_), .Y(new_n14836_));
  AOI21X1  g14644(.A0(new_n14836_), .A1(new_n14833_), .B0(new_n12447_), .Y(new_n14837_));
  NOR2X1   g14645(.A(new_n14837_), .B(\asqrt[21] ), .Y(new_n14838_));
  AOI21X1  g14646(.A0(new_n14838_), .A1(new_n14824_), .B0(new_n14827_), .Y(new_n14839_));
  OAI21X1  g14647(.A0(new_n14839_), .A1(new_n14823_), .B0(\asqrt[22] ), .Y(new_n14840_));
  AOI21X1  g14648(.A0(new_n14232_), .A1(new_n14225_), .B0(new_n14270_), .Y(new_n14841_));
  AND2X1   g14649(.A(new_n14841_), .B(new_n14268_), .Y(new_n14842_));
  AOI22X1  g14650(.A0(new_n14232_), .A1(new_n14225_), .B0(new_n14212_), .B1(\asqrt[21] ), .Y(new_n14843_));
  AOI21X1  g14651(.A0(new_n14843_), .A1(\asqrt[16] ), .B0(new_n14230_), .Y(new_n14844_));
  AOI21X1  g14652(.A0(new_n14842_), .A1(\asqrt[16] ), .B0(new_n14844_), .Y(new_n14845_));
  INVX1    g14653(.A(new_n14845_), .Y(new_n14846_));
  INVX1    g14654(.A(new_n14820_), .Y(new_n14847_));
  NAND3X1  g14655(.A(new_n14836_), .B(new_n14833_), .C(new_n12447_), .Y(new_n14848_));
  AOI21X1  g14656(.A0(new_n14848_), .A1(new_n14847_), .B0(new_n14837_), .Y(new_n14849_));
  OAI21X1  g14657(.A0(new_n14849_), .A1(new_n11896_), .B0(new_n11362_), .Y(new_n14850_));
  OAI21X1  g14658(.A0(new_n14850_), .A1(new_n14839_), .B0(new_n14846_), .Y(new_n14851_));
  AOI21X1  g14659(.A0(new_n14851_), .A1(new_n14840_), .B0(new_n10849_), .Y(new_n14852_));
  AND2X1   g14660(.A(new_n14274_), .B(new_n14272_), .Y(new_n14853_));
  NOR3X1   g14661(.A(new_n14853_), .B(new_n14240_), .C(new_n14273_), .Y(new_n14854_));
  NOR3X1   g14662(.A(new_n14754_), .B(new_n14853_), .C(new_n14273_), .Y(new_n14855_));
  NOR2X1   g14663(.A(new_n14855_), .B(new_n14239_), .Y(new_n14856_));
  AOI21X1  g14664(.A0(new_n14854_), .A1(\asqrt[16] ), .B0(new_n14856_), .Y(new_n14857_));
  INVX1    g14665(.A(new_n14857_), .Y(new_n14858_));
  NAND3X1  g14666(.A(new_n14851_), .B(new_n14840_), .C(new_n10849_), .Y(new_n14859_));
  AOI21X1  g14667(.A0(new_n14859_), .A1(new_n14858_), .B0(new_n14852_), .Y(new_n14860_));
  OR2X1    g14668(.A(new_n14860_), .B(new_n10332_), .Y(new_n14861_));
  OR2X1    g14669(.A(new_n14849_), .B(new_n11896_), .Y(new_n14862_));
  NOR2X1   g14670(.A(new_n14821_), .B(new_n14820_), .Y(new_n14863_));
  INVX1    g14671(.A(new_n14827_), .Y(new_n14864_));
  OR2X1    g14672(.A(new_n14837_), .B(\asqrt[21] ), .Y(new_n14865_));
  OAI21X1  g14673(.A0(new_n14865_), .A1(new_n14863_), .B0(new_n14864_), .Y(new_n14866_));
  AOI21X1  g14674(.A0(new_n14866_), .A1(new_n14862_), .B0(new_n11362_), .Y(new_n14867_));
  AOI21X1  g14675(.A0(new_n14822_), .A1(\asqrt[21] ), .B0(\asqrt[22] ), .Y(new_n14868_));
  AOI21X1  g14676(.A0(new_n14868_), .A1(new_n14866_), .B0(new_n14845_), .Y(new_n14869_));
  NOR3X1   g14677(.A(new_n14869_), .B(new_n14867_), .C(\asqrt[23] ), .Y(new_n14870_));
  NOR2X1   g14678(.A(new_n14870_), .B(new_n14857_), .Y(new_n14871_));
  NAND4X1  g14679(.A(\asqrt[16] ), .B(new_n14250_), .C(new_n14248_), .D(new_n14276_), .Y(new_n14872_));
  NAND2X1  g14680(.A(new_n14250_), .B(new_n14276_), .Y(new_n14873_));
  OAI21X1  g14681(.A0(new_n14873_), .A1(new_n14754_), .B0(new_n14249_), .Y(new_n14874_));
  AND2X1   g14682(.A(new_n14874_), .B(new_n14872_), .Y(new_n14875_));
  INVX1    g14683(.A(new_n14875_), .Y(new_n14876_));
  OAI21X1  g14684(.A0(new_n14869_), .A1(new_n14867_), .B0(\asqrt[23] ), .Y(new_n14877_));
  NAND2X1  g14685(.A(new_n14877_), .B(new_n10332_), .Y(new_n14878_));
  OAI21X1  g14686(.A0(new_n14878_), .A1(new_n14871_), .B0(new_n14876_), .Y(new_n14879_));
  AOI21X1  g14687(.A0(new_n14879_), .A1(new_n14861_), .B0(new_n9833_), .Y(new_n14880_));
  AND2X1   g14688(.A(new_n14292_), .B(new_n14291_), .Y(new_n14881_));
  NOR3X1   g14689(.A(new_n14881_), .B(new_n14259_), .C(new_n14290_), .Y(new_n14882_));
  NOR3X1   g14690(.A(new_n14754_), .B(new_n14881_), .C(new_n14290_), .Y(new_n14883_));
  NOR2X1   g14691(.A(new_n14883_), .B(new_n14258_), .Y(new_n14884_));
  AOI21X1  g14692(.A0(new_n14882_), .A1(\asqrt[16] ), .B0(new_n14884_), .Y(new_n14885_));
  OAI21X1  g14693(.A0(new_n14870_), .A1(new_n14857_), .B0(new_n14877_), .Y(new_n14886_));
  AOI21X1  g14694(.A0(new_n14886_), .A1(\asqrt[24] ), .B0(\asqrt[25] ), .Y(new_n14887_));
  AOI21X1  g14695(.A0(new_n14887_), .A1(new_n14879_), .B0(new_n14885_), .Y(new_n14888_));
  OAI21X1  g14696(.A0(new_n14888_), .A1(new_n14880_), .B0(\asqrt[26] ), .Y(new_n14889_));
  AND2X1   g14697(.A(new_n14279_), .B(new_n14261_), .Y(new_n14890_));
  NOR3X1   g14698(.A(new_n14890_), .B(new_n14295_), .C(new_n14262_), .Y(new_n14891_));
  NOR3X1   g14699(.A(new_n14754_), .B(new_n14890_), .C(new_n14262_), .Y(new_n14892_));
  NOR2X1   g14700(.A(new_n14892_), .B(new_n14267_), .Y(new_n14893_));
  AOI21X1  g14701(.A0(new_n14891_), .A1(\asqrt[16] ), .B0(new_n14893_), .Y(new_n14894_));
  NOR3X1   g14702(.A(new_n14888_), .B(new_n14880_), .C(\asqrt[26] ), .Y(new_n14895_));
  OAI21X1  g14703(.A0(new_n14895_), .A1(new_n14894_), .B0(new_n14889_), .Y(new_n14896_));
  AND2X1   g14704(.A(new_n14896_), .B(\asqrt[27] ), .Y(new_n14897_));
  OR2X1    g14705(.A(new_n14895_), .B(new_n14894_), .Y(new_n14898_));
  OR4X1    g14706(.A(new_n14754_), .B(new_n14286_), .C(new_n14289_), .D(new_n14305_), .Y(new_n14899_));
  NAND2X1  g14707(.A(new_n14298_), .B(new_n14281_), .Y(new_n14900_));
  OAI21X1  g14708(.A0(new_n14900_), .A1(new_n14754_), .B0(new_n14289_), .Y(new_n14901_));
  AND2X1   g14709(.A(new_n14901_), .B(new_n14899_), .Y(new_n14902_));
  AND2X1   g14710(.A(new_n14889_), .B(new_n8874_), .Y(new_n14903_));
  AOI21X1  g14711(.A0(new_n14903_), .A1(new_n14898_), .B0(new_n14902_), .Y(new_n14904_));
  OAI21X1  g14712(.A0(new_n14904_), .A1(new_n14897_), .B0(\asqrt[28] ), .Y(new_n14905_));
  AOI21X1  g14713(.A0(new_n14306_), .A1(new_n14299_), .B0(new_n14345_), .Y(new_n14906_));
  AND2X1   g14714(.A(new_n14906_), .B(new_n14343_), .Y(new_n14907_));
  AOI22X1  g14715(.A0(new_n14306_), .A1(new_n14299_), .B0(new_n14287_), .B1(\asqrt[27] ), .Y(new_n14908_));
  AOI21X1  g14716(.A0(new_n14908_), .A1(\asqrt[16] ), .B0(new_n14304_), .Y(new_n14909_));
  AOI21X1  g14717(.A0(new_n14907_), .A1(\asqrt[16] ), .B0(new_n14909_), .Y(new_n14910_));
  INVX1    g14718(.A(new_n14910_), .Y(new_n14911_));
  AND2X1   g14719(.A(new_n14886_), .B(\asqrt[24] ), .Y(new_n14912_));
  OR2X1    g14720(.A(new_n14870_), .B(new_n14857_), .Y(new_n14913_));
  AND2X1   g14721(.A(new_n14877_), .B(new_n10332_), .Y(new_n14914_));
  AOI21X1  g14722(.A0(new_n14914_), .A1(new_n14913_), .B0(new_n14875_), .Y(new_n14915_));
  OAI21X1  g14723(.A0(new_n14915_), .A1(new_n14912_), .B0(\asqrt[25] ), .Y(new_n14916_));
  INVX1    g14724(.A(new_n14885_), .Y(new_n14917_));
  OAI21X1  g14725(.A0(new_n14860_), .A1(new_n10332_), .B0(new_n9833_), .Y(new_n14918_));
  OAI21X1  g14726(.A0(new_n14918_), .A1(new_n14915_), .B0(new_n14917_), .Y(new_n14919_));
  AOI21X1  g14727(.A0(new_n14919_), .A1(new_n14916_), .B0(new_n9353_), .Y(new_n14920_));
  INVX1    g14728(.A(new_n14894_), .Y(new_n14921_));
  NAND3X1  g14729(.A(new_n14919_), .B(new_n14916_), .C(new_n9353_), .Y(new_n14922_));
  AOI21X1  g14730(.A0(new_n14922_), .A1(new_n14921_), .B0(new_n14920_), .Y(new_n14923_));
  OAI21X1  g14731(.A0(new_n14923_), .A1(new_n8874_), .B0(new_n8412_), .Y(new_n14924_));
  OAI21X1  g14732(.A0(new_n14924_), .A1(new_n14904_), .B0(new_n14911_), .Y(new_n14925_));
  AOI21X1  g14733(.A0(new_n14925_), .A1(new_n14905_), .B0(new_n7970_), .Y(new_n14926_));
  AND2X1   g14734(.A(new_n14349_), .B(new_n14347_), .Y(new_n14927_));
  NOR3X1   g14735(.A(new_n14927_), .B(new_n14314_), .C(new_n14348_), .Y(new_n14928_));
  NOR3X1   g14736(.A(new_n14754_), .B(new_n14927_), .C(new_n14348_), .Y(new_n14929_));
  NOR2X1   g14737(.A(new_n14929_), .B(new_n14313_), .Y(new_n14930_));
  AOI21X1  g14738(.A0(new_n14928_), .A1(\asqrt[16] ), .B0(new_n14930_), .Y(new_n14931_));
  INVX1    g14739(.A(new_n14931_), .Y(new_n14932_));
  NAND3X1  g14740(.A(new_n14925_), .B(new_n14905_), .C(new_n7970_), .Y(new_n14933_));
  AOI21X1  g14741(.A0(new_n14933_), .A1(new_n14932_), .B0(new_n14926_), .Y(new_n14934_));
  OR2X1    g14742(.A(new_n14934_), .B(new_n7527_), .Y(new_n14935_));
  AND2X1   g14743(.A(new_n14933_), .B(new_n14932_), .Y(new_n14936_));
  NAND4X1  g14744(.A(\asqrt[16] ), .B(new_n14324_), .C(new_n14322_), .D(new_n14351_), .Y(new_n14937_));
  NAND2X1  g14745(.A(new_n14324_), .B(new_n14351_), .Y(new_n14938_));
  OAI21X1  g14746(.A0(new_n14938_), .A1(new_n14754_), .B0(new_n14323_), .Y(new_n14939_));
  AND2X1   g14747(.A(new_n14939_), .B(new_n14937_), .Y(new_n14940_));
  INVX1    g14748(.A(new_n14940_), .Y(new_n14941_));
  OR2X1    g14749(.A(new_n14926_), .B(\asqrt[30] ), .Y(new_n14942_));
  OAI21X1  g14750(.A0(new_n14942_), .A1(new_n14936_), .B0(new_n14941_), .Y(new_n14943_));
  AOI21X1  g14751(.A0(new_n14943_), .A1(new_n14935_), .B0(new_n7103_), .Y(new_n14944_));
  AND2X1   g14752(.A(new_n14367_), .B(new_n14366_), .Y(new_n14945_));
  NOR3X1   g14753(.A(new_n14945_), .B(new_n14333_), .C(new_n14365_), .Y(new_n14946_));
  NOR3X1   g14754(.A(new_n14754_), .B(new_n14945_), .C(new_n14365_), .Y(new_n14947_));
  NOR2X1   g14755(.A(new_n14947_), .B(new_n14332_), .Y(new_n14948_));
  AOI21X1  g14756(.A0(new_n14946_), .A1(\asqrt[16] ), .B0(new_n14948_), .Y(new_n14949_));
  OR2X1    g14757(.A(new_n14923_), .B(new_n8874_), .Y(new_n14950_));
  NOR2X1   g14758(.A(new_n14895_), .B(new_n14894_), .Y(new_n14951_));
  INVX1    g14759(.A(new_n14902_), .Y(new_n14952_));
  NAND2X1  g14760(.A(new_n14889_), .B(new_n8874_), .Y(new_n14953_));
  OAI21X1  g14761(.A0(new_n14953_), .A1(new_n14951_), .B0(new_n14952_), .Y(new_n14954_));
  AOI21X1  g14762(.A0(new_n14954_), .A1(new_n14950_), .B0(new_n8412_), .Y(new_n14955_));
  AOI21X1  g14763(.A0(new_n14896_), .A1(\asqrt[27] ), .B0(\asqrt[28] ), .Y(new_n14956_));
  AOI21X1  g14764(.A0(new_n14956_), .A1(new_n14954_), .B0(new_n14910_), .Y(new_n14957_));
  OAI21X1  g14765(.A0(new_n14957_), .A1(new_n14955_), .B0(\asqrt[29] ), .Y(new_n14958_));
  NOR3X1   g14766(.A(new_n14957_), .B(new_n14955_), .C(\asqrt[29] ), .Y(new_n14959_));
  OAI21X1  g14767(.A0(new_n14959_), .A1(new_n14931_), .B0(new_n14958_), .Y(new_n14960_));
  AOI21X1  g14768(.A0(new_n14960_), .A1(\asqrt[30] ), .B0(\asqrt[31] ), .Y(new_n14961_));
  AOI21X1  g14769(.A0(new_n14961_), .A1(new_n14943_), .B0(new_n14949_), .Y(new_n14962_));
  OAI21X1  g14770(.A0(new_n14962_), .A1(new_n14944_), .B0(\asqrt[32] ), .Y(new_n14963_));
  AND2X1   g14771(.A(new_n14354_), .B(new_n14335_), .Y(new_n14964_));
  NOR3X1   g14772(.A(new_n14964_), .B(new_n14341_), .C(new_n14336_), .Y(new_n14965_));
  NOR3X1   g14773(.A(new_n14754_), .B(new_n14964_), .C(new_n14336_), .Y(new_n14966_));
  NOR2X1   g14774(.A(new_n14966_), .B(new_n14342_), .Y(new_n14967_));
  AOI21X1  g14775(.A0(new_n14965_), .A1(\asqrt[16] ), .B0(new_n14967_), .Y(new_n14968_));
  NOR3X1   g14776(.A(new_n14962_), .B(new_n14944_), .C(\asqrt[32] ), .Y(new_n14969_));
  OAI21X1  g14777(.A0(new_n14969_), .A1(new_n14968_), .B0(new_n14963_), .Y(new_n14970_));
  AND2X1   g14778(.A(new_n14970_), .B(\asqrt[33] ), .Y(new_n14971_));
  OR2X1    g14779(.A(new_n14969_), .B(new_n14968_), .Y(new_n14972_));
  NAND4X1  g14780(.A(\asqrt[16] ), .B(new_n14372_), .C(new_n14360_), .D(new_n14356_), .Y(new_n14973_));
  NAND2X1  g14781(.A(new_n14372_), .B(new_n14356_), .Y(new_n14974_));
  OAI21X1  g14782(.A0(new_n14974_), .A1(new_n14754_), .B0(new_n14364_), .Y(new_n14975_));
  AND2X1   g14783(.A(new_n14975_), .B(new_n14973_), .Y(new_n14976_));
  AND2X1   g14784(.A(new_n14960_), .B(\asqrt[30] ), .Y(new_n14977_));
  NAND2X1  g14785(.A(new_n14933_), .B(new_n14932_), .Y(new_n14978_));
  NOR2X1   g14786(.A(new_n14926_), .B(\asqrt[30] ), .Y(new_n14979_));
  AOI21X1  g14787(.A0(new_n14979_), .A1(new_n14978_), .B0(new_n14940_), .Y(new_n14980_));
  OAI21X1  g14788(.A0(new_n14980_), .A1(new_n14977_), .B0(\asqrt[31] ), .Y(new_n14981_));
  INVX1    g14789(.A(new_n14949_), .Y(new_n14982_));
  OAI21X1  g14790(.A0(new_n14934_), .A1(new_n7527_), .B0(new_n7103_), .Y(new_n14983_));
  OAI21X1  g14791(.A0(new_n14983_), .A1(new_n14980_), .B0(new_n14982_), .Y(new_n14984_));
  AOI21X1  g14792(.A0(new_n14984_), .A1(new_n14981_), .B0(new_n6699_), .Y(new_n14985_));
  NOR2X1   g14793(.A(new_n14985_), .B(\asqrt[33] ), .Y(new_n14986_));
  AOI21X1  g14794(.A0(new_n14986_), .A1(new_n14972_), .B0(new_n14976_), .Y(new_n14987_));
  OAI21X1  g14795(.A0(new_n14987_), .A1(new_n14971_), .B0(\asqrt[34] ), .Y(new_n14988_));
  AOI21X1  g14796(.A0(new_n14380_), .A1(new_n14373_), .B0(new_n14416_), .Y(new_n14989_));
  AND2X1   g14797(.A(new_n14989_), .B(new_n14414_), .Y(new_n14990_));
  AOI22X1  g14798(.A0(new_n14380_), .A1(new_n14373_), .B0(new_n14362_), .B1(\asqrt[33] ), .Y(new_n14991_));
  AOI21X1  g14799(.A0(new_n14991_), .A1(\asqrt[16] ), .B0(new_n14378_), .Y(new_n14992_));
  AOI21X1  g14800(.A0(new_n14990_), .A1(\asqrt[16] ), .B0(new_n14992_), .Y(new_n14993_));
  INVX1    g14801(.A(new_n14993_), .Y(new_n14994_));
  INVX1    g14802(.A(new_n14968_), .Y(new_n14995_));
  NAND3X1  g14803(.A(new_n14984_), .B(new_n14981_), .C(new_n6699_), .Y(new_n14996_));
  AOI21X1  g14804(.A0(new_n14996_), .A1(new_n14995_), .B0(new_n14985_), .Y(new_n14997_));
  OAI21X1  g14805(.A0(new_n14997_), .A1(new_n6294_), .B0(new_n5941_), .Y(new_n14998_));
  OAI21X1  g14806(.A0(new_n14998_), .A1(new_n14987_), .B0(new_n14994_), .Y(new_n14999_));
  AOI21X1  g14807(.A0(new_n14999_), .A1(new_n14988_), .B0(new_n5541_), .Y(new_n15000_));
  AND2X1   g14808(.A(new_n14420_), .B(new_n14418_), .Y(new_n15001_));
  NOR3X1   g14809(.A(new_n15001_), .B(new_n14388_), .C(new_n14419_), .Y(new_n15002_));
  NOR3X1   g14810(.A(new_n14754_), .B(new_n15001_), .C(new_n14419_), .Y(new_n15003_));
  NOR2X1   g14811(.A(new_n15003_), .B(new_n14387_), .Y(new_n15004_));
  AOI21X1  g14812(.A0(new_n15002_), .A1(\asqrt[16] ), .B0(new_n15004_), .Y(new_n15005_));
  INVX1    g14813(.A(new_n15005_), .Y(new_n15006_));
  NAND3X1  g14814(.A(new_n14999_), .B(new_n14988_), .C(new_n5541_), .Y(new_n15007_));
  AOI21X1  g14815(.A0(new_n15007_), .A1(new_n15006_), .B0(new_n15000_), .Y(new_n15008_));
  OR2X1    g14816(.A(new_n15008_), .B(new_n5176_), .Y(new_n15009_));
  OR2X1    g14817(.A(new_n14997_), .B(new_n6294_), .Y(new_n15010_));
  NOR2X1   g14818(.A(new_n14969_), .B(new_n14968_), .Y(new_n15011_));
  INVX1    g14819(.A(new_n14976_), .Y(new_n15012_));
  OR2X1    g14820(.A(new_n14985_), .B(\asqrt[33] ), .Y(new_n15013_));
  OAI21X1  g14821(.A0(new_n15013_), .A1(new_n15011_), .B0(new_n15012_), .Y(new_n15014_));
  AOI21X1  g14822(.A0(new_n15014_), .A1(new_n15010_), .B0(new_n5941_), .Y(new_n15015_));
  AOI21X1  g14823(.A0(new_n14970_), .A1(\asqrt[33] ), .B0(\asqrt[34] ), .Y(new_n15016_));
  AOI21X1  g14824(.A0(new_n15016_), .A1(new_n15014_), .B0(new_n14993_), .Y(new_n15017_));
  NOR3X1   g14825(.A(new_n15017_), .B(new_n15015_), .C(\asqrt[35] ), .Y(new_n15018_));
  NOR2X1   g14826(.A(new_n15018_), .B(new_n15005_), .Y(new_n15019_));
  OR4X1    g14827(.A(new_n14754_), .B(new_n14424_), .C(new_n14395_), .D(new_n14392_), .Y(new_n15020_));
  NAND2X1  g14828(.A(new_n14396_), .B(new_n14422_), .Y(new_n15021_));
  OAI21X1  g14829(.A0(new_n15021_), .A1(new_n14754_), .B0(new_n14395_), .Y(new_n15022_));
  AND2X1   g14830(.A(new_n15022_), .B(new_n15020_), .Y(new_n15023_));
  INVX1    g14831(.A(new_n15023_), .Y(new_n15024_));
  OAI21X1  g14832(.A0(new_n15017_), .A1(new_n15015_), .B0(\asqrt[35] ), .Y(new_n15025_));
  NAND2X1  g14833(.A(new_n15025_), .B(new_n5176_), .Y(new_n15026_));
  OAI21X1  g14834(.A0(new_n15026_), .A1(new_n15019_), .B0(new_n15024_), .Y(new_n15027_));
  AOI21X1  g14835(.A0(new_n15027_), .A1(new_n15009_), .B0(new_n4826_), .Y(new_n15028_));
  AND2X1   g14836(.A(new_n14452_), .B(new_n14451_), .Y(new_n15029_));
  NOR3X1   g14837(.A(new_n15029_), .B(new_n14405_), .C(new_n14450_), .Y(new_n15030_));
  NOR3X1   g14838(.A(new_n14754_), .B(new_n15029_), .C(new_n14450_), .Y(new_n15031_));
  NOR2X1   g14839(.A(new_n15031_), .B(new_n14404_), .Y(new_n15032_));
  AOI21X1  g14840(.A0(new_n15030_), .A1(\asqrt[16] ), .B0(new_n15032_), .Y(new_n15033_));
  OAI21X1  g14841(.A0(new_n15018_), .A1(new_n15005_), .B0(new_n15025_), .Y(new_n15034_));
  AOI21X1  g14842(.A0(new_n15034_), .A1(\asqrt[36] ), .B0(\asqrt[37] ), .Y(new_n15035_));
  AOI21X1  g14843(.A0(new_n15035_), .A1(new_n15027_), .B0(new_n15033_), .Y(new_n15036_));
  OAI21X1  g14844(.A0(new_n15036_), .A1(new_n15028_), .B0(\asqrt[38] ), .Y(new_n15037_));
  AND2X1   g14845(.A(new_n14426_), .B(new_n14407_), .Y(new_n15038_));
  NOR3X1   g14846(.A(new_n15038_), .B(new_n14455_), .C(new_n14408_), .Y(new_n15039_));
  NOR3X1   g14847(.A(new_n14754_), .B(new_n15038_), .C(new_n14408_), .Y(new_n15040_));
  NOR2X1   g14848(.A(new_n15040_), .B(new_n14413_), .Y(new_n15041_));
  AOI21X1  g14849(.A0(new_n15039_), .A1(\asqrt[16] ), .B0(new_n15041_), .Y(new_n15042_));
  NOR3X1   g14850(.A(new_n15036_), .B(new_n15028_), .C(\asqrt[38] ), .Y(new_n15043_));
  OAI21X1  g14851(.A0(new_n15043_), .A1(new_n15042_), .B0(new_n15037_), .Y(new_n15044_));
  AND2X1   g14852(.A(new_n15044_), .B(\asqrt[39] ), .Y(new_n15045_));
  OR2X1    g14853(.A(new_n15043_), .B(new_n15042_), .Y(new_n15046_));
  OR4X1    g14854(.A(new_n14754_), .B(new_n14433_), .C(new_n14459_), .D(new_n14458_), .Y(new_n15047_));
  OR2X1    g14855(.A(new_n14433_), .B(new_n14458_), .Y(new_n15048_));
  OAI21X1  g14856(.A0(new_n15048_), .A1(new_n14754_), .B0(new_n14459_), .Y(new_n15049_));
  AND2X1   g14857(.A(new_n15049_), .B(new_n15047_), .Y(new_n15050_));
  AND2X1   g14858(.A(new_n15037_), .B(new_n4165_), .Y(new_n15051_));
  AOI21X1  g14859(.A0(new_n15051_), .A1(new_n15046_), .B0(new_n15050_), .Y(new_n15052_));
  OAI21X1  g14860(.A0(new_n15052_), .A1(new_n15045_), .B0(\asqrt[40] ), .Y(new_n15053_));
  AOI21X1  g14861(.A0(new_n14442_), .A1(new_n14436_), .B0(new_n14475_), .Y(new_n15054_));
  AND2X1   g14862(.A(new_n15054_), .B(new_n14473_), .Y(new_n15055_));
  AOI22X1  g14863(.A0(new_n14442_), .A1(new_n14436_), .B0(new_n14434_), .B1(\asqrt[39] ), .Y(new_n15056_));
  AOI21X1  g14864(.A0(new_n15056_), .A1(\asqrt[16] ), .B0(new_n14441_), .Y(new_n15057_));
  AOI21X1  g14865(.A0(new_n15055_), .A1(\asqrt[16] ), .B0(new_n15057_), .Y(new_n15058_));
  INVX1    g14866(.A(new_n15058_), .Y(new_n15059_));
  AND2X1   g14867(.A(new_n15034_), .B(\asqrt[36] ), .Y(new_n15060_));
  OR2X1    g14868(.A(new_n15018_), .B(new_n15005_), .Y(new_n15061_));
  AND2X1   g14869(.A(new_n15025_), .B(new_n5176_), .Y(new_n15062_));
  AOI21X1  g14870(.A0(new_n15062_), .A1(new_n15061_), .B0(new_n15023_), .Y(new_n15063_));
  OAI21X1  g14871(.A0(new_n15063_), .A1(new_n15060_), .B0(\asqrt[37] ), .Y(new_n15064_));
  INVX1    g14872(.A(new_n15033_), .Y(new_n15065_));
  OAI21X1  g14873(.A0(new_n15008_), .A1(new_n5176_), .B0(new_n4826_), .Y(new_n15066_));
  OAI21X1  g14874(.A0(new_n15066_), .A1(new_n15063_), .B0(new_n15065_), .Y(new_n15067_));
  AOI21X1  g14875(.A0(new_n15067_), .A1(new_n15064_), .B0(new_n4493_), .Y(new_n15068_));
  INVX1    g14876(.A(new_n15042_), .Y(new_n15069_));
  NAND3X1  g14877(.A(new_n15067_), .B(new_n15064_), .C(new_n4493_), .Y(new_n15070_));
  AOI21X1  g14878(.A0(new_n15070_), .A1(new_n15069_), .B0(new_n15068_), .Y(new_n15071_));
  OAI21X1  g14879(.A0(new_n15071_), .A1(new_n4165_), .B0(new_n3863_), .Y(new_n15072_));
  OAI21X1  g14880(.A0(new_n15072_), .A1(new_n15052_), .B0(new_n15059_), .Y(new_n15073_));
  AOI21X1  g14881(.A0(new_n15073_), .A1(new_n15053_), .B0(new_n3564_), .Y(new_n15074_));
  AND2X1   g14882(.A(new_n14480_), .B(new_n14477_), .Y(new_n15075_));
  NOR3X1   g14883(.A(new_n15075_), .B(new_n14449_), .C(new_n14478_), .Y(new_n15076_));
  NOR3X1   g14884(.A(new_n14754_), .B(new_n15075_), .C(new_n14478_), .Y(new_n15077_));
  NOR2X1   g14885(.A(new_n15077_), .B(new_n14479_), .Y(new_n15078_));
  AOI21X1  g14886(.A0(new_n15076_), .A1(\asqrt[16] ), .B0(new_n15078_), .Y(new_n15079_));
  INVX1    g14887(.A(new_n15079_), .Y(new_n15080_));
  NAND3X1  g14888(.A(new_n15073_), .B(new_n15053_), .C(new_n3564_), .Y(new_n15081_));
  AOI21X1  g14889(.A0(new_n15081_), .A1(new_n15080_), .B0(new_n15074_), .Y(new_n15082_));
  OR2X1    g14890(.A(new_n15082_), .B(new_n3276_), .Y(new_n15083_));
  OR2X1    g14891(.A(new_n15071_), .B(new_n4165_), .Y(new_n15084_));
  NOR2X1   g14892(.A(new_n15043_), .B(new_n15042_), .Y(new_n15085_));
  INVX1    g14893(.A(new_n15050_), .Y(new_n15086_));
  NAND2X1  g14894(.A(new_n15037_), .B(new_n4165_), .Y(new_n15087_));
  OAI21X1  g14895(.A0(new_n15087_), .A1(new_n15085_), .B0(new_n15086_), .Y(new_n15088_));
  AOI21X1  g14896(.A0(new_n15088_), .A1(new_n15084_), .B0(new_n3863_), .Y(new_n15089_));
  AOI21X1  g14897(.A0(new_n15044_), .A1(\asqrt[39] ), .B0(\asqrt[40] ), .Y(new_n15090_));
  AOI21X1  g14898(.A0(new_n15090_), .A1(new_n15088_), .B0(new_n15058_), .Y(new_n15091_));
  NOR3X1   g14899(.A(new_n15091_), .B(new_n15089_), .C(\asqrt[41] ), .Y(new_n15092_));
  NOR2X1   g14900(.A(new_n15092_), .B(new_n15079_), .Y(new_n15093_));
  OR4X1    g14901(.A(new_n14754_), .B(new_n14482_), .C(new_n14469_), .D(new_n14464_), .Y(new_n15094_));
  OR2X1    g14902(.A(new_n14482_), .B(new_n14464_), .Y(new_n15095_));
  OAI21X1  g14903(.A0(new_n15095_), .A1(new_n14754_), .B0(new_n14469_), .Y(new_n15096_));
  AND2X1   g14904(.A(new_n15096_), .B(new_n15094_), .Y(new_n15097_));
  INVX1    g14905(.A(new_n15097_), .Y(new_n15098_));
  OAI21X1  g14906(.A0(new_n15091_), .A1(new_n15089_), .B0(\asqrt[41] ), .Y(new_n15099_));
  NAND2X1  g14907(.A(new_n15099_), .B(new_n3276_), .Y(new_n15100_));
  OAI21X1  g14908(.A0(new_n15100_), .A1(new_n15093_), .B0(new_n15098_), .Y(new_n15101_));
  AOI21X1  g14909(.A0(new_n15101_), .A1(new_n15083_), .B0(new_n3008_), .Y(new_n15102_));
  AND2X1   g14910(.A(new_n14512_), .B(new_n14511_), .Y(new_n15103_));
  NOR3X1   g14911(.A(new_n15103_), .B(new_n14489_), .C(new_n14510_), .Y(new_n15104_));
  NOR3X1   g14912(.A(new_n14754_), .B(new_n15103_), .C(new_n14510_), .Y(new_n15105_));
  NOR2X1   g14913(.A(new_n15105_), .B(new_n14488_), .Y(new_n15106_));
  AOI21X1  g14914(.A0(new_n15104_), .A1(\asqrt[16] ), .B0(new_n15106_), .Y(new_n15107_));
  OAI21X1  g14915(.A0(new_n15092_), .A1(new_n15079_), .B0(new_n15099_), .Y(new_n15108_));
  AOI21X1  g14916(.A0(new_n15108_), .A1(\asqrt[42] ), .B0(\asqrt[43] ), .Y(new_n15109_));
  AOI21X1  g14917(.A0(new_n15109_), .A1(new_n15101_), .B0(new_n15107_), .Y(new_n15110_));
  OAI21X1  g14918(.A0(new_n15110_), .A1(new_n15102_), .B0(\asqrt[44] ), .Y(new_n15111_));
  AND2X1   g14919(.A(new_n14500_), .B(new_n14492_), .Y(new_n15112_));
  NOR3X1   g14920(.A(new_n15112_), .B(new_n14515_), .C(new_n14493_), .Y(new_n15113_));
  NOR3X1   g14921(.A(new_n14754_), .B(new_n15112_), .C(new_n14493_), .Y(new_n15114_));
  NOR2X1   g14922(.A(new_n15114_), .B(new_n14498_), .Y(new_n15115_));
  AOI21X1  g14923(.A0(new_n15113_), .A1(\asqrt[16] ), .B0(new_n15115_), .Y(new_n15116_));
  NOR3X1   g14924(.A(new_n15110_), .B(new_n15102_), .C(\asqrt[44] ), .Y(new_n15117_));
  OAI21X1  g14925(.A0(new_n15117_), .A1(new_n15116_), .B0(new_n15111_), .Y(new_n15118_));
  AND2X1   g14926(.A(new_n15118_), .B(\asqrt[45] ), .Y(new_n15119_));
  OR2X1    g14927(.A(new_n15117_), .B(new_n15116_), .Y(new_n15120_));
  OR4X1    g14928(.A(new_n14754_), .B(new_n14507_), .C(new_n14505_), .D(new_n14533_), .Y(new_n15121_));
  OR2X1    g14929(.A(new_n14507_), .B(new_n14533_), .Y(new_n15122_));
  OAI21X1  g14930(.A0(new_n15122_), .A1(new_n14754_), .B0(new_n14505_), .Y(new_n15123_));
  AND2X1   g14931(.A(new_n15123_), .B(new_n15121_), .Y(new_n15124_));
  AND2X1   g14932(.A(new_n15111_), .B(new_n2570_), .Y(new_n15125_));
  AOI21X1  g14933(.A0(new_n15125_), .A1(new_n15120_), .B0(new_n15124_), .Y(new_n15126_));
  OAI21X1  g14934(.A0(new_n15126_), .A1(new_n15119_), .B0(\asqrt[46] ), .Y(new_n15127_));
  AOI21X1  g14935(.A0(new_n14525_), .A1(new_n14519_), .B0(new_n14548_), .Y(new_n15128_));
  AND2X1   g14936(.A(new_n15128_), .B(new_n14546_), .Y(new_n15129_));
  AOI22X1  g14937(.A0(new_n14525_), .A1(new_n14519_), .B0(new_n14508_), .B1(\asqrt[45] ), .Y(new_n15130_));
  AOI21X1  g14938(.A0(new_n15130_), .A1(\asqrt[16] ), .B0(new_n14524_), .Y(new_n15131_));
  AOI21X1  g14939(.A0(new_n15129_), .A1(\asqrt[16] ), .B0(new_n15131_), .Y(new_n15132_));
  INVX1    g14940(.A(new_n15132_), .Y(new_n15133_));
  AND2X1   g14941(.A(new_n15108_), .B(\asqrt[42] ), .Y(new_n15134_));
  OR2X1    g14942(.A(new_n15092_), .B(new_n15079_), .Y(new_n15135_));
  AND2X1   g14943(.A(new_n15099_), .B(new_n3276_), .Y(new_n15136_));
  AOI21X1  g14944(.A0(new_n15136_), .A1(new_n15135_), .B0(new_n15097_), .Y(new_n15137_));
  OAI21X1  g14945(.A0(new_n15137_), .A1(new_n15134_), .B0(\asqrt[43] ), .Y(new_n15138_));
  INVX1    g14946(.A(new_n15107_), .Y(new_n15139_));
  OAI21X1  g14947(.A0(new_n15082_), .A1(new_n3276_), .B0(new_n3008_), .Y(new_n15140_));
  OAI21X1  g14948(.A0(new_n15140_), .A1(new_n15137_), .B0(new_n15139_), .Y(new_n15141_));
  AOI21X1  g14949(.A0(new_n15141_), .A1(new_n15138_), .B0(new_n2769_), .Y(new_n15142_));
  INVX1    g14950(.A(new_n15116_), .Y(new_n15143_));
  NAND3X1  g14951(.A(new_n15141_), .B(new_n15138_), .C(new_n2769_), .Y(new_n15144_));
  AOI21X1  g14952(.A0(new_n15144_), .A1(new_n15143_), .B0(new_n15142_), .Y(new_n15145_));
  OAI21X1  g14953(.A0(new_n15145_), .A1(new_n2570_), .B0(new_n2263_), .Y(new_n15146_));
  OAI21X1  g14954(.A0(new_n15146_), .A1(new_n15126_), .B0(new_n15133_), .Y(new_n15147_));
  AOI21X1  g14955(.A0(new_n15147_), .A1(new_n15127_), .B0(new_n2040_), .Y(new_n15148_));
  AND2X1   g14956(.A(new_n14553_), .B(new_n14550_), .Y(new_n15149_));
  NOR3X1   g14957(.A(new_n15149_), .B(new_n14532_), .C(new_n14551_), .Y(new_n15150_));
  NOR3X1   g14958(.A(new_n14754_), .B(new_n15149_), .C(new_n14551_), .Y(new_n15151_));
  NOR2X1   g14959(.A(new_n15151_), .B(new_n14552_), .Y(new_n15152_));
  AOI21X1  g14960(.A0(new_n15150_), .A1(\asqrt[16] ), .B0(new_n15152_), .Y(new_n15153_));
  INVX1    g14961(.A(new_n15153_), .Y(new_n15154_));
  NAND3X1  g14962(.A(new_n15147_), .B(new_n15127_), .C(new_n2040_), .Y(new_n15155_));
  AOI21X1  g14963(.A0(new_n15155_), .A1(new_n15154_), .B0(new_n15148_), .Y(new_n15156_));
  OR2X1    g14964(.A(new_n15156_), .B(new_n1834_), .Y(new_n15157_));
  OR2X1    g14965(.A(new_n15145_), .B(new_n2570_), .Y(new_n15158_));
  NOR2X1   g14966(.A(new_n15117_), .B(new_n15116_), .Y(new_n15159_));
  INVX1    g14967(.A(new_n15124_), .Y(new_n15160_));
  NAND2X1  g14968(.A(new_n15111_), .B(new_n2570_), .Y(new_n15161_));
  OAI21X1  g14969(.A0(new_n15161_), .A1(new_n15159_), .B0(new_n15160_), .Y(new_n15162_));
  AOI21X1  g14970(.A0(new_n15162_), .A1(new_n15158_), .B0(new_n2263_), .Y(new_n15163_));
  AOI21X1  g14971(.A0(new_n15118_), .A1(\asqrt[45] ), .B0(\asqrt[46] ), .Y(new_n15164_));
  AOI21X1  g14972(.A0(new_n15164_), .A1(new_n15162_), .B0(new_n15132_), .Y(new_n15165_));
  NOR3X1   g14973(.A(new_n15165_), .B(new_n15163_), .C(\asqrt[47] ), .Y(new_n15166_));
  NOR2X1   g14974(.A(new_n15166_), .B(new_n15153_), .Y(new_n15167_));
  OR4X1    g14975(.A(new_n14754_), .B(new_n14555_), .C(new_n14542_), .D(new_n14537_), .Y(new_n15168_));
  OR2X1    g14976(.A(new_n14555_), .B(new_n14537_), .Y(new_n15169_));
  OAI21X1  g14977(.A0(new_n15169_), .A1(new_n14754_), .B0(new_n14542_), .Y(new_n15170_));
  AND2X1   g14978(.A(new_n15170_), .B(new_n15168_), .Y(new_n15171_));
  INVX1    g14979(.A(new_n15171_), .Y(new_n15172_));
  OAI21X1  g14980(.A0(new_n15165_), .A1(new_n15163_), .B0(\asqrt[47] ), .Y(new_n15173_));
  NAND2X1  g14981(.A(new_n15173_), .B(new_n1834_), .Y(new_n15174_));
  OAI21X1  g14982(.A0(new_n15174_), .A1(new_n15167_), .B0(new_n15172_), .Y(new_n15175_));
  AOI21X1  g14983(.A0(new_n15175_), .A1(new_n15157_), .B0(new_n1632_), .Y(new_n15176_));
  OAI21X1  g14984(.A0(new_n15166_), .A1(new_n15153_), .B0(new_n15173_), .Y(new_n15177_));
  AOI21X1  g14985(.A0(new_n15177_), .A1(\asqrt[48] ), .B0(\asqrt[49] ), .Y(new_n15178_));
  AND2X1   g14986(.A(new_n14599_), .B(new_n14598_), .Y(new_n15179_));
  NOR3X1   g14987(.A(new_n14564_), .B(new_n15179_), .C(new_n14597_), .Y(new_n15180_));
  NOR3X1   g14988(.A(new_n14754_), .B(new_n15179_), .C(new_n14597_), .Y(new_n15181_));
  NOR2X1   g14989(.A(new_n15181_), .B(new_n14563_), .Y(new_n15182_));
  AOI21X1  g14990(.A0(new_n15180_), .A1(\asqrt[16] ), .B0(new_n15182_), .Y(new_n15183_));
  AOI21X1  g14991(.A0(new_n15178_), .A1(new_n15175_), .B0(new_n15183_), .Y(new_n15184_));
  OAI21X1  g14992(.A0(new_n15184_), .A1(new_n15176_), .B0(\asqrt[50] ), .Y(new_n15185_));
  AND2X1   g14993(.A(new_n14573_), .B(new_n14565_), .Y(new_n15186_));
  NOR3X1   g14994(.A(new_n15186_), .B(new_n14602_), .C(new_n14566_), .Y(new_n15187_));
  NOR3X1   g14995(.A(new_n14754_), .B(new_n15186_), .C(new_n14566_), .Y(new_n15188_));
  NOR2X1   g14996(.A(new_n15188_), .B(new_n14571_), .Y(new_n15189_));
  AOI21X1  g14997(.A0(new_n15187_), .A1(\asqrt[16] ), .B0(new_n15189_), .Y(new_n15190_));
  NOR3X1   g14998(.A(new_n15184_), .B(new_n15176_), .C(\asqrt[50] ), .Y(new_n15191_));
  OAI21X1  g14999(.A0(new_n15191_), .A1(new_n15190_), .B0(new_n15185_), .Y(new_n15192_));
  AND2X1   g15000(.A(new_n15192_), .B(\asqrt[51] ), .Y(new_n15193_));
  OR2X1    g15001(.A(new_n15191_), .B(new_n15190_), .Y(new_n15194_));
  OR4X1    g15002(.A(new_n14754_), .B(new_n14580_), .C(new_n14606_), .D(new_n14605_), .Y(new_n15195_));
  OR2X1    g15003(.A(new_n14580_), .B(new_n14605_), .Y(new_n15196_));
  OAI21X1  g15004(.A0(new_n15196_), .A1(new_n14754_), .B0(new_n14606_), .Y(new_n15197_));
  AND2X1   g15005(.A(new_n15197_), .B(new_n15195_), .Y(new_n15198_));
  AND2X1   g15006(.A(new_n15185_), .B(new_n1277_), .Y(new_n15199_));
  AOI21X1  g15007(.A0(new_n15199_), .A1(new_n15194_), .B0(new_n15198_), .Y(new_n15200_));
  OAI21X1  g15008(.A0(new_n15200_), .A1(new_n15193_), .B0(\asqrt[52] ), .Y(new_n15201_));
  AOI21X1  g15009(.A0(new_n14589_), .A1(new_n14583_), .B0(new_n14622_), .Y(new_n15202_));
  AND2X1   g15010(.A(new_n15202_), .B(new_n14620_), .Y(new_n15203_));
  AOI22X1  g15011(.A0(new_n14589_), .A1(new_n14583_), .B0(new_n14581_), .B1(\asqrt[51] ), .Y(new_n15204_));
  AOI21X1  g15012(.A0(new_n15204_), .A1(\asqrt[16] ), .B0(new_n14588_), .Y(new_n15205_));
  AOI21X1  g15013(.A0(new_n15203_), .A1(\asqrt[16] ), .B0(new_n15205_), .Y(new_n15206_));
  INVX1    g15014(.A(new_n15206_), .Y(new_n15207_));
  AND2X1   g15015(.A(new_n15177_), .B(\asqrt[48] ), .Y(new_n15208_));
  OR2X1    g15016(.A(new_n15166_), .B(new_n15153_), .Y(new_n15209_));
  AND2X1   g15017(.A(new_n15173_), .B(new_n1834_), .Y(new_n15210_));
  AOI21X1  g15018(.A0(new_n15210_), .A1(new_n15209_), .B0(new_n15171_), .Y(new_n15211_));
  OAI21X1  g15019(.A0(new_n15211_), .A1(new_n15208_), .B0(\asqrt[49] ), .Y(new_n15212_));
  OAI21X1  g15020(.A0(new_n15156_), .A1(new_n1834_), .B0(new_n1632_), .Y(new_n15213_));
  INVX1    g15021(.A(new_n15183_), .Y(new_n15214_));
  OAI21X1  g15022(.A0(new_n15213_), .A1(new_n15211_), .B0(new_n15214_), .Y(new_n15215_));
  AOI21X1  g15023(.A0(new_n15215_), .A1(new_n15212_), .B0(new_n1469_), .Y(new_n15216_));
  INVX1    g15024(.A(new_n15190_), .Y(new_n15217_));
  NAND3X1  g15025(.A(new_n15215_), .B(new_n15212_), .C(new_n1469_), .Y(new_n15218_));
  AOI21X1  g15026(.A0(new_n15218_), .A1(new_n15217_), .B0(new_n15216_), .Y(new_n15219_));
  OAI21X1  g15027(.A0(new_n15219_), .A1(new_n1277_), .B0(new_n1111_), .Y(new_n15220_));
  OAI21X1  g15028(.A0(new_n15220_), .A1(new_n15200_), .B0(new_n15207_), .Y(new_n15221_));
  AOI21X1  g15029(.A0(new_n15221_), .A1(new_n15201_), .B0(new_n968_), .Y(new_n15222_));
  AND2X1   g15030(.A(new_n14627_), .B(new_n14624_), .Y(new_n15223_));
  NOR3X1   g15031(.A(new_n15223_), .B(new_n14596_), .C(new_n14625_), .Y(new_n15224_));
  NOR3X1   g15032(.A(new_n14754_), .B(new_n15223_), .C(new_n14625_), .Y(new_n15225_));
  NOR2X1   g15033(.A(new_n15225_), .B(new_n14626_), .Y(new_n15226_));
  AOI21X1  g15034(.A0(new_n15224_), .A1(\asqrt[16] ), .B0(new_n15226_), .Y(new_n15227_));
  INVX1    g15035(.A(new_n15227_), .Y(new_n15228_));
  NAND3X1  g15036(.A(new_n15221_), .B(new_n15201_), .C(new_n968_), .Y(new_n15229_));
  AOI21X1  g15037(.A0(new_n15229_), .A1(new_n15228_), .B0(new_n15222_), .Y(new_n15230_));
  OR2X1    g15038(.A(new_n15230_), .B(new_n902_), .Y(new_n15231_));
  OR2X1    g15039(.A(new_n15219_), .B(new_n1277_), .Y(new_n15232_));
  NOR2X1   g15040(.A(new_n15191_), .B(new_n15190_), .Y(new_n15233_));
  INVX1    g15041(.A(new_n15198_), .Y(new_n15234_));
  NAND2X1  g15042(.A(new_n15185_), .B(new_n1277_), .Y(new_n15235_));
  OAI21X1  g15043(.A0(new_n15235_), .A1(new_n15233_), .B0(new_n15234_), .Y(new_n15236_));
  AOI21X1  g15044(.A0(new_n15236_), .A1(new_n15232_), .B0(new_n1111_), .Y(new_n15237_));
  AOI21X1  g15045(.A0(new_n15192_), .A1(\asqrt[51] ), .B0(\asqrt[52] ), .Y(new_n15238_));
  AOI21X1  g15046(.A0(new_n15238_), .A1(new_n15236_), .B0(new_n15206_), .Y(new_n15239_));
  NOR3X1   g15047(.A(new_n15239_), .B(new_n15237_), .C(\asqrt[53] ), .Y(new_n15240_));
  NOR2X1   g15048(.A(new_n15240_), .B(new_n15227_), .Y(new_n15241_));
  OR4X1    g15049(.A(new_n14754_), .B(new_n14629_), .C(new_n14616_), .D(new_n14611_), .Y(new_n15242_));
  OR2X1    g15050(.A(new_n14629_), .B(new_n14611_), .Y(new_n15243_));
  OAI21X1  g15051(.A0(new_n15243_), .A1(new_n14754_), .B0(new_n14616_), .Y(new_n15244_));
  AND2X1   g15052(.A(new_n15244_), .B(new_n15242_), .Y(new_n15245_));
  INVX1    g15053(.A(new_n15245_), .Y(new_n15246_));
  OAI21X1  g15054(.A0(new_n15239_), .A1(new_n15237_), .B0(\asqrt[53] ), .Y(new_n15247_));
  NAND2X1  g15055(.A(new_n15247_), .B(new_n902_), .Y(new_n15248_));
  OAI21X1  g15056(.A0(new_n15248_), .A1(new_n15241_), .B0(new_n15246_), .Y(new_n15249_));
  AOI21X1  g15057(.A0(new_n15249_), .A1(new_n15231_), .B0(new_n697_), .Y(new_n15250_));
  AND2X1   g15058(.A(new_n14674_), .B(new_n14673_), .Y(new_n15251_));
  NOR3X1   g15059(.A(new_n15251_), .B(new_n14636_), .C(new_n14672_), .Y(new_n15252_));
  NOR3X1   g15060(.A(new_n14754_), .B(new_n15251_), .C(new_n14672_), .Y(new_n15253_));
  NOR2X1   g15061(.A(new_n15253_), .B(new_n14635_), .Y(new_n15254_));
  AOI21X1  g15062(.A0(new_n15252_), .A1(\asqrt[16] ), .B0(new_n15254_), .Y(new_n15255_));
  OAI21X1  g15063(.A0(new_n15240_), .A1(new_n15227_), .B0(new_n15247_), .Y(new_n15256_));
  AOI21X1  g15064(.A0(new_n15256_), .A1(\asqrt[54] ), .B0(\asqrt[55] ), .Y(new_n15257_));
  AOI21X1  g15065(.A0(new_n15257_), .A1(new_n15249_), .B0(new_n15255_), .Y(new_n15258_));
  OAI21X1  g15066(.A0(new_n15258_), .A1(new_n15250_), .B0(\asqrt[56] ), .Y(new_n15259_));
  AND2X1   g15067(.A(new_n14647_), .B(new_n14639_), .Y(new_n15260_));
  NOR3X1   g15068(.A(new_n15260_), .B(new_n14677_), .C(new_n14640_), .Y(new_n15261_));
  NOR3X1   g15069(.A(new_n14754_), .B(new_n15260_), .C(new_n14640_), .Y(new_n15262_));
  NOR2X1   g15070(.A(new_n15262_), .B(new_n14645_), .Y(new_n15263_));
  AOI21X1  g15071(.A0(new_n15261_), .A1(\asqrt[16] ), .B0(new_n15263_), .Y(new_n15264_));
  NOR3X1   g15072(.A(new_n15258_), .B(new_n15250_), .C(\asqrt[56] ), .Y(new_n15265_));
  OAI21X1  g15073(.A0(new_n15265_), .A1(new_n15264_), .B0(new_n15259_), .Y(new_n15266_));
  AND2X1   g15074(.A(new_n15266_), .B(\asqrt[57] ), .Y(new_n15267_));
  OR2X1    g15075(.A(new_n15265_), .B(new_n15264_), .Y(new_n15268_));
  OR4X1    g15076(.A(new_n14754_), .B(new_n14654_), .C(new_n14681_), .D(new_n14680_), .Y(new_n15269_));
  OR2X1    g15077(.A(new_n14654_), .B(new_n14680_), .Y(new_n15270_));
  OAI21X1  g15078(.A0(new_n15270_), .A1(new_n14754_), .B0(new_n14681_), .Y(new_n15271_));
  AND2X1   g15079(.A(new_n15271_), .B(new_n15269_), .Y(new_n15272_));
  AND2X1   g15080(.A(new_n15259_), .B(new_n481_), .Y(new_n15273_));
  AOI21X1  g15081(.A0(new_n15273_), .A1(new_n15268_), .B0(new_n15272_), .Y(new_n15274_));
  OAI21X1  g15082(.A0(new_n15274_), .A1(new_n15267_), .B0(\asqrt[58] ), .Y(new_n15275_));
  AOI21X1  g15083(.A0(new_n14663_), .A1(new_n14657_), .B0(new_n14697_), .Y(new_n15276_));
  AND2X1   g15084(.A(new_n15276_), .B(new_n14695_), .Y(new_n15277_));
  AOI22X1  g15085(.A0(new_n14663_), .A1(new_n14657_), .B0(new_n14655_), .B1(\asqrt[57] ), .Y(new_n15278_));
  AOI21X1  g15086(.A0(new_n15278_), .A1(\asqrt[16] ), .B0(new_n14662_), .Y(new_n15279_));
  AOI21X1  g15087(.A0(new_n15277_), .A1(\asqrt[16] ), .B0(new_n15279_), .Y(new_n15280_));
  INVX1    g15088(.A(new_n15280_), .Y(new_n15281_));
  AND2X1   g15089(.A(new_n15256_), .B(\asqrt[54] ), .Y(new_n15282_));
  OR2X1    g15090(.A(new_n15240_), .B(new_n15227_), .Y(new_n15283_));
  AND2X1   g15091(.A(new_n15247_), .B(new_n902_), .Y(new_n15284_));
  AOI21X1  g15092(.A0(new_n15284_), .A1(new_n15283_), .B0(new_n15245_), .Y(new_n15285_));
  OAI21X1  g15093(.A0(new_n15285_), .A1(new_n15282_), .B0(\asqrt[55] ), .Y(new_n15286_));
  INVX1    g15094(.A(new_n15255_), .Y(new_n15287_));
  OAI21X1  g15095(.A0(new_n15230_), .A1(new_n902_), .B0(new_n697_), .Y(new_n15288_));
  OAI21X1  g15096(.A0(new_n15288_), .A1(new_n15285_), .B0(new_n15287_), .Y(new_n15289_));
  AOI21X1  g15097(.A0(new_n15289_), .A1(new_n15286_), .B0(new_n582_), .Y(new_n15290_));
  INVX1    g15098(.A(new_n15264_), .Y(new_n15291_));
  NAND3X1  g15099(.A(new_n15289_), .B(new_n15286_), .C(new_n582_), .Y(new_n15292_));
  AOI21X1  g15100(.A0(new_n15292_), .A1(new_n15291_), .B0(new_n15290_), .Y(new_n15293_));
  OAI21X1  g15101(.A0(new_n15293_), .A1(new_n481_), .B0(new_n399_), .Y(new_n15294_));
  OAI21X1  g15102(.A0(new_n15294_), .A1(new_n15274_), .B0(new_n15281_), .Y(new_n15295_));
  AOI21X1  g15103(.A0(new_n15295_), .A1(new_n15275_), .B0(new_n328_), .Y(new_n15296_));
  AND2X1   g15104(.A(new_n14701_), .B(new_n14699_), .Y(new_n15297_));
  NOR3X1   g15105(.A(new_n15297_), .B(new_n14671_), .C(new_n14700_), .Y(new_n15298_));
  NOR3X1   g15106(.A(new_n14754_), .B(new_n15297_), .C(new_n14700_), .Y(new_n15299_));
  NOR2X1   g15107(.A(new_n15299_), .B(new_n14670_), .Y(new_n15300_));
  AOI21X1  g15108(.A0(new_n15298_), .A1(\asqrt[16] ), .B0(new_n15300_), .Y(new_n15301_));
  INVX1    g15109(.A(new_n15301_), .Y(new_n15302_));
  NAND3X1  g15110(.A(new_n15295_), .B(new_n15275_), .C(new_n328_), .Y(new_n15303_));
  AOI21X1  g15111(.A0(new_n15303_), .A1(new_n15302_), .B0(new_n15296_), .Y(new_n15304_));
  OR2X1    g15112(.A(new_n15304_), .B(new_n292_), .Y(new_n15305_));
  OR2X1    g15113(.A(new_n15293_), .B(new_n481_), .Y(new_n15306_));
  NOR2X1   g15114(.A(new_n15265_), .B(new_n15264_), .Y(new_n15307_));
  INVX1    g15115(.A(new_n15272_), .Y(new_n15308_));
  NAND2X1  g15116(.A(new_n15259_), .B(new_n481_), .Y(new_n15309_));
  OAI21X1  g15117(.A0(new_n15309_), .A1(new_n15307_), .B0(new_n15308_), .Y(new_n15310_));
  AOI21X1  g15118(.A0(new_n15310_), .A1(new_n15306_), .B0(new_n399_), .Y(new_n15311_));
  AOI21X1  g15119(.A0(new_n15266_), .A1(\asqrt[57] ), .B0(\asqrt[58] ), .Y(new_n15312_));
  AOI21X1  g15120(.A0(new_n15312_), .A1(new_n15310_), .B0(new_n15280_), .Y(new_n15313_));
  NOR3X1   g15121(.A(new_n15313_), .B(new_n15311_), .C(\asqrt[59] ), .Y(new_n15314_));
  NOR2X1   g15122(.A(new_n15314_), .B(new_n15301_), .Y(new_n15315_));
  OR4X1    g15123(.A(new_n14754_), .B(new_n14703_), .C(new_n14691_), .D(new_n14686_), .Y(new_n15316_));
  OR2X1    g15124(.A(new_n14703_), .B(new_n14686_), .Y(new_n15317_));
  OAI21X1  g15125(.A0(new_n15317_), .A1(new_n14754_), .B0(new_n14691_), .Y(new_n15318_));
  AND2X1   g15126(.A(new_n15318_), .B(new_n15316_), .Y(new_n15319_));
  INVX1    g15127(.A(new_n15319_), .Y(new_n15320_));
  OAI21X1  g15128(.A0(new_n15313_), .A1(new_n15311_), .B0(\asqrt[59] ), .Y(new_n15321_));
  NAND2X1  g15129(.A(new_n15321_), .B(new_n292_), .Y(new_n15322_));
  OAI21X1  g15130(.A0(new_n15322_), .A1(new_n15315_), .B0(new_n15320_), .Y(new_n15323_));
  AOI21X1  g15131(.A0(new_n15323_), .A1(new_n15305_), .B0(new_n217_), .Y(new_n15324_));
  AND2X1   g15132(.A(new_n14763_), .B(new_n14762_), .Y(new_n15325_));
  NOR3X1   g15133(.A(new_n15325_), .B(new_n14710_), .C(new_n14761_), .Y(new_n15326_));
  NOR3X1   g15134(.A(new_n14754_), .B(new_n15325_), .C(new_n14761_), .Y(new_n15327_));
  NOR2X1   g15135(.A(new_n15327_), .B(new_n14709_), .Y(new_n15328_));
  AOI21X1  g15136(.A0(new_n15326_), .A1(\asqrt[16] ), .B0(new_n15328_), .Y(new_n15329_));
  OAI21X1  g15137(.A0(new_n15314_), .A1(new_n15301_), .B0(new_n15321_), .Y(new_n15330_));
  AOI21X1  g15138(.A0(new_n15330_), .A1(\asqrt[60] ), .B0(\asqrt[61] ), .Y(new_n15331_));
  AOI21X1  g15139(.A0(new_n15331_), .A1(new_n15323_), .B0(new_n15329_), .Y(new_n15332_));
  OAI21X1  g15140(.A0(new_n15332_), .A1(new_n15324_), .B0(\asqrt[62] ), .Y(new_n15333_));
  AND2X1   g15141(.A(new_n14721_), .B(new_n14713_), .Y(new_n15334_));
  NOR3X1   g15142(.A(new_n15334_), .B(new_n14766_), .C(new_n14714_), .Y(new_n15335_));
  NOR3X1   g15143(.A(new_n14754_), .B(new_n15334_), .C(new_n14714_), .Y(new_n15336_));
  NOR2X1   g15144(.A(new_n15336_), .B(new_n14719_), .Y(new_n15337_));
  AOI21X1  g15145(.A0(new_n15335_), .A1(\asqrt[16] ), .B0(new_n15337_), .Y(new_n15338_));
  NOR3X1   g15146(.A(new_n15332_), .B(new_n15324_), .C(\asqrt[62] ), .Y(new_n15339_));
  OAI21X1  g15147(.A0(new_n15339_), .A1(new_n15338_), .B0(new_n15333_), .Y(new_n15340_));
  NOR4X1   g15148(.A(new_n14754_), .B(new_n14728_), .C(new_n14770_), .D(new_n14769_), .Y(new_n15341_));
  NOR3X1   g15149(.A(new_n14754_), .B(new_n14728_), .C(new_n14769_), .Y(new_n15342_));
  NOR2X1   g15150(.A(new_n15342_), .B(new_n14727_), .Y(new_n15343_));
  NOR2X1   g15151(.A(new_n15343_), .B(new_n15341_), .Y(new_n15344_));
  INVX1    g15152(.A(new_n15344_), .Y(new_n15345_));
  AND2X1   g15153(.A(new_n14736_), .B(new_n14729_), .Y(new_n15346_));
  AOI21X1  g15154(.A0(new_n15346_), .A1(\asqrt[16] ), .B0(new_n14790_), .Y(new_n15347_));
  AND2X1   g15155(.A(new_n15347_), .B(new_n15345_), .Y(new_n15348_));
  AOI21X1  g15156(.A0(new_n15348_), .A1(new_n15340_), .B0(\asqrt[63] ), .Y(new_n15349_));
  NOR2X1   g15157(.A(new_n15339_), .B(new_n15338_), .Y(new_n15350_));
  NAND2X1  g15158(.A(new_n15344_), .B(new_n15333_), .Y(new_n15351_));
  AOI21X1  g15159(.A0(new_n14778_), .A1(new_n14774_), .B0(new_n14735_), .Y(new_n15352_));
  AOI21X1  g15160(.A0(new_n14736_), .A1(new_n14729_), .B0(new_n193_), .Y(new_n15353_));
  OAI21X1  g15161(.A0(new_n15352_), .A1(new_n14729_), .B0(new_n15353_), .Y(new_n15354_));
  INVX1    g15162(.A(new_n14734_), .Y(new_n15355_));
  NOR4X1   g15163(.A(new_n14751_), .B(new_n14746_), .C(new_n15355_), .D(new_n14731_), .Y(new_n15356_));
  OAI21X1  g15164(.A0(new_n14743_), .A1(new_n14742_), .B0(new_n15356_), .Y(new_n15357_));
  NOR2X1   g15165(.A(new_n15357_), .B(new_n14741_), .Y(new_n15358_));
  INVX1    g15166(.A(new_n15358_), .Y(new_n15359_));
  AND2X1   g15167(.A(new_n15359_), .B(new_n15354_), .Y(new_n15360_));
  OAI21X1  g15168(.A0(new_n15351_), .A1(new_n15350_), .B0(new_n15360_), .Y(new_n15361_));
  NOR2X1   g15169(.A(new_n15361_), .B(new_n15349_), .Y(new_n15362_));
  OAI21X1  g15170(.A0(new_n15361_), .A1(new_n15349_), .B0(\a[30] ), .Y(new_n15363_));
  NOR3X1   g15171(.A(\a[30] ), .B(\a[29] ), .C(\a[28] ), .Y(new_n15364_));
  INVX1    g15172(.A(new_n15364_), .Y(new_n15365_));
  AOI21X1  g15173(.A0(new_n15365_), .A1(new_n15363_), .B0(new_n14754_), .Y(new_n15366_));
  OR2X1    g15174(.A(new_n15364_), .B(new_n14751_), .Y(new_n15367_));
  NOR4X1   g15175(.A(new_n15367_), .B(new_n14746_), .C(new_n14790_), .D(new_n14741_), .Y(new_n15368_));
  NAND2X1  g15176(.A(new_n15368_), .B(new_n15363_), .Y(new_n15369_));
  INVX1    g15177(.A(\a[30] ), .Y(new_n15370_));
  OAI21X1  g15178(.A0(new_n15361_), .A1(new_n15349_), .B0(new_n15370_), .Y(new_n15371_));
  INVX1    g15179(.A(new_n14758_), .Y(new_n15372_));
  AND2X1   g15180(.A(new_n15330_), .B(\asqrt[60] ), .Y(new_n15373_));
  OR2X1    g15181(.A(new_n15314_), .B(new_n15301_), .Y(new_n15374_));
  AND2X1   g15182(.A(new_n15321_), .B(new_n292_), .Y(new_n15375_));
  AOI21X1  g15183(.A0(new_n15375_), .A1(new_n15374_), .B0(new_n15319_), .Y(new_n15376_));
  OAI21X1  g15184(.A0(new_n15376_), .A1(new_n15373_), .B0(\asqrt[61] ), .Y(new_n15377_));
  INVX1    g15185(.A(new_n15329_), .Y(new_n15378_));
  OAI21X1  g15186(.A0(new_n15304_), .A1(new_n292_), .B0(new_n217_), .Y(new_n15379_));
  OAI21X1  g15187(.A0(new_n15379_), .A1(new_n15376_), .B0(new_n15378_), .Y(new_n15380_));
  AOI21X1  g15188(.A0(new_n15380_), .A1(new_n15377_), .B0(new_n199_), .Y(new_n15381_));
  INVX1    g15189(.A(new_n15338_), .Y(new_n15382_));
  NAND3X1  g15190(.A(new_n15380_), .B(new_n15377_), .C(new_n199_), .Y(new_n15383_));
  AOI21X1  g15191(.A0(new_n15383_), .A1(new_n15382_), .B0(new_n15381_), .Y(new_n15384_));
  INVX1    g15192(.A(new_n15348_), .Y(new_n15385_));
  OAI21X1  g15193(.A0(new_n15385_), .A1(new_n15384_), .B0(new_n193_), .Y(new_n15386_));
  OR2X1    g15194(.A(new_n15339_), .B(new_n15338_), .Y(new_n15387_));
  AND2X1   g15195(.A(new_n15344_), .B(new_n15333_), .Y(new_n15388_));
  INVX1    g15196(.A(new_n15360_), .Y(new_n15389_));
  AOI21X1  g15197(.A0(new_n15388_), .A1(new_n15387_), .B0(new_n15389_), .Y(new_n15390_));
  AOI21X1  g15198(.A0(new_n15390_), .A1(new_n15386_), .B0(new_n15372_), .Y(new_n15391_));
  AOI21X1  g15199(.A0(new_n15371_), .A1(\a[31] ), .B0(new_n15391_), .Y(new_n15392_));
  AOI21X1  g15200(.A0(new_n15392_), .A1(new_n15369_), .B0(new_n15366_), .Y(new_n15393_));
  OR2X1    g15201(.A(new_n15393_), .B(new_n14165_), .Y(new_n15394_));
  AND2X1   g15202(.A(new_n15392_), .B(new_n15369_), .Y(new_n15395_));
  OR2X1    g15203(.A(new_n15366_), .B(\asqrt[17] ), .Y(new_n15396_));
  OAI21X1  g15204(.A0(new_n15361_), .A1(new_n15349_), .B0(new_n14758_), .Y(new_n15397_));
  INVX1    g15205(.A(new_n15354_), .Y(new_n15398_));
  NOR3X1   g15206(.A(new_n15358_), .B(new_n15398_), .C(new_n14754_), .Y(new_n15399_));
  OAI21X1  g15207(.A0(new_n15351_), .A1(new_n15350_), .B0(new_n15399_), .Y(new_n15400_));
  OR2X1    g15208(.A(new_n15400_), .B(new_n15349_), .Y(new_n15401_));
  AOI21X1  g15209(.A0(new_n15401_), .A1(new_n15397_), .B0(new_n14757_), .Y(new_n15402_));
  OAI21X1  g15210(.A0(new_n15400_), .A1(new_n15349_), .B0(new_n14757_), .Y(new_n15403_));
  NOR2X1   g15211(.A(new_n15403_), .B(new_n15391_), .Y(new_n15404_));
  OR2X1    g15212(.A(new_n15404_), .B(new_n15402_), .Y(new_n15405_));
  OAI21X1  g15213(.A0(new_n15396_), .A1(new_n15395_), .B0(new_n15405_), .Y(new_n15406_));
  AOI21X1  g15214(.A0(new_n15406_), .A1(new_n15394_), .B0(new_n13571_), .Y(new_n15407_));
  NOR3X1   g15215(.A(new_n14784_), .B(new_n14806_), .C(new_n14760_), .Y(new_n15408_));
  OAI21X1  g15216(.A0(new_n15361_), .A1(new_n15349_), .B0(new_n15408_), .Y(new_n15409_));
  NOR2X1   g15217(.A(new_n14806_), .B(new_n14760_), .Y(new_n15410_));
  OAI21X1  g15218(.A0(new_n15361_), .A1(new_n15349_), .B0(new_n15410_), .Y(new_n15411_));
  NAND2X1  g15219(.A(new_n15411_), .B(new_n14784_), .Y(new_n15412_));
  AND2X1   g15220(.A(new_n15412_), .B(new_n15409_), .Y(new_n15413_));
  AOI21X1  g15221(.A0(new_n15390_), .A1(new_n15386_), .B0(new_n15370_), .Y(new_n15414_));
  OAI21X1  g15222(.A0(new_n15364_), .A1(new_n15414_), .B0(\asqrt[16] ), .Y(new_n15415_));
  AND2X1   g15223(.A(new_n15368_), .B(new_n15363_), .Y(new_n15416_));
  INVX1    g15224(.A(\a[31] ), .Y(new_n15417_));
  AOI21X1  g15225(.A0(new_n15390_), .A1(new_n15386_), .B0(\a[30] ), .Y(new_n15418_));
  OAI21X1  g15226(.A0(new_n15418_), .A1(new_n15417_), .B0(new_n15397_), .Y(new_n15419_));
  OAI21X1  g15227(.A0(new_n15419_), .A1(new_n15416_), .B0(new_n15415_), .Y(new_n15420_));
  AOI21X1  g15228(.A0(new_n15420_), .A1(\asqrt[17] ), .B0(\asqrt[18] ), .Y(new_n15421_));
  AOI21X1  g15229(.A0(new_n15421_), .A1(new_n15406_), .B0(new_n15413_), .Y(new_n15422_));
  OAI21X1  g15230(.A0(new_n15422_), .A1(new_n15407_), .B0(\asqrt[19] ), .Y(new_n15423_));
  AOI21X1  g15231(.A0(new_n14830_), .A1(new_n14829_), .B0(new_n14796_), .Y(new_n15424_));
  AND2X1   g15232(.A(new_n15424_), .B(new_n14786_), .Y(new_n15425_));
  OAI21X1  g15233(.A0(new_n15361_), .A1(new_n15349_), .B0(new_n15425_), .Y(new_n15426_));
  AOI22X1  g15234(.A0(new_n14830_), .A1(new_n14829_), .B0(new_n14810_), .B1(\asqrt[18] ), .Y(new_n15427_));
  OAI21X1  g15235(.A0(new_n15361_), .A1(new_n15349_), .B0(new_n15427_), .Y(new_n15428_));
  NAND2X1  g15236(.A(new_n15428_), .B(new_n14796_), .Y(new_n15429_));
  AND2X1   g15237(.A(new_n15429_), .B(new_n15426_), .Y(new_n15430_));
  NOR3X1   g15238(.A(new_n15422_), .B(new_n15407_), .C(\asqrt[19] ), .Y(new_n15431_));
  OAI21X1  g15239(.A0(new_n15431_), .A1(new_n15430_), .B0(new_n15423_), .Y(new_n15432_));
  AND2X1   g15240(.A(new_n15432_), .B(\asqrt[20] ), .Y(new_n15433_));
  OR2X1    g15241(.A(new_n15431_), .B(new_n15430_), .Y(new_n15434_));
  INVX1    g15242(.A(new_n15362_), .Y(\asqrt[15] ));
  AND2X1   g15243(.A(new_n14811_), .B(new_n14797_), .Y(new_n15436_));
  NOR3X1   g15244(.A(new_n15436_), .B(new_n14834_), .C(new_n14798_), .Y(new_n15437_));
  NOR2X1   g15245(.A(new_n15436_), .B(new_n14798_), .Y(new_n15438_));
  OAI21X1  g15246(.A0(new_n15361_), .A1(new_n15349_), .B0(new_n15438_), .Y(new_n15439_));
  AOI22X1  g15247(.A0(new_n15439_), .A1(new_n14834_), .B0(new_n15437_), .B1(\asqrt[15] ), .Y(new_n15440_));
  AND2X1   g15248(.A(new_n15423_), .B(new_n12447_), .Y(new_n15441_));
  AOI21X1  g15249(.A0(new_n15441_), .A1(new_n15434_), .B0(new_n15440_), .Y(new_n15442_));
  OAI21X1  g15250(.A0(new_n15442_), .A1(new_n15433_), .B0(\asqrt[21] ), .Y(new_n15443_));
  NAND4X1  g15251(.A(\asqrt[15] ), .B(new_n14848_), .C(new_n14820_), .D(new_n14813_), .Y(new_n15444_));
  NOR3X1   g15252(.A(new_n15362_), .B(new_n14821_), .C(new_n14837_), .Y(new_n15445_));
  OAI21X1  g15253(.A0(new_n15445_), .A1(new_n14820_), .B0(new_n15444_), .Y(new_n15446_));
  AND2X1   g15254(.A(new_n15420_), .B(\asqrt[17] ), .Y(new_n15447_));
  NAND2X1  g15255(.A(new_n15392_), .B(new_n15369_), .Y(new_n15448_));
  AND2X1   g15256(.A(new_n15415_), .B(new_n14165_), .Y(new_n15449_));
  NOR2X1   g15257(.A(new_n15404_), .B(new_n15402_), .Y(new_n15450_));
  AOI21X1  g15258(.A0(new_n15449_), .A1(new_n15448_), .B0(new_n15450_), .Y(new_n15451_));
  OAI21X1  g15259(.A0(new_n15451_), .A1(new_n15447_), .B0(\asqrt[18] ), .Y(new_n15452_));
  NAND2X1  g15260(.A(new_n15412_), .B(new_n15409_), .Y(new_n15453_));
  OAI21X1  g15261(.A0(new_n15393_), .A1(new_n14165_), .B0(new_n13571_), .Y(new_n15454_));
  OAI21X1  g15262(.A0(new_n15454_), .A1(new_n15451_), .B0(new_n15453_), .Y(new_n15455_));
  AOI21X1  g15263(.A0(new_n15455_), .A1(new_n15452_), .B0(new_n13000_), .Y(new_n15456_));
  INVX1    g15264(.A(new_n15430_), .Y(new_n15457_));
  NAND3X1  g15265(.A(new_n15455_), .B(new_n15452_), .C(new_n13000_), .Y(new_n15458_));
  AOI21X1  g15266(.A0(new_n15458_), .A1(new_n15457_), .B0(new_n15456_), .Y(new_n15459_));
  OAI21X1  g15267(.A0(new_n15459_), .A1(new_n12447_), .B0(new_n11896_), .Y(new_n15460_));
  OAI21X1  g15268(.A0(new_n15460_), .A1(new_n15442_), .B0(new_n15446_), .Y(new_n15461_));
  AOI21X1  g15269(.A0(new_n15461_), .A1(new_n15443_), .B0(new_n11362_), .Y(new_n15462_));
  AND2X1   g15270(.A(new_n14838_), .B(new_n14824_), .Y(new_n15463_));
  NOR3X1   g15271(.A(new_n15463_), .B(new_n14864_), .C(new_n14823_), .Y(new_n15464_));
  NOR3X1   g15272(.A(new_n15362_), .B(new_n15463_), .C(new_n14823_), .Y(new_n15465_));
  NOR2X1   g15273(.A(new_n15465_), .B(new_n14827_), .Y(new_n15466_));
  AOI21X1  g15274(.A0(new_n15464_), .A1(\asqrt[15] ), .B0(new_n15466_), .Y(new_n15467_));
  INVX1    g15275(.A(new_n15467_), .Y(new_n15468_));
  NAND3X1  g15276(.A(new_n15461_), .B(new_n15443_), .C(new_n11362_), .Y(new_n15469_));
  AOI21X1  g15277(.A0(new_n15469_), .A1(new_n15468_), .B0(new_n15462_), .Y(new_n15470_));
  OR2X1    g15278(.A(new_n15470_), .B(new_n10849_), .Y(new_n15471_));
  AND2X1   g15279(.A(new_n15469_), .B(new_n15468_), .Y(new_n15472_));
  AND2X1   g15280(.A(new_n14868_), .B(new_n14866_), .Y(new_n15473_));
  NOR3X1   g15281(.A(new_n15473_), .B(new_n14846_), .C(new_n14867_), .Y(new_n15474_));
  NOR3X1   g15282(.A(new_n15362_), .B(new_n15473_), .C(new_n14867_), .Y(new_n15475_));
  NOR2X1   g15283(.A(new_n15475_), .B(new_n14845_), .Y(new_n15476_));
  AOI21X1  g15284(.A0(new_n15474_), .A1(\asqrt[15] ), .B0(new_n15476_), .Y(new_n15477_));
  INVX1    g15285(.A(new_n15477_), .Y(new_n15478_));
  OR2X1    g15286(.A(new_n15459_), .B(new_n12447_), .Y(new_n15479_));
  NOR2X1   g15287(.A(new_n15431_), .B(new_n15430_), .Y(new_n15480_));
  INVX1    g15288(.A(new_n15440_), .Y(new_n15481_));
  NAND2X1  g15289(.A(new_n15423_), .B(new_n12447_), .Y(new_n15482_));
  OAI21X1  g15290(.A0(new_n15482_), .A1(new_n15480_), .B0(new_n15481_), .Y(new_n15483_));
  AOI21X1  g15291(.A0(new_n15483_), .A1(new_n15479_), .B0(new_n11896_), .Y(new_n15484_));
  INVX1    g15292(.A(new_n15446_), .Y(new_n15485_));
  AOI21X1  g15293(.A0(new_n15432_), .A1(\asqrt[20] ), .B0(\asqrt[21] ), .Y(new_n15486_));
  AOI21X1  g15294(.A0(new_n15486_), .A1(new_n15483_), .B0(new_n15485_), .Y(new_n15487_));
  OAI21X1  g15295(.A0(new_n15487_), .A1(new_n15484_), .B0(\asqrt[22] ), .Y(new_n15488_));
  NAND2X1  g15296(.A(new_n15488_), .B(new_n10849_), .Y(new_n15489_));
  OAI21X1  g15297(.A0(new_n15489_), .A1(new_n15472_), .B0(new_n15478_), .Y(new_n15490_));
  AOI21X1  g15298(.A0(new_n15490_), .A1(new_n15471_), .B0(new_n10332_), .Y(new_n15491_));
  OR4X1    g15299(.A(new_n15362_), .B(new_n14870_), .C(new_n14858_), .D(new_n14852_), .Y(new_n15492_));
  OR2X1    g15300(.A(new_n14870_), .B(new_n14852_), .Y(new_n15493_));
  OAI21X1  g15301(.A0(new_n15493_), .A1(new_n15362_), .B0(new_n14858_), .Y(new_n15494_));
  AND2X1   g15302(.A(new_n15494_), .B(new_n15492_), .Y(new_n15495_));
  NOR3X1   g15303(.A(new_n15487_), .B(new_n15484_), .C(\asqrt[22] ), .Y(new_n15496_));
  OAI21X1  g15304(.A0(new_n15496_), .A1(new_n15467_), .B0(new_n15488_), .Y(new_n15497_));
  AOI21X1  g15305(.A0(new_n15497_), .A1(\asqrt[23] ), .B0(\asqrt[24] ), .Y(new_n15498_));
  AOI21X1  g15306(.A0(new_n15498_), .A1(new_n15490_), .B0(new_n15495_), .Y(new_n15499_));
  OAI21X1  g15307(.A0(new_n15499_), .A1(new_n15491_), .B0(\asqrt[25] ), .Y(new_n15500_));
  AOI21X1  g15308(.A0(new_n14914_), .A1(new_n14913_), .B0(new_n14876_), .Y(new_n15501_));
  AND2X1   g15309(.A(new_n15501_), .B(new_n14861_), .Y(new_n15502_));
  AOI22X1  g15310(.A0(new_n14914_), .A1(new_n14913_), .B0(new_n14886_), .B1(\asqrt[24] ), .Y(new_n15503_));
  AOI21X1  g15311(.A0(new_n15503_), .A1(\asqrt[15] ), .B0(new_n14875_), .Y(new_n15504_));
  AOI21X1  g15312(.A0(new_n15502_), .A1(\asqrt[15] ), .B0(new_n15504_), .Y(new_n15505_));
  NOR3X1   g15313(.A(new_n15499_), .B(new_n15491_), .C(\asqrt[25] ), .Y(new_n15506_));
  OAI21X1  g15314(.A0(new_n15506_), .A1(new_n15505_), .B0(new_n15500_), .Y(new_n15507_));
  AND2X1   g15315(.A(new_n15507_), .B(\asqrt[26] ), .Y(new_n15508_));
  INVX1    g15316(.A(new_n15505_), .Y(new_n15509_));
  AND2X1   g15317(.A(new_n15497_), .B(\asqrt[23] ), .Y(new_n15510_));
  NAND2X1  g15318(.A(new_n15469_), .B(new_n15468_), .Y(new_n15511_));
  AND2X1   g15319(.A(new_n15488_), .B(new_n10849_), .Y(new_n15512_));
  AOI21X1  g15320(.A0(new_n15512_), .A1(new_n15511_), .B0(new_n15477_), .Y(new_n15513_));
  OAI21X1  g15321(.A0(new_n15513_), .A1(new_n15510_), .B0(\asqrt[24] ), .Y(new_n15514_));
  INVX1    g15322(.A(new_n15495_), .Y(new_n15515_));
  OAI21X1  g15323(.A0(new_n15470_), .A1(new_n10849_), .B0(new_n10332_), .Y(new_n15516_));
  OAI21X1  g15324(.A0(new_n15516_), .A1(new_n15513_), .B0(new_n15515_), .Y(new_n15517_));
  NAND3X1  g15325(.A(new_n15517_), .B(new_n15514_), .C(new_n9833_), .Y(new_n15518_));
  NAND2X1  g15326(.A(new_n15518_), .B(new_n15509_), .Y(new_n15519_));
  AND2X1   g15327(.A(new_n14887_), .B(new_n14879_), .Y(new_n15520_));
  NOR3X1   g15328(.A(new_n15520_), .B(new_n14917_), .C(new_n14880_), .Y(new_n15521_));
  NOR3X1   g15329(.A(new_n15362_), .B(new_n15520_), .C(new_n14880_), .Y(new_n15522_));
  NOR2X1   g15330(.A(new_n15522_), .B(new_n14885_), .Y(new_n15523_));
  AOI21X1  g15331(.A0(new_n15521_), .A1(\asqrt[15] ), .B0(new_n15523_), .Y(new_n15524_));
  AND2X1   g15332(.A(new_n15500_), .B(new_n9353_), .Y(new_n15525_));
  AOI21X1  g15333(.A0(new_n15525_), .A1(new_n15519_), .B0(new_n15524_), .Y(new_n15526_));
  OAI21X1  g15334(.A0(new_n15526_), .A1(new_n15508_), .B0(\asqrt[27] ), .Y(new_n15527_));
  OR4X1    g15335(.A(new_n15362_), .B(new_n14895_), .C(new_n14921_), .D(new_n14920_), .Y(new_n15528_));
  OR2X1    g15336(.A(new_n14895_), .B(new_n14920_), .Y(new_n15529_));
  OAI21X1  g15337(.A0(new_n15529_), .A1(new_n15362_), .B0(new_n14921_), .Y(new_n15530_));
  AND2X1   g15338(.A(new_n15530_), .B(new_n15528_), .Y(new_n15531_));
  INVX1    g15339(.A(new_n15531_), .Y(new_n15532_));
  AOI21X1  g15340(.A0(new_n15517_), .A1(new_n15514_), .B0(new_n9833_), .Y(new_n15533_));
  AOI21X1  g15341(.A0(new_n15518_), .A1(new_n15509_), .B0(new_n15533_), .Y(new_n15534_));
  OAI21X1  g15342(.A0(new_n15534_), .A1(new_n9353_), .B0(new_n8874_), .Y(new_n15535_));
  OAI21X1  g15343(.A0(new_n15535_), .A1(new_n15526_), .B0(new_n15532_), .Y(new_n15536_));
  AOI21X1  g15344(.A0(new_n15536_), .A1(new_n15527_), .B0(new_n8412_), .Y(new_n15537_));
  AND2X1   g15345(.A(new_n14903_), .B(new_n14898_), .Y(new_n15538_));
  NOR3X1   g15346(.A(new_n15538_), .B(new_n14952_), .C(new_n14897_), .Y(new_n15539_));
  NOR3X1   g15347(.A(new_n15362_), .B(new_n15538_), .C(new_n14897_), .Y(new_n15540_));
  NOR2X1   g15348(.A(new_n15540_), .B(new_n14902_), .Y(new_n15541_));
  AOI21X1  g15349(.A0(new_n15539_), .A1(\asqrt[15] ), .B0(new_n15541_), .Y(new_n15542_));
  INVX1    g15350(.A(new_n15542_), .Y(new_n15543_));
  NAND3X1  g15351(.A(new_n15536_), .B(new_n15527_), .C(new_n8412_), .Y(new_n15544_));
  AOI21X1  g15352(.A0(new_n15544_), .A1(new_n15543_), .B0(new_n15537_), .Y(new_n15545_));
  OR2X1    g15353(.A(new_n15545_), .B(new_n7970_), .Y(new_n15546_));
  AND2X1   g15354(.A(new_n15544_), .B(new_n15543_), .Y(new_n15547_));
  AND2X1   g15355(.A(new_n14956_), .B(new_n14954_), .Y(new_n15548_));
  NOR3X1   g15356(.A(new_n15548_), .B(new_n14911_), .C(new_n14955_), .Y(new_n15549_));
  NOR3X1   g15357(.A(new_n15362_), .B(new_n15548_), .C(new_n14955_), .Y(new_n15550_));
  NOR2X1   g15358(.A(new_n15550_), .B(new_n14910_), .Y(new_n15551_));
  AOI21X1  g15359(.A0(new_n15549_), .A1(\asqrt[15] ), .B0(new_n15551_), .Y(new_n15552_));
  INVX1    g15360(.A(new_n15552_), .Y(new_n15553_));
  OR2X1    g15361(.A(new_n15534_), .B(new_n9353_), .Y(new_n15554_));
  AND2X1   g15362(.A(new_n15518_), .B(new_n15509_), .Y(new_n15555_));
  INVX1    g15363(.A(new_n15524_), .Y(new_n15556_));
  NAND2X1  g15364(.A(new_n15500_), .B(new_n9353_), .Y(new_n15557_));
  OAI21X1  g15365(.A0(new_n15557_), .A1(new_n15555_), .B0(new_n15556_), .Y(new_n15558_));
  AOI21X1  g15366(.A0(new_n15558_), .A1(new_n15554_), .B0(new_n8874_), .Y(new_n15559_));
  AOI21X1  g15367(.A0(new_n15507_), .A1(\asqrt[26] ), .B0(\asqrt[27] ), .Y(new_n15560_));
  AOI21X1  g15368(.A0(new_n15560_), .A1(new_n15558_), .B0(new_n15531_), .Y(new_n15561_));
  OAI21X1  g15369(.A0(new_n15561_), .A1(new_n15559_), .B0(\asqrt[28] ), .Y(new_n15562_));
  NAND2X1  g15370(.A(new_n15562_), .B(new_n7970_), .Y(new_n15563_));
  OAI21X1  g15371(.A0(new_n15563_), .A1(new_n15547_), .B0(new_n15553_), .Y(new_n15564_));
  AOI21X1  g15372(.A0(new_n15564_), .A1(new_n15546_), .B0(new_n7527_), .Y(new_n15565_));
  NAND4X1  g15373(.A(\asqrt[15] ), .B(new_n14933_), .C(new_n14931_), .D(new_n14958_), .Y(new_n15566_));
  NAND2X1  g15374(.A(new_n14933_), .B(new_n14958_), .Y(new_n15567_));
  OAI21X1  g15375(.A0(new_n15567_), .A1(new_n15362_), .B0(new_n14932_), .Y(new_n15568_));
  AND2X1   g15376(.A(new_n15568_), .B(new_n15566_), .Y(new_n15569_));
  NOR3X1   g15377(.A(new_n15561_), .B(new_n15559_), .C(\asqrt[28] ), .Y(new_n15570_));
  OAI21X1  g15378(.A0(new_n15570_), .A1(new_n15542_), .B0(new_n15562_), .Y(new_n15571_));
  AOI21X1  g15379(.A0(new_n15571_), .A1(\asqrt[29] ), .B0(\asqrt[30] ), .Y(new_n15572_));
  AOI21X1  g15380(.A0(new_n15572_), .A1(new_n15564_), .B0(new_n15569_), .Y(new_n15573_));
  OAI21X1  g15381(.A0(new_n15573_), .A1(new_n15565_), .B0(\asqrt[31] ), .Y(new_n15574_));
  AOI21X1  g15382(.A0(new_n14979_), .A1(new_n14978_), .B0(new_n14941_), .Y(new_n15575_));
  AND2X1   g15383(.A(new_n15575_), .B(new_n14935_), .Y(new_n15576_));
  AOI22X1  g15384(.A0(new_n14979_), .A1(new_n14978_), .B0(new_n14960_), .B1(\asqrt[30] ), .Y(new_n15577_));
  AOI21X1  g15385(.A0(new_n15577_), .A1(\asqrt[15] ), .B0(new_n14940_), .Y(new_n15578_));
  AOI21X1  g15386(.A0(new_n15576_), .A1(\asqrt[15] ), .B0(new_n15578_), .Y(new_n15579_));
  NOR3X1   g15387(.A(new_n15573_), .B(new_n15565_), .C(\asqrt[31] ), .Y(new_n15580_));
  OAI21X1  g15388(.A0(new_n15580_), .A1(new_n15579_), .B0(new_n15574_), .Y(new_n15581_));
  AND2X1   g15389(.A(new_n15581_), .B(\asqrt[32] ), .Y(new_n15582_));
  INVX1    g15390(.A(new_n15579_), .Y(new_n15583_));
  AND2X1   g15391(.A(new_n15571_), .B(\asqrt[29] ), .Y(new_n15584_));
  NAND2X1  g15392(.A(new_n15544_), .B(new_n15543_), .Y(new_n15585_));
  AND2X1   g15393(.A(new_n15562_), .B(new_n7970_), .Y(new_n15586_));
  AOI21X1  g15394(.A0(new_n15586_), .A1(new_n15585_), .B0(new_n15552_), .Y(new_n15587_));
  OAI21X1  g15395(.A0(new_n15587_), .A1(new_n15584_), .B0(\asqrt[30] ), .Y(new_n15588_));
  INVX1    g15396(.A(new_n15569_), .Y(new_n15589_));
  OAI21X1  g15397(.A0(new_n15545_), .A1(new_n7970_), .B0(new_n7527_), .Y(new_n15590_));
  OAI21X1  g15398(.A0(new_n15590_), .A1(new_n15587_), .B0(new_n15589_), .Y(new_n15591_));
  NAND3X1  g15399(.A(new_n15591_), .B(new_n15588_), .C(new_n7103_), .Y(new_n15592_));
  NAND2X1  g15400(.A(new_n15592_), .B(new_n15583_), .Y(new_n15593_));
  AND2X1   g15401(.A(new_n14961_), .B(new_n14943_), .Y(new_n15594_));
  NOR3X1   g15402(.A(new_n15594_), .B(new_n14982_), .C(new_n14944_), .Y(new_n15595_));
  NOR3X1   g15403(.A(new_n15362_), .B(new_n15594_), .C(new_n14944_), .Y(new_n15596_));
  NOR2X1   g15404(.A(new_n15596_), .B(new_n14949_), .Y(new_n15597_));
  AOI21X1  g15405(.A0(new_n15595_), .A1(\asqrt[15] ), .B0(new_n15597_), .Y(new_n15598_));
  AND2X1   g15406(.A(new_n15574_), .B(new_n6699_), .Y(new_n15599_));
  AOI21X1  g15407(.A0(new_n15599_), .A1(new_n15593_), .B0(new_n15598_), .Y(new_n15600_));
  OAI21X1  g15408(.A0(new_n15600_), .A1(new_n15582_), .B0(\asqrt[33] ), .Y(new_n15601_));
  NAND4X1  g15409(.A(\asqrt[15] ), .B(new_n14996_), .C(new_n14968_), .D(new_n14963_), .Y(new_n15602_));
  NAND2X1  g15410(.A(new_n14996_), .B(new_n14963_), .Y(new_n15603_));
  OAI21X1  g15411(.A0(new_n15603_), .A1(new_n15362_), .B0(new_n14995_), .Y(new_n15604_));
  AND2X1   g15412(.A(new_n15604_), .B(new_n15602_), .Y(new_n15605_));
  INVX1    g15413(.A(new_n15605_), .Y(new_n15606_));
  AOI21X1  g15414(.A0(new_n15591_), .A1(new_n15588_), .B0(new_n7103_), .Y(new_n15607_));
  AOI21X1  g15415(.A0(new_n15592_), .A1(new_n15583_), .B0(new_n15607_), .Y(new_n15608_));
  OAI21X1  g15416(.A0(new_n15608_), .A1(new_n6699_), .B0(new_n6294_), .Y(new_n15609_));
  OAI21X1  g15417(.A0(new_n15609_), .A1(new_n15600_), .B0(new_n15606_), .Y(new_n15610_));
  AOI21X1  g15418(.A0(new_n15610_), .A1(new_n15601_), .B0(new_n5941_), .Y(new_n15611_));
  AND2X1   g15419(.A(new_n14986_), .B(new_n14972_), .Y(new_n15612_));
  NOR3X1   g15420(.A(new_n15612_), .B(new_n15012_), .C(new_n14971_), .Y(new_n15613_));
  NOR3X1   g15421(.A(new_n15362_), .B(new_n15612_), .C(new_n14971_), .Y(new_n15614_));
  NOR2X1   g15422(.A(new_n15614_), .B(new_n14976_), .Y(new_n15615_));
  AOI21X1  g15423(.A0(new_n15613_), .A1(\asqrt[15] ), .B0(new_n15615_), .Y(new_n15616_));
  INVX1    g15424(.A(new_n15616_), .Y(new_n15617_));
  NAND3X1  g15425(.A(new_n15610_), .B(new_n15601_), .C(new_n5941_), .Y(new_n15618_));
  AOI21X1  g15426(.A0(new_n15618_), .A1(new_n15617_), .B0(new_n15611_), .Y(new_n15619_));
  OR2X1    g15427(.A(new_n15619_), .B(new_n5541_), .Y(new_n15620_));
  AND2X1   g15428(.A(new_n15618_), .B(new_n15617_), .Y(new_n15621_));
  AND2X1   g15429(.A(new_n15016_), .B(new_n15014_), .Y(new_n15622_));
  NOR3X1   g15430(.A(new_n15622_), .B(new_n14994_), .C(new_n15015_), .Y(new_n15623_));
  NOR3X1   g15431(.A(new_n15362_), .B(new_n15622_), .C(new_n15015_), .Y(new_n15624_));
  NOR2X1   g15432(.A(new_n15624_), .B(new_n14993_), .Y(new_n15625_));
  AOI21X1  g15433(.A0(new_n15623_), .A1(\asqrt[15] ), .B0(new_n15625_), .Y(new_n15626_));
  INVX1    g15434(.A(new_n15626_), .Y(new_n15627_));
  OR2X1    g15435(.A(new_n15608_), .B(new_n6699_), .Y(new_n15628_));
  AND2X1   g15436(.A(new_n15592_), .B(new_n15583_), .Y(new_n15629_));
  INVX1    g15437(.A(new_n15598_), .Y(new_n15630_));
  NAND2X1  g15438(.A(new_n15574_), .B(new_n6699_), .Y(new_n15631_));
  OAI21X1  g15439(.A0(new_n15631_), .A1(new_n15629_), .B0(new_n15630_), .Y(new_n15632_));
  AOI21X1  g15440(.A0(new_n15632_), .A1(new_n15628_), .B0(new_n6294_), .Y(new_n15633_));
  AOI21X1  g15441(.A0(new_n15581_), .A1(\asqrt[32] ), .B0(\asqrt[33] ), .Y(new_n15634_));
  AOI21X1  g15442(.A0(new_n15634_), .A1(new_n15632_), .B0(new_n15605_), .Y(new_n15635_));
  OAI21X1  g15443(.A0(new_n15635_), .A1(new_n15633_), .B0(\asqrt[34] ), .Y(new_n15636_));
  NAND2X1  g15444(.A(new_n15636_), .B(new_n5541_), .Y(new_n15637_));
  OAI21X1  g15445(.A0(new_n15637_), .A1(new_n15621_), .B0(new_n15627_), .Y(new_n15638_));
  AOI21X1  g15446(.A0(new_n15638_), .A1(new_n15620_), .B0(new_n5176_), .Y(new_n15639_));
  NAND4X1  g15447(.A(\asqrt[15] ), .B(new_n15007_), .C(new_n15005_), .D(new_n15025_), .Y(new_n15640_));
  OR2X1    g15448(.A(new_n15018_), .B(new_n15000_), .Y(new_n15641_));
  OAI21X1  g15449(.A0(new_n15641_), .A1(new_n15362_), .B0(new_n15006_), .Y(new_n15642_));
  AND2X1   g15450(.A(new_n15642_), .B(new_n15640_), .Y(new_n15643_));
  NOR3X1   g15451(.A(new_n15635_), .B(new_n15633_), .C(\asqrt[34] ), .Y(new_n15644_));
  OAI21X1  g15452(.A0(new_n15644_), .A1(new_n15616_), .B0(new_n15636_), .Y(new_n15645_));
  AOI21X1  g15453(.A0(new_n15645_), .A1(\asqrt[35] ), .B0(\asqrt[36] ), .Y(new_n15646_));
  AOI21X1  g15454(.A0(new_n15646_), .A1(new_n15638_), .B0(new_n15643_), .Y(new_n15647_));
  OAI21X1  g15455(.A0(new_n15647_), .A1(new_n15639_), .B0(\asqrt[37] ), .Y(new_n15648_));
  AOI21X1  g15456(.A0(new_n15062_), .A1(new_n15061_), .B0(new_n15024_), .Y(new_n15649_));
  AND2X1   g15457(.A(new_n15649_), .B(new_n15009_), .Y(new_n15650_));
  AOI22X1  g15458(.A0(new_n15062_), .A1(new_n15061_), .B0(new_n15034_), .B1(\asqrt[36] ), .Y(new_n15651_));
  AOI21X1  g15459(.A0(new_n15651_), .A1(\asqrt[15] ), .B0(new_n15023_), .Y(new_n15652_));
  AOI21X1  g15460(.A0(new_n15650_), .A1(\asqrt[15] ), .B0(new_n15652_), .Y(new_n15653_));
  NOR3X1   g15461(.A(new_n15647_), .B(new_n15639_), .C(\asqrt[37] ), .Y(new_n15654_));
  OAI21X1  g15462(.A0(new_n15654_), .A1(new_n15653_), .B0(new_n15648_), .Y(new_n15655_));
  AND2X1   g15463(.A(new_n15655_), .B(\asqrt[38] ), .Y(new_n15656_));
  INVX1    g15464(.A(new_n15653_), .Y(new_n15657_));
  AND2X1   g15465(.A(new_n15645_), .B(\asqrt[35] ), .Y(new_n15658_));
  NAND2X1  g15466(.A(new_n15618_), .B(new_n15617_), .Y(new_n15659_));
  AND2X1   g15467(.A(new_n15636_), .B(new_n5541_), .Y(new_n15660_));
  AOI21X1  g15468(.A0(new_n15660_), .A1(new_n15659_), .B0(new_n15626_), .Y(new_n15661_));
  OAI21X1  g15469(.A0(new_n15661_), .A1(new_n15658_), .B0(\asqrt[36] ), .Y(new_n15662_));
  INVX1    g15470(.A(new_n15643_), .Y(new_n15663_));
  OAI21X1  g15471(.A0(new_n15619_), .A1(new_n5541_), .B0(new_n5176_), .Y(new_n15664_));
  OAI21X1  g15472(.A0(new_n15664_), .A1(new_n15661_), .B0(new_n15663_), .Y(new_n15665_));
  NAND3X1  g15473(.A(new_n15665_), .B(new_n15662_), .C(new_n4826_), .Y(new_n15666_));
  NAND2X1  g15474(.A(new_n15666_), .B(new_n15657_), .Y(new_n15667_));
  AND2X1   g15475(.A(new_n15035_), .B(new_n15027_), .Y(new_n15668_));
  NOR3X1   g15476(.A(new_n15668_), .B(new_n15065_), .C(new_n15028_), .Y(new_n15669_));
  NOR3X1   g15477(.A(new_n15362_), .B(new_n15668_), .C(new_n15028_), .Y(new_n15670_));
  NOR2X1   g15478(.A(new_n15670_), .B(new_n15033_), .Y(new_n15671_));
  AOI21X1  g15479(.A0(new_n15669_), .A1(\asqrt[15] ), .B0(new_n15671_), .Y(new_n15672_));
  AND2X1   g15480(.A(new_n15648_), .B(new_n4493_), .Y(new_n15673_));
  AOI21X1  g15481(.A0(new_n15673_), .A1(new_n15667_), .B0(new_n15672_), .Y(new_n15674_));
  OAI21X1  g15482(.A0(new_n15674_), .A1(new_n15656_), .B0(\asqrt[39] ), .Y(new_n15675_));
  NAND4X1  g15483(.A(\asqrt[15] ), .B(new_n15070_), .C(new_n15042_), .D(new_n15037_), .Y(new_n15676_));
  OR2X1    g15484(.A(new_n15043_), .B(new_n15068_), .Y(new_n15677_));
  OAI21X1  g15485(.A0(new_n15677_), .A1(new_n15362_), .B0(new_n15069_), .Y(new_n15678_));
  AND2X1   g15486(.A(new_n15678_), .B(new_n15676_), .Y(new_n15679_));
  INVX1    g15487(.A(new_n15679_), .Y(new_n15680_));
  AOI21X1  g15488(.A0(new_n15665_), .A1(new_n15662_), .B0(new_n4826_), .Y(new_n15681_));
  AOI21X1  g15489(.A0(new_n15666_), .A1(new_n15657_), .B0(new_n15681_), .Y(new_n15682_));
  OAI21X1  g15490(.A0(new_n15682_), .A1(new_n4493_), .B0(new_n4165_), .Y(new_n15683_));
  OAI21X1  g15491(.A0(new_n15683_), .A1(new_n15674_), .B0(new_n15680_), .Y(new_n15684_));
  AOI21X1  g15492(.A0(new_n15684_), .A1(new_n15675_), .B0(new_n3863_), .Y(new_n15685_));
  AND2X1   g15493(.A(new_n15051_), .B(new_n15046_), .Y(new_n15686_));
  NOR3X1   g15494(.A(new_n15686_), .B(new_n15086_), .C(new_n15045_), .Y(new_n15687_));
  NOR3X1   g15495(.A(new_n15362_), .B(new_n15686_), .C(new_n15045_), .Y(new_n15688_));
  NOR2X1   g15496(.A(new_n15688_), .B(new_n15050_), .Y(new_n15689_));
  AOI21X1  g15497(.A0(new_n15687_), .A1(\asqrt[15] ), .B0(new_n15689_), .Y(new_n15690_));
  INVX1    g15498(.A(new_n15690_), .Y(new_n15691_));
  NAND3X1  g15499(.A(new_n15684_), .B(new_n15675_), .C(new_n3863_), .Y(new_n15692_));
  AOI21X1  g15500(.A0(new_n15692_), .A1(new_n15691_), .B0(new_n15685_), .Y(new_n15693_));
  OR2X1    g15501(.A(new_n15693_), .B(new_n3564_), .Y(new_n15694_));
  AND2X1   g15502(.A(new_n15692_), .B(new_n15691_), .Y(new_n15695_));
  AND2X1   g15503(.A(new_n15090_), .B(new_n15088_), .Y(new_n15696_));
  NOR3X1   g15504(.A(new_n15696_), .B(new_n15059_), .C(new_n15089_), .Y(new_n15697_));
  NOR3X1   g15505(.A(new_n15362_), .B(new_n15696_), .C(new_n15089_), .Y(new_n15698_));
  NOR2X1   g15506(.A(new_n15698_), .B(new_n15058_), .Y(new_n15699_));
  AOI21X1  g15507(.A0(new_n15697_), .A1(\asqrt[15] ), .B0(new_n15699_), .Y(new_n15700_));
  INVX1    g15508(.A(new_n15700_), .Y(new_n15701_));
  OR2X1    g15509(.A(new_n15682_), .B(new_n4493_), .Y(new_n15702_));
  AND2X1   g15510(.A(new_n15666_), .B(new_n15657_), .Y(new_n15703_));
  INVX1    g15511(.A(new_n15672_), .Y(new_n15704_));
  NAND2X1  g15512(.A(new_n15648_), .B(new_n4493_), .Y(new_n15705_));
  OAI21X1  g15513(.A0(new_n15705_), .A1(new_n15703_), .B0(new_n15704_), .Y(new_n15706_));
  AOI21X1  g15514(.A0(new_n15706_), .A1(new_n15702_), .B0(new_n4165_), .Y(new_n15707_));
  AOI21X1  g15515(.A0(new_n15655_), .A1(\asqrt[38] ), .B0(\asqrt[39] ), .Y(new_n15708_));
  AOI21X1  g15516(.A0(new_n15708_), .A1(new_n15706_), .B0(new_n15679_), .Y(new_n15709_));
  OAI21X1  g15517(.A0(new_n15709_), .A1(new_n15707_), .B0(\asqrt[40] ), .Y(new_n15710_));
  NAND2X1  g15518(.A(new_n15710_), .B(new_n3564_), .Y(new_n15711_));
  OAI21X1  g15519(.A0(new_n15711_), .A1(new_n15695_), .B0(new_n15701_), .Y(new_n15712_));
  AOI21X1  g15520(.A0(new_n15712_), .A1(new_n15694_), .B0(new_n3276_), .Y(new_n15713_));
  NAND4X1  g15521(.A(\asqrt[15] ), .B(new_n15081_), .C(new_n15079_), .D(new_n15099_), .Y(new_n15714_));
  OR2X1    g15522(.A(new_n15092_), .B(new_n15074_), .Y(new_n15715_));
  OAI21X1  g15523(.A0(new_n15715_), .A1(new_n15362_), .B0(new_n15080_), .Y(new_n15716_));
  AND2X1   g15524(.A(new_n15716_), .B(new_n15714_), .Y(new_n15717_));
  NOR3X1   g15525(.A(new_n15709_), .B(new_n15707_), .C(\asqrt[40] ), .Y(new_n15718_));
  OAI21X1  g15526(.A0(new_n15718_), .A1(new_n15690_), .B0(new_n15710_), .Y(new_n15719_));
  AOI21X1  g15527(.A0(new_n15719_), .A1(\asqrt[41] ), .B0(\asqrt[42] ), .Y(new_n15720_));
  AOI21X1  g15528(.A0(new_n15720_), .A1(new_n15712_), .B0(new_n15717_), .Y(new_n15721_));
  OAI21X1  g15529(.A0(new_n15721_), .A1(new_n15713_), .B0(\asqrt[43] ), .Y(new_n15722_));
  AOI21X1  g15530(.A0(new_n15136_), .A1(new_n15135_), .B0(new_n15098_), .Y(new_n15723_));
  AND2X1   g15531(.A(new_n15723_), .B(new_n15083_), .Y(new_n15724_));
  AOI22X1  g15532(.A0(new_n15136_), .A1(new_n15135_), .B0(new_n15108_), .B1(\asqrt[42] ), .Y(new_n15725_));
  AOI21X1  g15533(.A0(new_n15725_), .A1(\asqrt[15] ), .B0(new_n15097_), .Y(new_n15726_));
  AOI21X1  g15534(.A0(new_n15724_), .A1(\asqrt[15] ), .B0(new_n15726_), .Y(new_n15727_));
  NOR3X1   g15535(.A(new_n15721_), .B(new_n15713_), .C(\asqrt[43] ), .Y(new_n15728_));
  OAI21X1  g15536(.A0(new_n15728_), .A1(new_n15727_), .B0(new_n15722_), .Y(new_n15729_));
  AND2X1   g15537(.A(new_n15729_), .B(\asqrt[44] ), .Y(new_n15730_));
  OR2X1    g15538(.A(new_n15728_), .B(new_n15727_), .Y(new_n15731_));
  AND2X1   g15539(.A(new_n15109_), .B(new_n15101_), .Y(new_n15732_));
  NOR3X1   g15540(.A(new_n15732_), .B(new_n15139_), .C(new_n15102_), .Y(new_n15733_));
  NOR3X1   g15541(.A(new_n15362_), .B(new_n15732_), .C(new_n15102_), .Y(new_n15734_));
  NOR2X1   g15542(.A(new_n15734_), .B(new_n15107_), .Y(new_n15735_));
  AOI21X1  g15543(.A0(new_n15733_), .A1(\asqrt[15] ), .B0(new_n15735_), .Y(new_n15736_));
  AND2X1   g15544(.A(new_n15722_), .B(new_n2769_), .Y(new_n15737_));
  AOI21X1  g15545(.A0(new_n15737_), .A1(new_n15731_), .B0(new_n15736_), .Y(new_n15738_));
  OAI21X1  g15546(.A0(new_n15738_), .A1(new_n15730_), .B0(\asqrt[45] ), .Y(new_n15739_));
  OR4X1    g15547(.A(new_n15362_), .B(new_n15117_), .C(new_n15143_), .D(new_n15142_), .Y(new_n15740_));
  OR2X1    g15548(.A(new_n15117_), .B(new_n15142_), .Y(new_n15741_));
  OAI21X1  g15549(.A0(new_n15741_), .A1(new_n15362_), .B0(new_n15143_), .Y(new_n15742_));
  AND2X1   g15550(.A(new_n15742_), .B(new_n15740_), .Y(new_n15743_));
  INVX1    g15551(.A(new_n15743_), .Y(new_n15744_));
  AND2X1   g15552(.A(new_n15719_), .B(\asqrt[41] ), .Y(new_n15745_));
  NAND2X1  g15553(.A(new_n15692_), .B(new_n15691_), .Y(new_n15746_));
  AND2X1   g15554(.A(new_n15710_), .B(new_n3564_), .Y(new_n15747_));
  AOI21X1  g15555(.A0(new_n15747_), .A1(new_n15746_), .B0(new_n15700_), .Y(new_n15748_));
  OAI21X1  g15556(.A0(new_n15748_), .A1(new_n15745_), .B0(\asqrt[42] ), .Y(new_n15749_));
  INVX1    g15557(.A(new_n15717_), .Y(new_n15750_));
  OAI21X1  g15558(.A0(new_n15693_), .A1(new_n3564_), .B0(new_n3276_), .Y(new_n15751_));
  OAI21X1  g15559(.A0(new_n15751_), .A1(new_n15748_), .B0(new_n15750_), .Y(new_n15752_));
  AOI21X1  g15560(.A0(new_n15752_), .A1(new_n15749_), .B0(new_n3008_), .Y(new_n15753_));
  INVX1    g15561(.A(new_n15727_), .Y(new_n15754_));
  NAND3X1  g15562(.A(new_n15752_), .B(new_n15749_), .C(new_n3008_), .Y(new_n15755_));
  AOI21X1  g15563(.A0(new_n15755_), .A1(new_n15754_), .B0(new_n15753_), .Y(new_n15756_));
  OAI21X1  g15564(.A0(new_n15756_), .A1(new_n2769_), .B0(new_n2570_), .Y(new_n15757_));
  OAI21X1  g15565(.A0(new_n15757_), .A1(new_n15738_), .B0(new_n15744_), .Y(new_n15758_));
  AOI21X1  g15566(.A0(new_n15758_), .A1(new_n15739_), .B0(new_n2263_), .Y(new_n15759_));
  AND2X1   g15567(.A(new_n15125_), .B(new_n15120_), .Y(new_n15760_));
  NOR3X1   g15568(.A(new_n15760_), .B(new_n15160_), .C(new_n15119_), .Y(new_n15761_));
  NOR3X1   g15569(.A(new_n15362_), .B(new_n15760_), .C(new_n15119_), .Y(new_n15762_));
  NOR2X1   g15570(.A(new_n15762_), .B(new_n15124_), .Y(new_n15763_));
  AOI21X1  g15571(.A0(new_n15761_), .A1(\asqrt[15] ), .B0(new_n15763_), .Y(new_n15764_));
  INVX1    g15572(.A(new_n15764_), .Y(new_n15765_));
  NAND3X1  g15573(.A(new_n15758_), .B(new_n15739_), .C(new_n2263_), .Y(new_n15766_));
  AOI21X1  g15574(.A0(new_n15766_), .A1(new_n15765_), .B0(new_n15759_), .Y(new_n15767_));
  OR2X1    g15575(.A(new_n15767_), .B(new_n2040_), .Y(new_n15768_));
  AND2X1   g15576(.A(new_n15766_), .B(new_n15765_), .Y(new_n15769_));
  AND2X1   g15577(.A(new_n15164_), .B(new_n15162_), .Y(new_n15770_));
  NOR3X1   g15578(.A(new_n15770_), .B(new_n15133_), .C(new_n15163_), .Y(new_n15771_));
  NOR3X1   g15579(.A(new_n15362_), .B(new_n15770_), .C(new_n15163_), .Y(new_n15772_));
  NOR2X1   g15580(.A(new_n15772_), .B(new_n15132_), .Y(new_n15773_));
  AOI21X1  g15581(.A0(new_n15771_), .A1(\asqrt[15] ), .B0(new_n15773_), .Y(new_n15774_));
  INVX1    g15582(.A(new_n15774_), .Y(new_n15775_));
  OR2X1    g15583(.A(new_n15756_), .B(new_n2769_), .Y(new_n15776_));
  NOR2X1   g15584(.A(new_n15728_), .B(new_n15727_), .Y(new_n15777_));
  INVX1    g15585(.A(new_n15736_), .Y(new_n15778_));
  NAND2X1  g15586(.A(new_n15722_), .B(new_n2769_), .Y(new_n15779_));
  OAI21X1  g15587(.A0(new_n15779_), .A1(new_n15777_), .B0(new_n15778_), .Y(new_n15780_));
  AOI21X1  g15588(.A0(new_n15780_), .A1(new_n15776_), .B0(new_n2570_), .Y(new_n15781_));
  AOI21X1  g15589(.A0(new_n15729_), .A1(\asqrt[44] ), .B0(\asqrt[45] ), .Y(new_n15782_));
  AOI21X1  g15590(.A0(new_n15782_), .A1(new_n15780_), .B0(new_n15743_), .Y(new_n15783_));
  OAI21X1  g15591(.A0(new_n15783_), .A1(new_n15781_), .B0(\asqrt[46] ), .Y(new_n15784_));
  NAND2X1  g15592(.A(new_n15784_), .B(new_n2040_), .Y(new_n15785_));
  OAI21X1  g15593(.A0(new_n15785_), .A1(new_n15769_), .B0(new_n15775_), .Y(new_n15786_));
  AOI21X1  g15594(.A0(new_n15786_), .A1(new_n15768_), .B0(new_n1834_), .Y(new_n15787_));
  NAND4X1  g15595(.A(\asqrt[15] ), .B(new_n15155_), .C(new_n15153_), .D(new_n15173_), .Y(new_n15788_));
  OR2X1    g15596(.A(new_n15166_), .B(new_n15148_), .Y(new_n15789_));
  OAI21X1  g15597(.A0(new_n15789_), .A1(new_n15362_), .B0(new_n15154_), .Y(new_n15790_));
  AND2X1   g15598(.A(new_n15790_), .B(new_n15788_), .Y(new_n15791_));
  NOR3X1   g15599(.A(new_n15783_), .B(new_n15781_), .C(\asqrt[46] ), .Y(new_n15792_));
  OAI21X1  g15600(.A0(new_n15792_), .A1(new_n15764_), .B0(new_n15784_), .Y(new_n15793_));
  AOI21X1  g15601(.A0(new_n15793_), .A1(\asqrt[47] ), .B0(\asqrt[48] ), .Y(new_n15794_));
  AOI21X1  g15602(.A0(new_n15794_), .A1(new_n15786_), .B0(new_n15791_), .Y(new_n15795_));
  OAI21X1  g15603(.A0(new_n15795_), .A1(new_n15787_), .B0(\asqrt[49] ), .Y(new_n15796_));
  AOI21X1  g15604(.A0(new_n15210_), .A1(new_n15209_), .B0(new_n15172_), .Y(new_n15797_));
  AND2X1   g15605(.A(new_n15797_), .B(new_n15157_), .Y(new_n15798_));
  AOI22X1  g15606(.A0(new_n15210_), .A1(new_n15209_), .B0(new_n15177_), .B1(\asqrt[48] ), .Y(new_n15799_));
  AOI21X1  g15607(.A0(new_n15799_), .A1(\asqrt[15] ), .B0(new_n15171_), .Y(new_n15800_));
  AOI21X1  g15608(.A0(new_n15798_), .A1(\asqrt[15] ), .B0(new_n15800_), .Y(new_n15801_));
  NOR3X1   g15609(.A(new_n15795_), .B(new_n15787_), .C(\asqrt[49] ), .Y(new_n15802_));
  OAI21X1  g15610(.A0(new_n15802_), .A1(new_n15801_), .B0(new_n15796_), .Y(new_n15803_));
  AND2X1   g15611(.A(new_n15803_), .B(\asqrt[50] ), .Y(new_n15804_));
  OR2X1    g15612(.A(new_n15802_), .B(new_n15801_), .Y(new_n15805_));
  AND2X1   g15613(.A(new_n15796_), .B(new_n1469_), .Y(new_n15806_));
  AND2X1   g15614(.A(new_n15178_), .B(new_n15175_), .Y(new_n15807_));
  NOR3X1   g15615(.A(new_n15214_), .B(new_n15807_), .C(new_n15176_), .Y(new_n15808_));
  NOR3X1   g15616(.A(new_n15362_), .B(new_n15807_), .C(new_n15176_), .Y(new_n15809_));
  NOR2X1   g15617(.A(new_n15809_), .B(new_n15183_), .Y(new_n15810_));
  AOI21X1  g15618(.A0(new_n15808_), .A1(\asqrt[15] ), .B0(new_n15810_), .Y(new_n15811_));
  AOI21X1  g15619(.A0(new_n15806_), .A1(new_n15805_), .B0(new_n15811_), .Y(new_n15812_));
  OAI21X1  g15620(.A0(new_n15812_), .A1(new_n15804_), .B0(\asqrt[51] ), .Y(new_n15813_));
  OR4X1    g15621(.A(new_n15362_), .B(new_n15191_), .C(new_n15217_), .D(new_n15216_), .Y(new_n15814_));
  OR2X1    g15622(.A(new_n15191_), .B(new_n15216_), .Y(new_n15815_));
  OAI21X1  g15623(.A0(new_n15815_), .A1(new_n15362_), .B0(new_n15217_), .Y(new_n15816_));
  AND2X1   g15624(.A(new_n15816_), .B(new_n15814_), .Y(new_n15817_));
  INVX1    g15625(.A(new_n15817_), .Y(new_n15818_));
  AND2X1   g15626(.A(new_n15793_), .B(\asqrt[47] ), .Y(new_n15819_));
  NAND2X1  g15627(.A(new_n15766_), .B(new_n15765_), .Y(new_n15820_));
  AND2X1   g15628(.A(new_n15784_), .B(new_n2040_), .Y(new_n15821_));
  AOI21X1  g15629(.A0(new_n15821_), .A1(new_n15820_), .B0(new_n15774_), .Y(new_n15822_));
  OAI21X1  g15630(.A0(new_n15822_), .A1(new_n15819_), .B0(\asqrt[48] ), .Y(new_n15823_));
  INVX1    g15631(.A(new_n15791_), .Y(new_n15824_));
  OAI21X1  g15632(.A0(new_n15767_), .A1(new_n2040_), .B0(new_n1834_), .Y(new_n15825_));
  OAI21X1  g15633(.A0(new_n15825_), .A1(new_n15822_), .B0(new_n15824_), .Y(new_n15826_));
  AOI21X1  g15634(.A0(new_n15826_), .A1(new_n15823_), .B0(new_n1632_), .Y(new_n15827_));
  INVX1    g15635(.A(new_n15801_), .Y(new_n15828_));
  NAND3X1  g15636(.A(new_n15826_), .B(new_n15823_), .C(new_n1632_), .Y(new_n15829_));
  AOI21X1  g15637(.A0(new_n15829_), .A1(new_n15828_), .B0(new_n15827_), .Y(new_n15830_));
  OAI21X1  g15638(.A0(new_n15830_), .A1(new_n1469_), .B0(new_n1277_), .Y(new_n15831_));
  OAI21X1  g15639(.A0(new_n15831_), .A1(new_n15812_), .B0(new_n15818_), .Y(new_n15832_));
  AOI21X1  g15640(.A0(new_n15832_), .A1(new_n15813_), .B0(new_n1111_), .Y(new_n15833_));
  AND2X1   g15641(.A(new_n15199_), .B(new_n15194_), .Y(new_n15834_));
  NOR3X1   g15642(.A(new_n15834_), .B(new_n15234_), .C(new_n15193_), .Y(new_n15835_));
  NOR3X1   g15643(.A(new_n15362_), .B(new_n15834_), .C(new_n15193_), .Y(new_n15836_));
  NOR2X1   g15644(.A(new_n15836_), .B(new_n15198_), .Y(new_n15837_));
  AOI21X1  g15645(.A0(new_n15835_), .A1(\asqrt[15] ), .B0(new_n15837_), .Y(new_n15838_));
  INVX1    g15646(.A(new_n15838_), .Y(new_n15839_));
  NAND3X1  g15647(.A(new_n15832_), .B(new_n15813_), .C(new_n1111_), .Y(new_n15840_));
  AOI21X1  g15648(.A0(new_n15840_), .A1(new_n15839_), .B0(new_n15833_), .Y(new_n15841_));
  OR2X1    g15649(.A(new_n15841_), .B(new_n968_), .Y(new_n15842_));
  OR2X1    g15650(.A(new_n15830_), .B(new_n1469_), .Y(new_n15843_));
  NOR2X1   g15651(.A(new_n15802_), .B(new_n15801_), .Y(new_n15844_));
  NAND2X1  g15652(.A(new_n15796_), .B(new_n1469_), .Y(new_n15845_));
  INVX1    g15653(.A(new_n15811_), .Y(new_n15846_));
  OAI21X1  g15654(.A0(new_n15845_), .A1(new_n15844_), .B0(new_n15846_), .Y(new_n15847_));
  AOI21X1  g15655(.A0(new_n15847_), .A1(new_n15843_), .B0(new_n1277_), .Y(new_n15848_));
  AOI21X1  g15656(.A0(new_n15803_), .A1(\asqrt[50] ), .B0(\asqrt[51] ), .Y(new_n15849_));
  AOI21X1  g15657(.A0(new_n15849_), .A1(new_n15847_), .B0(new_n15817_), .Y(new_n15850_));
  NOR3X1   g15658(.A(new_n15850_), .B(new_n15848_), .C(\asqrt[52] ), .Y(new_n15851_));
  NOR2X1   g15659(.A(new_n15851_), .B(new_n15838_), .Y(new_n15852_));
  AND2X1   g15660(.A(new_n15238_), .B(new_n15236_), .Y(new_n15853_));
  NOR3X1   g15661(.A(new_n15853_), .B(new_n15207_), .C(new_n15237_), .Y(new_n15854_));
  NOR3X1   g15662(.A(new_n15362_), .B(new_n15853_), .C(new_n15237_), .Y(new_n15855_));
  NOR2X1   g15663(.A(new_n15855_), .B(new_n15206_), .Y(new_n15856_));
  AOI21X1  g15664(.A0(new_n15854_), .A1(\asqrt[15] ), .B0(new_n15856_), .Y(new_n15857_));
  INVX1    g15665(.A(new_n15857_), .Y(new_n15858_));
  OAI21X1  g15666(.A0(new_n15850_), .A1(new_n15848_), .B0(\asqrt[52] ), .Y(new_n15859_));
  NAND2X1  g15667(.A(new_n15859_), .B(new_n968_), .Y(new_n15860_));
  OAI21X1  g15668(.A0(new_n15860_), .A1(new_n15852_), .B0(new_n15858_), .Y(new_n15861_));
  AOI21X1  g15669(.A0(new_n15861_), .A1(new_n15842_), .B0(new_n902_), .Y(new_n15862_));
  NAND4X1  g15670(.A(\asqrt[15] ), .B(new_n15229_), .C(new_n15227_), .D(new_n15247_), .Y(new_n15863_));
  OR2X1    g15671(.A(new_n15240_), .B(new_n15222_), .Y(new_n15864_));
  OAI21X1  g15672(.A0(new_n15864_), .A1(new_n15362_), .B0(new_n15228_), .Y(new_n15865_));
  AND2X1   g15673(.A(new_n15865_), .B(new_n15863_), .Y(new_n15866_));
  OAI21X1  g15674(.A0(new_n15851_), .A1(new_n15838_), .B0(new_n15859_), .Y(new_n15867_));
  AOI21X1  g15675(.A0(new_n15867_), .A1(\asqrt[53] ), .B0(\asqrt[54] ), .Y(new_n15868_));
  AOI21X1  g15676(.A0(new_n15868_), .A1(new_n15861_), .B0(new_n15866_), .Y(new_n15869_));
  OAI21X1  g15677(.A0(new_n15869_), .A1(new_n15862_), .B0(\asqrt[55] ), .Y(new_n15870_));
  AOI21X1  g15678(.A0(new_n15284_), .A1(new_n15283_), .B0(new_n15246_), .Y(new_n15871_));
  AND2X1   g15679(.A(new_n15871_), .B(new_n15231_), .Y(new_n15872_));
  AOI22X1  g15680(.A0(new_n15284_), .A1(new_n15283_), .B0(new_n15256_), .B1(\asqrt[54] ), .Y(new_n15873_));
  AOI21X1  g15681(.A0(new_n15873_), .A1(\asqrt[15] ), .B0(new_n15245_), .Y(new_n15874_));
  AOI21X1  g15682(.A0(new_n15872_), .A1(\asqrt[15] ), .B0(new_n15874_), .Y(new_n15875_));
  NOR3X1   g15683(.A(new_n15869_), .B(new_n15862_), .C(\asqrt[55] ), .Y(new_n15876_));
  OAI21X1  g15684(.A0(new_n15876_), .A1(new_n15875_), .B0(new_n15870_), .Y(new_n15877_));
  AND2X1   g15685(.A(new_n15877_), .B(\asqrt[56] ), .Y(new_n15878_));
  OR2X1    g15686(.A(new_n15876_), .B(new_n15875_), .Y(new_n15879_));
  AND2X1   g15687(.A(new_n15257_), .B(new_n15249_), .Y(new_n15880_));
  NOR3X1   g15688(.A(new_n15880_), .B(new_n15287_), .C(new_n15250_), .Y(new_n15881_));
  NOR3X1   g15689(.A(new_n15362_), .B(new_n15880_), .C(new_n15250_), .Y(new_n15882_));
  NOR2X1   g15690(.A(new_n15882_), .B(new_n15255_), .Y(new_n15883_));
  AOI21X1  g15691(.A0(new_n15881_), .A1(\asqrt[15] ), .B0(new_n15883_), .Y(new_n15884_));
  AND2X1   g15692(.A(new_n15870_), .B(new_n582_), .Y(new_n15885_));
  AOI21X1  g15693(.A0(new_n15885_), .A1(new_n15879_), .B0(new_n15884_), .Y(new_n15886_));
  OAI21X1  g15694(.A0(new_n15886_), .A1(new_n15878_), .B0(\asqrt[57] ), .Y(new_n15887_));
  OR4X1    g15695(.A(new_n15362_), .B(new_n15265_), .C(new_n15291_), .D(new_n15290_), .Y(new_n15888_));
  OR2X1    g15696(.A(new_n15265_), .B(new_n15290_), .Y(new_n15889_));
  OAI21X1  g15697(.A0(new_n15889_), .A1(new_n15362_), .B0(new_n15291_), .Y(new_n15890_));
  AND2X1   g15698(.A(new_n15890_), .B(new_n15888_), .Y(new_n15891_));
  INVX1    g15699(.A(new_n15891_), .Y(new_n15892_));
  AND2X1   g15700(.A(new_n15867_), .B(\asqrt[53] ), .Y(new_n15893_));
  OR2X1    g15701(.A(new_n15851_), .B(new_n15838_), .Y(new_n15894_));
  AND2X1   g15702(.A(new_n15859_), .B(new_n968_), .Y(new_n15895_));
  AOI21X1  g15703(.A0(new_n15895_), .A1(new_n15894_), .B0(new_n15857_), .Y(new_n15896_));
  OAI21X1  g15704(.A0(new_n15896_), .A1(new_n15893_), .B0(\asqrt[54] ), .Y(new_n15897_));
  INVX1    g15705(.A(new_n15866_), .Y(new_n15898_));
  OAI21X1  g15706(.A0(new_n15841_), .A1(new_n968_), .B0(new_n902_), .Y(new_n15899_));
  OAI21X1  g15707(.A0(new_n15899_), .A1(new_n15896_), .B0(new_n15898_), .Y(new_n15900_));
  AOI21X1  g15708(.A0(new_n15900_), .A1(new_n15897_), .B0(new_n697_), .Y(new_n15901_));
  INVX1    g15709(.A(new_n15875_), .Y(new_n15902_));
  NAND3X1  g15710(.A(new_n15900_), .B(new_n15897_), .C(new_n697_), .Y(new_n15903_));
  AOI21X1  g15711(.A0(new_n15903_), .A1(new_n15902_), .B0(new_n15901_), .Y(new_n15904_));
  OAI21X1  g15712(.A0(new_n15904_), .A1(new_n582_), .B0(new_n481_), .Y(new_n15905_));
  OAI21X1  g15713(.A0(new_n15905_), .A1(new_n15886_), .B0(new_n15892_), .Y(new_n15906_));
  AOI21X1  g15714(.A0(new_n15906_), .A1(new_n15887_), .B0(new_n399_), .Y(new_n15907_));
  AND2X1   g15715(.A(new_n15273_), .B(new_n15268_), .Y(new_n15908_));
  NOR3X1   g15716(.A(new_n15908_), .B(new_n15308_), .C(new_n15267_), .Y(new_n15909_));
  NOR3X1   g15717(.A(new_n15362_), .B(new_n15908_), .C(new_n15267_), .Y(new_n15910_));
  NOR2X1   g15718(.A(new_n15910_), .B(new_n15272_), .Y(new_n15911_));
  AOI21X1  g15719(.A0(new_n15909_), .A1(\asqrt[15] ), .B0(new_n15911_), .Y(new_n15912_));
  INVX1    g15720(.A(new_n15912_), .Y(new_n15913_));
  NAND3X1  g15721(.A(new_n15906_), .B(new_n15887_), .C(new_n399_), .Y(new_n15914_));
  AOI21X1  g15722(.A0(new_n15914_), .A1(new_n15913_), .B0(new_n15907_), .Y(new_n15915_));
  OR2X1    g15723(.A(new_n15915_), .B(new_n328_), .Y(new_n15916_));
  OR2X1    g15724(.A(new_n15904_), .B(new_n582_), .Y(new_n15917_));
  NOR2X1   g15725(.A(new_n15876_), .B(new_n15875_), .Y(new_n15918_));
  INVX1    g15726(.A(new_n15884_), .Y(new_n15919_));
  NAND2X1  g15727(.A(new_n15870_), .B(new_n582_), .Y(new_n15920_));
  OAI21X1  g15728(.A0(new_n15920_), .A1(new_n15918_), .B0(new_n15919_), .Y(new_n15921_));
  AOI21X1  g15729(.A0(new_n15921_), .A1(new_n15917_), .B0(new_n481_), .Y(new_n15922_));
  AOI21X1  g15730(.A0(new_n15877_), .A1(\asqrt[56] ), .B0(\asqrt[57] ), .Y(new_n15923_));
  AOI21X1  g15731(.A0(new_n15923_), .A1(new_n15921_), .B0(new_n15891_), .Y(new_n15924_));
  NOR3X1   g15732(.A(new_n15924_), .B(new_n15922_), .C(\asqrt[58] ), .Y(new_n15925_));
  NOR2X1   g15733(.A(new_n15925_), .B(new_n15912_), .Y(new_n15926_));
  AND2X1   g15734(.A(new_n15312_), .B(new_n15310_), .Y(new_n15927_));
  NOR3X1   g15735(.A(new_n15927_), .B(new_n15281_), .C(new_n15311_), .Y(new_n15928_));
  NOR3X1   g15736(.A(new_n15362_), .B(new_n15927_), .C(new_n15311_), .Y(new_n15929_));
  NOR2X1   g15737(.A(new_n15929_), .B(new_n15280_), .Y(new_n15930_));
  AOI21X1  g15738(.A0(new_n15928_), .A1(\asqrt[15] ), .B0(new_n15930_), .Y(new_n15931_));
  INVX1    g15739(.A(new_n15931_), .Y(new_n15932_));
  OAI21X1  g15740(.A0(new_n15924_), .A1(new_n15922_), .B0(\asqrt[58] ), .Y(new_n15933_));
  NAND2X1  g15741(.A(new_n15933_), .B(new_n328_), .Y(new_n15934_));
  OAI21X1  g15742(.A0(new_n15934_), .A1(new_n15926_), .B0(new_n15932_), .Y(new_n15935_));
  AOI21X1  g15743(.A0(new_n15935_), .A1(new_n15916_), .B0(new_n292_), .Y(new_n15936_));
  OR4X1    g15744(.A(new_n15362_), .B(new_n15314_), .C(new_n15302_), .D(new_n15296_), .Y(new_n15937_));
  OR2X1    g15745(.A(new_n15314_), .B(new_n15296_), .Y(new_n15938_));
  OAI21X1  g15746(.A0(new_n15938_), .A1(new_n15362_), .B0(new_n15302_), .Y(new_n15939_));
  AND2X1   g15747(.A(new_n15939_), .B(new_n15937_), .Y(new_n15940_));
  OAI21X1  g15748(.A0(new_n15925_), .A1(new_n15912_), .B0(new_n15933_), .Y(new_n15941_));
  AOI21X1  g15749(.A0(new_n15941_), .A1(\asqrt[59] ), .B0(\asqrt[60] ), .Y(new_n15942_));
  AOI21X1  g15750(.A0(new_n15942_), .A1(new_n15935_), .B0(new_n15940_), .Y(new_n15943_));
  OAI21X1  g15751(.A0(new_n15943_), .A1(new_n15936_), .B0(\asqrt[61] ), .Y(new_n15944_));
  AOI21X1  g15752(.A0(new_n15375_), .A1(new_n15374_), .B0(new_n15320_), .Y(new_n15945_));
  AND2X1   g15753(.A(new_n15945_), .B(new_n15305_), .Y(new_n15946_));
  AOI22X1  g15754(.A0(new_n15375_), .A1(new_n15374_), .B0(new_n15330_), .B1(\asqrt[60] ), .Y(new_n15947_));
  AOI21X1  g15755(.A0(new_n15947_), .A1(\asqrt[15] ), .B0(new_n15319_), .Y(new_n15948_));
  AOI21X1  g15756(.A0(new_n15946_), .A1(\asqrt[15] ), .B0(new_n15948_), .Y(new_n15949_));
  NOR3X1   g15757(.A(new_n15943_), .B(new_n15936_), .C(\asqrt[61] ), .Y(new_n15950_));
  OAI21X1  g15758(.A0(new_n15950_), .A1(new_n15949_), .B0(new_n15944_), .Y(new_n15951_));
  AND2X1   g15759(.A(new_n15951_), .B(\asqrt[62] ), .Y(new_n15952_));
  OR2X1    g15760(.A(new_n15950_), .B(new_n15949_), .Y(new_n15953_));
  AND2X1   g15761(.A(new_n15331_), .B(new_n15323_), .Y(new_n15954_));
  NOR3X1   g15762(.A(new_n15954_), .B(new_n15378_), .C(new_n15324_), .Y(new_n15955_));
  NOR3X1   g15763(.A(new_n15362_), .B(new_n15954_), .C(new_n15324_), .Y(new_n15956_));
  NOR2X1   g15764(.A(new_n15956_), .B(new_n15329_), .Y(new_n15957_));
  AOI21X1  g15765(.A0(new_n15955_), .A1(\asqrt[15] ), .B0(new_n15957_), .Y(new_n15958_));
  AND2X1   g15766(.A(new_n15944_), .B(new_n199_), .Y(new_n15959_));
  AOI21X1  g15767(.A0(new_n15959_), .A1(new_n15953_), .B0(new_n15958_), .Y(new_n15960_));
  NOR4X1   g15768(.A(new_n15362_), .B(new_n15339_), .C(new_n15382_), .D(new_n15381_), .Y(new_n15961_));
  NAND3X1  g15769(.A(\asqrt[15] ), .B(new_n15383_), .C(new_n15333_), .Y(new_n15962_));
  AOI21X1  g15770(.A0(new_n15962_), .A1(new_n15382_), .B0(new_n15961_), .Y(new_n15963_));
  INVX1    g15771(.A(new_n15963_), .Y(new_n15964_));
  NOR3X1   g15772(.A(new_n15362_), .B(new_n15344_), .C(new_n15384_), .Y(new_n15965_));
  AOI21X1  g15773(.A0(new_n15388_), .A1(new_n15387_), .B0(new_n15965_), .Y(new_n15966_));
  AND2X1   g15774(.A(new_n15966_), .B(new_n15964_), .Y(new_n15967_));
  OAI21X1  g15775(.A0(new_n15960_), .A1(new_n15952_), .B0(new_n15967_), .Y(new_n15968_));
  AND2X1   g15776(.A(new_n15941_), .B(\asqrt[59] ), .Y(new_n15969_));
  OR2X1    g15777(.A(new_n15925_), .B(new_n15912_), .Y(new_n15970_));
  AND2X1   g15778(.A(new_n15933_), .B(new_n328_), .Y(new_n15971_));
  AOI21X1  g15779(.A0(new_n15971_), .A1(new_n15970_), .B0(new_n15931_), .Y(new_n15972_));
  OAI21X1  g15780(.A0(new_n15972_), .A1(new_n15969_), .B0(\asqrt[60] ), .Y(new_n15973_));
  INVX1    g15781(.A(new_n15940_), .Y(new_n15974_));
  OAI21X1  g15782(.A0(new_n15915_), .A1(new_n328_), .B0(new_n292_), .Y(new_n15975_));
  OAI21X1  g15783(.A0(new_n15975_), .A1(new_n15972_), .B0(new_n15974_), .Y(new_n15976_));
  AOI21X1  g15784(.A0(new_n15976_), .A1(new_n15973_), .B0(new_n217_), .Y(new_n15977_));
  INVX1    g15785(.A(new_n15949_), .Y(new_n15978_));
  NAND3X1  g15786(.A(new_n15976_), .B(new_n15973_), .C(new_n217_), .Y(new_n15979_));
  AOI21X1  g15787(.A0(new_n15979_), .A1(new_n15978_), .B0(new_n15977_), .Y(new_n15980_));
  OAI21X1  g15788(.A0(new_n15980_), .A1(new_n199_), .B0(new_n15963_), .Y(new_n15981_));
  AOI21X1  g15789(.A0(new_n15390_), .A1(new_n15386_), .B0(new_n15344_), .Y(new_n15982_));
  AOI21X1  g15790(.A0(new_n15345_), .A1(new_n15340_), .B0(new_n193_), .Y(new_n15983_));
  OAI21X1  g15791(.A0(new_n15982_), .A1(new_n15340_), .B0(new_n15983_), .Y(new_n15984_));
  OR2X1    g15792(.A(new_n15351_), .B(new_n15350_), .Y(new_n15985_));
  NOR4X1   g15793(.A(new_n15358_), .B(new_n15398_), .C(new_n15343_), .D(new_n15341_), .Y(new_n15986_));
  NAND3X1  g15794(.A(new_n15986_), .B(new_n15985_), .C(new_n15386_), .Y(new_n15987_));
  AND2X1   g15795(.A(new_n15987_), .B(new_n15984_), .Y(new_n15988_));
  OAI21X1  g15796(.A0(new_n15981_), .A1(new_n15960_), .B0(new_n15988_), .Y(new_n15989_));
  AOI21X1  g15797(.A0(new_n15968_), .A1(new_n193_), .B0(new_n15989_), .Y(new_n15990_));
  OR2X1    g15798(.A(new_n15980_), .B(new_n199_), .Y(new_n15991_));
  NOR2X1   g15799(.A(new_n15950_), .B(new_n15949_), .Y(new_n15992_));
  INVX1    g15800(.A(new_n15958_), .Y(new_n15993_));
  NAND2X1  g15801(.A(new_n15944_), .B(new_n199_), .Y(new_n15994_));
  OAI21X1  g15802(.A0(new_n15994_), .A1(new_n15992_), .B0(new_n15993_), .Y(new_n15995_));
  INVX1    g15803(.A(new_n15967_), .Y(new_n15996_));
  AOI21X1  g15804(.A0(new_n15995_), .A1(new_n15991_), .B0(new_n15996_), .Y(new_n15997_));
  AOI21X1  g15805(.A0(new_n15951_), .A1(\asqrt[62] ), .B0(new_n15964_), .Y(new_n15998_));
  INVX1    g15806(.A(new_n15988_), .Y(new_n15999_));
  AOI21X1  g15807(.A0(new_n15998_), .A1(new_n15995_), .B0(new_n15999_), .Y(new_n16000_));
  OAI21X1  g15808(.A0(new_n15997_), .A1(\asqrt[63] ), .B0(new_n16000_), .Y(\asqrt[14] ));
  NOR2X1   g15809(.A(\a[27] ), .B(\a[26] ), .Y(new_n16002_));
  MX2X1    g15810(.A(new_n16002_), .B(\asqrt[14] ), .S0(\a[28] ), .Y(new_n16003_));
  AND2X1   g15811(.A(new_n16003_), .B(\asqrt[15] ), .Y(new_n16004_));
  NOR3X1   g15812(.A(\a[28] ), .B(\a[27] ), .C(\a[26] ), .Y(new_n16005_));
  NOR3X1   g15813(.A(new_n16005_), .B(new_n15358_), .C(new_n15398_), .Y(new_n16006_));
  NAND3X1  g15814(.A(new_n16006_), .B(new_n15985_), .C(new_n15386_), .Y(new_n16007_));
  AOI21X1  g15815(.A0(\asqrt[14] ), .A1(\a[28] ), .B0(new_n16007_), .Y(new_n16008_));
  INVX1    g15816(.A(\a[28] ), .Y(new_n16009_));
  INVX1    g15817(.A(\a[29] ), .Y(new_n16010_));
  AOI21X1  g15818(.A0(\asqrt[14] ), .A1(new_n16009_), .B0(new_n16010_), .Y(new_n16011_));
  NOR2X1   g15819(.A(\a[29] ), .B(\a[28] ), .Y(new_n16012_));
  AND2X1   g15820(.A(\asqrt[14] ), .B(new_n16012_), .Y(new_n16013_));
  NOR3X1   g15821(.A(new_n16013_), .B(new_n16011_), .C(new_n16008_), .Y(new_n16014_));
  OAI21X1  g15822(.A0(new_n16014_), .A1(new_n16004_), .B0(\asqrt[16] ), .Y(new_n16015_));
  INVX1    g15823(.A(new_n16002_), .Y(new_n16016_));
  MX2X1    g15824(.A(new_n16016_), .B(new_n15990_), .S0(\a[28] ), .Y(new_n16017_));
  OAI21X1  g15825(.A0(new_n16017_), .A1(new_n15362_), .B0(new_n14754_), .Y(new_n16018_));
  NAND3X1  g15826(.A(new_n15987_), .B(new_n15984_), .C(\asqrt[15] ), .Y(new_n16019_));
  INVX1    g15827(.A(new_n16019_), .Y(new_n16020_));
  OAI21X1  g15828(.A0(new_n15981_), .A1(new_n15960_), .B0(new_n16020_), .Y(new_n16021_));
  AOI21X1  g15829(.A0(new_n15968_), .A1(new_n193_), .B0(new_n16021_), .Y(new_n16022_));
  AOI21X1  g15830(.A0(\asqrt[14] ), .A1(new_n16012_), .B0(new_n16022_), .Y(new_n16023_));
  OR2X1    g15831(.A(new_n16022_), .B(\a[30] ), .Y(new_n16024_));
  OAI22X1  g15832(.A0(new_n16024_), .A1(new_n16013_), .B0(new_n16023_), .B1(new_n15370_), .Y(new_n16025_));
  OAI21X1  g15833(.A0(new_n16018_), .A1(new_n16014_), .B0(new_n16025_), .Y(new_n16026_));
  AOI21X1  g15834(.A0(new_n16026_), .A1(new_n16015_), .B0(new_n14165_), .Y(new_n16027_));
  NOR4X1   g15835(.A(new_n15990_), .B(new_n15392_), .C(new_n15416_), .D(new_n15366_), .Y(new_n16028_));
  AND2X1   g15836(.A(new_n15369_), .B(new_n15415_), .Y(new_n16029_));
  AOI21X1  g15837(.A0(new_n16029_), .A1(\asqrt[14] ), .B0(new_n15419_), .Y(new_n16030_));
  NOR2X1   g15838(.A(new_n16030_), .B(new_n16028_), .Y(new_n16031_));
  INVX1    g15839(.A(new_n16031_), .Y(new_n16032_));
  NAND3X1  g15840(.A(new_n16026_), .B(new_n16015_), .C(new_n14165_), .Y(new_n16033_));
  AOI21X1  g15841(.A0(new_n16033_), .A1(new_n16032_), .B0(new_n16027_), .Y(new_n16034_));
  OR2X1    g15842(.A(new_n16034_), .B(new_n13571_), .Y(new_n16035_));
  AND2X1   g15843(.A(new_n16033_), .B(new_n16032_), .Y(new_n16036_));
  AOI21X1  g15844(.A0(new_n15449_), .A1(new_n15448_), .B0(new_n15405_), .Y(new_n16037_));
  NAND3X1  g15845(.A(new_n16037_), .B(\asqrt[14] ), .C(new_n15394_), .Y(new_n16038_));
  OAI22X1  g15846(.A0(new_n15396_), .A1(new_n15395_), .B0(new_n15393_), .B1(new_n14165_), .Y(new_n16039_));
  OAI21X1  g15847(.A0(new_n16039_), .A1(new_n15990_), .B0(new_n15405_), .Y(new_n16040_));
  AND2X1   g15848(.A(new_n16040_), .B(new_n16038_), .Y(new_n16041_));
  INVX1    g15849(.A(new_n16041_), .Y(new_n16042_));
  OR2X1    g15850(.A(new_n16027_), .B(\asqrt[18] ), .Y(new_n16043_));
  OAI21X1  g15851(.A0(new_n16043_), .A1(new_n16036_), .B0(new_n16042_), .Y(new_n16044_));
  AOI21X1  g15852(.A0(new_n16044_), .A1(new_n16035_), .B0(new_n13000_), .Y(new_n16045_));
  OR2X1    g15853(.A(new_n15454_), .B(new_n15451_), .Y(new_n16046_));
  NAND4X1  g15854(.A(\asqrt[14] ), .B(new_n16046_), .C(new_n15413_), .D(new_n15452_), .Y(new_n16047_));
  NAND2X1  g15855(.A(new_n16046_), .B(new_n15452_), .Y(new_n16048_));
  OAI21X1  g15856(.A0(new_n16048_), .A1(new_n15990_), .B0(new_n15453_), .Y(new_n16049_));
  AND2X1   g15857(.A(new_n16049_), .B(new_n16047_), .Y(new_n16050_));
  OR2X1    g15858(.A(new_n16017_), .B(new_n15362_), .Y(new_n16051_));
  INVX1    g15859(.A(new_n16007_), .Y(new_n16052_));
  OAI21X1  g15860(.A0(new_n15990_), .A1(new_n16009_), .B0(new_n16052_), .Y(new_n16053_));
  OAI21X1  g15861(.A0(new_n15990_), .A1(\a[28] ), .B0(\a[29] ), .Y(new_n16054_));
  INVX1    g15862(.A(new_n16012_), .Y(new_n16055_));
  OR2X1    g15863(.A(new_n15990_), .B(new_n16055_), .Y(new_n16056_));
  NAND3X1  g15864(.A(new_n16056_), .B(new_n16054_), .C(new_n16053_), .Y(new_n16057_));
  AOI21X1  g15865(.A0(new_n16057_), .A1(new_n16051_), .B0(new_n14754_), .Y(new_n16058_));
  AOI21X1  g15866(.A0(new_n16003_), .A1(\asqrt[15] ), .B0(\asqrt[16] ), .Y(new_n16059_));
  OR2X1    g15867(.A(new_n16023_), .B(new_n15370_), .Y(new_n16060_));
  OR2X1    g15868(.A(new_n16024_), .B(new_n16013_), .Y(new_n16061_));
  AOI22X1  g15869(.A0(new_n16061_), .A1(new_n16060_), .B0(new_n16059_), .B1(new_n16057_), .Y(new_n16062_));
  OAI21X1  g15870(.A0(new_n16062_), .A1(new_n16058_), .B0(\asqrt[17] ), .Y(new_n16063_));
  NOR3X1   g15871(.A(new_n16062_), .B(new_n16058_), .C(\asqrt[17] ), .Y(new_n16064_));
  OAI21X1  g15872(.A0(new_n16064_), .A1(new_n16031_), .B0(new_n16063_), .Y(new_n16065_));
  AOI21X1  g15873(.A0(new_n16065_), .A1(\asqrt[18] ), .B0(\asqrt[19] ), .Y(new_n16066_));
  AOI21X1  g15874(.A0(new_n16066_), .A1(new_n16044_), .B0(new_n16050_), .Y(new_n16067_));
  OAI21X1  g15875(.A0(new_n16067_), .A1(new_n16045_), .B0(\asqrt[20] ), .Y(new_n16068_));
  OR4X1    g15876(.A(new_n15990_), .B(new_n15431_), .C(new_n15457_), .D(new_n15456_), .Y(new_n16069_));
  NAND2X1  g15877(.A(new_n15458_), .B(new_n15423_), .Y(new_n16070_));
  OAI21X1  g15878(.A0(new_n16070_), .A1(new_n15990_), .B0(new_n15457_), .Y(new_n16071_));
  AND2X1   g15879(.A(new_n16071_), .B(new_n16069_), .Y(new_n16072_));
  NOR3X1   g15880(.A(new_n16067_), .B(new_n16045_), .C(\asqrt[20] ), .Y(new_n16073_));
  OAI21X1  g15881(.A0(new_n16073_), .A1(new_n16072_), .B0(new_n16068_), .Y(new_n16074_));
  AND2X1   g15882(.A(new_n16074_), .B(\asqrt[21] ), .Y(new_n16075_));
  INVX1    g15883(.A(new_n16072_), .Y(new_n16076_));
  AND2X1   g15884(.A(new_n16065_), .B(\asqrt[18] ), .Y(new_n16077_));
  NAND2X1  g15885(.A(new_n16033_), .B(new_n16032_), .Y(new_n16078_));
  NOR2X1   g15886(.A(new_n16027_), .B(\asqrt[18] ), .Y(new_n16079_));
  AOI21X1  g15887(.A0(new_n16079_), .A1(new_n16078_), .B0(new_n16041_), .Y(new_n16080_));
  OAI21X1  g15888(.A0(new_n16080_), .A1(new_n16077_), .B0(\asqrt[19] ), .Y(new_n16081_));
  INVX1    g15889(.A(new_n16050_), .Y(new_n16082_));
  OAI21X1  g15890(.A0(new_n16034_), .A1(new_n13571_), .B0(new_n13000_), .Y(new_n16083_));
  OAI21X1  g15891(.A0(new_n16083_), .A1(new_n16080_), .B0(new_n16082_), .Y(new_n16084_));
  NAND3X1  g15892(.A(new_n16084_), .B(new_n16081_), .C(new_n12447_), .Y(new_n16085_));
  NAND2X1  g15893(.A(new_n16085_), .B(new_n16076_), .Y(new_n16086_));
  AND2X1   g15894(.A(new_n15441_), .B(new_n15434_), .Y(new_n16087_));
  NOR4X1   g15895(.A(new_n15990_), .B(new_n16087_), .C(new_n15481_), .D(new_n15433_), .Y(new_n16088_));
  AOI22X1  g15896(.A0(new_n15441_), .A1(new_n15434_), .B0(new_n15432_), .B1(\asqrt[20] ), .Y(new_n16089_));
  AOI21X1  g15897(.A0(new_n16089_), .A1(\asqrt[14] ), .B0(new_n15440_), .Y(new_n16090_));
  NOR2X1   g15898(.A(new_n16090_), .B(new_n16088_), .Y(new_n16091_));
  AOI21X1  g15899(.A0(new_n16084_), .A1(new_n16081_), .B0(new_n12447_), .Y(new_n16092_));
  NOR2X1   g15900(.A(new_n16092_), .B(\asqrt[21] ), .Y(new_n16093_));
  AOI21X1  g15901(.A0(new_n16093_), .A1(new_n16086_), .B0(new_n16091_), .Y(new_n16094_));
  OAI21X1  g15902(.A0(new_n16094_), .A1(new_n16075_), .B0(\asqrt[22] ), .Y(new_n16095_));
  AND2X1   g15903(.A(new_n15486_), .B(new_n15483_), .Y(new_n16096_));
  OR4X1    g15904(.A(new_n15990_), .B(new_n16096_), .C(new_n15446_), .D(new_n15484_), .Y(new_n16097_));
  OR2X1    g15905(.A(new_n16096_), .B(new_n15484_), .Y(new_n16098_));
  OAI21X1  g15906(.A0(new_n16098_), .A1(new_n15990_), .B0(new_n15446_), .Y(new_n16099_));
  AND2X1   g15907(.A(new_n16099_), .B(new_n16097_), .Y(new_n16100_));
  INVX1    g15908(.A(new_n16100_), .Y(new_n16101_));
  AOI21X1  g15909(.A0(new_n16085_), .A1(new_n16076_), .B0(new_n16092_), .Y(new_n16102_));
  OAI21X1  g15910(.A0(new_n16102_), .A1(new_n11896_), .B0(new_n11362_), .Y(new_n16103_));
  OAI21X1  g15911(.A0(new_n16103_), .A1(new_n16094_), .B0(new_n16101_), .Y(new_n16104_));
  AOI21X1  g15912(.A0(new_n16104_), .A1(new_n16095_), .B0(new_n10849_), .Y(new_n16105_));
  OR4X1    g15913(.A(new_n15990_), .B(new_n15496_), .C(new_n15468_), .D(new_n15462_), .Y(new_n16106_));
  NAND2X1  g15914(.A(new_n15469_), .B(new_n15488_), .Y(new_n16107_));
  OAI21X1  g15915(.A0(new_n16107_), .A1(new_n15990_), .B0(new_n15468_), .Y(new_n16108_));
  AND2X1   g15916(.A(new_n16108_), .B(new_n16106_), .Y(new_n16109_));
  INVX1    g15917(.A(new_n16109_), .Y(new_n16110_));
  NAND3X1  g15918(.A(new_n16104_), .B(new_n16095_), .C(new_n10849_), .Y(new_n16111_));
  AOI21X1  g15919(.A0(new_n16111_), .A1(new_n16110_), .B0(new_n16105_), .Y(new_n16112_));
  OR2X1    g15920(.A(new_n16112_), .B(new_n10332_), .Y(new_n16113_));
  AND2X1   g15921(.A(new_n16111_), .B(new_n16110_), .Y(new_n16114_));
  OAI21X1  g15922(.A0(new_n15489_), .A1(new_n15472_), .B0(new_n15477_), .Y(new_n16115_));
  NOR3X1   g15923(.A(new_n16115_), .B(new_n15990_), .C(new_n15510_), .Y(new_n16116_));
  AOI22X1  g15924(.A0(new_n15512_), .A1(new_n15511_), .B0(new_n15497_), .B1(\asqrt[23] ), .Y(new_n16117_));
  AOI21X1  g15925(.A0(new_n16117_), .A1(\asqrt[14] ), .B0(new_n15477_), .Y(new_n16118_));
  NOR2X1   g15926(.A(new_n16118_), .B(new_n16116_), .Y(new_n16119_));
  INVX1    g15927(.A(new_n16119_), .Y(new_n16120_));
  OR2X1    g15928(.A(new_n16105_), .B(\asqrt[24] ), .Y(new_n16121_));
  OAI21X1  g15929(.A0(new_n16121_), .A1(new_n16114_), .B0(new_n16120_), .Y(new_n16122_));
  AOI21X1  g15930(.A0(new_n16122_), .A1(new_n16113_), .B0(new_n9833_), .Y(new_n16123_));
  AND2X1   g15931(.A(new_n15498_), .B(new_n15490_), .Y(new_n16124_));
  OR4X1    g15932(.A(new_n15990_), .B(new_n16124_), .C(new_n15515_), .D(new_n15491_), .Y(new_n16125_));
  OR2X1    g15933(.A(new_n16124_), .B(new_n15491_), .Y(new_n16126_));
  OAI21X1  g15934(.A0(new_n16126_), .A1(new_n15990_), .B0(new_n15515_), .Y(new_n16127_));
  AND2X1   g15935(.A(new_n16127_), .B(new_n16125_), .Y(new_n16128_));
  OR2X1    g15936(.A(new_n16102_), .B(new_n11896_), .Y(new_n16129_));
  AND2X1   g15937(.A(new_n16085_), .B(new_n16076_), .Y(new_n16130_));
  INVX1    g15938(.A(new_n16091_), .Y(new_n16131_));
  OR2X1    g15939(.A(new_n16092_), .B(\asqrt[21] ), .Y(new_n16132_));
  OAI21X1  g15940(.A0(new_n16132_), .A1(new_n16130_), .B0(new_n16131_), .Y(new_n16133_));
  AOI21X1  g15941(.A0(new_n16133_), .A1(new_n16129_), .B0(new_n11362_), .Y(new_n16134_));
  AOI21X1  g15942(.A0(new_n16074_), .A1(\asqrt[21] ), .B0(\asqrt[22] ), .Y(new_n16135_));
  AOI21X1  g15943(.A0(new_n16135_), .A1(new_n16133_), .B0(new_n16100_), .Y(new_n16136_));
  OAI21X1  g15944(.A0(new_n16136_), .A1(new_n16134_), .B0(\asqrt[23] ), .Y(new_n16137_));
  NOR3X1   g15945(.A(new_n16136_), .B(new_n16134_), .C(\asqrt[23] ), .Y(new_n16138_));
  OAI21X1  g15946(.A0(new_n16138_), .A1(new_n16109_), .B0(new_n16137_), .Y(new_n16139_));
  AOI21X1  g15947(.A0(new_n16139_), .A1(\asqrt[24] ), .B0(\asqrt[25] ), .Y(new_n16140_));
  AOI21X1  g15948(.A0(new_n16140_), .A1(new_n16122_), .B0(new_n16128_), .Y(new_n16141_));
  OAI21X1  g15949(.A0(new_n16141_), .A1(new_n16123_), .B0(\asqrt[26] ), .Y(new_n16142_));
  OR4X1    g15950(.A(new_n15990_), .B(new_n15506_), .C(new_n15509_), .D(new_n15533_), .Y(new_n16143_));
  NAND2X1  g15951(.A(new_n15518_), .B(new_n15500_), .Y(new_n16144_));
  OAI21X1  g15952(.A0(new_n16144_), .A1(new_n15990_), .B0(new_n15509_), .Y(new_n16145_));
  AND2X1   g15953(.A(new_n16145_), .B(new_n16143_), .Y(new_n16146_));
  NOR3X1   g15954(.A(new_n16141_), .B(new_n16123_), .C(\asqrt[26] ), .Y(new_n16147_));
  OAI21X1  g15955(.A0(new_n16147_), .A1(new_n16146_), .B0(new_n16142_), .Y(new_n16148_));
  AND2X1   g15956(.A(new_n16148_), .B(\asqrt[27] ), .Y(new_n16149_));
  INVX1    g15957(.A(new_n16146_), .Y(new_n16150_));
  AND2X1   g15958(.A(new_n16139_), .B(\asqrt[24] ), .Y(new_n16151_));
  NAND2X1  g15959(.A(new_n16111_), .B(new_n16110_), .Y(new_n16152_));
  NOR2X1   g15960(.A(new_n16105_), .B(\asqrt[24] ), .Y(new_n16153_));
  AOI21X1  g15961(.A0(new_n16153_), .A1(new_n16152_), .B0(new_n16119_), .Y(new_n16154_));
  OAI21X1  g15962(.A0(new_n16154_), .A1(new_n16151_), .B0(\asqrt[25] ), .Y(new_n16155_));
  INVX1    g15963(.A(new_n16128_), .Y(new_n16156_));
  OAI21X1  g15964(.A0(new_n16112_), .A1(new_n10332_), .B0(new_n9833_), .Y(new_n16157_));
  OAI21X1  g15965(.A0(new_n16157_), .A1(new_n16154_), .B0(new_n16156_), .Y(new_n16158_));
  NAND3X1  g15966(.A(new_n16158_), .B(new_n16155_), .C(new_n9353_), .Y(new_n16159_));
  NAND2X1  g15967(.A(new_n16159_), .B(new_n16150_), .Y(new_n16160_));
  AND2X1   g15968(.A(new_n15525_), .B(new_n15519_), .Y(new_n16161_));
  NOR4X1   g15969(.A(new_n15990_), .B(new_n16161_), .C(new_n15556_), .D(new_n15508_), .Y(new_n16162_));
  AOI22X1  g15970(.A0(new_n15525_), .A1(new_n15519_), .B0(new_n15507_), .B1(\asqrt[26] ), .Y(new_n16163_));
  AOI21X1  g15971(.A0(new_n16163_), .A1(\asqrt[14] ), .B0(new_n15524_), .Y(new_n16164_));
  NOR2X1   g15972(.A(new_n16164_), .B(new_n16162_), .Y(new_n16165_));
  AOI21X1  g15973(.A0(new_n16158_), .A1(new_n16155_), .B0(new_n9353_), .Y(new_n16166_));
  NOR2X1   g15974(.A(new_n16166_), .B(\asqrt[27] ), .Y(new_n16167_));
  AOI21X1  g15975(.A0(new_n16167_), .A1(new_n16160_), .B0(new_n16165_), .Y(new_n16168_));
  OAI21X1  g15976(.A0(new_n16168_), .A1(new_n16149_), .B0(\asqrt[28] ), .Y(new_n16169_));
  AND2X1   g15977(.A(new_n15560_), .B(new_n15558_), .Y(new_n16170_));
  OR4X1    g15978(.A(new_n15990_), .B(new_n16170_), .C(new_n15532_), .D(new_n15559_), .Y(new_n16171_));
  OR2X1    g15979(.A(new_n16170_), .B(new_n15559_), .Y(new_n16172_));
  OAI21X1  g15980(.A0(new_n16172_), .A1(new_n15990_), .B0(new_n15532_), .Y(new_n16173_));
  AND2X1   g15981(.A(new_n16173_), .B(new_n16171_), .Y(new_n16174_));
  INVX1    g15982(.A(new_n16174_), .Y(new_n16175_));
  AOI21X1  g15983(.A0(new_n16159_), .A1(new_n16150_), .B0(new_n16166_), .Y(new_n16176_));
  OAI21X1  g15984(.A0(new_n16176_), .A1(new_n8874_), .B0(new_n8412_), .Y(new_n16177_));
  OAI21X1  g15985(.A0(new_n16177_), .A1(new_n16168_), .B0(new_n16175_), .Y(new_n16178_));
  AOI21X1  g15986(.A0(new_n16178_), .A1(new_n16169_), .B0(new_n7970_), .Y(new_n16179_));
  OR4X1    g15987(.A(new_n15990_), .B(new_n15570_), .C(new_n15543_), .D(new_n15537_), .Y(new_n16180_));
  NAND2X1  g15988(.A(new_n15544_), .B(new_n15562_), .Y(new_n16181_));
  OAI21X1  g15989(.A0(new_n16181_), .A1(new_n15990_), .B0(new_n15543_), .Y(new_n16182_));
  AND2X1   g15990(.A(new_n16182_), .B(new_n16180_), .Y(new_n16183_));
  INVX1    g15991(.A(new_n16183_), .Y(new_n16184_));
  NAND3X1  g15992(.A(new_n16178_), .B(new_n16169_), .C(new_n7970_), .Y(new_n16185_));
  AOI21X1  g15993(.A0(new_n16185_), .A1(new_n16184_), .B0(new_n16179_), .Y(new_n16186_));
  OR2X1    g15994(.A(new_n16186_), .B(new_n7527_), .Y(new_n16187_));
  AND2X1   g15995(.A(new_n16185_), .B(new_n16184_), .Y(new_n16188_));
  AOI21X1  g15996(.A0(new_n15586_), .A1(new_n15585_), .B0(new_n15553_), .Y(new_n16189_));
  AND2X1   g15997(.A(new_n16189_), .B(new_n15546_), .Y(new_n16190_));
  AOI22X1  g15998(.A0(new_n15586_), .A1(new_n15585_), .B0(new_n15571_), .B1(\asqrt[29] ), .Y(new_n16191_));
  AOI21X1  g15999(.A0(new_n16191_), .A1(\asqrt[14] ), .B0(new_n15552_), .Y(new_n16192_));
  AOI21X1  g16000(.A0(new_n16190_), .A1(\asqrt[14] ), .B0(new_n16192_), .Y(new_n16193_));
  INVX1    g16001(.A(new_n16193_), .Y(new_n16194_));
  OR2X1    g16002(.A(new_n16179_), .B(\asqrt[30] ), .Y(new_n16195_));
  OAI21X1  g16003(.A0(new_n16195_), .A1(new_n16188_), .B0(new_n16194_), .Y(new_n16196_));
  AOI21X1  g16004(.A0(new_n16196_), .A1(new_n16187_), .B0(new_n7103_), .Y(new_n16197_));
  AND2X1   g16005(.A(new_n15572_), .B(new_n15564_), .Y(new_n16198_));
  OR4X1    g16006(.A(new_n15990_), .B(new_n16198_), .C(new_n15589_), .D(new_n15565_), .Y(new_n16199_));
  OR2X1    g16007(.A(new_n16198_), .B(new_n15565_), .Y(new_n16200_));
  OAI21X1  g16008(.A0(new_n16200_), .A1(new_n15990_), .B0(new_n15589_), .Y(new_n16201_));
  AND2X1   g16009(.A(new_n16201_), .B(new_n16199_), .Y(new_n16202_));
  OR2X1    g16010(.A(new_n16176_), .B(new_n8874_), .Y(new_n16203_));
  AND2X1   g16011(.A(new_n16159_), .B(new_n16150_), .Y(new_n16204_));
  INVX1    g16012(.A(new_n16165_), .Y(new_n16205_));
  OR2X1    g16013(.A(new_n16166_), .B(\asqrt[27] ), .Y(new_n16206_));
  OAI21X1  g16014(.A0(new_n16206_), .A1(new_n16204_), .B0(new_n16205_), .Y(new_n16207_));
  AOI21X1  g16015(.A0(new_n16207_), .A1(new_n16203_), .B0(new_n8412_), .Y(new_n16208_));
  AOI21X1  g16016(.A0(new_n16148_), .A1(\asqrt[27] ), .B0(\asqrt[28] ), .Y(new_n16209_));
  AOI21X1  g16017(.A0(new_n16209_), .A1(new_n16207_), .B0(new_n16174_), .Y(new_n16210_));
  OAI21X1  g16018(.A0(new_n16210_), .A1(new_n16208_), .B0(\asqrt[29] ), .Y(new_n16211_));
  NOR3X1   g16019(.A(new_n16210_), .B(new_n16208_), .C(\asqrt[29] ), .Y(new_n16212_));
  OAI21X1  g16020(.A0(new_n16212_), .A1(new_n16183_), .B0(new_n16211_), .Y(new_n16213_));
  AOI21X1  g16021(.A0(new_n16213_), .A1(\asqrt[30] ), .B0(\asqrt[31] ), .Y(new_n16214_));
  AOI21X1  g16022(.A0(new_n16214_), .A1(new_n16196_), .B0(new_n16202_), .Y(new_n16215_));
  OAI21X1  g16023(.A0(new_n16215_), .A1(new_n16197_), .B0(\asqrt[32] ), .Y(new_n16216_));
  OR4X1    g16024(.A(new_n15990_), .B(new_n15580_), .C(new_n15583_), .D(new_n15607_), .Y(new_n16217_));
  NAND2X1  g16025(.A(new_n15592_), .B(new_n15574_), .Y(new_n16218_));
  OAI21X1  g16026(.A0(new_n16218_), .A1(new_n15990_), .B0(new_n15583_), .Y(new_n16219_));
  AND2X1   g16027(.A(new_n16219_), .B(new_n16217_), .Y(new_n16220_));
  NOR3X1   g16028(.A(new_n16215_), .B(new_n16197_), .C(\asqrt[32] ), .Y(new_n16221_));
  OAI21X1  g16029(.A0(new_n16221_), .A1(new_n16220_), .B0(new_n16216_), .Y(new_n16222_));
  AND2X1   g16030(.A(new_n16222_), .B(\asqrt[33] ), .Y(new_n16223_));
  OR2X1    g16031(.A(new_n16221_), .B(new_n16220_), .Y(new_n16224_));
  AND2X1   g16032(.A(new_n15599_), .B(new_n15593_), .Y(new_n16225_));
  NOR4X1   g16033(.A(new_n15990_), .B(new_n16225_), .C(new_n15630_), .D(new_n15582_), .Y(new_n16226_));
  AOI22X1  g16034(.A0(new_n15599_), .A1(new_n15593_), .B0(new_n15581_), .B1(\asqrt[32] ), .Y(new_n16227_));
  AOI21X1  g16035(.A0(new_n16227_), .A1(\asqrt[14] ), .B0(new_n15598_), .Y(new_n16228_));
  NOR2X1   g16036(.A(new_n16228_), .B(new_n16226_), .Y(new_n16229_));
  AND2X1   g16037(.A(new_n16216_), .B(new_n6294_), .Y(new_n16230_));
  AOI21X1  g16038(.A0(new_n16230_), .A1(new_n16224_), .B0(new_n16229_), .Y(new_n16231_));
  OAI21X1  g16039(.A0(new_n16231_), .A1(new_n16223_), .B0(\asqrt[34] ), .Y(new_n16232_));
  AND2X1   g16040(.A(new_n15634_), .B(new_n15632_), .Y(new_n16233_));
  OR4X1    g16041(.A(new_n15990_), .B(new_n16233_), .C(new_n15606_), .D(new_n15633_), .Y(new_n16234_));
  OR2X1    g16042(.A(new_n16233_), .B(new_n15633_), .Y(new_n16235_));
  OAI21X1  g16043(.A0(new_n16235_), .A1(new_n15990_), .B0(new_n15606_), .Y(new_n16236_));
  AND2X1   g16044(.A(new_n16236_), .B(new_n16234_), .Y(new_n16237_));
  INVX1    g16045(.A(new_n16237_), .Y(new_n16238_));
  AND2X1   g16046(.A(new_n16213_), .B(\asqrt[30] ), .Y(new_n16239_));
  NAND2X1  g16047(.A(new_n16185_), .B(new_n16184_), .Y(new_n16240_));
  NOR2X1   g16048(.A(new_n16179_), .B(\asqrt[30] ), .Y(new_n16241_));
  AOI21X1  g16049(.A0(new_n16241_), .A1(new_n16240_), .B0(new_n16193_), .Y(new_n16242_));
  OAI21X1  g16050(.A0(new_n16242_), .A1(new_n16239_), .B0(\asqrt[31] ), .Y(new_n16243_));
  INVX1    g16051(.A(new_n16202_), .Y(new_n16244_));
  OAI21X1  g16052(.A0(new_n16186_), .A1(new_n7527_), .B0(new_n7103_), .Y(new_n16245_));
  OAI21X1  g16053(.A0(new_n16245_), .A1(new_n16242_), .B0(new_n16244_), .Y(new_n16246_));
  AOI21X1  g16054(.A0(new_n16246_), .A1(new_n16243_), .B0(new_n6699_), .Y(new_n16247_));
  INVX1    g16055(.A(new_n16220_), .Y(new_n16248_));
  NAND3X1  g16056(.A(new_n16246_), .B(new_n16243_), .C(new_n6699_), .Y(new_n16249_));
  AOI21X1  g16057(.A0(new_n16249_), .A1(new_n16248_), .B0(new_n16247_), .Y(new_n16250_));
  OAI21X1  g16058(.A0(new_n16250_), .A1(new_n6294_), .B0(new_n5941_), .Y(new_n16251_));
  OAI21X1  g16059(.A0(new_n16251_), .A1(new_n16231_), .B0(new_n16238_), .Y(new_n16252_));
  AOI21X1  g16060(.A0(new_n16252_), .A1(new_n16232_), .B0(new_n5541_), .Y(new_n16253_));
  OR4X1    g16061(.A(new_n15990_), .B(new_n15644_), .C(new_n15617_), .D(new_n15611_), .Y(new_n16254_));
  NAND2X1  g16062(.A(new_n15618_), .B(new_n15636_), .Y(new_n16255_));
  OAI21X1  g16063(.A0(new_n16255_), .A1(new_n15990_), .B0(new_n15617_), .Y(new_n16256_));
  AND2X1   g16064(.A(new_n16256_), .B(new_n16254_), .Y(new_n16257_));
  INVX1    g16065(.A(new_n16257_), .Y(new_n16258_));
  NAND3X1  g16066(.A(new_n16252_), .B(new_n16232_), .C(new_n5541_), .Y(new_n16259_));
  AOI21X1  g16067(.A0(new_n16259_), .A1(new_n16258_), .B0(new_n16253_), .Y(new_n16260_));
  OR2X1    g16068(.A(new_n16260_), .B(new_n5176_), .Y(new_n16261_));
  OR2X1    g16069(.A(new_n16250_), .B(new_n6294_), .Y(new_n16262_));
  NOR2X1   g16070(.A(new_n16221_), .B(new_n16220_), .Y(new_n16263_));
  INVX1    g16071(.A(new_n16229_), .Y(new_n16264_));
  NAND2X1  g16072(.A(new_n16216_), .B(new_n6294_), .Y(new_n16265_));
  OAI21X1  g16073(.A0(new_n16265_), .A1(new_n16263_), .B0(new_n16264_), .Y(new_n16266_));
  AOI21X1  g16074(.A0(new_n16266_), .A1(new_n16262_), .B0(new_n5941_), .Y(new_n16267_));
  AOI21X1  g16075(.A0(new_n16222_), .A1(\asqrt[33] ), .B0(\asqrt[34] ), .Y(new_n16268_));
  AOI21X1  g16076(.A0(new_n16268_), .A1(new_n16266_), .B0(new_n16237_), .Y(new_n16269_));
  NOR3X1   g16077(.A(new_n16269_), .B(new_n16267_), .C(\asqrt[35] ), .Y(new_n16270_));
  NOR2X1   g16078(.A(new_n16270_), .B(new_n16257_), .Y(new_n16271_));
  OAI21X1  g16079(.A0(new_n15637_), .A1(new_n15621_), .B0(new_n15626_), .Y(new_n16272_));
  NOR3X1   g16080(.A(new_n16272_), .B(new_n15990_), .C(new_n15658_), .Y(new_n16273_));
  AOI22X1  g16081(.A0(new_n15660_), .A1(new_n15659_), .B0(new_n15645_), .B1(\asqrt[35] ), .Y(new_n16274_));
  AOI21X1  g16082(.A0(new_n16274_), .A1(\asqrt[14] ), .B0(new_n15626_), .Y(new_n16275_));
  NOR2X1   g16083(.A(new_n16275_), .B(new_n16273_), .Y(new_n16276_));
  INVX1    g16084(.A(new_n16276_), .Y(new_n16277_));
  OAI21X1  g16085(.A0(new_n16269_), .A1(new_n16267_), .B0(\asqrt[35] ), .Y(new_n16278_));
  NAND2X1  g16086(.A(new_n16278_), .B(new_n5176_), .Y(new_n16279_));
  OAI21X1  g16087(.A0(new_n16279_), .A1(new_n16271_), .B0(new_n16277_), .Y(new_n16280_));
  AOI21X1  g16088(.A0(new_n16280_), .A1(new_n16261_), .B0(new_n4826_), .Y(new_n16281_));
  AND2X1   g16089(.A(new_n15646_), .B(new_n15638_), .Y(new_n16282_));
  OR4X1    g16090(.A(new_n15990_), .B(new_n16282_), .C(new_n15663_), .D(new_n15639_), .Y(new_n16283_));
  OR2X1    g16091(.A(new_n16282_), .B(new_n15639_), .Y(new_n16284_));
  OAI21X1  g16092(.A0(new_n16284_), .A1(new_n15990_), .B0(new_n15663_), .Y(new_n16285_));
  AND2X1   g16093(.A(new_n16285_), .B(new_n16283_), .Y(new_n16286_));
  OAI21X1  g16094(.A0(new_n16270_), .A1(new_n16257_), .B0(new_n16278_), .Y(new_n16287_));
  AOI21X1  g16095(.A0(new_n16287_), .A1(\asqrt[36] ), .B0(\asqrt[37] ), .Y(new_n16288_));
  AOI21X1  g16096(.A0(new_n16288_), .A1(new_n16280_), .B0(new_n16286_), .Y(new_n16289_));
  OAI21X1  g16097(.A0(new_n16289_), .A1(new_n16281_), .B0(\asqrt[38] ), .Y(new_n16290_));
  OR4X1    g16098(.A(new_n15990_), .B(new_n15654_), .C(new_n15657_), .D(new_n15681_), .Y(new_n16291_));
  NAND2X1  g16099(.A(new_n15666_), .B(new_n15648_), .Y(new_n16292_));
  OAI21X1  g16100(.A0(new_n16292_), .A1(new_n15990_), .B0(new_n15657_), .Y(new_n16293_));
  AND2X1   g16101(.A(new_n16293_), .B(new_n16291_), .Y(new_n16294_));
  NOR3X1   g16102(.A(new_n16289_), .B(new_n16281_), .C(\asqrt[38] ), .Y(new_n16295_));
  OAI21X1  g16103(.A0(new_n16295_), .A1(new_n16294_), .B0(new_n16290_), .Y(new_n16296_));
  AND2X1   g16104(.A(new_n16296_), .B(\asqrt[39] ), .Y(new_n16297_));
  OR2X1    g16105(.A(new_n16295_), .B(new_n16294_), .Y(new_n16298_));
  AND2X1   g16106(.A(new_n15673_), .B(new_n15667_), .Y(new_n16299_));
  NOR4X1   g16107(.A(new_n15990_), .B(new_n16299_), .C(new_n15704_), .D(new_n15656_), .Y(new_n16300_));
  AOI22X1  g16108(.A0(new_n15673_), .A1(new_n15667_), .B0(new_n15655_), .B1(\asqrt[38] ), .Y(new_n16301_));
  AOI21X1  g16109(.A0(new_n16301_), .A1(\asqrt[14] ), .B0(new_n15672_), .Y(new_n16302_));
  NOR2X1   g16110(.A(new_n16302_), .B(new_n16300_), .Y(new_n16303_));
  AND2X1   g16111(.A(new_n16290_), .B(new_n4165_), .Y(new_n16304_));
  AOI21X1  g16112(.A0(new_n16304_), .A1(new_n16298_), .B0(new_n16303_), .Y(new_n16305_));
  OAI21X1  g16113(.A0(new_n16305_), .A1(new_n16297_), .B0(\asqrt[40] ), .Y(new_n16306_));
  AND2X1   g16114(.A(new_n15708_), .B(new_n15706_), .Y(new_n16307_));
  OR4X1    g16115(.A(new_n15990_), .B(new_n16307_), .C(new_n15680_), .D(new_n15707_), .Y(new_n16308_));
  OR2X1    g16116(.A(new_n16307_), .B(new_n15707_), .Y(new_n16309_));
  OAI21X1  g16117(.A0(new_n16309_), .A1(new_n15990_), .B0(new_n15680_), .Y(new_n16310_));
  AND2X1   g16118(.A(new_n16310_), .B(new_n16308_), .Y(new_n16311_));
  INVX1    g16119(.A(new_n16311_), .Y(new_n16312_));
  AND2X1   g16120(.A(new_n16287_), .B(\asqrt[36] ), .Y(new_n16313_));
  OR2X1    g16121(.A(new_n16270_), .B(new_n16257_), .Y(new_n16314_));
  AND2X1   g16122(.A(new_n16278_), .B(new_n5176_), .Y(new_n16315_));
  AOI21X1  g16123(.A0(new_n16315_), .A1(new_n16314_), .B0(new_n16276_), .Y(new_n16316_));
  OAI21X1  g16124(.A0(new_n16316_), .A1(new_n16313_), .B0(\asqrt[37] ), .Y(new_n16317_));
  INVX1    g16125(.A(new_n16286_), .Y(new_n16318_));
  OAI21X1  g16126(.A0(new_n16260_), .A1(new_n5176_), .B0(new_n4826_), .Y(new_n16319_));
  OAI21X1  g16127(.A0(new_n16319_), .A1(new_n16316_), .B0(new_n16318_), .Y(new_n16320_));
  AOI21X1  g16128(.A0(new_n16320_), .A1(new_n16317_), .B0(new_n4493_), .Y(new_n16321_));
  INVX1    g16129(.A(new_n16294_), .Y(new_n16322_));
  NAND3X1  g16130(.A(new_n16320_), .B(new_n16317_), .C(new_n4493_), .Y(new_n16323_));
  AOI21X1  g16131(.A0(new_n16323_), .A1(new_n16322_), .B0(new_n16321_), .Y(new_n16324_));
  OAI21X1  g16132(.A0(new_n16324_), .A1(new_n4165_), .B0(new_n3863_), .Y(new_n16325_));
  OAI21X1  g16133(.A0(new_n16325_), .A1(new_n16305_), .B0(new_n16312_), .Y(new_n16326_));
  AOI21X1  g16134(.A0(new_n16326_), .A1(new_n16306_), .B0(new_n3564_), .Y(new_n16327_));
  OR4X1    g16135(.A(new_n15990_), .B(new_n15718_), .C(new_n15691_), .D(new_n15685_), .Y(new_n16328_));
  NAND2X1  g16136(.A(new_n15692_), .B(new_n15710_), .Y(new_n16329_));
  OAI21X1  g16137(.A0(new_n16329_), .A1(new_n15990_), .B0(new_n15691_), .Y(new_n16330_));
  AND2X1   g16138(.A(new_n16330_), .B(new_n16328_), .Y(new_n16331_));
  INVX1    g16139(.A(new_n16331_), .Y(new_n16332_));
  NAND3X1  g16140(.A(new_n16326_), .B(new_n16306_), .C(new_n3564_), .Y(new_n16333_));
  AOI21X1  g16141(.A0(new_n16333_), .A1(new_n16332_), .B0(new_n16327_), .Y(new_n16334_));
  OR2X1    g16142(.A(new_n16334_), .B(new_n3276_), .Y(new_n16335_));
  OR2X1    g16143(.A(new_n16324_), .B(new_n4165_), .Y(new_n16336_));
  NOR2X1   g16144(.A(new_n16295_), .B(new_n16294_), .Y(new_n16337_));
  INVX1    g16145(.A(new_n16303_), .Y(new_n16338_));
  NAND2X1  g16146(.A(new_n16290_), .B(new_n4165_), .Y(new_n16339_));
  OAI21X1  g16147(.A0(new_n16339_), .A1(new_n16337_), .B0(new_n16338_), .Y(new_n16340_));
  AOI21X1  g16148(.A0(new_n16340_), .A1(new_n16336_), .B0(new_n3863_), .Y(new_n16341_));
  AOI21X1  g16149(.A0(new_n16296_), .A1(\asqrt[39] ), .B0(\asqrt[40] ), .Y(new_n16342_));
  AOI21X1  g16150(.A0(new_n16342_), .A1(new_n16340_), .B0(new_n16311_), .Y(new_n16343_));
  NOR3X1   g16151(.A(new_n16343_), .B(new_n16341_), .C(\asqrt[41] ), .Y(new_n16344_));
  NOR2X1   g16152(.A(new_n16344_), .B(new_n16331_), .Y(new_n16345_));
  OAI21X1  g16153(.A0(new_n15711_), .A1(new_n15695_), .B0(new_n15700_), .Y(new_n16346_));
  NOR3X1   g16154(.A(new_n16346_), .B(new_n15990_), .C(new_n15745_), .Y(new_n16347_));
  AOI22X1  g16155(.A0(new_n15747_), .A1(new_n15746_), .B0(new_n15719_), .B1(\asqrt[41] ), .Y(new_n16348_));
  AOI21X1  g16156(.A0(new_n16348_), .A1(\asqrt[14] ), .B0(new_n15700_), .Y(new_n16349_));
  NOR2X1   g16157(.A(new_n16349_), .B(new_n16347_), .Y(new_n16350_));
  INVX1    g16158(.A(new_n16350_), .Y(new_n16351_));
  OAI21X1  g16159(.A0(new_n16343_), .A1(new_n16341_), .B0(\asqrt[41] ), .Y(new_n16352_));
  NAND2X1  g16160(.A(new_n16352_), .B(new_n3276_), .Y(new_n16353_));
  OAI21X1  g16161(.A0(new_n16353_), .A1(new_n16345_), .B0(new_n16351_), .Y(new_n16354_));
  AOI21X1  g16162(.A0(new_n16354_), .A1(new_n16335_), .B0(new_n3008_), .Y(new_n16355_));
  AND2X1   g16163(.A(new_n15720_), .B(new_n15712_), .Y(new_n16356_));
  OR4X1    g16164(.A(new_n15990_), .B(new_n16356_), .C(new_n15750_), .D(new_n15713_), .Y(new_n16357_));
  OR2X1    g16165(.A(new_n16356_), .B(new_n15713_), .Y(new_n16358_));
  OAI21X1  g16166(.A0(new_n16358_), .A1(new_n15990_), .B0(new_n15750_), .Y(new_n16359_));
  AND2X1   g16167(.A(new_n16359_), .B(new_n16357_), .Y(new_n16360_));
  OAI21X1  g16168(.A0(new_n16344_), .A1(new_n16331_), .B0(new_n16352_), .Y(new_n16361_));
  AOI21X1  g16169(.A0(new_n16361_), .A1(\asqrt[42] ), .B0(\asqrt[43] ), .Y(new_n16362_));
  AOI21X1  g16170(.A0(new_n16362_), .A1(new_n16354_), .B0(new_n16360_), .Y(new_n16363_));
  OAI21X1  g16171(.A0(new_n16363_), .A1(new_n16355_), .B0(\asqrt[44] ), .Y(new_n16364_));
  OR4X1    g16172(.A(new_n15990_), .B(new_n15728_), .C(new_n15754_), .D(new_n15753_), .Y(new_n16365_));
  OR2X1    g16173(.A(new_n15728_), .B(new_n15753_), .Y(new_n16366_));
  OAI21X1  g16174(.A0(new_n16366_), .A1(new_n15990_), .B0(new_n15754_), .Y(new_n16367_));
  AND2X1   g16175(.A(new_n16367_), .B(new_n16365_), .Y(new_n16368_));
  NOR3X1   g16176(.A(new_n16363_), .B(new_n16355_), .C(\asqrt[44] ), .Y(new_n16369_));
  OAI21X1  g16177(.A0(new_n16369_), .A1(new_n16368_), .B0(new_n16364_), .Y(new_n16370_));
  AND2X1   g16178(.A(new_n16370_), .B(\asqrt[45] ), .Y(new_n16371_));
  OR2X1    g16179(.A(new_n16369_), .B(new_n16368_), .Y(new_n16372_));
  AND2X1   g16180(.A(new_n15737_), .B(new_n15731_), .Y(new_n16373_));
  NOR4X1   g16181(.A(new_n15990_), .B(new_n16373_), .C(new_n15778_), .D(new_n15730_), .Y(new_n16374_));
  AOI22X1  g16182(.A0(new_n15737_), .A1(new_n15731_), .B0(new_n15729_), .B1(\asqrt[44] ), .Y(new_n16375_));
  AOI21X1  g16183(.A0(new_n16375_), .A1(\asqrt[14] ), .B0(new_n15736_), .Y(new_n16376_));
  NOR2X1   g16184(.A(new_n16376_), .B(new_n16374_), .Y(new_n16377_));
  AND2X1   g16185(.A(new_n16364_), .B(new_n2570_), .Y(new_n16378_));
  AOI21X1  g16186(.A0(new_n16378_), .A1(new_n16372_), .B0(new_n16377_), .Y(new_n16379_));
  OAI21X1  g16187(.A0(new_n16379_), .A1(new_n16371_), .B0(\asqrt[46] ), .Y(new_n16380_));
  AND2X1   g16188(.A(new_n15782_), .B(new_n15780_), .Y(new_n16381_));
  OR4X1    g16189(.A(new_n15990_), .B(new_n16381_), .C(new_n15744_), .D(new_n15781_), .Y(new_n16382_));
  OR2X1    g16190(.A(new_n16381_), .B(new_n15781_), .Y(new_n16383_));
  OAI21X1  g16191(.A0(new_n16383_), .A1(new_n15990_), .B0(new_n15744_), .Y(new_n16384_));
  AND2X1   g16192(.A(new_n16384_), .B(new_n16382_), .Y(new_n16385_));
  INVX1    g16193(.A(new_n16385_), .Y(new_n16386_));
  AND2X1   g16194(.A(new_n16361_), .B(\asqrt[42] ), .Y(new_n16387_));
  OR2X1    g16195(.A(new_n16344_), .B(new_n16331_), .Y(new_n16388_));
  AND2X1   g16196(.A(new_n16352_), .B(new_n3276_), .Y(new_n16389_));
  AOI21X1  g16197(.A0(new_n16389_), .A1(new_n16388_), .B0(new_n16350_), .Y(new_n16390_));
  OAI21X1  g16198(.A0(new_n16390_), .A1(new_n16387_), .B0(\asqrt[43] ), .Y(new_n16391_));
  INVX1    g16199(.A(new_n16360_), .Y(new_n16392_));
  OAI21X1  g16200(.A0(new_n16334_), .A1(new_n3276_), .B0(new_n3008_), .Y(new_n16393_));
  OAI21X1  g16201(.A0(new_n16393_), .A1(new_n16390_), .B0(new_n16392_), .Y(new_n16394_));
  AOI21X1  g16202(.A0(new_n16394_), .A1(new_n16391_), .B0(new_n2769_), .Y(new_n16395_));
  INVX1    g16203(.A(new_n16368_), .Y(new_n16396_));
  NAND3X1  g16204(.A(new_n16394_), .B(new_n16391_), .C(new_n2769_), .Y(new_n16397_));
  AOI21X1  g16205(.A0(new_n16397_), .A1(new_n16396_), .B0(new_n16395_), .Y(new_n16398_));
  OAI21X1  g16206(.A0(new_n16398_), .A1(new_n2570_), .B0(new_n2263_), .Y(new_n16399_));
  OAI21X1  g16207(.A0(new_n16399_), .A1(new_n16379_), .B0(new_n16386_), .Y(new_n16400_));
  AOI21X1  g16208(.A0(new_n16400_), .A1(new_n16380_), .B0(new_n2040_), .Y(new_n16401_));
  OR4X1    g16209(.A(new_n15990_), .B(new_n15792_), .C(new_n15765_), .D(new_n15759_), .Y(new_n16402_));
  OR2X1    g16210(.A(new_n15792_), .B(new_n15759_), .Y(new_n16403_));
  OAI21X1  g16211(.A0(new_n16403_), .A1(new_n15990_), .B0(new_n15765_), .Y(new_n16404_));
  AND2X1   g16212(.A(new_n16404_), .B(new_n16402_), .Y(new_n16405_));
  INVX1    g16213(.A(new_n16405_), .Y(new_n16406_));
  NAND3X1  g16214(.A(new_n16400_), .B(new_n16380_), .C(new_n2040_), .Y(new_n16407_));
  AOI21X1  g16215(.A0(new_n16407_), .A1(new_n16406_), .B0(new_n16401_), .Y(new_n16408_));
  OR2X1    g16216(.A(new_n16408_), .B(new_n1834_), .Y(new_n16409_));
  OR2X1    g16217(.A(new_n16398_), .B(new_n2570_), .Y(new_n16410_));
  NOR2X1   g16218(.A(new_n16369_), .B(new_n16368_), .Y(new_n16411_));
  INVX1    g16219(.A(new_n16377_), .Y(new_n16412_));
  NAND2X1  g16220(.A(new_n16364_), .B(new_n2570_), .Y(new_n16413_));
  OAI21X1  g16221(.A0(new_n16413_), .A1(new_n16411_), .B0(new_n16412_), .Y(new_n16414_));
  AOI21X1  g16222(.A0(new_n16414_), .A1(new_n16410_), .B0(new_n2263_), .Y(new_n16415_));
  AOI21X1  g16223(.A0(new_n16370_), .A1(\asqrt[45] ), .B0(\asqrt[46] ), .Y(new_n16416_));
  AOI21X1  g16224(.A0(new_n16416_), .A1(new_n16414_), .B0(new_n16385_), .Y(new_n16417_));
  NOR3X1   g16225(.A(new_n16417_), .B(new_n16415_), .C(\asqrt[47] ), .Y(new_n16418_));
  NOR2X1   g16226(.A(new_n16418_), .B(new_n16405_), .Y(new_n16419_));
  AOI21X1  g16227(.A0(new_n15821_), .A1(new_n15820_), .B0(new_n15775_), .Y(new_n16420_));
  AND2X1   g16228(.A(new_n16420_), .B(new_n15768_), .Y(new_n16421_));
  AOI22X1  g16229(.A0(new_n15821_), .A1(new_n15820_), .B0(new_n15793_), .B1(\asqrt[47] ), .Y(new_n16422_));
  AOI21X1  g16230(.A0(new_n16422_), .A1(\asqrt[14] ), .B0(new_n15774_), .Y(new_n16423_));
  AOI21X1  g16231(.A0(new_n16421_), .A1(\asqrt[14] ), .B0(new_n16423_), .Y(new_n16424_));
  INVX1    g16232(.A(new_n16424_), .Y(new_n16425_));
  OAI21X1  g16233(.A0(new_n16417_), .A1(new_n16415_), .B0(\asqrt[47] ), .Y(new_n16426_));
  NAND2X1  g16234(.A(new_n16426_), .B(new_n1834_), .Y(new_n16427_));
  OAI21X1  g16235(.A0(new_n16427_), .A1(new_n16419_), .B0(new_n16425_), .Y(new_n16428_));
  AOI21X1  g16236(.A0(new_n16428_), .A1(new_n16409_), .B0(new_n1632_), .Y(new_n16429_));
  AND2X1   g16237(.A(new_n15794_), .B(new_n15786_), .Y(new_n16430_));
  OR4X1    g16238(.A(new_n15990_), .B(new_n16430_), .C(new_n15824_), .D(new_n15787_), .Y(new_n16431_));
  OR2X1    g16239(.A(new_n16430_), .B(new_n15787_), .Y(new_n16432_));
  OAI21X1  g16240(.A0(new_n16432_), .A1(new_n15990_), .B0(new_n15824_), .Y(new_n16433_));
  AND2X1   g16241(.A(new_n16433_), .B(new_n16431_), .Y(new_n16434_));
  OAI21X1  g16242(.A0(new_n16418_), .A1(new_n16405_), .B0(new_n16426_), .Y(new_n16435_));
  AOI21X1  g16243(.A0(new_n16435_), .A1(\asqrt[48] ), .B0(\asqrt[49] ), .Y(new_n16436_));
  AOI21X1  g16244(.A0(new_n16436_), .A1(new_n16428_), .B0(new_n16434_), .Y(new_n16437_));
  OAI21X1  g16245(.A0(new_n16437_), .A1(new_n16429_), .B0(\asqrt[50] ), .Y(new_n16438_));
  OR4X1    g16246(.A(new_n15990_), .B(new_n15802_), .C(new_n15828_), .D(new_n15827_), .Y(new_n16439_));
  OR2X1    g16247(.A(new_n15802_), .B(new_n15827_), .Y(new_n16440_));
  OAI21X1  g16248(.A0(new_n16440_), .A1(new_n15990_), .B0(new_n15828_), .Y(new_n16441_));
  AND2X1   g16249(.A(new_n16441_), .B(new_n16439_), .Y(new_n16442_));
  NOR3X1   g16250(.A(new_n16437_), .B(new_n16429_), .C(\asqrt[50] ), .Y(new_n16443_));
  OAI21X1  g16251(.A0(new_n16443_), .A1(new_n16442_), .B0(new_n16438_), .Y(new_n16444_));
  AND2X1   g16252(.A(new_n16444_), .B(\asqrt[51] ), .Y(new_n16445_));
  OR2X1    g16253(.A(new_n16443_), .B(new_n16442_), .Y(new_n16446_));
  AND2X1   g16254(.A(new_n16438_), .B(new_n1277_), .Y(new_n16447_));
  AND2X1   g16255(.A(new_n15806_), .B(new_n15805_), .Y(new_n16448_));
  NOR3X1   g16256(.A(new_n15846_), .B(new_n16448_), .C(new_n15804_), .Y(new_n16449_));
  AOI22X1  g16257(.A0(new_n15806_), .A1(new_n15805_), .B0(new_n15803_), .B1(\asqrt[50] ), .Y(new_n16450_));
  AOI21X1  g16258(.A0(new_n16450_), .A1(\asqrt[14] ), .B0(new_n15811_), .Y(new_n16451_));
  AOI21X1  g16259(.A0(new_n16449_), .A1(\asqrt[14] ), .B0(new_n16451_), .Y(new_n16452_));
  AOI21X1  g16260(.A0(new_n16447_), .A1(new_n16446_), .B0(new_n16452_), .Y(new_n16453_));
  OAI21X1  g16261(.A0(new_n16453_), .A1(new_n16445_), .B0(\asqrt[52] ), .Y(new_n16454_));
  AND2X1   g16262(.A(new_n15849_), .B(new_n15847_), .Y(new_n16455_));
  OR4X1    g16263(.A(new_n15990_), .B(new_n16455_), .C(new_n15818_), .D(new_n15848_), .Y(new_n16456_));
  OR2X1    g16264(.A(new_n16455_), .B(new_n15848_), .Y(new_n16457_));
  OAI21X1  g16265(.A0(new_n16457_), .A1(new_n15990_), .B0(new_n15818_), .Y(new_n16458_));
  AND2X1   g16266(.A(new_n16458_), .B(new_n16456_), .Y(new_n16459_));
  INVX1    g16267(.A(new_n16459_), .Y(new_n16460_));
  AND2X1   g16268(.A(new_n16435_), .B(\asqrt[48] ), .Y(new_n16461_));
  OR2X1    g16269(.A(new_n16418_), .B(new_n16405_), .Y(new_n16462_));
  AND2X1   g16270(.A(new_n16426_), .B(new_n1834_), .Y(new_n16463_));
  AOI21X1  g16271(.A0(new_n16463_), .A1(new_n16462_), .B0(new_n16424_), .Y(new_n16464_));
  OAI21X1  g16272(.A0(new_n16464_), .A1(new_n16461_), .B0(\asqrt[49] ), .Y(new_n16465_));
  INVX1    g16273(.A(new_n16434_), .Y(new_n16466_));
  OAI21X1  g16274(.A0(new_n16408_), .A1(new_n1834_), .B0(new_n1632_), .Y(new_n16467_));
  OAI21X1  g16275(.A0(new_n16467_), .A1(new_n16464_), .B0(new_n16466_), .Y(new_n16468_));
  AOI21X1  g16276(.A0(new_n16468_), .A1(new_n16465_), .B0(new_n1469_), .Y(new_n16469_));
  INVX1    g16277(.A(new_n16442_), .Y(new_n16470_));
  NAND3X1  g16278(.A(new_n16468_), .B(new_n16465_), .C(new_n1469_), .Y(new_n16471_));
  AOI21X1  g16279(.A0(new_n16471_), .A1(new_n16470_), .B0(new_n16469_), .Y(new_n16472_));
  OAI21X1  g16280(.A0(new_n16472_), .A1(new_n1277_), .B0(new_n1111_), .Y(new_n16473_));
  OAI21X1  g16281(.A0(new_n16473_), .A1(new_n16453_), .B0(new_n16460_), .Y(new_n16474_));
  AOI21X1  g16282(.A0(new_n16474_), .A1(new_n16454_), .B0(new_n968_), .Y(new_n16475_));
  OR4X1    g16283(.A(new_n15990_), .B(new_n15851_), .C(new_n15839_), .D(new_n15833_), .Y(new_n16476_));
  OR2X1    g16284(.A(new_n15851_), .B(new_n15833_), .Y(new_n16477_));
  OAI21X1  g16285(.A0(new_n16477_), .A1(new_n15990_), .B0(new_n15839_), .Y(new_n16478_));
  AND2X1   g16286(.A(new_n16478_), .B(new_n16476_), .Y(new_n16479_));
  INVX1    g16287(.A(new_n16479_), .Y(new_n16480_));
  NAND3X1  g16288(.A(new_n16474_), .B(new_n16454_), .C(new_n968_), .Y(new_n16481_));
  AOI21X1  g16289(.A0(new_n16481_), .A1(new_n16480_), .B0(new_n16475_), .Y(new_n16482_));
  OR2X1    g16290(.A(new_n16482_), .B(new_n902_), .Y(new_n16483_));
  OR2X1    g16291(.A(new_n16472_), .B(new_n1277_), .Y(new_n16484_));
  NOR2X1   g16292(.A(new_n16443_), .B(new_n16442_), .Y(new_n16485_));
  NAND2X1  g16293(.A(new_n16438_), .B(new_n1277_), .Y(new_n16486_));
  INVX1    g16294(.A(new_n16452_), .Y(new_n16487_));
  OAI21X1  g16295(.A0(new_n16486_), .A1(new_n16485_), .B0(new_n16487_), .Y(new_n16488_));
  AOI21X1  g16296(.A0(new_n16488_), .A1(new_n16484_), .B0(new_n1111_), .Y(new_n16489_));
  AOI21X1  g16297(.A0(new_n16444_), .A1(\asqrt[51] ), .B0(\asqrt[52] ), .Y(new_n16490_));
  AOI21X1  g16298(.A0(new_n16490_), .A1(new_n16488_), .B0(new_n16459_), .Y(new_n16491_));
  NOR3X1   g16299(.A(new_n16491_), .B(new_n16489_), .C(\asqrt[53] ), .Y(new_n16492_));
  NOR2X1   g16300(.A(new_n16492_), .B(new_n16479_), .Y(new_n16493_));
  OAI21X1  g16301(.A0(new_n15860_), .A1(new_n15852_), .B0(new_n15857_), .Y(new_n16494_));
  NOR3X1   g16302(.A(new_n16494_), .B(new_n15990_), .C(new_n15893_), .Y(new_n16495_));
  AOI22X1  g16303(.A0(new_n15895_), .A1(new_n15894_), .B0(new_n15867_), .B1(\asqrt[53] ), .Y(new_n16496_));
  AOI21X1  g16304(.A0(new_n16496_), .A1(\asqrt[14] ), .B0(new_n15857_), .Y(new_n16497_));
  NOR2X1   g16305(.A(new_n16497_), .B(new_n16495_), .Y(new_n16498_));
  INVX1    g16306(.A(new_n16498_), .Y(new_n16499_));
  OAI21X1  g16307(.A0(new_n16491_), .A1(new_n16489_), .B0(\asqrt[53] ), .Y(new_n16500_));
  NAND2X1  g16308(.A(new_n16500_), .B(new_n902_), .Y(new_n16501_));
  OAI21X1  g16309(.A0(new_n16501_), .A1(new_n16493_), .B0(new_n16499_), .Y(new_n16502_));
  AOI21X1  g16310(.A0(new_n16502_), .A1(new_n16483_), .B0(new_n697_), .Y(new_n16503_));
  AND2X1   g16311(.A(new_n15868_), .B(new_n15861_), .Y(new_n16504_));
  OR4X1    g16312(.A(new_n15990_), .B(new_n16504_), .C(new_n15898_), .D(new_n15862_), .Y(new_n16505_));
  OR2X1    g16313(.A(new_n16504_), .B(new_n15862_), .Y(new_n16506_));
  OAI21X1  g16314(.A0(new_n16506_), .A1(new_n15990_), .B0(new_n15898_), .Y(new_n16507_));
  AND2X1   g16315(.A(new_n16507_), .B(new_n16505_), .Y(new_n16508_));
  OAI21X1  g16316(.A0(new_n16492_), .A1(new_n16479_), .B0(new_n16500_), .Y(new_n16509_));
  AOI21X1  g16317(.A0(new_n16509_), .A1(\asqrt[54] ), .B0(\asqrt[55] ), .Y(new_n16510_));
  AOI21X1  g16318(.A0(new_n16510_), .A1(new_n16502_), .B0(new_n16508_), .Y(new_n16511_));
  OAI21X1  g16319(.A0(new_n16511_), .A1(new_n16503_), .B0(\asqrt[56] ), .Y(new_n16512_));
  NAND3X1  g16320(.A(new_n15903_), .B(new_n15875_), .C(new_n15870_), .Y(new_n16513_));
  NOR3X1   g16321(.A(new_n15990_), .B(new_n15876_), .C(new_n15901_), .Y(new_n16514_));
  OAI22X1  g16322(.A0(new_n16514_), .A1(new_n15875_), .B0(new_n16513_), .B1(new_n15990_), .Y(new_n16515_));
  INVX1    g16323(.A(new_n16515_), .Y(new_n16516_));
  NOR3X1   g16324(.A(new_n16511_), .B(new_n16503_), .C(\asqrt[56] ), .Y(new_n16517_));
  OAI21X1  g16325(.A0(new_n16517_), .A1(new_n16516_), .B0(new_n16512_), .Y(new_n16518_));
  AND2X1   g16326(.A(new_n16518_), .B(\asqrt[57] ), .Y(new_n16519_));
  OR2X1    g16327(.A(new_n16517_), .B(new_n16516_), .Y(new_n16520_));
  AND2X1   g16328(.A(new_n15885_), .B(new_n15879_), .Y(new_n16521_));
  NOR4X1   g16329(.A(new_n15990_), .B(new_n16521_), .C(new_n15919_), .D(new_n15878_), .Y(new_n16522_));
  AOI22X1  g16330(.A0(new_n15885_), .A1(new_n15879_), .B0(new_n15877_), .B1(\asqrt[56] ), .Y(new_n16523_));
  AOI21X1  g16331(.A0(new_n16523_), .A1(\asqrt[14] ), .B0(new_n15884_), .Y(new_n16524_));
  NOR2X1   g16332(.A(new_n16524_), .B(new_n16522_), .Y(new_n16525_));
  AND2X1   g16333(.A(new_n16512_), .B(new_n481_), .Y(new_n16526_));
  AOI21X1  g16334(.A0(new_n16526_), .A1(new_n16520_), .B0(new_n16525_), .Y(new_n16527_));
  OAI21X1  g16335(.A0(new_n16527_), .A1(new_n16519_), .B0(\asqrt[58] ), .Y(new_n16528_));
  AND2X1   g16336(.A(new_n15923_), .B(new_n15921_), .Y(new_n16529_));
  NOR3X1   g16337(.A(new_n16529_), .B(new_n15892_), .C(new_n15922_), .Y(new_n16530_));
  NOR2X1   g16338(.A(new_n16529_), .B(new_n15922_), .Y(new_n16531_));
  AOI21X1  g16339(.A0(new_n16531_), .A1(\asqrt[14] ), .B0(new_n15891_), .Y(new_n16532_));
  AOI21X1  g16340(.A0(new_n16530_), .A1(\asqrt[14] ), .B0(new_n16532_), .Y(new_n16533_));
  INVX1    g16341(.A(new_n16533_), .Y(new_n16534_));
  AND2X1   g16342(.A(new_n16509_), .B(\asqrt[54] ), .Y(new_n16535_));
  OR2X1    g16343(.A(new_n16492_), .B(new_n16479_), .Y(new_n16536_));
  AND2X1   g16344(.A(new_n16500_), .B(new_n902_), .Y(new_n16537_));
  AOI21X1  g16345(.A0(new_n16537_), .A1(new_n16536_), .B0(new_n16498_), .Y(new_n16538_));
  OAI21X1  g16346(.A0(new_n16538_), .A1(new_n16535_), .B0(\asqrt[55] ), .Y(new_n16539_));
  INVX1    g16347(.A(new_n16508_), .Y(new_n16540_));
  OAI21X1  g16348(.A0(new_n16482_), .A1(new_n902_), .B0(new_n697_), .Y(new_n16541_));
  OAI21X1  g16349(.A0(new_n16541_), .A1(new_n16538_), .B0(new_n16540_), .Y(new_n16542_));
  AOI21X1  g16350(.A0(new_n16542_), .A1(new_n16539_), .B0(new_n582_), .Y(new_n16543_));
  NAND3X1  g16351(.A(new_n16542_), .B(new_n16539_), .C(new_n582_), .Y(new_n16544_));
  AOI21X1  g16352(.A0(new_n16544_), .A1(new_n16515_), .B0(new_n16543_), .Y(new_n16545_));
  OAI21X1  g16353(.A0(new_n16545_), .A1(new_n481_), .B0(new_n399_), .Y(new_n16546_));
  OAI21X1  g16354(.A0(new_n16546_), .A1(new_n16527_), .B0(new_n16534_), .Y(new_n16547_));
  AOI21X1  g16355(.A0(new_n16547_), .A1(new_n16528_), .B0(new_n328_), .Y(new_n16548_));
  OR4X1    g16356(.A(new_n15990_), .B(new_n15925_), .C(new_n15913_), .D(new_n15907_), .Y(new_n16549_));
  OR2X1    g16357(.A(new_n15925_), .B(new_n15907_), .Y(new_n16550_));
  OAI21X1  g16358(.A0(new_n16550_), .A1(new_n15990_), .B0(new_n15913_), .Y(new_n16551_));
  AND2X1   g16359(.A(new_n16551_), .B(new_n16549_), .Y(new_n16552_));
  INVX1    g16360(.A(new_n16552_), .Y(new_n16553_));
  NAND3X1  g16361(.A(new_n16547_), .B(new_n16528_), .C(new_n328_), .Y(new_n16554_));
  AOI21X1  g16362(.A0(new_n16554_), .A1(new_n16553_), .B0(new_n16548_), .Y(new_n16555_));
  OR2X1    g16363(.A(new_n16555_), .B(new_n292_), .Y(new_n16556_));
  AND2X1   g16364(.A(new_n16554_), .B(new_n16553_), .Y(new_n16557_));
  OAI21X1  g16365(.A0(new_n15934_), .A1(new_n15926_), .B0(new_n15931_), .Y(new_n16558_));
  NOR3X1   g16366(.A(new_n16558_), .B(new_n15990_), .C(new_n15969_), .Y(new_n16559_));
  AOI22X1  g16367(.A0(new_n15971_), .A1(new_n15970_), .B0(new_n15941_), .B1(\asqrt[59] ), .Y(new_n16560_));
  AOI21X1  g16368(.A0(new_n16560_), .A1(\asqrt[14] ), .B0(new_n15931_), .Y(new_n16561_));
  NOR2X1   g16369(.A(new_n16561_), .B(new_n16559_), .Y(new_n16562_));
  INVX1    g16370(.A(new_n16562_), .Y(new_n16563_));
  OR2X1    g16371(.A(new_n16548_), .B(\asqrt[60] ), .Y(new_n16564_));
  OAI21X1  g16372(.A0(new_n16564_), .A1(new_n16557_), .B0(new_n16563_), .Y(new_n16565_));
  AOI21X1  g16373(.A0(new_n16565_), .A1(new_n16556_), .B0(new_n217_), .Y(new_n16566_));
  AND2X1   g16374(.A(new_n15942_), .B(new_n15935_), .Y(new_n16567_));
  OR4X1    g16375(.A(new_n15990_), .B(new_n16567_), .C(new_n15974_), .D(new_n15936_), .Y(new_n16568_));
  OR2X1    g16376(.A(new_n16567_), .B(new_n15936_), .Y(new_n16569_));
  OAI21X1  g16377(.A0(new_n16569_), .A1(new_n15990_), .B0(new_n15974_), .Y(new_n16570_));
  AND2X1   g16378(.A(new_n16570_), .B(new_n16568_), .Y(new_n16571_));
  OR2X1    g16379(.A(new_n16545_), .B(new_n481_), .Y(new_n16572_));
  NOR2X1   g16380(.A(new_n16517_), .B(new_n16516_), .Y(new_n16573_));
  INVX1    g16381(.A(new_n16525_), .Y(new_n16574_));
  NAND2X1  g16382(.A(new_n16512_), .B(new_n481_), .Y(new_n16575_));
  OAI21X1  g16383(.A0(new_n16575_), .A1(new_n16573_), .B0(new_n16574_), .Y(new_n16576_));
  AOI21X1  g16384(.A0(new_n16576_), .A1(new_n16572_), .B0(new_n399_), .Y(new_n16577_));
  AOI21X1  g16385(.A0(new_n16518_), .A1(\asqrt[57] ), .B0(\asqrt[58] ), .Y(new_n16578_));
  AOI21X1  g16386(.A0(new_n16578_), .A1(new_n16576_), .B0(new_n16533_), .Y(new_n16579_));
  OAI21X1  g16387(.A0(new_n16579_), .A1(new_n16577_), .B0(\asqrt[59] ), .Y(new_n16580_));
  NOR3X1   g16388(.A(new_n16579_), .B(new_n16577_), .C(\asqrt[59] ), .Y(new_n16581_));
  OAI21X1  g16389(.A0(new_n16581_), .A1(new_n16552_), .B0(new_n16580_), .Y(new_n16582_));
  AOI21X1  g16390(.A0(new_n16582_), .A1(\asqrt[60] ), .B0(\asqrt[61] ), .Y(new_n16583_));
  AOI21X1  g16391(.A0(new_n16583_), .A1(new_n16565_), .B0(new_n16571_), .Y(new_n16584_));
  OAI21X1  g16392(.A0(new_n16584_), .A1(new_n16566_), .B0(\asqrt[62] ), .Y(new_n16585_));
  OR4X1    g16393(.A(new_n15990_), .B(new_n15950_), .C(new_n15978_), .D(new_n15977_), .Y(new_n16586_));
  OR2X1    g16394(.A(new_n15950_), .B(new_n15977_), .Y(new_n16587_));
  OAI21X1  g16395(.A0(new_n16587_), .A1(new_n15990_), .B0(new_n15978_), .Y(new_n16588_));
  AND2X1   g16396(.A(new_n16588_), .B(new_n16586_), .Y(new_n16589_));
  NOR3X1   g16397(.A(new_n16584_), .B(new_n16566_), .C(\asqrt[62] ), .Y(new_n16590_));
  OAI21X1  g16398(.A0(new_n16590_), .A1(new_n16589_), .B0(new_n16585_), .Y(new_n16591_));
  AND2X1   g16399(.A(new_n15959_), .B(new_n15953_), .Y(new_n16592_));
  NOR4X1   g16400(.A(new_n15990_), .B(new_n16592_), .C(new_n15993_), .D(new_n15952_), .Y(new_n16593_));
  INVX1    g16401(.A(new_n16593_), .Y(new_n16594_));
  OAI22X1  g16402(.A0(new_n15994_), .A1(new_n15992_), .B0(new_n15980_), .B1(new_n199_), .Y(new_n16595_));
  OAI21X1  g16403(.A0(new_n16595_), .A1(new_n15990_), .B0(new_n15993_), .Y(new_n16596_));
  AND2X1   g16404(.A(new_n16596_), .B(new_n16594_), .Y(new_n16597_));
  INVX1    g16405(.A(new_n16597_), .Y(new_n16598_));
  AND2X1   g16406(.A(new_n15998_), .B(new_n15995_), .Y(new_n16599_));
  AOI21X1  g16407(.A0(new_n15995_), .A1(new_n15991_), .B0(new_n15963_), .Y(new_n16600_));
  AOI21X1  g16408(.A0(new_n16600_), .A1(\asqrt[14] ), .B0(new_n16599_), .Y(new_n16601_));
  AND2X1   g16409(.A(new_n16601_), .B(new_n16598_), .Y(new_n16602_));
  AOI21X1  g16410(.A0(new_n16602_), .A1(new_n16591_), .B0(\asqrt[63] ), .Y(new_n16603_));
  NOR2X1   g16411(.A(new_n16590_), .B(new_n16589_), .Y(new_n16604_));
  NAND2X1  g16412(.A(new_n16597_), .B(new_n16585_), .Y(new_n16605_));
  NAND2X1  g16413(.A(new_n15995_), .B(new_n15991_), .Y(new_n16606_));
  AOI21X1  g16414(.A0(\asqrt[14] ), .A1(new_n15964_), .B0(new_n16606_), .Y(new_n16607_));
  NOR3X1   g16415(.A(new_n16607_), .B(new_n16600_), .C(new_n193_), .Y(new_n16608_));
  AND2X1   g16416(.A(new_n15968_), .B(new_n193_), .Y(new_n16609_));
  INVX1    g16417(.A(new_n15987_), .Y(new_n16610_));
  OR2X1    g16418(.A(new_n16610_), .B(new_n15961_), .Y(new_n16611_));
  AOI21X1  g16419(.A0(new_n15962_), .A1(new_n15382_), .B0(new_n16611_), .Y(new_n16612_));
  NAND2X1  g16420(.A(new_n16612_), .B(new_n15984_), .Y(new_n16613_));
  NOR3X1   g16421(.A(new_n16613_), .B(new_n16599_), .C(new_n16609_), .Y(new_n16614_));
  NOR2X1   g16422(.A(new_n16614_), .B(new_n16608_), .Y(new_n16615_));
  OAI21X1  g16423(.A0(new_n16605_), .A1(new_n16604_), .B0(new_n16615_), .Y(new_n16616_));
  NOR2X1   g16424(.A(new_n16616_), .B(new_n16603_), .Y(new_n16617_));
  INVX1    g16425(.A(new_n16617_), .Y(\asqrt[13] ));
  OAI21X1  g16426(.A0(new_n16616_), .A1(new_n16603_), .B0(\a[26] ), .Y(new_n16619_));
  INVX1    g16427(.A(\a[26] ), .Y(new_n16620_));
  NOR2X1   g16428(.A(\a[25] ), .B(\a[24] ), .Y(new_n16621_));
  NAND2X1  g16429(.A(new_n16621_), .B(new_n16620_), .Y(new_n16622_));
  AND2X1   g16430(.A(new_n16622_), .B(new_n16619_), .Y(new_n16623_));
  AND2X1   g16431(.A(new_n16582_), .B(\asqrt[60] ), .Y(new_n16624_));
  NAND2X1  g16432(.A(new_n16554_), .B(new_n16553_), .Y(new_n16625_));
  NOR2X1   g16433(.A(new_n16548_), .B(\asqrt[60] ), .Y(new_n16626_));
  AOI21X1  g16434(.A0(new_n16626_), .A1(new_n16625_), .B0(new_n16562_), .Y(new_n16627_));
  OAI21X1  g16435(.A0(new_n16627_), .A1(new_n16624_), .B0(\asqrt[61] ), .Y(new_n16628_));
  INVX1    g16436(.A(new_n16571_), .Y(new_n16629_));
  OAI21X1  g16437(.A0(new_n16555_), .A1(new_n292_), .B0(new_n217_), .Y(new_n16630_));
  OAI21X1  g16438(.A0(new_n16630_), .A1(new_n16627_), .B0(new_n16629_), .Y(new_n16631_));
  AOI21X1  g16439(.A0(new_n16631_), .A1(new_n16628_), .B0(new_n199_), .Y(new_n16632_));
  INVX1    g16440(.A(new_n16589_), .Y(new_n16633_));
  NAND3X1  g16441(.A(new_n16631_), .B(new_n16628_), .C(new_n199_), .Y(new_n16634_));
  AOI21X1  g16442(.A0(new_n16634_), .A1(new_n16633_), .B0(new_n16632_), .Y(new_n16635_));
  INVX1    g16443(.A(new_n16602_), .Y(new_n16636_));
  OAI21X1  g16444(.A0(new_n16636_), .A1(new_n16635_), .B0(new_n193_), .Y(new_n16637_));
  OR2X1    g16445(.A(new_n16590_), .B(new_n16589_), .Y(new_n16638_));
  AND2X1   g16446(.A(new_n16597_), .B(new_n16585_), .Y(new_n16639_));
  INVX1    g16447(.A(new_n16615_), .Y(new_n16640_));
  AOI21X1  g16448(.A0(new_n16639_), .A1(new_n16638_), .B0(new_n16640_), .Y(new_n16641_));
  AOI21X1  g16449(.A0(new_n16641_), .A1(new_n16637_), .B0(new_n16620_), .Y(new_n16642_));
  NAND3X1  g16450(.A(new_n16622_), .B(new_n15987_), .C(new_n15984_), .Y(new_n16643_));
  NOR4X1   g16451(.A(new_n16643_), .B(new_n16642_), .C(new_n16599_), .D(new_n16609_), .Y(new_n16644_));
  INVX1    g16452(.A(\a[27] ), .Y(new_n16645_));
  AOI21X1  g16453(.A0(new_n16641_), .A1(new_n16637_), .B0(\a[26] ), .Y(new_n16646_));
  OAI21X1  g16454(.A0(new_n16616_), .A1(new_n16603_), .B0(new_n16002_), .Y(new_n16647_));
  OAI21X1  g16455(.A0(new_n16646_), .A1(new_n16645_), .B0(new_n16647_), .Y(new_n16648_));
  OAI22X1  g16456(.A0(new_n16648_), .A1(new_n16644_), .B0(new_n16623_), .B1(new_n15990_), .Y(new_n16649_));
  AND2X1   g16457(.A(new_n16649_), .B(\asqrt[15] ), .Y(new_n16650_));
  OR4X1    g16458(.A(new_n16643_), .B(new_n16642_), .C(new_n16599_), .D(new_n16609_), .Y(new_n16651_));
  OAI21X1  g16459(.A0(new_n16616_), .A1(new_n16603_), .B0(new_n16620_), .Y(new_n16652_));
  AOI21X1  g16460(.A0(new_n16641_), .A1(new_n16637_), .B0(new_n16016_), .Y(new_n16653_));
  AOI21X1  g16461(.A0(new_n16652_), .A1(\a[27] ), .B0(new_n16653_), .Y(new_n16654_));
  NAND2X1  g16462(.A(new_n16654_), .B(new_n16651_), .Y(new_n16655_));
  AOI21X1  g16463(.A0(new_n16622_), .A1(new_n16619_), .B0(new_n15990_), .Y(new_n16656_));
  NOR2X1   g16464(.A(new_n16656_), .B(\asqrt[15] ), .Y(new_n16657_));
  AND2X1   g16465(.A(new_n16639_), .B(new_n16638_), .Y(new_n16658_));
  OR2X1    g16466(.A(new_n16614_), .B(new_n15990_), .Y(new_n16659_));
  OR4X1    g16467(.A(new_n16659_), .B(new_n16608_), .C(new_n16658_), .D(new_n16603_), .Y(new_n16660_));
  AOI21X1  g16468(.A0(new_n16660_), .A1(new_n16647_), .B0(new_n16009_), .Y(new_n16661_));
  NOR4X1   g16469(.A(new_n16659_), .B(new_n16608_), .C(new_n16658_), .D(new_n16603_), .Y(new_n16662_));
  NOR3X1   g16470(.A(new_n16662_), .B(new_n16653_), .C(\a[28] ), .Y(new_n16663_));
  NOR2X1   g16471(.A(new_n16663_), .B(new_n16661_), .Y(new_n16664_));
  AOI21X1  g16472(.A0(new_n16657_), .A1(new_n16655_), .B0(new_n16664_), .Y(new_n16665_));
  OAI21X1  g16473(.A0(new_n16665_), .A1(new_n16650_), .B0(\asqrt[16] ), .Y(new_n16666_));
  AND2X1   g16474(.A(new_n16056_), .B(new_n16054_), .Y(new_n16667_));
  NOR3X1   g16475(.A(new_n16667_), .B(new_n16008_), .C(new_n16004_), .Y(new_n16668_));
  OAI21X1  g16476(.A0(new_n16616_), .A1(new_n16603_), .B0(new_n16668_), .Y(new_n16669_));
  AOI21X1  g16477(.A0(new_n16003_), .A1(\asqrt[15] ), .B0(new_n16008_), .Y(new_n16670_));
  OAI21X1  g16478(.A0(new_n16616_), .A1(new_n16603_), .B0(new_n16670_), .Y(new_n16671_));
  NAND2X1  g16479(.A(new_n16671_), .B(new_n16667_), .Y(new_n16672_));
  NAND2X1  g16480(.A(new_n16672_), .B(new_n16669_), .Y(new_n16673_));
  AOI21X1  g16481(.A0(new_n16654_), .A1(new_n16651_), .B0(new_n16656_), .Y(new_n16674_));
  OAI21X1  g16482(.A0(new_n16674_), .A1(new_n15362_), .B0(new_n14754_), .Y(new_n16675_));
  OAI21X1  g16483(.A0(new_n16675_), .A1(new_n16665_), .B0(new_n16673_), .Y(new_n16676_));
  AOI21X1  g16484(.A0(new_n16676_), .A1(new_n16666_), .B0(new_n14165_), .Y(new_n16677_));
  AND2X1   g16485(.A(new_n16059_), .B(new_n16057_), .Y(new_n16678_));
  NOR3X1   g16486(.A(new_n16025_), .B(new_n16678_), .C(new_n16058_), .Y(new_n16679_));
  OAI21X1  g16487(.A0(new_n16616_), .A1(new_n16603_), .B0(new_n16679_), .Y(new_n16680_));
  NOR2X1   g16488(.A(new_n16678_), .B(new_n16058_), .Y(new_n16681_));
  OAI21X1  g16489(.A0(new_n16616_), .A1(new_n16603_), .B0(new_n16681_), .Y(new_n16682_));
  NAND2X1  g16490(.A(new_n16682_), .B(new_n16025_), .Y(new_n16683_));
  AND2X1   g16491(.A(new_n16683_), .B(new_n16680_), .Y(new_n16684_));
  INVX1    g16492(.A(new_n16684_), .Y(new_n16685_));
  NAND3X1  g16493(.A(new_n16676_), .B(new_n16666_), .C(new_n14165_), .Y(new_n16686_));
  AOI21X1  g16494(.A0(new_n16686_), .A1(new_n16685_), .B0(new_n16677_), .Y(new_n16687_));
  OR2X1    g16495(.A(new_n16687_), .B(new_n13571_), .Y(new_n16688_));
  OR2X1    g16496(.A(new_n16674_), .B(new_n15362_), .Y(new_n16689_));
  AND2X1   g16497(.A(new_n16654_), .B(new_n16651_), .Y(new_n16690_));
  OR2X1    g16498(.A(new_n16656_), .B(\asqrt[15] ), .Y(new_n16691_));
  OR2X1    g16499(.A(new_n16663_), .B(new_n16661_), .Y(new_n16692_));
  OAI21X1  g16500(.A0(new_n16691_), .A1(new_n16690_), .B0(new_n16692_), .Y(new_n16693_));
  AOI21X1  g16501(.A0(new_n16693_), .A1(new_n16689_), .B0(new_n14754_), .Y(new_n16694_));
  AOI21X1  g16502(.A0(new_n16649_), .A1(\asqrt[15] ), .B0(\asqrt[16] ), .Y(new_n16695_));
  AOI22X1  g16503(.A0(new_n16695_), .A1(new_n16693_), .B0(new_n16672_), .B1(new_n16669_), .Y(new_n16696_));
  NOR3X1   g16504(.A(new_n16696_), .B(new_n16694_), .C(\asqrt[17] ), .Y(new_n16697_));
  NOR2X1   g16505(.A(new_n16697_), .B(new_n16684_), .Y(new_n16698_));
  NOR3X1   g16506(.A(new_n16064_), .B(new_n16032_), .C(new_n16027_), .Y(new_n16699_));
  NAND3X1  g16507(.A(\asqrt[13] ), .B(new_n16033_), .C(new_n16063_), .Y(new_n16700_));
  AOI22X1  g16508(.A0(new_n16700_), .A1(new_n16032_), .B0(new_n16699_), .B1(\asqrt[13] ), .Y(new_n16701_));
  INVX1    g16509(.A(new_n16701_), .Y(new_n16702_));
  OR2X1    g16510(.A(new_n16677_), .B(\asqrt[18] ), .Y(new_n16703_));
  OAI21X1  g16511(.A0(new_n16703_), .A1(new_n16698_), .B0(new_n16702_), .Y(new_n16704_));
  AOI21X1  g16512(.A0(new_n16704_), .A1(new_n16688_), .B0(new_n13000_), .Y(new_n16705_));
  AOI21X1  g16513(.A0(new_n16079_), .A1(new_n16078_), .B0(new_n16042_), .Y(new_n16706_));
  AND2X1   g16514(.A(new_n16706_), .B(new_n16035_), .Y(new_n16707_));
  AOI22X1  g16515(.A0(new_n16079_), .A1(new_n16078_), .B0(new_n16065_), .B1(\asqrt[18] ), .Y(new_n16708_));
  AOI21X1  g16516(.A0(new_n16708_), .A1(\asqrt[13] ), .B0(new_n16041_), .Y(new_n16709_));
  AOI21X1  g16517(.A0(new_n16707_), .A1(\asqrt[13] ), .B0(new_n16709_), .Y(new_n16710_));
  OAI21X1  g16518(.A0(new_n16696_), .A1(new_n16694_), .B0(\asqrt[17] ), .Y(new_n16711_));
  OAI21X1  g16519(.A0(new_n16697_), .A1(new_n16684_), .B0(new_n16711_), .Y(new_n16712_));
  AOI21X1  g16520(.A0(new_n16712_), .A1(\asqrt[18] ), .B0(\asqrt[19] ), .Y(new_n16713_));
  AOI21X1  g16521(.A0(new_n16713_), .A1(new_n16704_), .B0(new_n16710_), .Y(new_n16714_));
  OAI21X1  g16522(.A0(new_n16714_), .A1(new_n16705_), .B0(\asqrt[20] ), .Y(new_n16715_));
  AND2X1   g16523(.A(new_n16066_), .B(new_n16044_), .Y(new_n16716_));
  NOR3X1   g16524(.A(new_n16716_), .B(new_n16082_), .C(new_n16045_), .Y(new_n16717_));
  NOR3X1   g16525(.A(new_n16617_), .B(new_n16716_), .C(new_n16045_), .Y(new_n16718_));
  NOR2X1   g16526(.A(new_n16718_), .B(new_n16050_), .Y(new_n16719_));
  AOI21X1  g16527(.A0(new_n16717_), .A1(\asqrt[13] ), .B0(new_n16719_), .Y(new_n16720_));
  NOR3X1   g16528(.A(new_n16714_), .B(new_n16705_), .C(\asqrt[20] ), .Y(new_n16721_));
  OAI21X1  g16529(.A0(new_n16721_), .A1(new_n16720_), .B0(new_n16715_), .Y(new_n16722_));
  AND2X1   g16530(.A(new_n16722_), .B(\asqrt[21] ), .Y(new_n16723_));
  OR2X1    g16531(.A(new_n16721_), .B(new_n16720_), .Y(new_n16724_));
  NOR3X1   g16532(.A(new_n16073_), .B(new_n16076_), .C(new_n16092_), .Y(new_n16725_));
  NOR3X1   g16533(.A(new_n16617_), .B(new_n16073_), .C(new_n16092_), .Y(new_n16726_));
  NOR2X1   g16534(.A(new_n16726_), .B(new_n16072_), .Y(new_n16727_));
  AOI21X1  g16535(.A0(new_n16725_), .A1(\asqrt[13] ), .B0(new_n16727_), .Y(new_n16728_));
  AND2X1   g16536(.A(new_n16715_), .B(new_n11896_), .Y(new_n16729_));
  AOI21X1  g16537(.A0(new_n16729_), .A1(new_n16724_), .B0(new_n16728_), .Y(new_n16730_));
  OAI21X1  g16538(.A0(new_n16730_), .A1(new_n16723_), .B0(\asqrt[22] ), .Y(new_n16731_));
  AND2X1   g16539(.A(new_n16093_), .B(new_n16086_), .Y(new_n16732_));
  NOR3X1   g16540(.A(new_n16732_), .B(new_n16131_), .C(new_n16075_), .Y(new_n16733_));
  NOR3X1   g16541(.A(new_n16617_), .B(new_n16732_), .C(new_n16075_), .Y(new_n16734_));
  NOR2X1   g16542(.A(new_n16734_), .B(new_n16091_), .Y(new_n16735_));
  AOI21X1  g16543(.A0(new_n16733_), .A1(\asqrt[13] ), .B0(new_n16735_), .Y(new_n16736_));
  INVX1    g16544(.A(new_n16736_), .Y(new_n16737_));
  AND2X1   g16545(.A(new_n16712_), .B(\asqrt[18] ), .Y(new_n16738_));
  OR2X1    g16546(.A(new_n16697_), .B(new_n16684_), .Y(new_n16739_));
  NOR2X1   g16547(.A(new_n16677_), .B(\asqrt[18] ), .Y(new_n16740_));
  AOI21X1  g16548(.A0(new_n16740_), .A1(new_n16739_), .B0(new_n16701_), .Y(new_n16741_));
  OAI21X1  g16549(.A0(new_n16741_), .A1(new_n16738_), .B0(\asqrt[19] ), .Y(new_n16742_));
  INVX1    g16550(.A(new_n16710_), .Y(new_n16743_));
  OAI21X1  g16551(.A0(new_n16687_), .A1(new_n13571_), .B0(new_n13000_), .Y(new_n16744_));
  OAI21X1  g16552(.A0(new_n16744_), .A1(new_n16741_), .B0(new_n16743_), .Y(new_n16745_));
  AOI21X1  g16553(.A0(new_n16745_), .A1(new_n16742_), .B0(new_n12447_), .Y(new_n16746_));
  INVX1    g16554(.A(new_n16720_), .Y(new_n16747_));
  NAND3X1  g16555(.A(new_n16745_), .B(new_n16742_), .C(new_n12447_), .Y(new_n16748_));
  AOI21X1  g16556(.A0(new_n16748_), .A1(new_n16747_), .B0(new_n16746_), .Y(new_n16749_));
  OAI21X1  g16557(.A0(new_n16749_), .A1(new_n11896_), .B0(new_n11362_), .Y(new_n16750_));
  OAI21X1  g16558(.A0(new_n16750_), .A1(new_n16730_), .B0(new_n16737_), .Y(new_n16751_));
  AOI21X1  g16559(.A0(new_n16751_), .A1(new_n16731_), .B0(new_n10849_), .Y(new_n16752_));
  AND2X1   g16560(.A(new_n16135_), .B(new_n16133_), .Y(new_n16753_));
  NOR3X1   g16561(.A(new_n16753_), .B(new_n16101_), .C(new_n16134_), .Y(new_n16754_));
  NOR3X1   g16562(.A(new_n16617_), .B(new_n16753_), .C(new_n16134_), .Y(new_n16755_));
  NOR2X1   g16563(.A(new_n16755_), .B(new_n16100_), .Y(new_n16756_));
  AOI21X1  g16564(.A0(new_n16754_), .A1(\asqrt[13] ), .B0(new_n16756_), .Y(new_n16757_));
  INVX1    g16565(.A(new_n16757_), .Y(new_n16758_));
  NAND3X1  g16566(.A(new_n16751_), .B(new_n16731_), .C(new_n10849_), .Y(new_n16759_));
  AOI21X1  g16567(.A0(new_n16759_), .A1(new_n16758_), .B0(new_n16752_), .Y(new_n16760_));
  OR2X1    g16568(.A(new_n16760_), .B(new_n10332_), .Y(new_n16761_));
  OR2X1    g16569(.A(new_n16749_), .B(new_n11896_), .Y(new_n16762_));
  NOR2X1   g16570(.A(new_n16721_), .B(new_n16720_), .Y(new_n16763_));
  INVX1    g16571(.A(new_n16728_), .Y(new_n16764_));
  NAND2X1  g16572(.A(new_n16715_), .B(new_n11896_), .Y(new_n16765_));
  OAI21X1  g16573(.A0(new_n16765_), .A1(new_n16763_), .B0(new_n16764_), .Y(new_n16766_));
  AOI21X1  g16574(.A0(new_n16766_), .A1(new_n16762_), .B0(new_n11362_), .Y(new_n16767_));
  AOI21X1  g16575(.A0(new_n16722_), .A1(\asqrt[21] ), .B0(\asqrt[22] ), .Y(new_n16768_));
  AOI21X1  g16576(.A0(new_n16768_), .A1(new_n16766_), .B0(new_n16736_), .Y(new_n16769_));
  NOR3X1   g16577(.A(new_n16769_), .B(new_n16767_), .C(\asqrt[23] ), .Y(new_n16770_));
  NOR2X1   g16578(.A(new_n16770_), .B(new_n16757_), .Y(new_n16771_));
  NAND4X1  g16579(.A(\asqrt[13] ), .B(new_n16111_), .C(new_n16109_), .D(new_n16137_), .Y(new_n16772_));
  NAND2X1  g16580(.A(new_n16111_), .B(new_n16137_), .Y(new_n16773_));
  OAI21X1  g16581(.A0(new_n16773_), .A1(new_n16617_), .B0(new_n16110_), .Y(new_n16774_));
  AND2X1   g16582(.A(new_n16774_), .B(new_n16772_), .Y(new_n16775_));
  INVX1    g16583(.A(new_n16775_), .Y(new_n16776_));
  OAI21X1  g16584(.A0(new_n16769_), .A1(new_n16767_), .B0(\asqrt[23] ), .Y(new_n16777_));
  NAND2X1  g16585(.A(new_n16777_), .B(new_n10332_), .Y(new_n16778_));
  OAI21X1  g16586(.A0(new_n16778_), .A1(new_n16771_), .B0(new_n16776_), .Y(new_n16779_));
  AOI21X1  g16587(.A0(new_n16779_), .A1(new_n16761_), .B0(new_n9833_), .Y(new_n16780_));
  AOI21X1  g16588(.A0(new_n16153_), .A1(new_n16152_), .B0(new_n16120_), .Y(new_n16781_));
  AND2X1   g16589(.A(new_n16781_), .B(new_n16113_), .Y(new_n16782_));
  AOI22X1  g16590(.A0(new_n16153_), .A1(new_n16152_), .B0(new_n16139_), .B1(\asqrt[24] ), .Y(new_n16783_));
  AOI21X1  g16591(.A0(new_n16783_), .A1(\asqrt[13] ), .B0(new_n16119_), .Y(new_n16784_));
  AOI21X1  g16592(.A0(new_n16782_), .A1(\asqrt[13] ), .B0(new_n16784_), .Y(new_n16785_));
  OAI21X1  g16593(.A0(new_n16770_), .A1(new_n16757_), .B0(new_n16777_), .Y(new_n16786_));
  AOI21X1  g16594(.A0(new_n16786_), .A1(\asqrt[24] ), .B0(\asqrt[25] ), .Y(new_n16787_));
  AOI21X1  g16595(.A0(new_n16787_), .A1(new_n16779_), .B0(new_n16785_), .Y(new_n16788_));
  OAI21X1  g16596(.A0(new_n16788_), .A1(new_n16780_), .B0(\asqrt[26] ), .Y(new_n16789_));
  AND2X1   g16597(.A(new_n16140_), .B(new_n16122_), .Y(new_n16790_));
  NOR3X1   g16598(.A(new_n16790_), .B(new_n16156_), .C(new_n16123_), .Y(new_n16791_));
  NOR3X1   g16599(.A(new_n16617_), .B(new_n16790_), .C(new_n16123_), .Y(new_n16792_));
  NOR2X1   g16600(.A(new_n16792_), .B(new_n16128_), .Y(new_n16793_));
  AOI21X1  g16601(.A0(new_n16791_), .A1(\asqrt[13] ), .B0(new_n16793_), .Y(new_n16794_));
  NOR3X1   g16602(.A(new_n16788_), .B(new_n16780_), .C(\asqrt[26] ), .Y(new_n16795_));
  OAI21X1  g16603(.A0(new_n16795_), .A1(new_n16794_), .B0(new_n16789_), .Y(new_n16796_));
  AND2X1   g16604(.A(new_n16796_), .B(\asqrt[27] ), .Y(new_n16797_));
  INVX1    g16605(.A(new_n16794_), .Y(new_n16798_));
  AND2X1   g16606(.A(new_n16786_), .B(\asqrt[24] ), .Y(new_n16799_));
  OR2X1    g16607(.A(new_n16770_), .B(new_n16757_), .Y(new_n16800_));
  AND2X1   g16608(.A(new_n16777_), .B(new_n10332_), .Y(new_n16801_));
  AOI21X1  g16609(.A0(new_n16801_), .A1(new_n16800_), .B0(new_n16775_), .Y(new_n16802_));
  OAI21X1  g16610(.A0(new_n16802_), .A1(new_n16799_), .B0(\asqrt[25] ), .Y(new_n16803_));
  INVX1    g16611(.A(new_n16785_), .Y(new_n16804_));
  OAI21X1  g16612(.A0(new_n16760_), .A1(new_n10332_), .B0(new_n9833_), .Y(new_n16805_));
  OAI21X1  g16613(.A0(new_n16805_), .A1(new_n16802_), .B0(new_n16804_), .Y(new_n16806_));
  NAND3X1  g16614(.A(new_n16806_), .B(new_n16803_), .C(new_n9353_), .Y(new_n16807_));
  NAND2X1  g16615(.A(new_n16807_), .B(new_n16798_), .Y(new_n16808_));
  NAND4X1  g16616(.A(\asqrt[13] ), .B(new_n16159_), .C(new_n16146_), .D(new_n16142_), .Y(new_n16809_));
  NAND2X1  g16617(.A(new_n16159_), .B(new_n16142_), .Y(new_n16810_));
  OAI21X1  g16618(.A0(new_n16810_), .A1(new_n16617_), .B0(new_n16150_), .Y(new_n16811_));
  AND2X1   g16619(.A(new_n16811_), .B(new_n16809_), .Y(new_n16812_));
  AOI21X1  g16620(.A0(new_n16806_), .A1(new_n16803_), .B0(new_n9353_), .Y(new_n16813_));
  NOR2X1   g16621(.A(new_n16813_), .B(\asqrt[27] ), .Y(new_n16814_));
  AOI21X1  g16622(.A0(new_n16814_), .A1(new_n16808_), .B0(new_n16812_), .Y(new_n16815_));
  OAI21X1  g16623(.A0(new_n16815_), .A1(new_n16797_), .B0(\asqrt[28] ), .Y(new_n16816_));
  AND2X1   g16624(.A(new_n16167_), .B(new_n16160_), .Y(new_n16817_));
  NOR3X1   g16625(.A(new_n16817_), .B(new_n16205_), .C(new_n16149_), .Y(new_n16818_));
  NOR3X1   g16626(.A(new_n16617_), .B(new_n16817_), .C(new_n16149_), .Y(new_n16819_));
  NOR2X1   g16627(.A(new_n16819_), .B(new_n16165_), .Y(new_n16820_));
  AOI21X1  g16628(.A0(new_n16818_), .A1(\asqrt[13] ), .B0(new_n16820_), .Y(new_n16821_));
  INVX1    g16629(.A(new_n16821_), .Y(new_n16822_));
  AOI21X1  g16630(.A0(new_n16807_), .A1(new_n16798_), .B0(new_n16813_), .Y(new_n16823_));
  OAI21X1  g16631(.A0(new_n16823_), .A1(new_n8874_), .B0(new_n8412_), .Y(new_n16824_));
  OAI21X1  g16632(.A0(new_n16824_), .A1(new_n16815_), .B0(new_n16822_), .Y(new_n16825_));
  AOI21X1  g16633(.A0(new_n16825_), .A1(new_n16816_), .B0(new_n7970_), .Y(new_n16826_));
  AND2X1   g16634(.A(new_n16209_), .B(new_n16207_), .Y(new_n16827_));
  NOR3X1   g16635(.A(new_n16827_), .B(new_n16175_), .C(new_n16208_), .Y(new_n16828_));
  NOR3X1   g16636(.A(new_n16617_), .B(new_n16827_), .C(new_n16208_), .Y(new_n16829_));
  NOR2X1   g16637(.A(new_n16829_), .B(new_n16174_), .Y(new_n16830_));
  AOI21X1  g16638(.A0(new_n16828_), .A1(\asqrt[13] ), .B0(new_n16830_), .Y(new_n16831_));
  INVX1    g16639(.A(new_n16831_), .Y(new_n16832_));
  NAND3X1  g16640(.A(new_n16825_), .B(new_n16816_), .C(new_n7970_), .Y(new_n16833_));
  AOI21X1  g16641(.A0(new_n16833_), .A1(new_n16832_), .B0(new_n16826_), .Y(new_n16834_));
  OR2X1    g16642(.A(new_n16834_), .B(new_n7527_), .Y(new_n16835_));
  AND2X1   g16643(.A(new_n16833_), .B(new_n16832_), .Y(new_n16836_));
  NAND4X1  g16644(.A(\asqrt[13] ), .B(new_n16185_), .C(new_n16183_), .D(new_n16211_), .Y(new_n16837_));
  NAND2X1  g16645(.A(new_n16185_), .B(new_n16211_), .Y(new_n16838_));
  OAI21X1  g16646(.A0(new_n16838_), .A1(new_n16617_), .B0(new_n16184_), .Y(new_n16839_));
  AND2X1   g16647(.A(new_n16839_), .B(new_n16837_), .Y(new_n16840_));
  INVX1    g16648(.A(new_n16840_), .Y(new_n16841_));
  OR2X1    g16649(.A(new_n16826_), .B(\asqrt[30] ), .Y(new_n16842_));
  OAI21X1  g16650(.A0(new_n16842_), .A1(new_n16836_), .B0(new_n16841_), .Y(new_n16843_));
  AOI21X1  g16651(.A0(new_n16843_), .A1(new_n16835_), .B0(new_n7103_), .Y(new_n16844_));
  AOI21X1  g16652(.A0(new_n16241_), .A1(new_n16240_), .B0(new_n16194_), .Y(new_n16845_));
  AND2X1   g16653(.A(new_n16845_), .B(new_n16187_), .Y(new_n16846_));
  AOI22X1  g16654(.A0(new_n16241_), .A1(new_n16240_), .B0(new_n16213_), .B1(\asqrt[30] ), .Y(new_n16847_));
  AOI21X1  g16655(.A0(new_n16847_), .A1(\asqrt[13] ), .B0(new_n16193_), .Y(new_n16848_));
  AOI21X1  g16656(.A0(new_n16846_), .A1(\asqrt[13] ), .B0(new_n16848_), .Y(new_n16849_));
  OR2X1    g16657(.A(new_n16823_), .B(new_n8874_), .Y(new_n16850_));
  AND2X1   g16658(.A(new_n16807_), .B(new_n16798_), .Y(new_n16851_));
  INVX1    g16659(.A(new_n16812_), .Y(new_n16852_));
  OR2X1    g16660(.A(new_n16813_), .B(\asqrt[27] ), .Y(new_n16853_));
  OAI21X1  g16661(.A0(new_n16853_), .A1(new_n16851_), .B0(new_n16852_), .Y(new_n16854_));
  AOI21X1  g16662(.A0(new_n16854_), .A1(new_n16850_), .B0(new_n8412_), .Y(new_n16855_));
  AOI21X1  g16663(.A0(new_n16796_), .A1(\asqrt[27] ), .B0(\asqrt[28] ), .Y(new_n16856_));
  AOI21X1  g16664(.A0(new_n16856_), .A1(new_n16854_), .B0(new_n16821_), .Y(new_n16857_));
  OAI21X1  g16665(.A0(new_n16857_), .A1(new_n16855_), .B0(\asqrt[29] ), .Y(new_n16858_));
  NOR3X1   g16666(.A(new_n16857_), .B(new_n16855_), .C(\asqrt[29] ), .Y(new_n16859_));
  OAI21X1  g16667(.A0(new_n16859_), .A1(new_n16831_), .B0(new_n16858_), .Y(new_n16860_));
  AOI21X1  g16668(.A0(new_n16860_), .A1(\asqrt[30] ), .B0(\asqrt[31] ), .Y(new_n16861_));
  AOI21X1  g16669(.A0(new_n16861_), .A1(new_n16843_), .B0(new_n16849_), .Y(new_n16862_));
  OAI21X1  g16670(.A0(new_n16862_), .A1(new_n16844_), .B0(\asqrt[32] ), .Y(new_n16863_));
  AND2X1   g16671(.A(new_n16214_), .B(new_n16196_), .Y(new_n16864_));
  NOR3X1   g16672(.A(new_n16864_), .B(new_n16244_), .C(new_n16197_), .Y(new_n16865_));
  NOR3X1   g16673(.A(new_n16617_), .B(new_n16864_), .C(new_n16197_), .Y(new_n16866_));
  NOR2X1   g16674(.A(new_n16866_), .B(new_n16202_), .Y(new_n16867_));
  AOI21X1  g16675(.A0(new_n16865_), .A1(\asqrt[13] ), .B0(new_n16867_), .Y(new_n16868_));
  NOR3X1   g16676(.A(new_n16862_), .B(new_n16844_), .C(\asqrt[32] ), .Y(new_n16869_));
  OAI21X1  g16677(.A0(new_n16869_), .A1(new_n16868_), .B0(new_n16863_), .Y(new_n16870_));
  AND2X1   g16678(.A(new_n16870_), .B(\asqrt[33] ), .Y(new_n16871_));
  OR2X1    g16679(.A(new_n16869_), .B(new_n16868_), .Y(new_n16872_));
  OR4X1    g16680(.A(new_n16617_), .B(new_n16221_), .C(new_n16248_), .D(new_n16247_), .Y(new_n16873_));
  OR2X1    g16681(.A(new_n16221_), .B(new_n16247_), .Y(new_n16874_));
  OAI21X1  g16682(.A0(new_n16874_), .A1(new_n16617_), .B0(new_n16248_), .Y(new_n16875_));
  AND2X1   g16683(.A(new_n16875_), .B(new_n16873_), .Y(new_n16876_));
  AND2X1   g16684(.A(new_n16863_), .B(new_n6294_), .Y(new_n16877_));
  AOI21X1  g16685(.A0(new_n16877_), .A1(new_n16872_), .B0(new_n16876_), .Y(new_n16878_));
  OAI21X1  g16686(.A0(new_n16878_), .A1(new_n16871_), .B0(\asqrt[34] ), .Y(new_n16879_));
  AND2X1   g16687(.A(new_n16230_), .B(new_n16224_), .Y(new_n16880_));
  NOR3X1   g16688(.A(new_n16880_), .B(new_n16264_), .C(new_n16223_), .Y(new_n16881_));
  NOR3X1   g16689(.A(new_n16617_), .B(new_n16880_), .C(new_n16223_), .Y(new_n16882_));
  NOR2X1   g16690(.A(new_n16882_), .B(new_n16229_), .Y(new_n16883_));
  AOI21X1  g16691(.A0(new_n16881_), .A1(\asqrt[13] ), .B0(new_n16883_), .Y(new_n16884_));
  INVX1    g16692(.A(new_n16884_), .Y(new_n16885_));
  AND2X1   g16693(.A(new_n16860_), .B(\asqrt[30] ), .Y(new_n16886_));
  NAND2X1  g16694(.A(new_n16833_), .B(new_n16832_), .Y(new_n16887_));
  NOR2X1   g16695(.A(new_n16826_), .B(\asqrt[30] ), .Y(new_n16888_));
  AOI21X1  g16696(.A0(new_n16888_), .A1(new_n16887_), .B0(new_n16840_), .Y(new_n16889_));
  OAI21X1  g16697(.A0(new_n16889_), .A1(new_n16886_), .B0(\asqrt[31] ), .Y(new_n16890_));
  INVX1    g16698(.A(new_n16849_), .Y(new_n16891_));
  OAI21X1  g16699(.A0(new_n16834_), .A1(new_n7527_), .B0(new_n7103_), .Y(new_n16892_));
  OAI21X1  g16700(.A0(new_n16892_), .A1(new_n16889_), .B0(new_n16891_), .Y(new_n16893_));
  AOI21X1  g16701(.A0(new_n16893_), .A1(new_n16890_), .B0(new_n6699_), .Y(new_n16894_));
  INVX1    g16702(.A(new_n16868_), .Y(new_n16895_));
  NAND3X1  g16703(.A(new_n16893_), .B(new_n16890_), .C(new_n6699_), .Y(new_n16896_));
  AOI21X1  g16704(.A0(new_n16896_), .A1(new_n16895_), .B0(new_n16894_), .Y(new_n16897_));
  OAI21X1  g16705(.A0(new_n16897_), .A1(new_n6294_), .B0(new_n5941_), .Y(new_n16898_));
  OAI21X1  g16706(.A0(new_n16898_), .A1(new_n16878_), .B0(new_n16885_), .Y(new_n16899_));
  AOI21X1  g16707(.A0(new_n16899_), .A1(new_n16879_), .B0(new_n5541_), .Y(new_n16900_));
  AND2X1   g16708(.A(new_n16268_), .B(new_n16266_), .Y(new_n16901_));
  NOR3X1   g16709(.A(new_n16901_), .B(new_n16238_), .C(new_n16267_), .Y(new_n16902_));
  NOR3X1   g16710(.A(new_n16617_), .B(new_n16901_), .C(new_n16267_), .Y(new_n16903_));
  NOR2X1   g16711(.A(new_n16903_), .B(new_n16237_), .Y(new_n16904_));
  AOI21X1  g16712(.A0(new_n16902_), .A1(\asqrt[13] ), .B0(new_n16904_), .Y(new_n16905_));
  INVX1    g16713(.A(new_n16905_), .Y(new_n16906_));
  NAND3X1  g16714(.A(new_n16899_), .B(new_n16879_), .C(new_n5541_), .Y(new_n16907_));
  AOI21X1  g16715(.A0(new_n16907_), .A1(new_n16906_), .B0(new_n16900_), .Y(new_n16908_));
  OR2X1    g16716(.A(new_n16908_), .B(new_n5176_), .Y(new_n16909_));
  OR2X1    g16717(.A(new_n16897_), .B(new_n6294_), .Y(new_n16910_));
  NOR2X1   g16718(.A(new_n16869_), .B(new_n16868_), .Y(new_n16911_));
  INVX1    g16719(.A(new_n16876_), .Y(new_n16912_));
  NAND2X1  g16720(.A(new_n16863_), .B(new_n6294_), .Y(new_n16913_));
  OAI21X1  g16721(.A0(new_n16913_), .A1(new_n16911_), .B0(new_n16912_), .Y(new_n16914_));
  AOI21X1  g16722(.A0(new_n16914_), .A1(new_n16910_), .B0(new_n5941_), .Y(new_n16915_));
  AOI21X1  g16723(.A0(new_n16870_), .A1(\asqrt[33] ), .B0(\asqrt[34] ), .Y(new_n16916_));
  AOI21X1  g16724(.A0(new_n16916_), .A1(new_n16914_), .B0(new_n16884_), .Y(new_n16917_));
  NOR3X1   g16725(.A(new_n16917_), .B(new_n16915_), .C(\asqrt[35] ), .Y(new_n16918_));
  NOR2X1   g16726(.A(new_n16918_), .B(new_n16905_), .Y(new_n16919_));
  OR4X1    g16727(.A(new_n16617_), .B(new_n16270_), .C(new_n16258_), .D(new_n16253_), .Y(new_n16920_));
  OR2X1    g16728(.A(new_n16270_), .B(new_n16253_), .Y(new_n16921_));
  OAI21X1  g16729(.A0(new_n16921_), .A1(new_n16617_), .B0(new_n16258_), .Y(new_n16922_));
  AND2X1   g16730(.A(new_n16922_), .B(new_n16920_), .Y(new_n16923_));
  INVX1    g16731(.A(new_n16923_), .Y(new_n16924_));
  OAI21X1  g16732(.A0(new_n16917_), .A1(new_n16915_), .B0(\asqrt[35] ), .Y(new_n16925_));
  NAND2X1  g16733(.A(new_n16925_), .B(new_n5176_), .Y(new_n16926_));
  OAI21X1  g16734(.A0(new_n16926_), .A1(new_n16919_), .B0(new_n16924_), .Y(new_n16927_));
  AOI21X1  g16735(.A0(new_n16927_), .A1(new_n16909_), .B0(new_n4826_), .Y(new_n16928_));
  AOI21X1  g16736(.A0(new_n16315_), .A1(new_n16314_), .B0(new_n16277_), .Y(new_n16929_));
  AND2X1   g16737(.A(new_n16929_), .B(new_n16261_), .Y(new_n16930_));
  AOI22X1  g16738(.A0(new_n16315_), .A1(new_n16314_), .B0(new_n16287_), .B1(\asqrt[36] ), .Y(new_n16931_));
  AOI21X1  g16739(.A0(new_n16931_), .A1(\asqrt[13] ), .B0(new_n16276_), .Y(new_n16932_));
  AOI21X1  g16740(.A0(new_n16930_), .A1(\asqrt[13] ), .B0(new_n16932_), .Y(new_n16933_));
  OAI21X1  g16741(.A0(new_n16918_), .A1(new_n16905_), .B0(new_n16925_), .Y(new_n16934_));
  AOI21X1  g16742(.A0(new_n16934_), .A1(\asqrt[36] ), .B0(\asqrt[37] ), .Y(new_n16935_));
  AOI21X1  g16743(.A0(new_n16935_), .A1(new_n16927_), .B0(new_n16933_), .Y(new_n16936_));
  OAI21X1  g16744(.A0(new_n16936_), .A1(new_n16928_), .B0(\asqrt[38] ), .Y(new_n16937_));
  AND2X1   g16745(.A(new_n16288_), .B(new_n16280_), .Y(new_n16938_));
  NOR3X1   g16746(.A(new_n16938_), .B(new_n16318_), .C(new_n16281_), .Y(new_n16939_));
  NOR3X1   g16747(.A(new_n16617_), .B(new_n16938_), .C(new_n16281_), .Y(new_n16940_));
  NOR2X1   g16748(.A(new_n16940_), .B(new_n16286_), .Y(new_n16941_));
  AOI21X1  g16749(.A0(new_n16939_), .A1(\asqrt[13] ), .B0(new_n16941_), .Y(new_n16942_));
  NOR3X1   g16750(.A(new_n16936_), .B(new_n16928_), .C(\asqrt[38] ), .Y(new_n16943_));
  OAI21X1  g16751(.A0(new_n16943_), .A1(new_n16942_), .B0(new_n16937_), .Y(new_n16944_));
  AND2X1   g16752(.A(new_n16944_), .B(\asqrt[39] ), .Y(new_n16945_));
  OR2X1    g16753(.A(new_n16943_), .B(new_n16942_), .Y(new_n16946_));
  OR4X1    g16754(.A(new_n16617_), .B(new_n16295_), .C(new_n16322_), .D(new_n16321_), .Y(new_n16947_));
  OR2X1    g16755(.A(new_n16295_), .B(new_n16321_), .Y(new_n16948_));
  OAI21X1  g16756(.A0(new_n16948_), .A1(new_n16617_), .B0(new_n16322_), .Y(new_n16949_));
  AND2X1   g16757(.A(new_n16949_), .B(new_n16947_), .Y(new_n16950_));
  AND2X1   g16758(.A(new_n16937_), .B(new_n4165_), .Y(new_n16951_));
  AOI21X1  g16759(.A0(new_n16951_), .A1(new_n16946_), .B0(new_n16950_), .Y(new_n16952_));
  OAI21X1  g16760(.A0(new_n16952_), .A1(new_n16945_), .B0(\asqrt[40] ), .Y(new_n16953_));
  AND2X1   g16761(.A(new_n16304_), .B(new_n16298_), .Y(new_n16954_));
  NOR3X1   g16762(.A(new_n16954_), .B(new_n16338_), .C(new_n16297_), .Y(new_n16955_));
  NOR3X1   g16763(.A(new_n16617_), .B(new_n16954_), .C(new_n16297_), .Y(new_n16956_));
  NOR2X1   g16764(.A(new_n16956_), .B(new_n16303_), .Y(new_n16957_));
  AOI21X1  g16765(.A0(new_n16955_), .A1(\asqrt[13] ), .B0(new_n16957_), .Y(new_n16958_));
  INVX1    g16766(.A(new_n16958_), .Y(new_n16959_));
  AND2X1   g16767(.A(new_n16934_), .B(\asqrt[36] ), .Y(new_n16960_));
  OR2X1    g16768(.A(new_n16918_), .B(new_n16905_), .Y(new_n16961_));
  AND2X1   g16769(.A(new_n16925_), .B(new_n5176_), .Y(new_n16962_));
  AOI21X1  g16770(.A0(new_n16962_), .A1(new_n16961_), .B0(new_n16923_), .Y(new_n16963_));
  OAI21X1  g16771(.A0(new_n16963_), .A1(new_n16960_), .B0(\asqrt[37] ), .Y(new_n16964_));
  INVX1    g16772(.A(new_n16933_), .Y(new_n16965_));
  OAI21X1  g16773(.A0(new_n16908_), .A1(new_n5176_), .B0(new_n4826_), .Y(new_n16966_));
  OAI21X1  g16774(.A0(new_n16966_), .A1(new_n16963_), .B0(new_n16965_), .Y(new_n16967_));
  AOI21X1  g16775(.A0(new_n16967_), .A1(new_n16964_), .B0(new_n4493_), .Y(new_n16968_));
  INVX1    g16776(.A(new_n16942_), .Y(new_n16969_));
  NAND3X1  g16777(.A(new_n16967_), .B(new_n16964_), .C(new_n4493_), .Y(new_n16970_));
  AOI21X1  g16778(.A0(new_n16970_), .A1(new_n16969_), .B0(new_n16968_), .Y(new_n16971_));
  OAI21X1  g16779(.A0(new_n16971_), .A1(new_n4165_), .B0(new_n3863_), .Y(new_n16972_));
  OAI21X1  g16780(.A0(new_n16972_), .A1(new_n16952_), .B0(new_n16959_), .Y(new_n16973_));
  AOI21X1  g16781(.A0(new_n16973_), .A1(new_n16953_), .B0(new_n3564_), .Y(new_n16974_));
  AND2X1   g16782(.A(new_n16342_), .B(new_n16340_), .Y(new_n16975_));
  NOR3X1   g16783(.A(new_n16975_), .B(new_n16312_), .C(new_n16341_), .Y(new_n16976_));
  NOR3X1   g16784(.A(new_n16617_), .B(new_n16975_), .C(new_n16341_), .Y(new_n16977_));
  NOR2X1   g16785(.A(new_n16977_), .B(new_n16311_), .Y(new_n16978_));
  AOI21X1  g16786(.A0(new_n16976_), .A1(\asqrt[13] ), .B0(new_n16978_), .Y(new_n16979_));
  INVX1    g16787(.A(new_n16979_), .Y(new_n16980_));
  NAND3X1  g16788(.A(new_n16973_), .B(new_n16953_), .C(new_n3564_), .Y(new_n16981_));
  AOI21X1  g16789(.A0(new_n16981_), .A1(new_n16980_), .B0(new_n16974_), .Y(new_n16982_));
  OR2X1    g16790(.A(new_n16982_), .B(new_n3276_), .Y(new_n16983_));
  OR2X1    g16791(.A(new_n16971_), .B(new_n4165_), .Y(new_n16984_));
  NOR2X1   g16792(.A(new_n16943_), .B(new_n16942_), .Y(new_n16985_));
  INVX1    g16793(.A(new_n16950_), .Y(new_n16986_));
  NAND2X1  g16794(.A(new_n16937_), .B(new_n4165_), .Y(new_n16987_));
  OAI21X1  g16795(.A0(new_n16987_), .A1(new_n16985_), .B0(new_n16986_), .Y(new_n16988_));
  AOI21X1  g16796(.A0(new_n16988_), .A1(new_n16984_), .B0(new_n3863_), .Y(new_n16989_));
  AOI21X1  g16797(.A0(new_n16944_), .A1(\asqrt[39] ), .B0(\asqrt[40] ), .Y(new_n16990_));
  AOI21X1  g16798(.A0(new_n16990_), .A1(new_n16988_), .B0(new_n16958_), .Y(new_n16991_));
  NOR3X1   g16799(.A(new_n16991_), .B(new_n16989_), .C(\asqrt[41] ), .Y(new_n16992_));
  NOR2X1   g16800(.A(new_n16992_), .B(new_n16979_), .Y(new_n16993_));
  OR4X1    g16801(.A(new_n16617_), .B(new_n16344_), .C(new_n16332_), .D(new_n16327_), .Y(new_n16994_));
  OR2X1    g16802(.A(new_n16344_), .B(new_n16327_), .Y(new_n16995_));
  OAI21X1  g16803(.A0(new_n16995_), .A1(new_n16617_), .B0(new_n16332_), .Y(new_n16996_));
  AND2X1   g16804(.A(new_n16996_), .B(new_n16994_), .Y(new_n16997_));
  INVX1    g16805(.A(new_n16997_), .Y(new_n16998_));
  OAI21X1  g16806(.A0(new_n16991_), .A1(new_n16989_), .B0(\asqrt[41] ), .Y(new_n16999_));
  NAND2X1  g16807(.A(new_n16999_), .B(new_n3276_), .Y(new_n17000_));
  OAI21X1  g16808(.A0(new_n17000_), .A1(new_n16993_), .B0(new_n16998_), .Y(new_n17001_));
  AOI21X1  g16809(.A0(new_n17001_), .A1(new_n16983_), .B0(new_n3008_), .Y(new_n17002_));
  AOI21X1  g16810(.A0(new_n16389_), .A1(new_n16388_), .B0(new_n16351_), .Y(new_n17003_));
  AND2X1   g16811(.A(new_n17003_), .B(new_n16335_), .Y(new_n17004_));
  AOI22X1  g16812(.A0(new_n16389_), .A1(new_n16388_), .B0(new_n16361_), .B1(\asqrt[42] ), .Y(new_n17005_));
  AOI21X1  g16813(.A0(new_n17005_), .A1(\asqrt[13] ), .B0(new_n16350_), .Y(new_n17006_));
  AOI21X1  g16814(.A0(new_n17004_), .A1(\asqrt[13] ), .B0(new_n17006_), .Y(new_n17007_));
  OAI21X1  g16815(.A0(new_n16992_), .A1(new_n16979_), .B0(new_n16999_), .Y(new_n17008_));
  AOI21X1  g16816(.A0(new_n17008_), .A1(\asqrt[42] ), .B0(\asqrt[43] ), .Y(new_n17009_));
  AOI21X1  g16817(.A0(new_n17009_), .A1(new_n17001_), .B0(new_n17007_), .Y(new_n17010_));
  OAI21X1  g16818(.A0(new_n17010_), .A1(new_n17002_), .B0(\asqrt[44] ), .Y(new_n17011_));
  AND2X1   g16819(.A(new_n16362_), .B(new_n16354_), .Y(new_n17012_));
  NOR3X1   g16820(.A(new_n17012_), .B(new_n16392_), .C(new_n16355_), .Y(new_n17013_));
  NOR3X1   g16821(.A(new_n16617_), .B(new_n17012_), .C(new_n16355_), .Y(new_n17014_));
  NOR2X1   g16822(.A(new_n17014_), .B(new_n16360_), .Y(new_n17015_));
  AOI21X1  g16823(.A0(new_n17013_), .A1(\asqrt[13] ), .B0(new_n17015_), .Y(new_n17016_));
  NOR3X1   g16824(.A(new_n17010_), .B(new_n17002_), .C(\asqrt[44] ), .Y(new_n17017_));
  OAI21X1  g16825(.A0(new_n17017_), .A1(new_n17016_), .B0(new_n17011_), .Y(new_n17018_));
  AND2X1   g16826(.A(new_n17018_), .B(\asqrt[45] ), .Y(new_n17019_));
  OR2X1    g16827(.A(new_n17017_), .B(new_n17016_), .Y(new_n17020_));
  OR4X1    g16828(.A(new_n16617_), .B(new_n16369_), .C(new_n16396_), .D(new_n16395_), .Y(new_n17021_));
  OR2X1    g16829(.A(new_n16369_), .B(new_n16395_), .Y(new_n17022_));
  OAI21X1  g16830(.A0(new_n17022_), .A1(new_n16617_), .B0(new_n16396_), .Y(new_n17023_));
  AND2X1   g16831(.A(new_n17023_), .B(new_n17021_), .Y(new_n17024_));
  AND2X1   g16832(.A(new_n17011_), .B(new_n2570_), .Y(new_n17025_));
  AOI21X1  g16833(.A0(new_n17025_), .A1(new_n17020_), .B0(new_n17024_), .Y(new_n17026_));
  OAI21X1  g16834(.A0(new_n17026_), .A1(new_n17019_), .B0(\asqrt[46] ), .Y(new_n17027_));
  AND2X1   g16835(.A(new_n16378_), .B(new_n16372_), .Y(new_n17028_));
  NOR3X1   g16836(.A(new_n17028_), .B(new_n16412_), .C(new_n16371_), .Y(new_n17029_));
  NOR3X1   g16837(.A(new_n16617_), .B(new_n17028_), .C(new_n16371_), .Y(new_n17030_));
  NOR2X1   g16838(.A(new_n17030_), .B(new_n16377_), .Y(new_n17031_));
  AOI21X1  g16839(.A0(new_n17029_), .A1(\asqrt[13] ), .B0(new_n17031_), .Y(new_n17032_));
  INVX1    g16840(.A(new_n17032_), .Y(new_n17033_));
  AND2X1   g16841(.A(new_n17008_), .B(\asqrt[42] ), .Y(new_n17034_));
  OR2X1    g16842(.A(new_n16992_), .B(new_n16979_), .Y(new_n17035_));
  AND2X1   g16843(.A(new_n16999_), .B(new_n3276_), .Y(new_n17036_));
  AOI21X1  g16844(.A0(new_n17036_), .A1(new_n17035_), .B0(new_n16997_), .Y(new_n17037_));
  OAI21X1  g16845(.A0(new_n17037_), .A1(new_n17034_), .B0(\asqrt[43] ), .Y(new_n17038_));
  INVX1    g16846(.A(new_n17007_), .Y(new_n17039_));
  OAI21X1  g16847(.A0(new_n16982_), .A1(new_n3276_), .B0(new_n3008_), .Y(new_n17040_));
  OAI21X1  g16848(.A0(new_n17040_), .A1(new_n17037_), .B0(new_n17039_), .Y(new_n17041_));
  AOI21X1  g16849(.A0(new_n17041_), .A1(new_n17038_), .B0(new_n2769_), .Y(new_n17042_));
  INVX1    g16850(.A(new_n17016_), .Y(new_n17043_));
  NAND3X1  g16851(.A(new_n17041_), .B(new_n17038_), .C(new_n2769_), .Y(new_n17044_));
  AOI21X1  g16852(.A0(new_n17044_), .A1(new_n17043_), .B0(new_n17042_), .Y(new_n17045_));
  OAI21X1  g16853(.A0(new_n17045_), .A1(new_n2570_), .B0(new_n2263_), .Y(new_n17046_));
  OAI21X1  g16854(.A0(new_n17046_), .A1(new_n17026_), .B0(new_n17033_), .Y(new_n17047_));
  AOI21X1  g16855(.A0(new_n17047_), .A1(new_n17027_), .B0(new_n2040_), .Y(new_n17048_));
  AND2X1   g16856(.A(new_n16416_), .B(new_n16414_), .Y(new_n17049_));
  NOR3X1   g16857(.A(new_n17049_), .B(new_n16386_), .C(new_n16415_), .Y(new_n17050_));
  NOR3X1   g16858(.A(new_n16617_), .B(new_n17049_), .C(new_n16415_), .Y(new_n17051_));
  NOR2X1   g16859(.A(new_n17051_), .B(new_n16385_), .Y(new_n17052_));
  AOI21X1  g16860(.A0(new_n17050_), .A1(\asqrt[13] ), .B0(new_n17052_), .Y(new_n17053_));
  INVX1    g16861(.A(new_n17053_), .Y(new_n17054_));
  NAND3X1  g16862(.A(new_n17047_), .B(new_n17027_), .C(new_n2040_), .Y(new_n17055_));
  AOI21X1  g16863(.A0(new_n17055_), .A1(new_n17054_), .B0(new_n17048_), .Y(new_n17056_));
  OR2X1    g16864(.A(new_n17056_), .B(new_n1834_), .Y(new_n17057_));
  OR2X1    g16865(.A(new_n17045_), .B(new_n2570_), .Y(new_n17058_));
  NOR2X1   g16866(.A(new_n17017_), .B(new_n17016_), .Y(new_n17059_));
  INVX1    g16867(.A(new_n17024_), .Y(new_n17060_));
  NAND2X1  g16868(.A(new_n17011_), .B(new_n2570_), .Y(new_n17061_));
  OAI21X1  g16869(.A0(new_n17061_), .A1(new_n17059_), .B0(new_n17060_), .Y(new_n17062_));
  AOI21X1  g16870(.A0(new_n17062_), .A1(new_n17058_), .B0(new_n2263_), .Y(new_n17063_));
  AOI21X1  g16871(.A0(new_n17018_), .A1(\asqrt[45] ), .B0(\asqrt[46] ), .Y(new_n17064_));
  AOI21X1  g16872(.A0(new_n17064_), .A1(new_n17062_), .B0(new_n17032_), .Y(new_n17065_));
  NOR3X1   g16873(.A(new_n17065_), .B(new_n17063_), .C(\asqrt[47] ), .Y(new_n17066_));
  NOR2X1   g16874(.A(new_n17066_), .B(new_n17053_), .Y(new_n17067_));
  OR4X1    g16875(.A(new_n16617_), .B(new_n16418_), .C(new_n16406_), .D(new_n16401_), .Y(new_n17068_));
  OR2X1    g16876(.A(new_n16418_), .B(new_n16401_), .Y(new_n17069_));
  OAI21X1  g16877(.A0(new_n17069_), .A1(new_n16617_), .B0(new_n16406_), .Y(new_n17070_));
  AND2X1   g16878(.A(new_n17070_), .B(new_n17068_), .Y(new_n17071_));
  INVX1    g16879(.A(new_n17071_), .Y(new_n17072_));
  OAI21X1  g16880(.A0(new_n17065_), .A1(new_n17063_), .B0(\asqrt[47] ), .Y(new_n17073_));
  NAND2X1  g16881(.A(new_n17073_), .B(new_n1834_), .Y(new_n17074_));
  OAI21X1  g16882(.A0(new_n17074_), .A1(new_n17067_), .B0(new_n17072_), .Y(new_n17075_));
  AOI21X1  g16883(.A0(new_n17075_), .A1(new_n17057_), .B0(new_n1632_), .Y(new_n17076_));
  AOI21X1  g16884(.A0(new_n16463_), .A1(new_n16462_), .B0(new_n16425_), .Y(new_n17077_));
  AND2X1   g16885(.A(new_n17077_), .B(new_n16409_), .Y(new_n17078_));
  AOI22X1  g16886(.A0(new_n16463_), .A1(new_n16462_), .B0(new_n16435_), .B1(\asqrt[48] ), .Y(new_n17079_));
  AOI21X1  g16887(.A0(new_n17079_), .A1(\asqrt[13] ), .B0(new_n16424_), .Y(new_n17080_));
  AOI21X1  g16888(.A0(new_n17078_), .A1(\asqrt[13] ), .B0(new_n17080_), .Y(new_n17081_));
  OAI21X1  g16889(.A0(new_n17066_), .A1(new_n17053_), .B0(new_n17073_), .Y(new_n17082_));
  AOI21X1  g16890(.A0(new_n17082_), .A1(\asqrt[48] ), .B0(\asqrt[49] ), .Y(new_n17083_));
  AOI21X1  g16891(.A0(new_n17083_), .A1(new_n17075_), .B0(new_n17081_), .Y(new_n17084_));
  OAI21X1  g16892(.A0(new_n17084_), .A1(new_n17076_), .B0(\asqrt[50] ), .Y(new_n17085_));
  AND2X1   g16893(.A(new_n16436_), .B(new_n16428_), .Y(new_n17086_));
  NOR3X1   g16894(.A(new_n17086_), .B(new_n16466_), .C(new_n16429_), .Y(new_n17087_));
  NOR3X1   g16895(.A(new_n16617_), .B(new_n17086_), .C(new_n16429_), .Y(new_n17088_));
  NOR2X1   g16896(.A(new_n17088_), .B(new_n16434_), .Y(new_n17089_));
  AOI21X1  g16897(.A0(new_n17087_), .A1(\asqrt[13] ), .B0(new_n17089_), .Y(new_n17090_));
  NOR3X1   g16898(.A(new_n17084_), .B(new_n17076_), .C(\asqrt[50] ), .Y(new_n17091_));
  OAI21X1  g16899(.A0(new_n17091_), .A1(new_n17090_), .B0(new_n17085_), .Y(new_n17092_));
  AND2X1   g16900(.A(new_n17092_), .B(\asqrt[51] ), .Y(new_n17093_));
  OR2X1    g16901(.A(new_n17091_), .B(new_n17090_), .Y(new_n17094_));
  OR4X1    g16902(.A(new_n16617_), .B(new_n16443_), .C(new_n16470_), .D(new_n16469_), .Y(new_n17095_));
  OR2X1    g16903(.A(new_n16443_), .B(new_n16469_), .Y(new_n17096_));
  OAI21X1  g16904(.A0(new_n17096_), .A1(new_n16617_), .B0(new_n16470_), .Y(new_n17097_));
  AND2X1   g16905(.A(new_n17097_), .B(new_n17095_), .Y(new_n17098_));
  AND2X1   g16906(.A(new_n17085_), .B(new_n1277_), .Y(new_n17099_));
  AOI21X1  g16907(.A0(new_n17099_), .A1(new_n17094_), .B0(new_n17098_), .Y(new_n17100_));
  OAI21X1  g16908(.A0(new_n17100_), .A1(new_n17093_), .B0(\asqrt[52] ), .Y(new_n17101_));
  AND2X1   g16909(.A(new_n17082_), .B(\asqrt[48] ), .Y(new_n17102_));
  OR2X1    g16910(.A(new_n17066_), .B(new_n17053_), .Y(new_n17103_));
  AND2X1   g16911(.A(new_n17073_), .B(new_n1834_), .Y(new_n17104_));
  AOI21X1  g16912(.A0(new_n17104_), .A1(new_n17103_), .B0(new_n17071_), .Y(new_n17105_));
  OAI21X1  g16913(.A0(new_n17105_), .A1(new_n17102_), .B0(\asqrt[49] ), .Y(new_n17106_));
  INVX1    g16914(.A(new_n17081_), .Y(new_n17107_));
  OAI21X1  g16915(.A0(new_n17056_), .A1(new_n1834_), .B0(new_n1632_), .Y(new_n17108_));
  OAI21X1  g16916(.A0(new_n17108_), .A1(new_n17105_), .B0(new_n17107_), .Y(new_n17109_));
  AOI21X1  g16917(.A0(new_n17109_), .A1(new_n17106_), .B0(new_n1469_), .Y(new_n17110_));
  INVX1    g16918(.A(new_n17090_), .Y(new_n17111_));
  NAND3X1  g16919(.A(new_n17109_), .B(new_n17106_), .C(new_n1469_), .Y(new_n17112_));
  AOI21X1  g16920(.A0(new_n17112_), .A1(new_n17111_), .B0(new_n17110_), .Y(new_n17113_));
  OAI21X1  g16921(.A0(new_n17113_), .A1(new_n1277_), .B0(new_n1111_), .Y(new_n17114_));
  AND2X1   g16922(.A(new_n16447_), .B(new_n16446_), .Y(new_n17115_));
  NOR3X1   g16923(.A(new_n16487_), .B(new_n17115_), .C(new_n16445_), .Y(new_n17116_));
  NOR3X1   g16924(.A(new_n16617_), .B(new_n17115_), .C(new_n16445_), .Y(new_n17117_));
  NOR2X1   g16925(.A(new_n17117_), .B(new_n16452_), .Y(new_n17118_));
  AOI21X1  g16926(.A0(new_n17116_), .A1(\asqrt[13] ), .B0(new_n17118_), .Y(new_n17119_));
  INVX1    g16927(.A(new_n17119_), .Y(new_n17120_));
  OAI21X1  g16928(.A0(new_n17114_), .A1(new_n17100_), .B0(new_n17120_), .Y(new_n17121_));
  AOI21X1  g16929(.A0(new_n17121_), .A1(new_n17101_), .B0(new_n968_), .Y(new_n17122_));
  AND2X1   g16930(.A(new_n16490_), .B(new_n16488_), .Y(new_n17123_));
  NOR3X1   g16931(.A(new_n17123_), .B(new_n16460_), .C(new_n16489_), .Y(new_n17124_));
  NOR3X1   g16932(.A(new_n16617_), .B(new_n17123_), .C(new_n16489_), .Y(new_n17125_));
  NOR2X1   g16933(.A(new_n17125_), .B(new_n16459_), .Y(new_n17126_));
  AOI21X1  g16934(.A0(new_n17124_), .A1(\asqrt[13] ), .B0(new_n17126_), .Y(new_n17127_));
  INVX1    g16935(.A(new_n17127_), .Y(new_n17128_));
  NAND3X1  g16936(.A(new_n17121_), .B(new_n17101_), .C(new_n968_), .Y(new_n17129_));
  AOI21X1  g16937(.A0(new_n17129_), .A1(new_n17128_), .B0(new_n17122_), .Y(new_n17130_));
  OR2X1    g16938(.A(new_n17130_), .B(new_n902_), .Y(new_n17131_));
  OR2X1    g16939(.A(new_n17113_), .B(new_n1277_), .Y(new_n17132_));
  NOR2X1   g16940(.A(new_n17091_), .B(new_n17090_), .Y(new_n17133_));
  INVX1    g16941(.A(new_n17098_), .Y(new_n17134_));
  NAND2X1  g16942(.A(new_n17085_), .B(new_n1277_), .Y(new_n17135_));
  OAI21X1  g16943(.A0(new_n17135_), .A1(new_n17133_), .B0(new_n17134_), .Y(new_n17136_));
  AOI21X1  g16944(.A0(new_n17136_), .A1(new_n17132_), .B0(new_n1111_), .Y(new_n17137_));
  AOI21X1  g16945(.A0(new_n17092_), .A1(\asqrt[51] ), .B0(\asqrt[52] ), .Y(new_n17138_));
  AOI21X1  g16946(.A0(new_n17138_), .A1(new_n17136_), .B0(new_n17119_), .Y(new_n17139_));
  NOR3X1   g16947(.A(new_n17139_), .B(new_n17137_), .C(\asqrt[53] ), .Y(new_n17140_));
  NOR2X1   g16948(.A(new_n17140_), .B(new_n17127_), .Y(new_n17141_));
  OR4X1    g16949(.A(new_n16617_), .B(new_n16492_), .C(new_n16480_), .D(new_n16475_), .Y(new_n17142_));
  OR2X1    g16950(.A(new_n16492_), .B(new_n16475_), .Y(new_n17143_));
  OAI21X1  g16951(.A0(new_n17143_), .A1(new_n16617_), .B0(new_n16480_), .Y(new_n17144_));
  AND2X1   g16952(.A(new_n17144_), .B(new_n17142_), .Y(new_n17145_));
  INVX1    g16953(.A(new_n17145_), .Y(new_n17146_));
  OAI21X1  g16954(.A0(new_n17139_), .A1(new_n17137_), .B0(\asqrt[53] ), .Y(new_n17147_));
  NAND2X1  g16955(.A(new_n17147_), .B(new_n902_), .Y(new_n17148_));
  OAI21X1  g16956(.A0(new_n17148_), .A1(new_n17141_), .B0(new_n17146_), .Y(new_n17149_));
  AOI21X1  g16957(.A0(new_n17149_), .A1(new_n17131_), .B0(new_n697_), .Y(new_n17150_));
  AOI21X1  g16958(.A0(new_n16537_), .A1(new_n16536_), .B0(new_n16499_), .Y(new_n17151_));
  AND2X1   g16959(.A(new_n17151_), .B(new_n16483_), .Y(new_n17152_));
  AOI22X1  g16960(.A0(new_n16537_), .A1(new_n16536_), .B0(new_n16509_), .B1(\asqrt[54] ), .Y(new_n17153_));
  AOI21X1  g16961(.A0(new_n17153_), .A1(\asqrt[13] ), .B0(new_n16498_), .Y(new_n17154_));
  AOI21X1  g16962(.A0(new_n17152_), .A1(\asqrt[13] ), .B0(new_n17154_), .Y(new_n17155_));
  OAI21X1  g16963(.A0(new_n17140_), .A1(new_n17127_), .B0(new_n17147_), .Y(new_n17156_));
  AOI21X1  g16964(.A0(new_n17156_), .A1(\asqrt[54] ), .B0(\asqrt[55] ), .Y(new_n17157_));
  AOI21X1  g16965(.A0(new_n17157_), .A1(new_n17149_), .B0(new_n17155_), .Y(new_n17158_));
  OAI21X1  g16966(.A0(new_n17158_), .A1(new_n17150_), .B0(\asqrt[56] ), .Y(new_n17159_));
  AND2X1   g16967(.A(new_n16510_), .B(new_n16502_), .Y(new_n17160_));
  NOR3X1   g16968(.A(new_n17160_), .B(new_n16540_), .C(new_n16503_), .Y(new_n17161_));
  NOR3X1   g16969(.A(new_n16617_), .B(new_n17160_), .C(new_n16503_), .Y(new_n17162_));
  NOR2X1   g16970(.A(new_n17162_), .B(new_n16508_), .Y(new_n17163_));
  AOI21X1  g16971(.A0(new_n17161_), .A1(\asqrt[13] ), .B0(new_n17163_), .Y(new_n17164_));
  NOR3X1   g16972(.A(new_n17158_), .B(new_n17150_), .C(\asqrt[56] ), .Y(new_n17165_));
  OAI21X1  g16973(.A0(new_n17165_), .A1(new_n17164_), .B0(new_n17159_), .Y(new_n17166_));
  AND2X1   g16974(.A(new_n17166_), .B(\asqrt[57] ), .Y(new_n17167_));
  OR2X1    g16975(.A(new_n17165_), .B(new_n17164_), .Y(new_n17168_));
  OR4X1    g16976(.A(new_n16617_), .B(new_n16517_), .C(new_n16515_), .D(new_n16543_), .Y(new_n17169_));
  OR2X1    g16977(.A(new_n16517_), .B(new_n16543_), .Y(new_n17170_));
  OAI21X1  g16978(.A0(new_n17170_), .A1(new_n16617_), .B0(new_n16515_), .Y(new_n17171_));
  AND2X1   g16979(.A(new_n17171_), .B(new_n17169_), .Y(new_n17172_));
  AND2X1   g16980(.A(new_n17159_), .B(new_n481_), .Y(new_n17173_));
  AOI21X1  g16981(.A0(new_n17173_), .A1(new_n17168_), .B0(new_n17172_), .Y(new_n17174_));
  OAI21X1  g16982(.A0(new_n17174_), .A1(new_n17167_), .B0(\asqrt[58] ), .Y(new_n17175_));
  AND2X1   g16983(.A(new_n16526_), .B(new_n16520_), .Y(new_n17176_));
  NOR3X1   g16984(.A(new_n17176_), .B(new_n16574_), .C(new_n16519_), .Y(new_n17177_));
  NOR3X1   g16985(.A(new_n16617_), .B(new_n17176_), .C(new_n16519_), .Y(new_n17178_));
  NOR2X1   g16986(.A(new_n17178_), .B(new_n16525_), .Y(new_n17179_));
  AOI21X1  g16987(.A0(new_n17177_), .A1(\asqrt[13] ), .B0(new_n17179_), .Y(new_n17180_));
  INVX1    g16988(.A(new_n17180_), .Y(new_n17181_));
  AND2X1   g16989(.A(new_n17156_), .B(\asqrt[54] ), .Y(new_n17182_));
  OR2X1    g16990(.A(new_n17140_), .B(new_n17127_), .Y(new_n17183_));
  AND2X1   g16991(.A(new_n17147_), .B(new_n902_), .Y(new_n17184_));
  AOI21X1  g16992(.A0(new_n17184_), .A1(new_n17183_), .B0(new_n17145_), .Y(new_n17185_));
  OAI21X1  g16993(.A0(new_n17185_), .A1(new_n17182_), .B0(\asqrt[55] ), .Y(new_n17186_));
  INVX1    g16994(.A(new_n17155_), .Y(new_n17187_));
  OAI21X1  g16995(.A0(new_n17130_), .A1(new_n902_), .B0(new_n697_), .Y(new_n17188_));
  OAI21X1  g16996(.A0(new_n17188_), .A1(new_n17185_), .B0(new_n17187_), .Y(new_n17189_));
  AOI21X1  g16997(.A0(new_n17189_), .A1(new_n17186_), .B0(new_n582_), .Y(new_n17190_));
  INVX1    g16998(.A(new_n17164_), .Y(new_n17191_));
  NAND3X1  g16999(.A(new_n17189_), .B(new_n17186_), .C(new_n582_), .Y(new_n17192_));
  AOI21X1  g17000(.A0(new_n17192_), .A1(new_n17191_), .B0(new_n17190_), .Y(new_n17193_));
  OAI21X1  g17001(.A0(new_n17193_), .A1(new_n481_), .B0(new_n399_), .Y(new_n17194_));
  OAI21X1  g17002(.A0(new_n17194_), .A1(new_n17174_), .B0(new_n17181_), .Y(new_n17195_));
  AOI21X1  g17003(.A0(new_n17195_), .A1(new_n17175_), .B0(new_n328_), .Y(new_n17196_));
  AND2X1   g17004(.A(new_n16578_), .B(new_n16576_), .Y(new_n17197_));
  NOR3X1   g17005(.A(new_n17197_), .B(new_n16534_), .C(new_n16577_), .Y(new_n17198_));
  NOR3X1   g17006(.A(new_n16617_), .B(new_n17197_), .C(new_n16577_), .Y(new_n17199_));
  NOR2X1   g17007(.A(new_n17199_), .B(new_n16533_), .Y(new_n17200_));
  AOI21X1  g17008(.A0(new_n17198_), .A1(\asqrt[13] ), .B0(new_n17200_), .Y(new_n17201_));
  INVX1    g17009(.A(new_n17201_), .Y(new_n17202_));
  NAND3X1  g17010(.A(new_n17195_), .B(new_n17175_), .C(new_n328_), .Y(new_n17203_));
  AOI21X1  g17011(.A0(new_n17203_), .A1(new_n17202_), .B0(new_n17196_), .Y(new_n17204_));
  OR2X1    g17012(.A(new_n17204_), .B(new_n292_), .Y(new_n17205_));
  OR2X1    g17013(.A(new_n17193_), .B(new_n481_), .Y(new_n17206_));
  NOR2X1   g17014(.A(new_n17165_), .B(new_n17164_), .Y(new_n17207_));
  INVX1    g17015(.A(new_n17172_), .Y(new_n17208_));
  NAND2X1  g17016(.A(new_n17159_), .B(new_n481_), .Y(new_n17209_));
  OAI21X1  g17017(.A0(new_n17209_), .A1(new_n17207_), .B0(new_n17208_), .Y(new_n17210_));
  AOI21X1  g17018(.A0(new_n17210_), .A1(new_n17206_), .B0(new_n399_), .Y(new_n17211_));
  AOI21X1  g17019(.A0(new_n17166_), .A1(\asqrt[57] ), .B0(\asqrt[58] ), .Y(new_n17212_));
  AOI21X1  g17020(.A0(new_n17212_), .A1(new_n17210_), .B0(new_n17180_), .Y(new_n17213_));
  NOR3X1   g17021(.A(new_n17213_), .B(new_n17211_), .C(\asqrt[59] ), .Y(new_n17214_));
  NOR2X1   g17022(.A(new_n17214_), .B(new_n17201_), .Y(new_n17215_));
  NAND4X1  g17023(.A(\asqrt[13] ), .B(new_n16554_), .C(new_n16552_), .D(new_n16580_), .Y(new_n17216_));
  NAND2X1  g17024(.A(new_n16554_), .B(new_n16580_), .Y(new_n17217_));
  OAI21X1  g17025(.A0(new_n17217_), .A1(new_n16617_), .B0(new_n16553_), .Y(new_n17218_));
  AND2X1   g17026(.A(new_n17218_), .B(new_n17216_), .Y(new_n17219_));
  INVX1    g17027(.A(new_n17219_), .Y(new_n17220_));
  OAI21X1  g17028(.A0(new_n17213_), .A1(new_n17211_), .B0(\asqrt[59] ), .Y(new_n17221_));
  NAND2X1  g17029(.A(new_n17221_), .B(new_n292_), .Y(new_n17222_));
  OAI21X1  g17030(.A0(new_n17222_), .A1(new_n17215_), .B0(new_n17220_), .Y(new_n17223_));
  AOI21X1  g17031(.A0(new_n17223_), .A1(new_n17205_), .B0(new_n217_), .Y(new_n17224_));
  AOI21X1  g17032(.A0(new_n16626_), .A1(new_n16625_), .B0(new_n16563_), .Y(new_n17225_));
  AND2X1   g17033(.A(new_n17225_), .B(new_n16556_), .Y(new_n17226_));
  AOI22X1  g17034(.A0(new_n16626_), .A1(new_n16625_), .B0(new_n16582_), .B1(\asqrt[60] ), .Y(new_n17227_));
  AOI21X1  g17035(.A0(new_n17227_), .A1(\asqrt[13] ), .B0(new_n16562_), .Y(new_n17228_));
  AOI21X1  g17036(.A0(new_n17226_), .A1(\asqrt[13] ), .B0(new_n17228_), .Y(new_n17229_));
  OAI21X1  g17037(.A0(new_n17214_), .A1(new_n17201_), .B0(new_n17221_), .Y(new_n17230_));
  AOI21X1  g17038(.A0(new_n17230_), .A1(\asqrt[60] ), .B0(\asqrt[61] ), .Y(new_n17231_));
  AOI21X1  g17039(.A0(new_n17231_), .A1(new_n17223_), .B0(new_n17229_), .Y(new_n17232_));
  OAI21X1  g17040(.A0(new_n17232_), .A1(new_n17224_), .B0(\asqrt[62] ), .Y(new_n17233_));
  AND2X1   g17041(.A(new_n16583_), .B(new_n16565_), .Y(new_n17234_));
  NOR3X1   g17042(.A(new_n17234_), .B(new_n16629_), .C(new_n16566_), .Y(new_n17235_));
  NOR3X1   g17043(.A(new_n16617_), .B(new_n17234_), .C(new_n16566_), .Y(new_n17236_));
  NOR2X1   g17044(.A(new_n17236_), .B(new_n16571_), .Y(new_n17237_));
  AOI21X1  g17045(.A0(new_n17235_), .A1(\asqrt[13] ), .B0(new_n17237_), .Y(new_n17238_));
  NOR3X1   g17046(.A(new_n17232_), .B(new_n17224_), .C(\asqrt[62] ), .Y(new_n17239_));
  OAI21X1  g17047(.A0(new_n17239_), .A1(new_n17238_), .B0(new_n17233_), .Y(new_n17240_));
  NOR4X1   g17048(.A(new_n16617_), .B(new_n16590_), .C(new_n16633_), .D(new_n16632_), .Y(new_n17241_));
  NOR3X1   g17049(.A(new_n16617_), .B(new_n16590_), .C(new_n16632_), .Y(new_n17242_));
  NOR2X1   g17050(.A(new_n17242_), .B(new_n16589_), .Y(new_n17243_));
  NOR2X1   g17051(.A(new_n17243_), .B(new_n17241_), .Y(new_n17244_));
  INVX1    g17052(.A(new_n17244_), .Y(new_n17245_));
  AND2X1   g17053(.A(new_n16598_), .B(new_n16591_), .Y(new_n17246_));
  AOI21X1  g17054(.A0(new_n17246_), .A1(\asqrt[13] ), .B0(new_n16658_), .Y(new_n17247_));
  AND2X1   g17055(.A(new_n17247_), .B(new_n17245_), .Y(new_n17248_));
  AOI21X1  g17056(.A0(new_n17248_), .A1(new_n17240_), .B0(\asqrt[63] ), .Y(new_n17249_));
  NOR2X1   g17057(.A(new_n17239_), .B(new_n17238_), .Y(new_n17250_));
  NAND2X1  g17058(.A(new_n17244_), .B(new_n17233_), .Y(new_n17251_));
  AOI21X1  g17059(.A0(new_n16641_), .A1(new_n16637_), .B0(new_n16597_), .Y(new_n17252_));
  AOI21X1  g17060(.A0(new_n16598_), .A1(new_n16591_), .B0(new_n193_), .Y(new_n17253_));
  OAI21X1  g17061(.A0(new_n17252_), .A1(new_n16591_), .B0(new_n17253_), .Y(new_n17254_));
  INVX1    g17062(.A(new_n16596_), .Y(new_n17255_));
  NOR4X1   g17063(.A(new_n16614_), .B(new_n16608_), .C(new_n17255_), .D(new_n16593_), .Y(new_n17256_));
  OAI21X1  g17064(.A0(new_n16605_), .A1(new_n16604_), .B0(new_n17256_), .Y(new_n17257_));
  NOR2X1   g17065(.A(new_n17257_), .B(new_n16603_), .Y(new_n17258_));
  INVX1    g17066(.A(new_n17258_), .Y(new_n17259_));
  AND2X1   g17067(.A(new_n17259_), .B(new_n17254_), .Y(new_n17260_));
  OAI21X1  g17068(.A0(new_n17251_), .A1(new_n17250_), .B0(new_n17260_), .Y(new_n17261_));
  NOR2X1   g17069(.A(new_n17261_), .B(new_n17249_), .Y(new_n17262_));
  INVX1    g17070(.A(\a[24] ), .Y(new_n17263_));
  AND2X1   g17071(.A(new_n17230_), .B(\asqrt[60] ), .Y(new_n17264_));
  OR2X1    g17072(.A(new_n17214_), .B(new_n17201_), .Y(new_n17265_));
  AND2X1   g17073(.A(new_n17221_), .B(new_n292_), .Y(new_n17266_));
  AOI21X1  g17074(.A0(new_n17266_), .A1(new_n17265_), .B0(new_n17219_), .Y(new_n17267_));
  OAI21X1  g17075(.A0(new_n17267_), .A1(new_n17264_), .B0(\asqrt[61] ), .Y(new_n17268_));
  INVX1    g17076(.A(new_n17229_), .Y(new_n17269_));
  OAI21X1  g17077(.A0(new_n17204_), .A1(new_n292_), .B0(new_n217_), .Y(new_n17270_));
  OAI21X1  g17078(.A0(new_n17270_), .A1(new_n17267_), .B0(new_n17269_), .Y(new_n17271_));
  AOI21X1  g17079(.A0(new_n17271_), .A1(new_n17268_), .B0(new_n199_), .Y(new_n17272_));
  INVX1    g17080(.A(new_n17238_), .Y(new_n17273_));
  NAND3X1  g17081(.A(new_n17271_), .B(new_n17268_), .C(new_n199_), .Y(new_n17274_));
  AOI21X1  g17082(.A0(new_n17274_), .A1(new_n17273_), .B0(new_n17272_), .Y(new_n17275_));
  INVX1    g17083(.A(new_n17248_), .Y(new_n17276_));
  OAI21X1  g17084(.A0(new_n17276_), .A1(new_n17275_), .B0(new_n193_), .Y(new_n17277_));
  OR2X1    g17085(.A(new_n17239_), .B(new_n17238_), .Y(new_n17278_));
  AND2X1   g17086(.A(new_n17244_), .B(new_n17233_), .Y(new_n17279_));
  INVX1    g17087(.A(new_n17260_), .Y(new_n17280_));
  AOI21X1  g17088(.A0(new_n17279_), .A1(new_n17278_), .B0(new_n17280_), .Y(new_n17281_));
  AOI21X1  g17089(.A0(new_n17281_), .A1(new_n17277_), .B0(new_n17263_), .Y(new_n17282_));
  NOR3X1   g17090(.A(\a[24] ), .B(\a[23] ), .C(\a[22] ), .Y(new_n17283_));
  OAI21X1  g17091(.A0(new_n17283_), .A1(new_n17282_), .B0(\asqrt[13] ), .Y(new_n17284_));
  OAI21X1  g17092(.A0(new_n17261_), .A1(new_n17249_), .B0(\a[24] ), .Y(new_n17285_));
  OR2X1    g17093(.A(new_n17283_), .B(new_n16614_), .Y(new_n17286_));
  NOR4X1   g17094(.A(new_n17286_), .B(new_n16608_), .C(new_n16658_), .D(new_n16603_), .Y(new_n17287_));
  AND2X1   g17095(.A(new_n17287_), .B(new_n17285_), .Y(new_n17288_));
  INVX1    g17096(.A(\a[25] ), .Y(new_n17289_));
  AOI21X1  g17097(.A0(new_n17281_), .A1(new_n17277_), .B0(\a[24] ), .Y(new_n17290_));
  OAI21X1  g17098(.A0(new_n17261_), .A1(new_n17249_), .B0(new_n16621_), .Y(new_n17291_));
  OAI21X1  g17099(.A0(new_n17290_), .A1(new_n17289_), .B0(new_n17291_), .Y(new_n17292_));
  OAI21X1  g17100(.A0(new_n17292_), .A1(new_n17288_), .B0(new_n17284_), .Y(new_n17293_));
  AND2X1   g17101(.A(new_n17293_), .B(\asqrt[14] ), .Y(new_n17294_));
  NAND2X1  g17102(.A(new_n17287_), .B(new_n17285_), .Y(new_n17295_));
  OAI21X1  g17103(.A0(new_n17261_), .A1(new_n17249_), .B0(new_n17263_), .Y(new_n17296_));
  INVX1    g17104(.A(new_n16621_), .Y(new_n17297_));
  AOI21X1  g17105(.A0(new_n17281_), .A1(new_n17277_), .B0(new_n17297_), .Y(new_n17298_));
  AOI21X1  g17106(.A0(new_n17296_), .A1(\a[25] ), .B0(new_n17298_), .Y(new_n17299_));
  NAND2X1  g17107(.A(new_n17299_), .B(new_n17295_), .Y(new_n17300_));
  AND2X1   g17108(.A(new_n17284_), .B(new_n15990_), .Y(new_n17301_));
  INVX1    g17109(.A(new_n17254_), .Y(new_n17302_));
  NOR3X1   g17110(.A(new_n17258_), .B(new_n17302_), .C(new_n16617_), .Y(new_n17303_));
  OAI21X1  g17111(.A0(new_n17251_), .A1(new_n17250_), .B0(new_n17303_), .Y(new_n17304_));
  OR2X1    g17112(.A(new_n17304_), .B(new_n17249_), .Y(new_n17305_));
  AOI21X1  g17113(.A0(new_n17305_), .A1(new_n17291_), .B0(new_n16620_), .Y(new_n17306_));
  OAI21X1  g17114(.A0(new_n17304_), .A1(new_n17249_), .B0(new_n16620_), .Y(new_n17307_));
  NOR2X1   g17115(.A(new_n17307_), .B(new_n17298_), .Y(new_n17308_));
  NOR2X1   g17116(.A(new_n17308_), .B(new_n17306_), .Y(new_n17309_));
  AOI21X1  g17117(.A0(new_n17301_), .A1(new_n17300_), .B0(new_n17309_), .Y(new_n17310_));
  OAI21X1  g17118(.A0(new_n17310_), .A1(new_n17294_), .B0(\asqrt[15] ), .Y(new_n17311_));
  OR4X1    g17119(.A(new_n17262_), .B(new_n16654_), .C(new_n16644_), .D(new_n16656_), .Y(new_n17312_));
  NOR3X1   g17120(.A(new_n17262_), .B(new_n16644_), .C(new_n16656_), .Y(new_n17313_));
  OAI21X1  g17121(.A0(new_n17313_), .A1(new_n16648_), .B0(new_n17312_), .Y(new_n17314_));
  INVX1    g17122(.A(new_n17283_), .Y(new_n17315_));
  AOI21X1  g17123(.A0(new_n17315_), .A1(new_n17285_), .B0(new_n16617_), .Y(new_n17316_));
  AOI21X1  g17124(.A0(new_n17299_), .A1(new_n17295_), .B0(new_n17316_), .Y(new_n17317_));
  OAI21X1  g17125(.A0(new_n17317_), .A1(new_n15990_), .B0(new_n15362_), .Y(new_n17318_));
  OAI21X1  g17126(.A0(new_n17318_), .A1(new_n17310_), .B0(new_n17314_), .Y(new_n17319_));
  AOI21X1  g17127(.A0(new_n17319_), .A1(new_n17311_), .B0(new_n14754_), .Y(new_n17320_));
  AOI21X1  g17128(.A0(new_n16657_), .A1(new_n16655_), .B0(new_n16692_), .Y(new_n17321_));
  AND2X1   g17129(.A(new_n17321_), .B(new_n16689_), .Y(new_n17322_));
  OAI21X1  g17130(.A0(new_n17261_), .A1(new_n17249_), .B0(new_n17322_), .Y(new_n17323_));
  AOI22X1  g17131(.A0(new_n16657_), .A1(new_n16655_), .B0(new_n16649_), .B1(\asqrt[15] ), .Y(new_n17324_));
  OAI21X1  g17132(.A0(new_n17261_), .A1(new_n17249_), .B0(new_n17324_), .Y(new_n17325_));
  NAND2X1  g17133(.A(new_n17325_), .B(new_n16692_), .Y(new_n17326_));
  AND2X1   g17134(.A(new_n17326_), .B(new_n17323_), .Y(new_n17327_));
  INVX1    g17135(.A(new_n17327_), .Y(new_n17328_));
  NAND3X1  g17136(.A(new_n17319_), .B(new_n17311_), .C(new_n14754_), .Y(new_n17329_));
  AOI21X1  g17137(.A0(new_n17329_), .A1(new_n17328_), .B0(new_n17320_), .Y(new_n17330_));
  OR2X1    g17138(.A(new_n17330_), .B(new_n14165_), .Y(new_n17331_));
  OR2X1    g17139(.A(new_n17317_), .B(new_n15990_), .Y(new_n17332_));
  AND2X1   g17140(.A(new_n17299_), .B(new_n17295_), .Y(new_n17333_));
  OR2X1    g17141(.A(new_n17316_), .B(\asqrt[14] ), .Y(new_n17334_));
  OR2X1    g17142(.A(new_n17308_), .B(new_n17306_), .Y(new_n17335_));
  OAI21X1  g17143(.A0(new_n17334_), .A1(new_n17333_), .B0(new_n17335_), .Y(new_n17336_));
  AOI21X1  g17144(.A0(new_n17336_), .A1(new_n17332_), .B0(new_n15362_), .Y(new_n17337_));
  OR2X1    g17145(.A(new_n17313_), .B(new_n16648_), .Y(new_n17338_));
  AOI21X1  g17146(.A0(new_n17293_), .A1(\asqrt[14] ), .B0(\asqrt[15] ), .Y(new_n17339_));
  AOI22X1  g17147(.A0(new_n17339_), .A1(new_n17336_), .B0(new_n17338_), .B1(new_n17312_), .Y(new_n17340_));
  NOR3X1   g17148(.A(new_n17340_), .B(new_n17337_), .C(\asqrt[16] ), .Y(new_n17341_));
  NOR2X1   g17149(.A(new_n17341_), .B(new_n17327_), .Y(new_n17342_));
  INVX1    g17150(.A(new_n17262_), .Y(\asqrt[12] ));
  AND2X1   g17151(.A(new_n16695_), .B(new_n16693_), .Y(new_n17344_));
  NOR3X1   g17152(.A(new_n17344_), .B(new_n16673_), .C(new_n16694_), .Y(new_n17345_));
  NOR2X1   g17153(.A(new_n17344_), .B(new_n16694_), .Y(new_n17346_));
  OAI21X1  g17154(.A0(new_n17261_), .A1(new_n17249_), .B0(new_n17346_), .Y(new_n17347_));
  AOI22X1  g17155(.A0(new_n17347_), .A1(new_n16673_), .B0(new_n17345_), .B1(\asqrt[12] ), .Y(new_n17348_));
  INVX1    g17156(.A(new_n17348_), .Y(new_n17349_));
  OAI21X1  g17157(.A0(new_n17340_), .A1(new_n17337_), .B0(\asqrt[16] ), .Y(new_n17350_));
  NAND2X1  g17158(.A(new_n17350_), .B(new_n14165_), .Y(new_n17351_));
  OAI21X1  g17159(.A0(new_n17351_), .A1(new_n17342_), .B0(new_n17349_), .Y(new_n17352_));
  AOI21X1  g17160(.A0(new_n17352_), .A1(new_n17331_), .B0(new_n13571_), .Y(new_n17353_));
  NAND4X1  g17161(.A(\asqrt[12] ), .B(new_n16686_), .C(new_n16684_), .D(new_n16711_), .Y(new_n17354_));
  NOR3X1   g17162(.A(new_n17262_), .B(new_n16697_), .C(new_n16677_), .Y(new_n17355_));
  OAI21X1  g17163(.A0(new_n17355_), .A1(new_n16684_), .B0(new_n17354_), .Y(new_n17356_));
  INVX1    g17164(.A(new_n17356_), .Y(new_n17357_));
  OAI21X1  g17165(.A0(new_n17341_), .A1(new_n17327_), .B0(new_n17350_), .Y(new_n17358_));
  AOI21X1  g17166(.A0(new_n17358_), .A1(\asqrt[17] ), .B0(\asqrt[18] ), .Y(new_n17359_));
  AOI21X1  g17167(.A0(new_n17359_), .A1(new_n17352_), .B0(new_n17357_), .Y(new_n17360_));
  OAI21X1  g17168(.A0(new_n17360_), .A1(new_n17353_), .B0(\asqrt[19] ), .Y(new_n17361_));
  AND2X1   g17169(.A(new_n16740_), .B(new_n16739_), .Y(new_n17362_));
  NOR3X1   g17170(.A(new_n17362_), .B(new_n16702_), .C(new_n16738_), .Y(new_n17363_));
  NOR3X1   g17171(.A(new_n17262_), .B(new_n17362_), .C(new_n16738_), .Y(new_n17364_));
  NOR2X1   g17172(.A(new_n17364_), .B(new_n16701_), .Y(new_n17365_));
  AOI21X1  g17173(.A0(new_n17363_), .A1(\asqrt[12] ), .B0(new_n17365_), .Y(new_n17366_));
  NOR3X1   g17174(.A(new_n17360_), .B(new_n17353_), .C(\asqrt[19] ), .Y(new_n17367_));
  OAI21X1  g17175(.A0(new_n17367_), .A1(new_n17366_), .B0(new_n17361_), .Y(new_n17368_));
  AND2X1   g17176(.A(new_n17368_), .B(\asqrt[20] ), .Y(new_n17369_));
  INVX1    g17177(.A(new_n17366_), .Y(new_n17370_));
  AND2X1   g17178(.A(new_n17358_), .B(\asqrt[17] ), .Y(new_n17371_));
  OR2X1    g17179(.A(new_n17341_), .B(new_n17327_), .Y(new_n17372_));
  AND2X1   g17180(.A(new_n17350_), .B(new_n14165_), .Y(new_n17373_));
  AOI21X1  g17181(.A0(new_n17373_), .A1(new_n17372_), .B0(new_n17348_), .Y(new_n17374_));
  OAI21X1  g17182(.A0(new_n17374_), .A1(new_n17371_), .B0(\asqrt[18] ), .Y(new_n17375_));
  OAI21X1  g17183(.A0(new_n17330_), .A1(new_n14165_), .B0(new_n13571_), .Y(new_n17376_));
  OAI21X1  g17184(.A0(new_n17376_), .A1(new_n17374_), .B0(new_n17356_), .Y(new_n17377_));
  NAND3X1  g17185(.A(new_n17377_), .B(new_n17375_), .C(new_n13000_), .Y(new_n17378_));
  NAND2X1  g17186(.A(new_n17378_), .B(new_n17370_), .Y(new_n17379_));
  AND2X1   g17187(.A(new_n16713_), .B(new_n16704_), .Y(new_n17380_));
  NOR3X1   g17188(.A(new_n17380_), .B(new_n16743_), .C(new_n16705_), .Y(new_n17381_));
  NOR3X1   g17189(.A(new_n17262_), .B(new_n17380_), .C(new_n16705_), .Y(new_n17382_));
  NOR2X1   g17190(.A(new_n17382_), .B(new_n16710_), .Y(new_n17383_));
  AOI21X1  g17191(.A0(new_n17381_), .A1(\asqrt[12] ), .B0(new_n17383_), .Y(new_n17384_));
  AND2X1   g17192(.A(new_n17361_), .B(new_n12447_), .Y(new_n17385_));
  AOI21X1  g17193(.A0(new_n17385_), .A1(new_n17379_), .B0(new_n17384_), .Y(new_n17386_));
  OAI21X1  g17194(.A0(new_n17386_), .A1(new_n17369_), .B0(\asqrt[21] ), .Y(new_n17387_));
  OR4X1    g17195(.A(new_n17262_), .B(new_n16721_), .C(new_n16747_), .D(new_n16746_), .Y(new_n17388_));
  OR2X1    g17196(.A(new_n16721_), .B(new_n16746_), .Y(new_n17389_));
  OAI21X1  g17197(.A0(new_n17389_), .A1(new_n17262_), .B0(new_n16747_), .Y(new_n17390_));
  AND2X1   g17198(.A(new_n17390_), .B(new_n17388_), .Y(new_n17391_));
  INVX1    g17199(.A(new_n17391_), .Y(new_n17392_));
  AOI21X1  g17200(.A0(new_n17377_), .A1(new_n17375_), .B0(new_n13000_), .Y(new_n17393_));
  AOI21X1  g17201(.A0(new_n17378_), .A1(new_n17370_), .B0(new_n17393_), .Y(new_n17394_));
  OAI21X1  g17202(.A0(new_n17394_), .A1(new_n12447_), .B0(new_n11896_), .Y(new_n17395_));
  OAI21X1  g17203(.A0(new_n17395_), .A1(new_n17386_), .B0(new_n17392_), .Y(new_n17396_));
  AOI21X1  g17204(.A0(new_n17396_), .A1(new_n17387_), .B0(new_n11362_), .Y(new_n17397_));
  OAI21X1  g17205(.A0(new_n16765_), .A1(new_n16763_), .B0(new_n16728_), .Y(new_n17398_));
  NOR2X1   g17206(.A(new_n17398_), .B(new_n16723_), .Y(new_n17399_));
  AOI22X1  g17207(.A0(new_n16729_), .A1(new_n16724_), .B0(new_n16722_), .B1(\asqrt[21] ), .Y(new_n17400_));
  AOI21X1  g17208(.A0(new_n17400_), .A1(\asqrt[12] ), .B0(new_n16728_), .Y(new_n17401_));
  AOI21X1  g17209(.A0(new_n17399_), .A1(\asqrt[12] ), .B0(new_n17401_), .Y(new_n17402_));
  INVX1    g17210(.A(new_n17402_), .Y(new_n17403_));
  NAND3X1  g17211(.A(new_n17396_), .B(new_n17387_), .C(new_n11362_), .Y(new_n17404_));
  AOI21X1  g17212(.A0(new_n17404_), .A1(new_n17403_), .B0(new_n17397_), .Y(new_n17405_));
  OR2X1    g17213(.A(new_n17405_), .B(new_n10849_), .Y(new_n17406_));
  AND2X1   g17214(.A(new_n17404_), .B(new_n17403_), .Y(new_n17407_));
  AND2X1   g17215(.A(new_n16768_), .B(new_n16766_), .Y(new_n17408_));
  NOR3X1   g17216(.A(new_n17408_), .B(new_n16737_), .C(new_n16767_), .Y(new_n17409_));
  NOR3X1   g17217(.A(new_n17262_), .B(new_n17408_), .C(new_n16767_), .Y(new_n17410_));
  NOR2X1   g17218(.A(new_n17410_), .B(new_n16736_), .Y(new_n17411_));
  AOI21X1  g17219(.A0(new_n17409_), .A1(\asqrt[12] ), .B0(new_n17411_), .Y(new_n17412_));
  INVX1    g17220(.A(new_n17412_), .Y(new_n17413_));
  OR2X1    g17221(.A(new_n17394_), .B(new_n12447_), .Y(new_n17414_));
  AND2X1   g17222(.A(new_n17378_), .B(new_n17370_), .Y(new_n17415_));
  INVX1    g17223(.A(new_n17384_), .Y(new_n17416_));
  NAND2X1  g17224(.A(new_n17361_), .B(new_n12447_), .Y(new_n17417_));
  OAI21X1  g17225(.A0(new_n17417_), .A1(new_n17415_), .B0(new_n17416_), .Y(new_n17418_));
  AOI21X1  g17226(.A0(new_n17418_), .A1(new_n17414_), .B0(new_n11896_), .Y(new_n17419_));
  AOI21X1  g17227(.A0(new_n17368_), .A1(\asqrt[20] ), .B0(\asqrt[21] ), .Y(new_n17420_));
  AOI21X1  g17228(.A0(new_n17420_), .A1(new_n17418_), .B0(new_n17391_), .Y(new_n17421_));
  OAI21X1  g17229(.A0(new_n17421_), .A1(new_n17419_), .B0(\asqrt[22] ), .Y(new_n17422_));
  NAND2X1  g17230(.A(new_n17422_), .B(new_n10849_), .Y(new_n17423_));
  OAI21X1  g17231(.A0(new_n17423_), .A1(new_n17407_), .B0(new_n17413_), .Y(new_n17424_));
  AOI21X1  g17232(.A0(new_n17424_), .A1(new_n17406_), .B0(new_n10332_), .Y(new_n17425_));
  OR4X1    g17233(.A(new_n17262_), .B(new_n16770_), .C(new_n16758_), .D(new_n16752_), .Y(new_n17426_));
  OR2X1    g17234(.A(new_n16770_), .B(new_n16752_), .Y(new_n17427_));
  OAI21X1  g17235(.A0(new_n17427_), .A1(new_n17262_), .B0(new_n16758_), .Y(new_n17428_));
  AND2X1   g17236(.A(new_n17428_), .B(new_n17426_), .Y(new_n17429_));
  NOR3X1   g17237(.A(new_n17421_), .B(new_n17419_), .C(\asqrt[22] ), .Y(new_n17430_));
  OAI21X1  g17238(.A0(new_n17430_), .A1(new_n17402_), .B0(new_n17422_), .Y(new_n17431_));
  AOI21X1  g17239(.A0(new_n17431_), .A1(\asqrt[23] ), .B0(\asqrt[24] ), .Y(new_n17432_));
  AOI21X1  g17240(.A0(new_n17432_), .A1(new_n17424_), .B0(new_n17429_), .Y(new_n17433_));
  OAI21X1  g17241(.A0(new_n17433_), .A1(new_n17425_), .B0(\asqrt[25] ), .Y(new_n17434_));
  AND2X1   g17242(.A(new_n16801_), .B(new_n16800_), .Y(new_n17435_));
  NOR3X1   g17243(.A(new_n17435_), .B(new_n16776_), .C(new_n16799_), .Y(new_n17436_));
  NOR3X1   g17244(.A(new_n17262_), .B(new_n17435_), .C(new_n16799_), .Y(new_n17437_));
  NOR2X1   g17245(.A(new_n17437_), .B(new_n16775_), .Y(new_n17438_));
  AOI21X1  g17246(.A0(new_n17436_), .A1(\asqrt[12] ), .B0(new_n17438_), .Y(new_n17439_));
  NOR3X1   g17247(.A(new_n17433_), .B(new_n17425_), .C(\asqrt[25] ), .Y(new_n17440_));
  OAI21X1  g17248(.A0(new_n17440_), .A1(new_n17439_), .B0(new_n17434_), .Y(new_n17441_));
  AND2X1   g17249(.A(new_n17441_), .B(\asqrt[26] ), .Y(new_n17442_));
  INVX1    g17250(.A(new_n17439_), .Y(new_n17443_));
  AND2X1   g17251(.A(new_n17431_), .B(\asqrt[23] ), .Y(new_n17444_));
  NAND2X1  g17252(.A(new_n17404_), .B(new_n17403_), .Y(new_n17445_));
  AND2X1   g17253(.A(new_n17422_), .B(new_n10849_), .Y(new_n17446_));
  AOI21X1  g17254(.A0(new_n17446_), .A1(new_n17445_), .B0(new_n17412_), .Y(new_n17447_));
  OAI21X1  g17255(.A0(new_n17447_), .A1(new_n17444_), .B0(\asqrt[24] ), .Y(new_n17448_));
  INVX1    g17256(.A(new_n17429_), .Y(new_n17449_));
  OAI21X1  g17257(.A0(new_n17405_), .A1(new_n10849_), .B0(new_n10332_), .Y(new_n17450_));
  OAI21X1  g17258(.A0(new_n17450_), .A1(new_n17447_), .B0(new_n17449_), .Y(new_n17451_));
  NAND3X1  g17259(.A(new_n17451_), .B(new_n17448_), .C(new_n9833_), .Y(new_n17452_));
  NAND2X1  g17260(.A(new_n17452_), .B(new_n17443_), .Y(new_n17453_));
  AND2X1   g17261(.A(new_n16787_), .B(new_n16779_), .Y(new_n17454_));
  NOR3X1   g17262(.A(new_n17454_), .B(new_n16804_), .C(new_n16780_), .Y(new_n17455_));
  NOR3X1   g17263(.A(new_n17262_), .B(new_n17454_), .C(new_n16780_), .Y(new_n17456_));
  NOR2X1   g17264(.A(new_n17456_), .B(new_n16785_), .Y(new_n17457_));
  AOI21X1  g17265(.A0(new_n17455_), .A1(\asqrt[12] ), .B0(new_n17457_), .Y(new_n17458_));
  AND2X1   g17266(.A(new_n17434_), .B(new_n9353_), .Y(new_n17459_));
  AOI21X1  g17267(.A0(new_n17459_), .A1(new_n17453_), .B0(new_n17458_), .Y(new_n17460_));
  OAI21X1  g17268(.A0(new_n17460_), .A1(new_n17442_), .B0(\asqrt[27] ), .Y(new_n17461_));
  NAND4X1  g17269(.A(\asqrt[12] ), .B(new_n16807_), .C(new_n16794_), .D(new_n16789_), .Y(new_n17462_));
  NAND2X1  g17270(.A(new_n16807_), .B(new_n16789_), .Y(new_n17463_));
  OAI21X1  g17271(.A0(new_n17463_), .A1(new_n17262_), .B0(new_n16798_), .Y(new_n17464_));
  AND2X1   g17272(.A(new_n17464_), .B(new_n17462_), .Y(new_n17465_));
  INVX1    g17273(.A(new_n17465_), .Y(new_n17466_));
  AOI21X1  g17274(.A0(new_n17451_), .A1(new_n17448_), .B0(new_n9833_), .Y(new_n17467_));
  AOI21X1  g17275(.A0(new_n17452_), .A1(new_n17443_), .B0(new_n17467_), .Y(new_n17468_));
  OAI21X1  g17276(.A0(new_n17468_), .A1(new_n9353_), .B0(new_n8874_), .Y(new_n17469_));
  OAI21X1  g17277(.A0(new_n17469_), .A1(new_n17460_), .B0(new_n17466_), .Y(new_n17470_));
  AOI21X1  g17278(.A0(new_n17470_), .A1(new_n17461_), .B0(new_n8412_), .Y(new_n17471_));
  AOI21X1  g17279(.A0(new_n16814_), .A1(new_n16808_), .B0(new_n16852_), .Y(new_n17472_));
  AND2X1   g17280(.A(new_n17472_), .B(new_n16850_), .Y(new_n17473_));
  AOI22X1  g17281(.A0(new_n16814_), .A1(new_n16808_), .B0(new_n16796_), .B1(\asqrt[27] ), .Y(new_n17474_));
  AOI21X1  g17282(.A0(new_n17474_), .A1(\asqrt[12] ), .B0(new_n16812_), .Y(new_n17475_));
  AOI21X1  g17283(.A0(new_n17473_), .A1(\asqrt[12] ), .B0(new_n17475_), .Y(new_n17476_));
  INVX1    g17284(.A(new_n17476_), .Y(new_n17477_));
  NAND3X1  g17285(.A(new_n17470_), .B(new_n17461_), .C(new_n8412_), .Y(new_n17478_));
  AOI21X1  g17286(.A0(new_n17478_), .A1(new_n17477_), .B0(new_n17471_), .Y(new_n17479_));
  OR2X1    g17287(.A(new_n17479_), .B(new_n7970_), .Y(new_n17480_));
  AND2X1   g17288(.A(new_n17478_), .B(new_n17477_), .Y(new_n17481_));
  AND2X1   g17289(.A(new_n16856_), .B(new_n16854_), .Y(new_n17482_));
  NOR3X1   g17290(.A(new_n17482_), .B(new_n16822_), .C(new_n16855_), .Y(new_n17483_));
  NOR3X1   g17291(.A(new_n17262_), .B(new_n17482_), .C(new_n16855_), .Y(new_n17484_));
  NOR2X1   g17292(.A(new_n17484_), .B(new_n16821_), .Y(new_n17485_));
  AOI21X1  g17293(.A0(new_n17483_), .A1(\asqrt[12] ), .B0(new_n17485_), .Y(new_n17486_));
  INVX1    g17294(.A(new_n17486_), .Y(new_n17487_));
  OR2X1    g17295(.A(new_n17468_), .B(new_n9353_), .Y(new_n17488_));
  AND2X1   g17296(.A(new_n17452_), .B(new_n17443_), .Y(new_n17489_));
  INVX1    g17297(.A(new_n17458_), .Y(new_n17490_));
  NAND2X1  g17298(.A(new_n17434_), .B(new_n9353_), .Y(new_n17491_));
  OAI21X1  g17299(.A0(new_n17491_), .A1(new_n17489_), .B0(new_n17490_), .Y(new_n17492_));
  AOI21X1  g17300(.A0(new_n17492_), .A1(new_n17488_), .B0(new_n8874_), .Y(new_n17493_));
  AOI21X1  g17301(.A0(new_n17441_), .A1(\asqrt[26] ), .B0(\asqrt[27] ), .Y(new_n17494_));
  AOI21X1  g17302(.A0(new_n17494_), .A1(new_n17492_), .B0(new_n17465_), .Y(new_n17495_));
  OAI21X1  g17303(.A0(new_n17495_), .A1(new_n17493_), .B0(\asqrt[28] ), .Y(new_n17496_));
  NAND2X1  g17304(.A(new_n17496_), .B(new_n7970_), .Y(new_n17497_));
  OAI21X1  g17305(.A0(new_n17497_), .A1(new_n17481_), .B0(new_n17487_), .Y(new_n17498_));
  AOI21X1  g17306(.A0(new_n17498_), .A1(new_n17480_), .B0(new_n7527_), .Y(new_n17499_));
  NAND4X1  g17307(.A(\asqrt[12] ), .B(new_n16833_), .C(new_n16831_), .D(new_n16858_), .Y(new_n17500_));
  NAND2X1  g17308(.A(new_n16833_), .B(new_n16858_), .Y(new_n17501_));
  OAI21X1  g17309(.A0(new_n17501_), .A1(new_n17262_), .B0(new_n16832_), .Y(new_n17502_));
  AND2X1   g17310(.A(new_n17502_), .B(new_n17500_), .Y(new_n17503_));
  NOR3X1   g17311(.A(new_n17495_), .B(new_n17493_), .C(\asqrt[28] ), .Y(new_n17504_));
  OAI21X1  g17312(.A0(new_n17504_), .A1(new_n17476_), .B0(new_n17496_), .Y(new_n17505_));
  AOI21X1  g17313(.A0(new_n17505_), .A1(\asqrt[29] ), .B0(\asqrt[30] ), .Y(new_n17506_));
  AOI21X1  g17314(.A0(new_n17506_), .A1(new_n17498_), .B0(new_n17503_), .Y(new_n17507_));
  OAI21X1  g17315(.A0(new_n17507_), .A1(new_n17499_), .B0(\asqrt[31] ), .Y(new_n17508_));
  AND2X1   g17316(.A(new_n16888_), .B(new_n16887_), .Y(new_n17509_));
  NOR3X1   g17317(.A(new_n17509_), .B(new_n16841_), .C(new_n16886_), .Y(new_n17510_));
  NOR3X1   g17318(.A(new_n17262_), .B(new_n17509_), .C(new_n16886_), .Y(new_n17511_));
  NOR2X1   g17319(.A(new_n17511_), .B(new_n16840_), .Y(new_n17512_));
  AOI21X1  g17320(.A0(new_n17510_), .A1(\asqrt[12] ), .B0(new_n17512_), .Y(new_n17513_));
  NOR3X1   g17321(.A(new_n17507_), .B(new_n17499_), .C(\asqrt[31] ), .Y(new_n17514_));
  OAI21X1  g17322(.A0(new_n17514_), .A1(new_n17513_), .B0(new_n17508_), .Y(new_n17515_));
  AND2X1   g17323(.A(new_n17515_), .B(\asqrt[32] ), .Y(new_n17516_));
  INVX1    g17324(.A(new_n17513_), .Y(new_n17517_));
  AND2X1   g17325(.A(new_n17505_), .B(\asqrt[29] ), .Y(new_n17518_));
  NAND2X1  g17326(.A(new_n17478_), .B(new_n17477_), .Y(new_n17519_));
  AND2X1   g17327(.A(new_n17496_), .B(new_n7970_), .Y(new_n17520_));
  AOI21X1  g17328(.A0(new_n17520_), .A1(new_n17519_), .B0(new_n17486_), .Y(new_n17521_));
  OAI21X1  g17329(.A0(new_n17521_), .A1(new_n17518_), .B0(\asqrt[30] ), .Y(new_n17522_));
  INVX1    g17330(.A(new_n17503_), .Y(new_n17523_));
  OAI21X1  g17331(.A0(new_n17479_), .A1(new_n7970_), .B0(new_n7527_), .Y(new_n17524_));
  OAI21X1  g17332(.A0(new_n17524_), .A1(new_n17521_), .B0(new_n17523_), .Y(new_n17525_));
  NAND3X1  g17333(.A(new_n17525_), .B(new_n17522_), .C(new_n7103_), .Y(new_n17526_));
  NAND2X1  g17334(.A(new_n17526_), .B(new_n17517_), .Y(new_n17527_));
  AND2X1   g17335(.A(new_n16861_), .B(new_n16843_), .Y(new_n17528_));
  NOR3X1   g17336(.A(new_n17528_), .B(new_n16891_), .C(new_n16844_), .Y(new_n17529_));
  NOR3X1   g17337(.A(new_n17262_), .B(new_n17528_), .C(new_n16844_), .Y(new_n17530_));
  NOR2X1   g17338(.A(new_n17530_), .B(new_n16849_), .Y(new_n17531_));
  AOI21X1  g17339(.A0(new_n17529_), .A1(\asqrt[12] ), .B0(new_n17531_), .Y(new_n17532_));
  AND2X1   g17340(.A(new_n17508_), .B(new_n6699_), .Y(new_n17533_));
  AOI21X1  g17341(.A0(new_n17533_), .A1(new_n17527_), .B0(new_n17532_), .Y(new_n17534_));
  OAI21X1  g17342(.A0(new_n17534_), .A1(new_n17516_), .B0(\asqrt[33] ), .Y(new_n17535_));
  OR4X1    g17343(.A(new_n17262_), .B(new_n16869_), .C(new_n16895_), .D(new_n16894_), .Y(new_n17536_));
  OR2X1    g17344(.A(new_n16869_), .B(new_n16894_), .Y(new_n17537_));
  OAI21X1  g17345(.A0(new_n17537_), .A1(new_n17262_), .B0(new_n16895_), .Y(new_n17538_));
  AND2X1   g17346(.A(new_n17538_), .B(new_n17536_), .Y(new_n17539_));
  INVX1    g17347(.A(new_n17539_), .Y(new_n17540_));
  AOI21X1  g17348(.A0(new_n17525_), .A1(new_n17522_), .B0(new_n7103_), .Y(new_n17541_));
  AOI21X1  g17349(.A0(new_n17526_), .A1(new_n17517_), .B0(new_n17541_), .Y(new_n17542_));
  OAI21X1  g17350(.A0(new_n17542_), .A1(new_n6699_), .B0(new_n6294_), .Y(new_n17543_));
  OAI21X1  g17351(.A0(new_n17543_), .A1(new_n17534_), .B0(new_n17540_), .Y(new_n17544_));
  AOI21X1  g17352(.A0(new_n17544_), .A1(new_n17535_), .B0(new_n5941_), .Y(new_n17545_));
  AOI21X1  g17353(.A0(new_n16877_), .A1(new_n16872_), .B0(new_n16912_), .Y(new_n17546_));
  AND2X1   g17354(.A(new_n17546_), .B(new_n16910_), .Y(new_n17547_));
  AOI22X1  g17355(.A0(new_n16877_), .A1(new_n16872_), .B0(new_n16870_), .B1(\asqrt[33] ), .Y(new_n17548_));
  AOI21X1  g17356(.A0(new_n17548_), .A1(\asqrt[12] ), .B0(new_n16876_), .Y(new_n17549_));
  AOI21X1  g17357(.A0(new_n17547_), .A1(\asqrt[12] ), .B0(new_n17549_), .Y(new_n17550_));
  INVX1    g17358(.A(new_n17550_), .Y(new_n17551_));
  NAND3X1  g17359(.A(new_n17544_), .B(new_n17535_), .C(new_n5941_), .Y(new_n17552_));
  AOI21X1  g17360(.A0(new_n17552_), .A1(new_n17551_), .B0(new_n17545_), .Y(new_n17553_));
  OR2X1    g17361(.A(new_n17553_), .B(new_n5541_), .Y(new_n17554_));
  OR2X1    g17362(.A(new_n17542_), .B(new_n6699_), .Y(new_n17555_));
  AND2X1   g17363(.A(new_n17526_), .B(new_n17517_), .Y(new_n17556_));
  INVX1    g17364(.A(new_n17532_), .Y(new_n17557_));
  NAND2X1  g17365(.A(new_n17508_), .B(new_n6699_), .Y(new_n17558_));
  OAI21X1  g17366(.A0(new_n17558_), .A1(new_n17556_), .B0(new_n17557_), .Y(new_n17559_));
  AOI21X1  g17367(.A0(new_n17559_), .A1(new_n17555_), .B0(new_n6294_), .Y(new_n17560_));
  AOI21X1  g17368(.A0(new_n17515_), .A1(\asqrt[32] ), .B0(\asqrt[33] ), .Y(new_n17561_));
  AOI21X1  g17369(.A0(new_n17561_), .A1(new_n17559_), .B0(new_n17539_), .Y(new_n17562_));
  NOR3X1   g17370(.A(new_n17562_), .B(new_n17560_), .C(\asqrt[34] ), .Y(new_n17563_));
  NOR2X1   g17371(.A(new_n17563_), .B(new_n17550_), .Y(new_n17564_));
  AND2X1   g17372(.A(new_n16916_), .B(new_n16914_), .Y(new_n17565_));
  NOR3X1   g17373(.A(new_n17565_), .B(new_n16885_), .C(new_n16915_), .Y(new_n17566_));
  NOR3X1   g17374(.A(new_n17262_), .B(new_n17565_), .C(new_n16915_), .Y(new_n17567_));
  NOR2X1   g17375(.A(new_n17567_), .B(new_n16884_), .Y(new_n17568_));
  AOI21X1  g17376(.A0(new_n17566_), .A1(\asqrt[12] ), .B0(new_n17568_), .Y(new_n17569_));
  INVX1    g17377(.A(new_n17569_), .Y(new_n17570_));
  OAI21X1  g17378(.A0(new_n17562_), .A1(new_n17560_), .B0(\asqrt[34] ), .Y(new_n17571_));
  NAND2X1  g17379(.A(new_n17571_), .B(new_n5541_), .Y(new_n17572_));
  OAI21X1  g17380(.A0(new_n17572_), .A1(new_n17564_), .B0(new_n17570_), .Y(new_n17573_));
  AOI21X1  g17381(.A0(new_n17573_), .A1(new_n17554_), .B0(new_n5176_), .Y(new_n17574_));
  OR4X1    g17382(.A(new_n17262_), .B(new_n16918_), .C(new_n16906_), .D(new_n16900_), .Y(new_n17575_));
  OR2X1    g17383(.A(new_n16918_), .B(new_n16900_), .Y(new_n17576_));
  OAI21X1  g17384(.A0(new_n17576_), .A1(new_n17262_), .B0(new_n16906_), .Y(new_n17577_));
  AND2X1   g17385(.A(new_n17577_), .B(new_n17575_), .Y(new_n17578_));
  OAI21X1  g17386(.A0(new_n17563_), .A1(new_n17550_), .B0(new_n17571_), .Y(new_n17579_));
  AOI21X1  g17387(.A0(new_n17579_), .A1(\asqrt[35] ), .B0(\asqrt[36] ), .Y(new_n17580_));
  AOI21X1  g17388(.A0(new_n17580_), .A1(new_n17573_), .B0(new_n17578_), .Y(new_n17581_));
  OAI21X1  g17389(.A0(new_n17581_), .A1(new_n17574_), .B0(\asqrt[37] ), .Y(new_n17582_));
  AND2X1   g17390(.A(new_n16962_), .B(new_n16961_), .Y(new_n17583_));
  NOR3X1   g17391(.A(new_n17583_), .B(new_n16924_), .C(new_n16960_), .Y(new_n17584_));
  NOR3X1   g17392(.A(new_n17262_), .B(new_n17583_), .C(new_n16960_), .Y(new_n17585_));
  NOR2X1   g17393(.A(new_n17585_), .B(new_n16923_), .Y(new_n17586_));
  AOI21X1  g17394(.A0(new_n17584_), .A1(\asqrt[12] ), .B0(new_n17586_), .Y(new_n17587_));
  NOR3X1   g17395(.A(new_n17581_), .B(new_n17574_), .C(\asqrt[37] ), .Y(new_n17588_));
  OAI21X1  g17396(.A0(new_n17588_), .A1(new_n17587_), .B0(new_n17582_), .Y(new_n17589_));
  AND2X1   g17397(.A(new_n17589_), .B(\asqrt[38] ), .Y(new_n17590_));
  OR2X1    g17398(.A(new_n17588_), .B(new_n17587_), .Y(new_n17591_));
  AND2X1   g17399(.A(new_n16935_), .B(new_n16927_), .Y(new_n17592_));
  NOR3X1   g17400(.A(new_n17592_), .B(new_n16965_), .C(new_n16928_), .Y(new_n17593_));
  NOR3X1   g17401(.A(new_n17262_), .B(new_n17592_), .C(new_n16928_), .Y(new_n17594_));
  NOR2X1   g17402(.A(new_n17594_), .B(new_n16933_), .Y(new_n17595_));
  AOI21X1  g17403(.A0(new_n17593_), .A1(\asqrt[12] ), .B0(new_n17595_), .Y(new_n17596_));
  AND2X1   g17404(.A(new_n17582_), .B(new_n4493_), .Y(new_n17597_));
  AOI21X1  g17405(.A0(new_n17597_), .A1(new_n17591_), .B0(new_n17596_), .Y(new_n17598_));
  OAI21X1  g17406(.A0(new_n17598_), .A1(new_n17590_), .B0(\asqrt[39] ), .Y(new_n17599_));
  OR4X1    g17407(.A(new_n17262_), .B(new_n16943_), .C(new_n16969_), .D(new_n16968_), .Y(new_n17600_));
  OR2X1    g17408(.A(new_n16943_), .B(new_n16968_), .Y(new_n17601_));
  OAI21X1  g17409(.A0(new_n17601_), .A1(new_n17262_), .B0(new_n16969_), .Y(new_n17602_));
  AND2X1   g17410(.A(new_n17602_), .B(new_n17600_), .Y(new_n17603_));
  INVX1    g17411(.A(new_n17603_), .Y(new_n17604_));
  AND2X1   g17412(.A(new_n17579_), .B(\asqrt[35] ), .Y(new_n17605_));
  OR2X1    g17413(.A(new_n17563_), .B(new_n17550_), .Y(new_n17606_));
  AND2X1   g17414(.A(new_n17571_), .B(new_n5541_), .Y(new_n17607_));
  AOI21X1  g17415(.A0(new_n17607_), .A1(new_n17606_), .B0(new_n17569_), .Y(new_n17608_));
  OAI21X1  g17416(.A0(new_n17608_), .A1(new_n17605_), .B0(\asqrt[36] ), .Y(new_n17609_));
  INVX1    g17417(.A(new_n17578_), .Y(new_n17610_));
  OAI21X1  g17418(.A0(new_n17553_), .A1(new_n5541_), .B0(new_n5176_), .Y(new_n17611_));
  OAI21X1  g17419(.A0(new_n17611_), .A1(new_n17608_), .B0(new_n17610_), .Y(new_n17612_));
  AOI21X1  g17420(.A0(new_n17612_), .A1(new_n17609_), .B0(new_n4826_), .Y(new_n17613_));
  INVX1    g17421(.A(new_n17587_), .Y(new_n17614_));
  NAND3X1  g17422(.A(new_n17612_), .B(new_n17609_), .C(new_n4826_), .Y(new_n17615_));
  AOI21X1  g17423(.A0(new_n17615_), .A1(new_n17614_), .B0(new_n17613_), .Y(new_n17616_));
  OAI21X1  g17424(.A0(new_n17616_), .A1(new_n4493_), .B0(new_n4165_), .Y(new_n17617_));
  OAI21X1  g17425(.A0(new_n17617_), .A1(new_n17598_), .B0(new_n17604_), .Y(new_n17618_));
  AOI21X1  g17426(.A0(new_n17618_), .A1(new_n17599_), .B0(new_n3863_), .Y(new_n17619_));
  AOI21X1  g17427(.A0(new_n16951_), .A1(new_n16946_), .B0(new_n16986_), .Y(new_n17620_));
  AND2X1   g17428(.A(new_n17620_), .B(new_n16984_), .Y(new_n17621_));
  AOI22X1  g17429(.A0(new_n16951_), .A1(new_n16946_), .B0(new_n16944_), .B1(\asqrt[39] ), .Y(new_n17622_));
  AOI21X1  g17430(.A0(new_n17622_), .A1(\asqrt[12] ), .B0(new_n16950_), .Y(new_n17623_));
  AOI21X1  g17431(.A0(new_n17621_), .A1(\asqrt[12] ), .B0(new_n17623_), .Y(new_n17624_));
  INVX1    g17432(.A(new_n17624_), .Y(new_n17625_));
  NAND3X1  g17433(.A(new_n17618_), .B(new_n17599_), .C(new_n3863_), .Y(new_n17626_));
  AOI21X1  g17434(.A0(new_n17626_), .A1(new_n17625_), .B0(new_n17619_), .Y(new_n17627_));
  OR2X1    g17435(.A(new_n17627_), .B(new_n3564_), .Y(new_n17628_));
  OR2X1    g17436(.A(new_n17616_), .B(new_n4493_), .Y(new_n17629_));
  NOR2X1   g17437(.A(new_n17588_), .B(new_n17587_), .Y(new_n17630_));
  INVX1    g17438(.A(new_n17596_), .Y(new_n17631_));
  NAND2X1  g17439(.A(new_n17582_), .B(new_n4493_), .Y(new_n17632_));
  OAI21X1  g17440(.A0(new_n17632_), .A1(new_n17630_), .B0(new_n17631_), .Y(new_n17633_));
  AOI21X1  g17441(.A0(new_n17633_), .A1(new_n17629_), .B0(new_n4165_), .Y(new_n17634_));
  AOI21X1  g17442(.A0(new_n17589_), .A1(\asqrt[38] ), .B0(\asqrt[39] ), .Y(new_n17635_));
  AOI21X1  g17443(.A0(new_n17635_), .A1(new_n17633_), .B0(new_n17603_), .Y(new_n17636_));
  NOR3X1   g17444(.A(new_n17636_), .B(new_n17634_), .C(\asqrt[40] ), .Y(new_n17637_));
  NOR2X1   g17445(.A(new_n17637_), .B(new_n17624_), .Y(new_n17638_));
  AND2X1   g17446(.A(new_n16990_), .B(new_n16988_), .Y(new_n17639_));
  NOR3X1   g17447(.A(new_n17639_), .B(new_n16959_), .C(new_n16989_), .Y(new_n17640_));
  NOR3X1   g17448(.A(new_n17262_), .B(new_n17639_), .C(new_n16989_), .Y(new_n17641_));
  NOR2X1   g17449(.A(new_n17641_), .B(new_n16958_), .Y(new_n17642_));
  AOI21X1  g17450(.A0(new_n17640_), .A1(\asqrt[12] ), .B0(new_n17642_), .Y(new_n17643_));
  INVX1    g17451(.A(new_n17643_), .Y(new_n17644_));
  OAI21X1  g17452(.A0(new_n17636_), .A1(new_n17634_), .B0(\asqrt[40] ), .Y(new_n17645_));
  NAND2X1  g17453(.A(new_n17645_), .B(new_n3564_), .Y(new_n17646_));
  OAI21X1  g17454(.A0(new_n17646_), .A1(new_n17638_), .B0(new_n17644_), .Y(new_n17647_));
  AOI21X1  g17455(.A0(new_n17647_), .A1(new_n17628_), .B0(new_n3276_), .Y(new_n17648_));
  OR4X1    g17456(.A(new_n17262_), .B(new_n16992_), .C(new_n16980_), .D(new_n16974_), .Y(new_n17649_));
  OR2X1    g17457(.A(new_n16992_), .B(new_n16974_), .Y(new_n17650_));
  OAI21X1  g17458(.A0(new_n17650_), .A1(new_n17262_), .B0(new_n16980_), .Y(new_n17651_));
  AND2X1   g17459(.A(new_n17651_), .B(new_n17649_), .Y(new_n17652_));
  OAI21X1  g17460(.A0(new_n17637_), .A1(new_n17624_), .B0(new_n17645_), .Y(new_n17653_));
  AOI21X1  g17461(.A0(new_n17653_), .A1(\asqrt[41] ), .B0(\asqrt[42] ), .Y(new_n17654_));
  AOI21X1  g17462(.A0(new_n17654_), .A1(new_n17647_), .B0(new_n17652_), .Y(new_n17655_));
  OAI21X1  g17463(.A0(new_n17655_), .A1(new_n17648_), .B0(\asqrt[43] ), .Y(new_n17656_));
  AND2X1   g17464(.A(new_n17036_), .B(new_n17035_), .Y(new_n17657_));
  NOR3X1   g17465(.A(new_n17657_), .B(new_n16998_), .C(new_n17034_), .Y(new_n17658_));
  NOR3X1   g17466(.A(new_n17262_), .B(new_n17657_), .C(new_n17034_), .Y(new_n17659_));
  NOR2X1   g17467(.A(new_n17659_), .B(new_n16997_), .Y(new_n17660_));
  AOI21X1  g17468(.A0(new_n17658_), .A1(\asqrt[12] ), .B0(new_n17660_), .Y(new_n17661_));
  NOR3X1   g17469(.A(new_n17655_), .B(new_n17648_), .C(\asqrt[43] ), .Y(new_n17662_));
  OAI21X1  g17470(.A0(new_n17662_), .A1(new_n17661_), .B0(new_n17656_), .Y(new_n17663_));
  AND2X1   g17471(.A(new_n17663_), .B(\asqrt[44] ), .Y(new_n17664_));
  OR2X1    g17472(.A(new_n17662_), .B(new_n17661_), .Y(new_n17665_));
  AND2X1   g17473(.A(new_n17009_), .B(new_n17001_), .Y(new_n17666_));
  NOR3X1   g17474(.A(new_n17666_), .B(new_n17039_), .C(new_n17002_), .Y(new_n17667_));
  NOR3X1   g17475(.A(new_n17262_), .B(new_n17666_), .C(new_n17002_), .Y(new_n17668_));
  NOR2X1   g17476(.A(new_n17668_), .B(new_n17007_), .Y(new_n17669_));
  AOI21X1  g17477(.A0(new_n17667_), .A1(\asqrt[12] ), .B0(new_n17669_), .Y(new_n17670_));
  AND2X1   g17478(.A(new_n17656_), .B(new_n2769_), .Y(new_n17671_));
  AOI21X1  g17479(.A0(new_n17671_), .A1(new_n17665_), .B0(new_n17670_), .Y(new_n17672_));
  OAI21X1  g17480(.A0(new_n17672_), .A1(new_n17664_), .B0(\asqrt[45] ), .Y(new_n17673_));
  OR4X1    g17481(.A(new_n17262_), .B(new_n17017_), .C(new_n17043_), .D(new_n17042_), .Y(new_n17674_));
  OR2X1    g17482(.A(new_n17017_), .B(new_n17042_), .Y(new_n17675_));
  OAI21X1  g17483(.A0(new_n17675_), .A1(new_n17262_), .B0(new_n17043_), .Y(new_n17676_));
  AND2X1   g17484(.A(new_n17676_), .B(new_n17674_), .Y(new_n17677_));
  INVX1    g17485(.A(new_n17677_), .Y(new_n17678_));
  AND2X1   g17486(.A(new_n17653_), .B(\asqrt[41] ), .Y(new_n17679_));
  OR2X1    g17487(.A(new_n17637_), .B(new_n17624_), .Y(new_n17680_));
  AND2X1   g17488(.A(new_n17645_), .B(new_n3564_), .Y(new_n17681_));
  AOI21X1  g17489(.A0(new_n17681_), .A1(new_n17680_), .B0(new_n17643_), .Y(new_n17682_));
  OAI21X1  g17490(.A0(new_n17682_), .A1(new_n17679_), .B0(\asqrt[42] ), .Y(new_n17683_));
  INVX1    g17491(.A(new_n17652_), .Y(new_n17684_));
  OAI21X1  g17492(.A0(new_n17627_), .A1(new_n3564_), .B0(new_n3276_), .Y(new_n17685_));
  OAI21X1  g17493(.A0(new_n17685_), .A1(new_n17682_), .B0(new_n17684_), .Y(new_n17686_));
  AOI21X1  g17494(.A0(new_n17686_), .A1(new_n17683_), .B0(new_n3008_), .Y(new_n17687_));
  INVX1    g17495(.A(new_n17661_), .Y(new_n17688_));
  NAND3X1  g17496(.A(new_n17686_), .B(new_n17683_), .C(new_n3008_), .Y(new_n17689_));
  AOI21X1  g17497(.A0(new_n17689_), .A1(new_n17688_), .B0(new_n17687_), .Y(new_n17690_));
  OAI21X1  g17498(.A0(new_n17690_), .A1(new_n2769_), .B0(new_n2570_), .Y(new_n17691_));
  OAI21X1  g17499(.A0(new_n17691_), .A1(new_n17672_), .B0(new_n17678_), .Y(new_n17692_));
  AOI21X1  g17500(.A0(new_n17692_), .A1(new_n17673_), .B0(new_n2263_), .Y(new_n17693_));
  AOI21X1  g17501(.A0(new_n17025_), .A1(new_n17020_), .B0(new_n17060_), .Y(new_n17694_));
  AND2X1   g17502(.A(new_n17694_), .B(new_n17058_), .Y(new_n17695_));
  AOI22X1  g17503(.A0(new_n17025_), .A1(new_n17020_), .B0(new_n17018_), .B1(\asqrt[45] ), .Y(new_n17696_));
  AOI21X1  g17504(.A0(new_n17696_), .A1(\asqrt[12] ), .B0(new_n17024_), .Y(new_n17697_));
  AOI21X1  g17505(.A0(new_n17695_), .A1(\asqrt[12] ), .B0(new_n17697_), .Y(new_n17698_));
  INVX1    g17506(.A(new_n17698_), .Y(new_n17699_));
  NAND3X1  g17507(.A(new_n17692_), .B(new_n17673_), .C(new_n2263_), .Y(new_n17700_));
  AOI21X1  g17508(.A0(new_n17700_), .A1(new_n17699_), .B0(new_n17693_), .Y(new_n17701_));
  OR2X1    g17509(.A(new_n17701_), .B(new_n2040_), .Y(new_n17702_));
  OR2X1    g17510(.A(new_n17690_), .B(new_n2769_), .Y(new_n17703_));
  NOR2X1   g17511(.A(new_n17662_), .B(new_n17661_), .Y(new_n17704_));
  INVX1    g17512(.A(new_n17670_), .Y(new_n17705_));
  NAND2X1  g17513(.A(new_n17656_), .B(new_n2769_), .Y(new_n17706_));
  OAI21X1  g17514(.A0(new_n17706_), .A1(new_n17704_), .B0(new_n17705_), .Y(new_n17707_));
  AOI21X1  g17515(.A0(new_n17707_), .A1(new_n17703_), .B0(new_n2570_), .Y(new_n17708_));
  AOI21X1  g17516(.A0(new_n17663_), .A1(\asqrt[44] ), .B0(\asqrt[45] ), .Y(new_n17709_));
  AOI21X1  g17517(.A0(new_n17709_), .A1(new_n17707_), .B0(new_n17677_), .Y(new_n17710_));
  NOR3X1   g17518(.A(new_n17710_), .B(new_n17708_), .C(\asqrt[46] ), .Y(new_n17711_));
  NOR2X1   g17519(.A(new_n17711_), .B(new_n17698_), .Y(new_n17712_));
  AND2X1   g17520(.A(new_n17064_), .B(new_n17062_), .Y(new_n17713_));
  NOR3X1   g17521(.A(new_n17713_), .B(new_n17033_), .C(new_n17063_), .Y(new_n17714_));
  NOR3X1   g17522(.A(new_n17262_), .B(new_n17713_), .C(new_n17063_), .Y(new_n17715_));
  NOR2X1   g17523(.A(new_n17715_), .B(new_n17032_), .Y(new_n17716_));
  AOI21X1  g17524(.A0(new_n17714_), .A1(\asqrt[12] ), .B0(new_n17716_), .Y(new_n17717_));
  INVX1    g17525(.A(new_n17717_), .Y(new_n17718_));
  OAI21X1  g17526(.A0(new_n17710_), .A1(new_n17708_), .B0(\asqrt[46] ), .Y(new_n17719_));
  NAND2X1  g17527(.A(new_n17719_), .B(new_n2040_), .Y(new_n17720_));
  OAI21X1  g17528(.A0(new_n17720_), .A1(new_n17712_), .B0(new_n17718_), .Y(new_n17721_));
  AOI21X1  g17529(.A0(new_n17721_), .A1(new_n17702_), .B0(new_n1834_), .Y(new_n17722_));
  OR4X1    g17530(.A(new_n17262_), .B(new_n17066_), .C(new_n17054_), .D(new_n17048_), .Y(new_n17723_));
  OR2X1    g17531(.A(new_n17066_), .B(new_n17048_), .Y(new_n17724_));
  OAI21X1  g17532(.A0(new_n17724_), .A1(new_n17262_), .B0(new_n17054_), .Y(new_n17725_));
  AND2X1   g17533(.A(new_n17725_), .B(new_n17723_), .Y(new_n17726_));
  OAI21X1  g17534(.A0(new_n17711_), .A1(new_n17698_), .B0(new_n17719_), .Y(new_n17727_));
  AOI21X1  g17535(.A0(new_n17727_), .A1(\asqrt[47] ), .B0(\asqrt[48] ), .Y(new_n17728_));
  AOI21X1  g17536(.A0(new_n17728_), .A1(new_n17721_), .B0(new_n17726_), .Y(new_n17729_));
  OAI21X1  g17537(.A0(new_n17729_), .A1(new_n17722_), .B0(\asqrt[49] ), .Y(new_n17730_));
  AND2X1   g17538(.A(new_n17104_), .B(new_n17103_), .Y(new_n17731_));
  NOR3X1   g17539(.A(new_n17731_), .B(new_n17072_), .C(new_n17102_), .Y(new_n17732_));
  NOR3X1   g17540(.A(new_n17262_), .B(new_n17731_), .C(new_n17102_), .Y(new_n17733_));
  NOR2X1   g17541(.A(new_n17733_), .B(new_n17071_), .Y(new_n17734_));
  AOI21X1  g17542(.A0(new_n17732_), .A1(\asqrt[12] ), .B0(new_n17734_), .Y(new_n17735_));
  NOR3X1   g17543(.A(new_n17729_), .B(new_n17722_), .C(\asqrt[49] ), .Y(new_n17736_));
  OAI21X1  g17544(.A0(new_n17736_), .A1(new_n17735_), .B0(new_n17730_), .Y(new_n17737_));
  AND2X1   g17545(.A(new_n17737_), .B(\asqrt[50] ), .Y(new_n17738_));
  OR2X1    g17546(.A(new_n17736_), .B(new_n17735_), .Y(new_n17739_));
  AND2X1   g17547(.A(new_n17083_), .B(new_n17075_), .Y(new_n17740_));
  NOR3X1   g17548(.A(new_n17740_), .B(new_n17107_), .C(new_n17076_), .Y(new_n17741_));
  NOR3X1   g17549(.A(new_n17262_), .B(new_n17740_), .C(new_n17076_), .Y(new_n17742_));
  NOR2X1   g17550(.A(new_n17742_), .B(new_n17081_), .Y(new_n17743_));
  AOI21X1  g17551(.A0(new_n17741_), .A1(\asqrt[12] ), .B0(new_n17743_), .Y(new_n17744_));
  AND2X1   g17552(.A(new_n17730_), .B(new_n1469_), .Y(new_n17745_));
  AOI21X1  g17553(.A0(new_n17745_), .A1(new_n17739_), .B0(new_n17744_), .Y(new_n17746_));
  OAI21X1  g17554(.A0(new_n17746_), .A1(new_n17738_), .B0(\asqrt[51] ), .Y(new_n17747_));
  OR4X1    g17555(.A(new_n17262_), .B(new_n17091_), .C(new_n17111_), .D(new_n17110_), .Y(new_n17748_));
  OR2X1    g17556(.A(new_n17091_), .B(new_n17110_), .Y(new_n17749_));
  OAI21X1  g17557(.A0(new_n17749_), .A1(new_n17262_), .B0(new_n17111_), .Y(new_n17750_));
  AND2X1   g17558(.A(new_n17750_), .B(new_n17748_), .Y(new_n17751_));
  INVX1    g17559(.A(new_n17751_), .Y(new_n17752_));
  AND2X1   g17560(.A(new_n17727_), .B(\asqrt[47] ), .Y(new_n17753_));
  OR2X1    g17561(.A(new_n17711_), .B(new_n17698_), .Y(new_n17754_));
  AND2X1   g17562(.A(new_n17719_), .B(new_n2040_), .Y(new_n17755_));
  AOI21X1  g17563(.A0(new_n17755_), .A1(new_n17754_), .B0(new_n17717_), .Y(new_n17756_));
  OAI21X1  g17564(.A0(new_n17756_), .A1(new_n17753_), .B0(\asqrt[48] ), .Y(new_n17757_));
  INVX1    g17565(.A(new_n17726_), .Y(new_n17758_));
  OAI21X1  g17566(.A0(new_n17701_), .A1(new_n2040_), .B0(new_n1834_), .Y(new_n17759_));
  OAI21X1  g17567(.A0(new_n17759_), .A1(new_n17756_), .B0(new_n17758_), .Y(new_n17760_));
  AOI21X1  g17568(.A0(new_n17760_), .A1(new_n17757_), .B0(new_n1632_), .Y(new_n17761_));
  INVX1    g17569(.A(new_n17735_), .Y(new_n17762_));
  NAND3X1  g17570(.A(new_n17760_), .B(new_n17757_), .C(new_n1632_), .Y(new_n17763_));
  AOI21X1  g17571(.A0(new_n17763_), .A1(new_n17762_), .B0(new_n17761_), .Y(new_n17764_));
  OAI21X1  g17572(.A0(new_n17764_), .A1(new_n1469_), .B0(new_n1277_), .Y(new_n17765_));
  OAI21X1  g17573(.A0(new_n17765_), .A1(new_n17746_), .B0(new_n17752_), .Y(new_n17766_));
  AOI21X1  g17574(.A0(new_n17766_), .A1(new_n17747_), .B0(new_n1111_), .Y(new_n17767_));
  AOI21X1  g17575(.A0(new_n17099_), .A1(new_n17094_), .B0(new_n17134_), .Y(new_n17768_));
  AND2X1   g17576(.A(new_n17768_), .B(new_n17132_), .Y(new_n17769_));
  AOI22X1  g17577(.A0(new_n17099_), .A1(new_n17094_), .B0(new_n17092_), .B1(\asqrt[51] ), .Y(new_n17770_));
  AOI21X1  g17578(.A0(new_n17770_), .A1(\asqrt[12] ), .B0(new_n17098_), .Y(new_n17771_));
  AOI21X1  g17579(.A0(new_n17769_), .A1(\asqrt[12] ), .B0(new_n17771_), .Y(new_n17772_));
  INVX1    g17580(.A(new_n17772_), .Y(new_n17773_));
  NAND3X1  g17581(.A(new_n17766_), .B(new_n17747_), .C(new_n1111_), .Y(new_n17774_));
  AOI21X1  g17582(.A0(new_n17774_), .A1(new_n17773_), .B0(new_n17767_), .Y(new_n17775_));
  OR2X1    g17583(.A(new_n17775_), .B(new_n968_), .Y(new_n17776_));
  OR2X1    g17584(.A(new_n17764_), .B(new_n1469_), .Y(new_n17777_));
  NOR2X1   g17585(.A(new_n17736_), .B(new_n17735_), .Y(new_n17778_));
  INVX1    g17586(.A(new_n17744_), .Y(new_n17779_));
  NAND2X1  g17587(.A(new_n17730_), .B(new_n1469_), .Y(new_n17780_));
  OAI21X1  g17588(.A0(new_n17780_), .A1(new_n17778_), .B0(new_n17779_), .Y(new_n17781_));
  AOI21X1  g17589(.A0(new_n17781_), .A1(new_n17777_), .B0(new_n1277_), .Y(new_n17782_));
  AOI21X1  g17590(.A0(new_n17737_), .A1(\asqrt[50] ), .B0(\asqrt[51] ), .Y(new_n17783_));
  AOI21X1  g17591(.A0(new_n17783_), .A1(new_n17781_), .B0(new_n17751_), .Y(new_n17784_));
  NOR3X1   g17592(.A(new_n17784_), .B(new_n17782_), .C(\asqrt[52] ), .Y(new_n17785_));
  NOR2X1   g17593(.A(new_n17785_), .B(new_n17772_), .Y(new_n17786_));
  OAI21X1  g17594(.A0(new_n17784_), .A1(new_n17782_), .B0(\asqrt[52] ), .Y(new_n17787_));
  NAND2X1  g17595(.A(new_n17787_), .B(new_n968_), .Y(new_n17788_));
  AND2X1   g17596(.A(new_n17138_), .B(new_n17136_), .Y(new_n17789_));
  NOR3X1   g17597(.A(new_n17120_), .B(new_n17789_), .C(new_n17137_), .Y(new_n17790_));
  NOR3X1   g17598(.A(new_n17262_), .B(new_n17789_), .C(new_n17137_), .Y(new_n17791_));
  NOR2X1   g17599(.A(new_n17791_), .B(new_n17119_), .Y(new_n17792_));
  AOI21X1  g17600(.A0(new_n17790_), .A1(\asqrt[12] ), .B0(new_n17792_), .Y(new_n17793_));
  INVX1    g17601(.A(new_n17793_), .Y(new_n17794_));
  OAI21X1  g17602(.A0(new_n17788_), .A1(new_n17786_), .B0(new_n17794_), .Y(new_n17795_));
  AOI21X1  g17603(.A0(new_n17795_), .A1(new_n17776_), .B0(new_n902_), .Y(new_n17796_));
  OR4X1    g17604(.A(new_n17262_), .B(new_n17140_), .C(new_n17128_), .D(new_n17122_), .Y(new_n17797_));
  OR2X1    g17605(.A(new_n17140_), .B(new_n17122_), .Y(new_n17798_));
  OAI21X1  g17606(.A0(new_n17798_), .A1(new_n17262_), .B0(new_n17128_), .Y(new_n17799_));
  AND2X1   g17607(.A(new_n17799_), .B(new_n17797_), .Y(new_n17800_));
  OAI21X1  g17608(.A0(new_n17785_), .A1(new_n17772_), .B0(new_n17787_), .Y(new_n17801_));
  AOI21X1  g17609(.A0(new_n17801_), .A1(\asqrt[53] ), .B0(\asqrt[54] ), .Y(new_n17802_));
  AOI21X1  g17610(.A0(new_n17802_), .A1(new_n17795_), .B0(new_n17800_), .Y(new_n17803_));
  OAI21X1  g17611(.A0(new_n17803_), .A1(new_n17796_), .B0(\asqrt[55] ), .Y(new_n17804_));
  AND2X1   g17612(.A(new_n17184_), .B(new_n17183_), .Y(new_n17805_));
  NOR3X1   g17613(.A(new_n17805_), .B(new_n17146_), .C(new_n17182_), .Y(new_n17806_));
  NOR3X1   g17614(.A(new_n17262_), .B(new_n17805_), .C(new_n17182_), .Y(new_n17807_));
  NOR2X1   g17615(.A(new_n17807_), .B(new_n17145_), .Y(new_n17808_));
  AOI21X1  g17616(.A0(new_n17806_), .A1(\asqrt[12] ), .B0(new_n17808_), .Y(new_n17809_));
  NOR3X1   g17617(.A(new_n17803_), .B(new_n17796_), .C(\asqrt[55] ), .Y(new_n17810_));
  OAI21X1  g17618(.A0(new_n17810_), .A1(new_n17809_), .B0(new_n17804_), .Y(new_n17811_));
  AND2X1   g17619(.A(new_n17811_), .B(\asqrt[56] ), .Y(new_n17812_));
  OR2X1    g17620(.A(new_n17810_), .B(new_n17809_), .Y(new_n17813_));
  AND2X1   g17621(.A(new_n17157_), .B(new_n17149_), .Y(new_n17814_));
  NOR3X1   g17622(.A(new_n17814_), .B(new_n17187_), .C(new_n17150_), .Y(new_n17815_));
  NOR3X1   g17623(.A(new_n17262_), .B(new_n17814_), .C(new_n17150_), .Y(new_n17816_));
  NOR2X1   g17624(.A(new_n17816_), .B(new_n17155_), .Y(new_n17817_));
  AOI21X1  g17625(.A0(new_n17815_), .A1(\asqrt[12] ), .B0(new_n17817_), .Y(new_n17818_));
  AND2X1   g17626(.A(new_n17804_), .B(new_n582_), .Y(new_n17819_));
  AOI21X1  g17627(.A0(new_n17819_), .A1(new_n17813_), .B0(new_n17818_), .Y(new_n17820_));
  OAI21X1  g17628(.A0(new_n17820_), .A1(new_n17812_), .B0(\asqrt[57] ), .Y(new_n17821_));
  OR4X1    g17629(.A(new_n17262_), .B(new_n17165_), .C(new_n17191_), .D(new_n17190_), .Y(new_n17822_));
  OR2X1    g17630(.A(new_n17165_), .B(new_n17190_), .Y(new_n17823_));
  OAI21X1  g17631(.A0(new_n17823_), .A1(new_n17262_), .B0(new_n17191_), .Y(new_n17824_));
  AND2X1   g17632(.A(new_n17824_), .B(new_n17822_), .Y(new_n17825_));
  INVX1    g17633(.A(new_n17825_), .Y(new_n17826_));
  AND2X1   g17634(.A(new_n17801_), .B(\asqrt[53] ), .Y(new_n17827_));
  OR2X1    g17635(.A(new_n17785_), .B(new_n17772_), .Y(new_n17828_));
  AND2X1   g17636(.A(new_n17787_), .B(new_n968_), .Y(new_n17829_));
  AOI21X1  g17637(.A0(new_n17829_), .A1(new_n17828_), .B0(new_n17793_), .Y(new_n17830_));
  OAI21X1  g17638(.A0(new_n17830_), .A1(new_n17827_), .B0(\asqrt[54] ), .Y(new_n17831_));
  INVX1    g17639(.A(new_n17800_), .Y(new_n17832_));
  OAI21X1  g17640(.A0(new_n17775_), .A1(new_n968_), .B0(new_n902_), .Y(new_n17833_));
  OAI21X1  g17641(.A0(new_n17833_), .A1(new_n17830_), .B0(new_n17832_), .Y(new_n17834_));
  AOI21X1  g17642(.A0(new_n17834_), .A1(new_n17831_), .B0(new_n697_), .Y(new_n17835_));
  INVX1    g17643(.A(new_n17809_), .Y(new_n17836_));
  NAND3X1  g17644(.A(new_n17834_), .B(new_n17831_), .C(new_n697_), .Y(new_n17837_));
  AOI21X1  g17645(.A0(new_n17837_), .A1(new_n17836_), .B0(new_n17835_), .Y(new_n17838_));
  OAI21X1  g17646(.A0(new_n17838_), .A1(new_n582_), .B0(new_n481_), .Y(new_n17839_));
  OAI21X1  g17647(.A0(new_n17839_), .A1(new_n17820_), .B0(new_n17826_), .Y(new_n17840_));
  AOI21X1  g17648(.A0(new_n17840_), .A1(new_n17821_), .B0(new_n399_), .Y(new_n17841_));
  AOI21X1  g17649(.A0(new_n17173_), .A1(new_n17168_), .B0(new_n17208_), .Y(new_n17842_));
  AND2X1   g17650(.A(new_n17842_), .B(new_n17206_), .Y(new_n17843_));
  AOI22X1  g17651(.A0(new_n17173_), .A1(new_n17168_), .B0(new_n17166_), .B1(\asqrt[57] ), .Y(new_n17844_));
  AOI21X1  g17652(.A0(new_n17844_), .A1(\asqrt[12] ), .B0(new_n17172_), .Y(new_n17845_));
  AOI21X1  g17653(.A0(new_n17843_), .A1(\asqrt[12] ), .B0(new_n17845_), .Y(new_n17846_));
  INVX1    g17654(.A(new_n17846_), .Y(new_n17847_));
  NAND3X1  g17655(.A(new_n17840_), .B(new_n17821_), .C(new_n399_), .Y(new_n17848_));
  AOI21X1  g17656(.A0(new_n17848_), .A1(new_n17847_), .B0(new_n17841_), .Y(new_n17849_));
  OR2X1    g17657(.A(new_n17849_), .B(new_n328_), .Y(new_n17850_));
  OR2X1    g17658(.A(new_n17838_), .B(new_n582_), .Y(new_n17851_));
  NOR2X1   g17659(.A(new_n17810_), .B(new_n17809_), .Y(new_n17852_));
  INVX1    g17660(.A(new_n17818_), .Y(new_n17853_));
  NAND2X1  g17661(.A(new_n17804_), .B(new_n582_), .Y(new_n17854_));
  OAI21X1  g17662(.A0(new_n17854_), .A1(new_n17852_), .B0(new_n17853_), .Y(new_n17855_));
  AOI21X1  g17663(.A0(new_n17855_), .A1(new_n17851_), .B0(new_n481_), .Y(new_n17856_));
  AOI21X1  g17664(.A0(new_n17811_), .A1(\asqrt[56] ), .B0(\asqrt[57] ), .Y(new_n17857_));
  AOI21X1  g17665(.A0(new_n17857_), .A1(new_n17855_), .B0(new_n17825_), .Y(new_n17858_));
  NOR3X1   g17666(.A(new_n17858_), .B(new_n17856_), .C(\asqrt[58] ), .Y(new_n17859_));
  NOR2X1   g17667(.A(new_n17859_), .B(new_n17846_), .Y(new_n17860_));
  AND2X1   g17668(.A(new_n17212_), .B(new_n17210_), .Y(new_n17861_));
  NOR3X1   g17669(.A(new_n17861_), .B(new_n17181_), .C(new_n17211_), .Y(new_n17862_));
  NOR3X1   g17670(.A(new_n17262_), .B(new_n17861_), .C(new_n17211_), .Y(new_n17863_));
  NOR2X1   g17671(.A(new_n17863_), .B(new_n17180_), .Y(new_n17864_));
  AOI21X1  g17672(.A0(new_n17862_), .A1(\asqrt[12] ), .B0(new_n17864_), .Y(new_n17865_));
  INVX1    g17673(.A(new_n17865_), .Y(new_n17866_));
  OAI21X1  g17674(.A0(new_n17858_), .A1(new_n17856_), .B0(\asqrt[58] ), .Y(new_n17867_));
  NAND2X1  g17675(.A(new_n17867_), .B(new_n328_), .Y(new_n17868_));
  OAI21X1  g17676(.A0(new_n17868_), .A1(new_n17860_), .B0(new_n17866_), .Y(new_n17869_));
  AOI21X1  g17677(.A0(new_n17869_), .A1(new_n17850_), .B0(new_n292_), .Y(new_n17870_));
  NAND4X1  g17678(.A(\asqrt[12] ), .B(new_n17203_), .C(new_n17201_), .D(new_n17221_), .Y(new_n17871_));
  OR2X1    g17679(.A(new_n17214_), .B(new_n17196_), .Y(new_n17872_));
  OAI21X1  g17680(.A0(new_n17872_), .A1(new_n17262_), .B0(new_n17202_), .Y(new_n17873_));
  AND2X1   g17681(.A(new_n17873_), .B(new_n17871_), .Y(new_n17874_));
  OAI21X1  g17682(.A0(new_n17859_), .A1(new_n17846_), .B0(new_n17867_), .Y(new_n17875_));
  AOI21X1  g17683(.A0(new_n17875_), .A1(\asqrt[59] ), .B0(\asqrt[60] ), .Y(new_n17876_));
  AOI21X1  g17684(.A0(new_n17876_), .A1(new_n17869_), .B0(new_n17874_), .Y(new_n17877_));
  OAI21X1  g17685(.A0(new_n17877_), .A1(new_n17870_), .B0(\asqrt[61] ), .Y(new_n17878_));
  AND2X1   g17686(.A(new_n17266_), .B(new_n17265_), .Y(new_n17879_));
  NOR3X1   g17687(.A(new_n17879_), .B(new_n17220_), .C(new_n17264_), .Y(new_n17880_));
  NOR3X1   g17688(.A(new_n17262_), .B(new_n17879_), .C(new_n17264_), .Y(new_n17881_));
  NOR2X1   g17689(.A(new_n17881_), .B(new_n17219_), .Y(new_n17882_));
  AOI21X1  g17690(.A0(new_n17880_), .A1(\asqrt[12] ), .B0(new_n17882_), .Y(new_n17883_));
  NOR3X1   g17691(.A(new_n17877_), .B(new_n17870_), .C(\asqrt[61] ), .Y(new_n17884_));
  OAI21X1  g17692(.A0(new_n17884_), .A1(new_n17883_), .B0(new_n17878_), .Y(new_n17885_));
  AND2X1   g17693(.A(new_n17885_), .B(\asqrt[62] ), .Y(new_n17886_));
  INVX1    g17694(.A(new_n17883_), .Y(new_n17887_));
  AND2X1   g17695(.A(new_n17875_), .B(\asqrt[59] ), .Y(new_n17888_));
  OR2X1    g17696(.A(new_n17859_), .B(new_n17846_), .Y(new_n17889_));
  AND2X1   g17697(.A(new_n17867_), .B(new_n328_), .Y(new_n17890_));
  AOI21X1  g17698(.A0(new_n17890_), .A1(new_n17889_), .B0(new_n17865_), .Y(new_n17891_));
  OAI21X1  g17699(.A0(new_n17891_), .A1(new_n17888_), .B0(\asqrt[60] ), .Y(new_n17892_));
  INVX1    g17700(.A(new_n17874_), .Y(new_n17893_));
  OAI21X1  g17701(.A0(new_n17849_), .A1(new_n328_), .B0(new_n292_), .Y(new_n17894_));
  OAI21X1  g17702(.A0(new_n17894_), .A1(new_n17891_), .B0(new_n17893_), .Y(new_n17895_));
  NAND3X1  g17703(.A(new_n17895_), .B(new_n17892_), .C(new_n217_), .Y(new_n17896_));
  NAND2X1  g17704(.A(new_n17896_), .B(new_n17887_), .Y(new_n17897_));
  AND2X1   g17705(.A(new_n17231_), .B(new_n17223_), .Y(new_n17898_));
  NOR3X1   g17706(.A(new_n17898_), .B(new_n17269_), .C(new_n17224_), .Y(new_n17899_));
  NOR3X1   g17707(.A(new_n17262_), .B(new_n17898_), .C(new_n17224_), .Y(new_n17900_));
  NOR2X1   g17708(.A(new_n17900_), .B(new_n17229_), .Y(new_n17901_));
  AOI21X1  g17709(.A0(new_n17899_), .A1(\asqrt[12] ), .B0(new_n17901_), .Y(new_n17902_));
  AOI21X1  g17710(.A0(new_n17895_), .A1(new_n17892_), .B0(new_n217_), .Y(new_n17903_));
  NOR2X1   g17711(.A(new_n17903_), .B(\asqrt[62] ), .Y(new_n17904_));
  AOI21X1  g17712(.A0(new_n17904_), .A1(new_n17897_), .B0(new_n17902_), .Y(new_n17905_));
  NOR4X1   g17713(.A(new_n17262_), .B(new_n17239_), .C(new_n17273_), .D(new_n17272_), .Y(new_n17906_));
  NAND3X1  g17714(.A(\asqrt[12] ), .B(new_n17274_), .C(new_n17233_), .Y(new_n17907_));
  AOI21X1  g17715(.A0(new_n17907_), .A1(new_n17273_), .B0(new_n17906_), .Y(new_n17908_));
  INVX1    g17716(.A(new_n17908_), .Y(new_n17909_));
  OR2X1    g17717(.A(new_n17251_), .B(new_n17250_), .Y(new_n17910_));
  INVX1    g17718(.A(new_n17910_), .Y(new_n17911_));
  AND2X1   g17719(.A(new_n17245_), .B(new_n17240_), .Y(new_n17912_));
  AOI21X1  g17720(.A0(new_n17912_), .A1(\asqrt[12] ), .B0(new_n17911_), .Y(new_n17913_));
  AND2X1   g17721(.A(new_n17913_), .B(new_n17909_), .Y(new_n17914_));
  OAI21X1  g17722(.A0(new_n17905_), .A1(new_n17886_), .B0(new_n17914_), .Y(new_n17915_));
  AOI21X1  g17723(.A0(new_n17896_), .A1(new_n17887_), .B0(new_n17903_), .Y(new_n17916_));
  OAI21X1  g17724(.A0(new_n17916_), .A1(new_n199_), .B0(new_n17908_), .Y(new_n17917_));
  AOI21X1  g17725(.A0(new_n17281_), .A1(new_n17277_), .B0(new_n17244_), .Y(new_n17918_));
  AOI21X1  g17726(.A0(new_n17245_), .A1(new_n17240_), .B0(new_n193_), .Y(new_n17919_));
  OAI21X1  g17727(.A0(new_n17918_), .A1(new_n17240_), .B0(new_n17919_), .Y(new_n17920_));
  OR2X1    g17728(.A(new_n17258_), .B(new_n17241_), .Y(new_n17921_));
  OR2X1    g17729(.A(new_n17921_), .B(new_n17243_), .Y(new_n17922_));
  NOR4X1   g17730(.A(new_n17922_), .B(new_n17302_), .C(new_n17911_), .D(new_n17249_), .Y(new_n17923_));
  INVX1    g17731(.A(new_n17923_), .Y(new_n17924_));
  AND2X1   g17732(.A(new_n17924_), .B(new_n17920_), .Y(new_n17925_));
  OAI21X1  g17733(.A0(new_n17917_), .A1(new_n17905_), .B0(new_n17925_), .Y(new_n17926_));
  AOI21X1  g17734(.A0(new_n17915_), .A1(new_n193_), .B0(new_n17926_), .Y(new_n17927_));
  NOR2X1   g17735(.A(\a[21] ), .B(\a[20] ), .Y(new_n17928_));
  INVX1    g17736(.A(new_n17928_), .Y(new_n17929_));
  MX2X1    g17737(.A(new_n17929_), .B(new_n17927_), .S0(\a[22] ), .Y(new_n17930_));
  OR2X1    g17738(.A(new_n17930_), .B(new_n17262_), .Y(new_n17931_));
  INVX1    g17739(.A(\a[22] ), .Y(new_n17932_));
  NOR3X1   g17740(.A(\a[22] ), .B(\a[21] ), .C(\a[20] ), .Y(new_n17933_));
  NOR3X1   g17741(.A(new_n17933_), .B(new_n17258_), .C(new_n17302_), .Y(new_n17934_));
  NAND3X1  g17742(.A(new_n17934_), .B(new_n17910_), .C(new_n17277_), .Y(new_n17935_));
  INVX1    g17743(.A(new_n17935_), .Y(new_n17936_));
  OAI21X1  g17744(.A0(new_n17927_), .A1(new_n17932_), .B0(new_n17936_), .Y(new_n17937_));
  OAI21X1  g17745(.A0(new_n17927_), .A1(\a[22] ), .B0(\a[23] ), .Y(new_n17938_));
  NOR2X1   g17746(.A(\a[23] ), .B(\a[22] ), .Y(new_n17939_));
  INVX1    g17747(.A(new_n17939_), .Y(new_n17940_));
  OR2X1    g17748(.A(new_n17927_), .B(new_n17940_), .Y(new_n17941_));
  NAND3X1  g17749(.A(new_n17941_), .B(new_n17938_), .C(new_n17937_), .Y(new_n17942_));
  AOI21X1  g17750(.A0(new_n17942_), .A1(new_n17931_), .B0(new_n16617_), .Y(new_n17943_));
  OR2X1    g17751(.A(new_n17916_), .B(new_n199_), .Y(new_n17944_));
  AND2X1   g17752(.A(new_n17896_), .B(new_n17887_), .Y(new_n17945_));
  INVX1    g17753(.A(new_n17902_), .Y(new_n17946_));
  OR2X1    g17754(.A(new_n17903_), .B(\asqrt[62] ), .Y(new_n17947_));
  OAI21X1  g17755(.A0(new_n17947_), .A1(new_n17945_), .B0(new_n17946_), .Y(new_n17948_));
  INVX1    g17756(.A(new_n17914_), .Y(new_n17949_));
  AOI21X1  g17757(.A0(new_n17948_), .A1(new_n17944_), .B0(new_n17949_), .Y(new_n17950_));
  AOI21X1  g17758(.A0(new_n17885_), .A1(\asqrt[62] ), .B0(new_n17909_), .Y(new_n17951_));
  INVX1    g17759(.A(new_n17925_), .Y(new_n17952_));
  AOI21X1  g17760(.A0(new_n17951_), .A1(new_n17948_), .B0(new_n17952_), .Y(new_n17953_));
  OAI21X1  g17761(.A0(new_n17950_), .A1(\asqrt[63] ), .B0(new_n17953_), .Y(\asqrt[11] ));
  MX2X1    g17762(.A(new_n17928_), .B(\asqrt[11] ), .S0(\a[22] ), .Y(new_n17955_));
  AOI21X1  g17763(.A0(new_n17955_), .A1(\asqrt[12] ), .B0(\asqrt[13] ), .Y(new_n17956_));
  NAND3X1  g17764(.A(new_n17924_), .B(new_n17920_), .C(\asqrt[12] ), .Y(new_n17957_));
  INVX1    g17765(.A(new_n17957_), .Y(new_n17958_));
  OAI21X1  g17766(.A0(new_n17917_), .A1(new_n17905_), .B0(new_n17958_), .Y(new_n17959_));
  AOI21X1  g17767(.A0(new_n17915_), .A1(new_n193_), .B0(new_n17959_), .Y(new_n17960_));
  AOI21X1  g17768(.A0(\asqrt[11] ), .A1(new_n17939_), .B0(new_n17960_), .Y(new_n17961_));
  OR2X1    g17769(.A(new_n17961_), .B(new_n17263_), .Y(new_n17962_));
  AND2X1   g17770(.A(\asqrt[11] ), .B(new_n17939_), .Y(new_n17963_));
  OR2X1    g17771(.A(new_n17960_), .B(\a[24] ), .Y(new_n17964_));
  OR2X1    g17772(.A(new_n17964_), .B(new_n17963_), .Y(new_n17965_));
  AOI22X1  g17773(.A0(new_n17965_), .A1(new_n17962_), .B0(new_n17956_), .B1(new_n17942_), .Y(new_n17966_));
  OAI21X1  g17774(.A0(new_n17966_), .A1(new_n17943_), .B0(\asqrt[14] ), .Y(new_n17967_));
  AND2X1   g17775(.A(new_n17295_), .B(new_n17284_), .Y(new_n17968_));
  NAND3X1  g17776(.A(new_n17968_), .B(\asqrt[11] ), .C(new_n17292_), .Y(new_n17969_));
  INVX1    g17777(.A(new_n17968_), .Y(new_n17970_));
  OAI21X1  g17778(.A0(new_n17970_), .A1(new_n17927_), .B0(new_n17299_), .Y(new_n17971_));
  AND2X1   g17779(.A(new_n17971_), .B(new_n17969_), .Y(new_n17972_));
  NOR3X1   g17780(.A(new_n17966_), .B(new_n17943_), .C(\asqrt[14] ), .Y(new_n17973_));
  OAI21X1  g17781(.A0(new_n17973_), .A1(new_n17972_), .B0(new_n17967_), .Y(new_n17974_));
  AND2X1   g17782(.A(new_n17974_), .B(\asqrt[15] ), .Y(new_n17975_));
  INVX1    g17783(.A(new_n17972_), .Y(new_n17976_));
  AND2X1   g17784(.A(new_n17955_), .B(\asqrt[12] ), .Y(new_n17977_));
  AOI21X1  g17785(.A0(\asqrt[11] ), .A1(\a[22] ), .B0(new_n17935_), .Y(new_n17978_));
  INVX1    g17786(.A(\a[23] ), .Y(new_n17979_));
  AOI21X1  g17787(.A0(\asqrt[11] ), .A1(new_n17932_), .B0(new_n17979_), .Y(new_n17980_));
  NOR3X1   g17788(.A(new_n17963_), .B(new_n17980_), .C(new_n17978_), .Y(new_n17981_));
  OAI21X1  g17789(.A0(new_n17981_), .A1(new_n17977_), .B0(\asqrt[13] ), .Y(new_n17982_));
  OAI21X1  g17790(.A0(new_n17930_), .A1(new_n17262_), .B0(new_n16617_), .Y(new_n17983_));
  OAI22X1  g17791(.A0(new_n17964_), .A1(new_n17963_), .B0(new_n17961_), .B1(new_n17263_), .Y(new_n17984_));
  OAI21X1  g17792(.A0(new_n17983_), .A1(new_n17981_), .B0(new_n17984_), .Y(new_n17985_));
  NAND3X1  g17793(.A(new_n17985_), .B(new_n17982_), .C(new_n15990_), .Y(new_n17986_));
  NAND2X1  g17794(.A(new_n17986_), .B(new_n17976_), .Y(new_n17987_));
  AOI21X1  g17795(.A0(new_n17301_), .A1(new_n17300_), .B0(new_n17335_), .Y(new_n17988_));
  AND2X1   g17796(.A(new_n17988_), .B(new_n17332_), .Y(new_n17989_));
  INVX1    g17797(.A(new_n17989_), .Y(new_n17990_));
  OR2X1    g17798(.A(new_n17990_), .B(new_n17927_), .Y(new_n17991_));
  OAI22X1  g17799(.A0(new_n17334_), .A1(new_n17333_), .B0(new_n17317_), .B1(new_n15990_), .Y(new_n17992_));
  OAI21X1  g17800(.A0(new_n17992_), .A1(new_n17927_), .B0(new_n17335_), .Y(new_n17993_));
  AND2X1   g17801(.A(new_n17993_), .B(new_n17991_), .Y(new_n17994_));
  AOI21X1  g17802(.A0(new_n17985_), .A1(new_n17982_), .B0(new_n15990_), .Y(new_n17995_));
  NOR2X1   g17803(.A(new_n17995_), .B(\asqrt[15] ), .Y(new_n17996_));
  AOI21X1  g17804(.A0(new_n17996_), .A1(new_n17987_), .B0(new_n17994_), .Y(new_n17997_));
  OAI21X1  g17805(.A0(new_n17997_), .A1(new_n17975_), .B0(\asqrt[16] ), .Y(new_n17998_));
  AND2X1   g17806(.A(new_n17339_), .B(new_n17336_), .Y(new_n17999_));
  OR4X1    g17807(.A(new_n17927_), .B(new_n17999_), .C(new_n17314_), .D(new_n17337_), .Y(new_n18000_));
  OR2X1    g17808(.A(new_n17999_), .B(new_n17337_), .Y(new_n18001_));
  OAI21X1  g17809(.A0(new_n18001_), .A1(new_n17927_), .B0(new_n17314_), .Y(new_n18002_));
  AND2X1   g17810(.A(new_n18002_), .B(new_n18000_), .Y(new_n18003_));
  INVX1    g17811(.A(new_n18003_), .Y(new_n18004_));
  AOI21X1  g17812(.A0(new_n17986_), .A1(new_n17976_), .B0(new_n17995_), .Y(new_n18005_));
  OAI21X1  g17813(.A0(new_n18005_), .A1(new_n15362_), .B0(new_n14754_), .Y(new_n18006_));
  OAI21X1  g17814(.A0(new_n18006_), .A1(new_n17997_), .B0(new_n18004_), .Y(new_n18007_));
  AOI21X1  g17815(.A0(new_n18007_), .A1(new_n17998_), .B0(new_n14165_), .Y(new_n18008_));
  NAND3X1  g17816(.A(new_n17329_), .B(new_n17327_), .C(new_n17350_), .Y(new_n18009_));
  NOR3X1   g17817(.A(new_n17927_), .B(new_n17341_), .C(new_n17320_), .Y(new_n18010_));
  OAI22X1  g17818(.A0(new_n18010_), .A1(new_n17327_), .B0(new_n18009_), .B1(new_n17927_), .Y(new_n18011_));
  NAND3X1  g17819(.A(new_n18007_), .B(new_n17998_), .C(new_n14165_), .Y(new_n18012_));
  AOI21X1  g17820(.A0(new_n18012_), .A1(new_n18011_), .B0(new_n18008_), .Y(new_n18013_));
  OR2X1    g17821(.A(new_n18013_), .B(new_n13571_), .Y(new_n18014_));
  AND2X1   g17822(.A(new_n18012_), .B(new_n18011_), .Y(new_n18015_));
  AND2X1   g17823(.A(new_n17373_), .B(new_n17372_), .Y(new_n18016_));
  NOR4X1   g17824(.A(new_n17927_), .B(new_n18016_), .C(new_n17349_), .D(new_n17371_), .Y(new_n18017_));
  AOI22X1  g17825(.A0(new_n17373_), .A1(new_n17372_), .B0(new_n17358_), .B1(\asqrt[17] ), .Y(new_n18018_));
  AOI21X1  g17826(.A0(new_n18018_), .A1(\asqrt[11] ), .B0(new_n17348_), .Y(new_n18019_));
  NOR2X1   g17827(.A(new_n18019_), .B(new_n18017_), .Y(new_n18020_));
  INVX1    g17828(.A(new_n18020_), .Y(new_n18021_));
  OR2X1    g17829(.A(new_n18008_), .B(\asqrt[18] ), .Y(new_n18022_));
  OAI21X1  g17830(.A0(new_n18022_), .A1(new_n18015_), .B0(new_n18021_), .Y(new_n18023_));
  AOI21X1  g17831(.A0(new_n18023_), .A1(new_n18014_), .B0(new_n13000_), .Y(new_n18024_));
  AND2X1   g17832(.A(new_n17359_), .B(new_n17352_), .Y(new_n18025_));
  OR4X1    g17833(.A(new_n17927_), .B(new_n18025_), .C(new_n17356_), .D(new_n17353_), .Y(new_n18026_));
  OR2X1    g17834(.A(new_n18025_), .B(new_n17353_), .Y(new_n18027_));
  OAI21X1  g17835(.A0(new_n18027_), .A1(new_n17927_), .B0(new_n17356_), .Y(new_n18028_));
  AND2X1   g17836(.A(new_n18028_), .B(new_n18026_), .Y(new_n18029_));
  OR2X1    g17837(.A(new_n18005_), .B(new_n15362_), .Y(new_n18030_));
  AND2X1   g17838(.A(new_n17986_), .B(new_n17976_), .Y(new_n18031_));
  INVX1    g17839(.A(new_n17994_), .Y(new_n18032_));
  OR2X1    g17840(.A(new_n17995_), .B(\asqrt[15] ), .Y(new_n18033_));
  OAI21X1  g17841(.A0(new_n18033_), .A1(new_n18031_), .B0(new_n18032_), .Y(new_n18034_));
  AOI21X1  g17842(.A0(new_n18034_), .A1(new_n18030_), .B0(new_n14754_), .Y(new_n18035_));
  AOI21X1  g17843(.A0(new_n17974_), .A1(\asqrt[15] ), .B0(\asqrt[16] ), .Y(new_n18036_));
  AOI21X1  g17844(.A0(new_n18036_), .A1(new_n18034_), .B0(new_n18003_), .Y(new_n18037_));
  OAI21X1  g17845(.A0(new_n18037_), .A1(new_n18035_), .B0(\asqrt[17] ), .Y(new_n18038_));
  INVX1    g17846(.A(new_n18011_), .Y(new_n18039_));
  NOR3X1   g17847(.A(new_n18037_), .B(new_n18035_), .C(\asqrt[17] ), .Y(new_n18040_));
  OAI21X1  g17848(.A0(new_n18040_), .A1(new_n18039_), .B0(new_n18038_), .Y(new_n18041_));
  AOI21X1  g17849(.A0(new_n18041_), .A1(\asqrt[18] ), .B0(\asqrt[19] ), .Y(new_n18042_));
  AOI21X1  g17850(.A0(new_n18042_), .A1(new_n18023_), .B0(new_n18029_), .Y(new_n18043_));
  OAI21X1  g17851(.A0(new_n18043_), .A1(new_n18024_), .B0(\asqrt[20] ), .Y(new_n18044_));
  OR4X1    g17852(.A(new_n17927_), .B(new_n17367_), .C(new_n17370_), .D(new_n17393_), .Y(new_n18045_));
  NAND2X1  g17853(.A(new_n17378_), .B(new_n17361_), .Y(new_n18046_));
  OAI21X1  g17854(.A0(new_n18046_), .A1(new_n17927_), .B0(new_n17370_), .Y(new_n18047_));
  AND2X1   g17855(.A(new_n18047_), .B(new_n18045_), .Y(new_n18048_));
  NOR3X1   g17856(.A(new_n18043_), .B(new_n18024_), .C(\asqrt[20] ), .Y(new_n18049_));
  OAI21X1  g17857(.A0(new_n18049_), .A1(new_n18048_), .B0(new_n18044_), .Y(new_n18050_));
  AND2X1   g17858(.A(new_n18050_), .B(\asqrt[21] ), .Y(new_n18051_));
  INVX1    g17859(.A(new_n18048_), .Y(new_n18052_));
  AND2X1   g17860(.A(new_n18041_), .B(\asqrt[18] ), .Y(new_n18053_));
  NAND2X1  g17861(.A(new_n18012_), .B(new_n18011_), .Y(new_n18054_));
  NOR2X1   g17862(.A(new_n18008_), .B(\asqrt[18] ), .Y(new_n18055_));
  AOI21X1  g17863(.A0(new_n18055_), .A1(new_n18054_), .B0(new_n18020_), .Y(new_n18056_));
  OAI21X1  g17864(.A0(new_n18056_), .A1(new_n18053_), .B0(\asqrt[19] ), .Y(new_n18057_));
  INVX1    g17865(.A(new_n18029_), .Y(new_n18058_));
  OAI21X1  g17866(.A0(new_n18013_), .A1(new_n13571_), .B0(new_n13000_), .Y(new_n18059_));
  OAI21X1  g17867(.A0(new_n18059_), .A1(new_n18056_), .B0(new_n18058_), .Y(new_n18060_));
  NAND3X1  g17868(.A(new_n18060_), .B(new_n18057_), .C(new_n12447_), .Y(new_n18061_));
  NAND2X1  g17869(.A(new_n18061_), .B(new_n18052_), .Y(new_n18062_));
  OAI21X1  g17870(.A0(new_n17417_), .A1(new_n17415_), .B0(new_n17384_), .Y(new_n18063_));
  NOR3X1   g17871(.A(new_n18063_), .B(new_n17927_), .C(new_n17369_), .Y(new_n18064_));
  AOI22X1  g17872(.A0(new_n17385_), .A1(new_n17379_), .B0(new_n17368_), .B1(\asqrt[20] ), .Y(new_n18065_));
  AOI21X1  g17873(.A0(new_n18065_), .A1(\asqrt[11] ), .B0(new_n17384_), .Y(new_n18066_));
  NOR2X1   g17874(.A(new_n18066_), .B(new_n18064_), .Y(new_n18067_));
  AOI21X1  g17875(.A0(new_n18060_), .A1(new_n18057_), .B0(new_n12447_), .Y(new_n18068_));
  NOR2X1   g17876(.A(new_n18068_), .B(\asqrt[21] ), .Y(new_n18069_));
  AOI21X1  g17877(.A0(new_n18069_), .A1(new_n18062_), .B0(new_n18067_), .Y(new_n18070_));
  OAI21X1  g17878(.A0(new_n18070_), .A1(new_n18051_), .B0(\asqrt[22] ), .Y(new_n18071_));
  AND2X1   g17879(.A(new_n17420_), .B(new_n17418_), .Y(new_n18072_));
  OR4X1    g17880(.A(new_n17927_), .B(new_n18072_), .C(new_n17392_), .D(new_n17419_), .Y(new_n18073_));
  OR2X1    g17881(.A(new_n18072_), .B(new_n17419_), .Y(new_n18074_));
  OAI21X1  g17882(.A0(new_n18074_), .A1(new_n17927_), .B0(new_n17392_), .Y(new_n18075_));
  AND2X1   g17883(.A(new_n18075_), .B(new_n18073_), .Y(new_n18076_));
  INVX1    g17884(.A(new_n18076_), .Y(new_n18077_));
  AOI21X1  g17885(.A0(new_n18061_), .A1(new_n18052_), .B0(new_n18068_), .Y(new_n18078_));
  OAI21X1  g17886(.A0(new_n18078_), .A1(new_n11896_), .B0(new_n11362_), .Y(new_n18079_));
  OAI21X1  g17887(.A0(new_n18079_), .A1(new_n18070_), .B0(new_n18077_), .Y(new_n18080_));
  AOI21X1  g17888(.A0(new_n18080_), .A1(new_n18071_), .B0(new_n10849_), .Y(new_n18081_));
  NAND3X1  g17889(.A(new_n17404_), .B(new_n17402_), .C(new_n17422_), .Y(new_n18082_));
  NOR3X1   g17890(.A(new_n17927_), .B(new_n17430_), .C(new_n17397_), .Y(new_n18083_));
  OAI22X1  g17891(.A0(new_n18083_), .A1(new_n17402_), .B0(new_n18082_), .B1(new_n17927_), .Y(new_n18084_));
  NAND3X1  g17892(.A(new_n18080_), .B(new_n18071_), .C(new_n10849_), .Y(new_n18085_));
  AOI21X1  g17893(.A0(new_n18085_), .A1(new_n18084_), .B0(new_n18081_), .Y(new_n18086_));
  OR2X1    g17894(.A(new_n18086_), .B(new_n10332_), .Y(new_n18087_));
  AND2X1   g17895(.A(new_n18085_), .B(new_n18084_), .Y(new_n18088_));
  AND2X1   g17896(.A(new_n17446_), .B(new_n17445_), .Y(new_n18089_));
  NOR4X1   g17897(.A(new_n17927_), .B(new_n18089_), .C(new_n17413_), .D(new_n17444_), .Y(new_n18090_));
  AOI22X1  g17898(.A0(new_n17446_), .A1(new_n17445_), .B0(new_n17431_), .B1(\asqrt[23] ), .Y(new_n18091_));
  AOI21X1  g17899(.A0(new_n18091_), .A1(\asqrt[11] ), .B0(new_n17412_), .Y(new_n18092_));
  NOR2X1   g17900(.A(new_n18092_), .B(new_n18090_), .Y(new_n18093_));
  INVX1    g17901(.A(new_n18093_), .Y(new_n18094_));
  OR2X1    g17902(.A(new_n18081_), .B(\asqrt[24] ), .Y(new_n18095_));
  OAI21X1  g17903(.A0(new_n18095_), .A1(new_n18088_), .B0(new_n18094_), .Y(new_n18096_));
  AOI21X1  g17904(.A0(new_n18096_), .A1(new_n18087_), .B0(new_n9833_), .Y(new_n18097_));
  OAI21X1  g17905(.A0(new_n17450_), .A1(new_n17447_), .B0(new_n17429_), .Y(new_n18098_));
  OR2X1    g17906(.A(new_n18098_), .B(new_n17425_), .Y(new_n18099_));
  AND2X1   g17907(.A(new_n17432_), .B(new_n17424_), .Y(new_n18100_));
  NOR3X1   g17908(.A(new_n17927_), .B(new_n18100_), .C(new_n17425_), .Y(new_n18101_));
  OAI22X1  g17909(.A0(new_n18101_), .A1(new_n17429_), .B0(new_n18099_), .B1(new_n17927_), .Y(new_n18102_));
  INVX1    g17910(.A(new_n18102_), .Y(new_n18103_));
  OR2X1    g17911(.A(new_n18078_), .B(new_n11896_), .Y(new_n18104_));
  AND2X1   g17912(.A(new_n18061_), .B(new_n18052_), .Y(new_n18105_));
  INVX1    g17913(.A(new_n18067_), .Y(new_n18106_));
  OR2X1    g17914(.A(new_n18068_), .B(\asqrt[21] ), .Y(new_n18107_));
  OAI21X1  g17915(.A0(new_n18107_), .A1(new_n18105_), .B0(new_n18106_), .Y(new_n18108_));
  AOI21X1  g17916(.A0(new_n18108_), .A1(new_n18104_), .B0(new_n11362_), .Y(new_n18109_));
  AOI21X1  g17917(.A0(new_n18050_), .A1(\asqrt[21] ), .B0(\asqrt[22] ), .Y(new_n18110_));
  AOI21X1  g17918(.A0(new_n18110_), .A1(new_n18108_), .B0(new_n18076_), .Y(new_n18111_));
  OAI21X1  g17919(.A0(new_n18111_), .A1(new_n18109_), .B0(\asqrt[23] ), .Y(new_n18112_));
  INVX1    g17920(.A(new_n18084_), .Y(new_n18113_));
  NOR3X1   g17921(.A(new_n18111_), .B(new_n18109_), .C(\asqrt[23] ), .Y(new_n18114_));
  OAI21X1  g17922(.A0(new_n18114_), .A1(new_n18113_), .B0(new_n18112_), .Y(new_n18115_));
  AOI21X1  g17923(.A0(new_n18115_), .A1(\asqrt[24] ), .B0(\asqrt[25] ), .Y(new_n18116_));
  AOI21X1  g17924(.A0(new_n18116_), .A1(new_n18096_), .B0(new_n18103_), .Y(new_n18117_));
  OAI21X1  g17925(.A0(new_n18117_), .A1(new_n18097_), .B0(\asqrt[26] ), .Y(new_n18118_));
  OR4X1    g17926(.A(new_n17927_), .B(new_n17440_), .C(new_n17443_), .D(new_n17467_), .Y(new_n18119_));
  NAND2X1  g17927(.A(new_n17452_), .B(new_n17434_), .Y(new_n18120_));
  OAI21X1  g17928(.A0(new_n18120_), .A1(new_n17927_), .B0(new_n17443_), .Y(new_n18121_));
  AND2X1   g17929(.A(new_n18121_), .B(new_n18119_), .Y(new_n18122_));
  NOR3X1   g17930(.A(new_n18117_), .B(new_n18097_), .C(\asqrt[26] ), .Y(new_n18123_));
  OAI21X1  g17931(.A0(new_n18123_), .A1(new_n18122_), .B0(new_n18118_), .Y(new_n18124_));
  AND2X1   g17932(.A(new_n18124_), .B(\asqrt[27] ), .Y(new_n18125_));
  INVX1    g17933(.A(new_n18122_), .Y(new_n18126_));
  AND2X1   g17934(.A(new_n18115_), .B(\asqrt[24] ), .Y(new_n18127_));
  NAND2X1  g17935(.A(new_n18085_), .B(new_n18084_), .Y(new_n18128_));
  NOR2X1   g17936(.A(new_n18081_), .B(\asqrt[24] ), .Y(new_n18129_));
  AOI21X1  g17937(.A0(new_n18129_), .A1(new_n18128_), .B0(new_n18093_), .Y(new_n18130_));
  OAI21X1  g17938(.A0(new_n18130_), .A1(new_n18127_), .B0(\asqrt[25] ), .Y(new_n18131_));
  OAI21X1  g17939(.A0(new_n18086_), .A1(new_n10332_), .B0(new_n9833_), .Y(new_n18132_));
  OAI21X1  g17940(.A0(new_n18132_), .A1(new_n18130_), .B0(new_n18102_), .Y(new_n18133_));
  NAND3X1  g17941(.A(new_n18133_), .B(new_n18131_), .C(new_n9353_), .Y(new_n18134_));
  NAND2X1  g17942(.A(new_n18134_), .B(new_n18126_), .Y(new_n18135_));
  OAI21X1  g17943(.A0(new_n17491_), .A1(new_n17489_), .B0(new_n17458_), .Y(new_n18136_));
  NOR3X1   g17944(.A(new_n18136_), .B(new_n17927_), .C(new_n17442_), .Y(new_n18137_));
  AOI22X1  g17945(.A0(new_n17459_), .A1(new_n17453_), .B0(new_n17441_), .B1(\asqrt[26] ), .Y(new_n18138_));
  AOI21X1  g17946(.A0(new_n18138_), .A1(\asqrt[11] ), .B0(new_n17458_), .Y(new_n18139_));
  NOR2X1   g17947(.A(new_n18139_), .B(new_n18137_), .Y(new_n18140_));
  AOI21X1  g17948(.A0(new_n18133_), .A1(new_n18131_), .B0(new_n9353_), .Y(new_n18141_));
  NOR2X1   g17949(.A(new_n18141_), .B(\asqrt[27] ), .Y(new_n18142_));
  AOI21X1  g17950(.A0(new_n18142_), .A1(new_n18135_), .B0(new_n18140_), .Y(new_n18143_));
  OAI21X1  g17951(.A0(new_n18143_), .A1(new_n18125_), .B0(\asqrt[28] ), .Y(new_n18144_));
  AND2X1   g17952(.A(new_n17494_), .B(new_n17492_), .Y(new_n18145_));
  OR2X1    g17953(.A(new_n17466_), .B(new_n17493_), .Y(new_n18146_));
  OR2X1    g17954(.A(new_n18146_), .B(new_n18145_), .Y(new_n18147_));
  NOR3X1   g17955(.A(new_n17927_), .B(new_n18145_), .C(new_n17493_), .Y(new_n18148_));
  OAI22X1  g17956(.A0(new_n18148_), .A1(new_n17465_), .B0(new_n18147_), .B1(new_n17927_), .Y(new_n18149_));
  AOI21X1  g17957(.A0(new_n18134_), .A1(new_n18126_), .B0(new_n18141_), .Y(new_n18150_));
  OAI21X1  g17958(.A0(new_n18150_), .A1(new_n8874_), .B0(new_n8412_), .Y(new_n18151_));
  OAI21X1  g17959(.A0(new_n18151_), .A1(new_n18143_), .B0(new_n18149_), .Y(new_n18152_));
  AOI21X1  g17960(.A0(new_n18152_), .A1(new_n18144_), .B0(new_n7970_), .Y(new_n18153_));
  OR4X1    g17961(.A(new_n17927_), .B(new_n17504_), .C(new_n17477_), .D(new_n17471_), .Y(new_n18154_));
  NAND2X1  g17962(.A(new_n17478_), .B(new_n17496_), .Y(new_n18155_));
  OAI21X1  g17963(.A0(new_n18155_), .A1(new_n17927_), .B0(new_n17477_), .Y(new_n18156_));
  AND2X1   g17964(.A(new_n18156_), .B(new_n18154_), .Y(new_n18157_));
  INVX1    g17965(.A(new_n18157_), .Y(new_n18158_));
  NAND3X1  g17966(.A(new_n18152_), .B(new_n18144_), .C(new_n7970_), .Y(new_n18159_));
  AOI21X1  g17967(.A0(new_n18159_), .A1(new_n18158_), .B0(new_n18153_), .Y(new_n18160_));
  OR2X1    g17968(.A(new_n18160_), .B(new_n7527_), .Y(new_n18161_));
  AND2X1   g17969(.A(new_n18159_), .B(new_n18158_), .Y(new_n18162_));
  AND2X1   g17970(.A(new_n17520_), .B(new_n17519_), .Y(new_n18163_));
  NOR4X1   g17971(.A(new_n17927_), .B(new_n18163_), .C(new_n17487_), .D(new_n17518_), .Y(new_n18164_));
  AOI22X1  g17972(.A0(new_n17520_), .A1(new_n17519_), .B0(new_n17505_), .B1(\asqrt[29] ), .Y(new_n18165_));
  AOI21X1  g17973(.A0(new_n18165_), .A1(\asqrt[11] ), .B0(new_n17486_), .Y(new_n18166_));
  NOR2X1   g17974(.A(new_n18166_), .B(new_n18164_), .Y(new_n18167_));
  INVX1    g17975(.A(new_n18167_), .Y(new_n18168_));
  OR2X1    g17976(.A(new_n18153_), .B(\asqrt[30] ), .Y(new_n18169_));
  OAI21X1  g17977(.A0(new_n18169_), .A1(new_n18162_), .B0(new_n18168_), .Y(new_n18170_));
  AOI21X1  g17978(.A0(new_n18170_), .A1(new_n18161_), .B0(new_n7103_), .Y(new_n18171_));
  AND2X1   g17979(.A(new_n17506_), .B(new_n17498_), .Y(new_n18172_));
  OR4X1    g17980(.A(new_n17927_), .B(new_n18172_), .C(new_n17523_), .D(new_n17499_), .Y(new_n18173_));
  OR2X1    g17981(.A(new_n18172_), .B(new_n17499_), .Y(new_n18174_));
  OAI21X1  g17982(.A0(new_n18174_), .A1(new_n17927_), .B0(new_n17523_), .Y(new_n18175_));
  AND2X1   g17983(.A(new_n18175_), .B(new_n18173_), .Y(new_n18176_));
  OR2X1    g17984(.A(new_n18150_), .B(new_n8874_), .Y(new_n18177_));
  AND2X1   g17985(.A(new_n18134_), .B(new_n18126_), .Y(new_n18178_));
  INVX1    g17986(.A(new_n18140_), .Y(new_n18179_));
  OR2X1    g17987(.A(new_n18141_), .B(\asqrt[27] ), .Y(new_n18180_));
  OAI21X1  g17988(.A0(new_n18180_), .A1(new_n18178_), .B0(new_n18179_), .Y(new_n18181_));
  AOI21X1  g17989(.A0(new_n18181_), .A1(new_n18177_), .B0(new_n8412_), .Y(new_n18182_));
  INVX1    g17990(.A(new_n18149_), .Y(new_n18183_));
  AOI21X1  g17991(.A0(new_n18124_), .A1(\asqrt[27] ), .B0(\asqrt[28] ), .Y(new_n18184_));
  AOI21X1  g17992(.A0(new_n18184_), .A1(new_n18181_), .B0(new_n18183_), .Y(new_n18185_));
  OAI21X1  g17993(.A0(new_n18185_), .A1(new_n18182_), .B0(\asqrt[29] ), .Y(new_n18186_));
  NOR3X1   g17994(.A(new_n18185_), .B(new_n18182_), .C(\asqrt[29] ), .Y(new_n18187_));
  OAI21X1  g17995(.A0(new_n18187_), .A1(new_n18157_), .B0(new_n18186_), .Y(new_n18188_));
  AOI21X1  g17996(.A0(new_n18188_), .A1(\asqrt[30] ), .B0(\asqrt[31] ), .Y(new_n18189_));
  AOI21X1  g17997(.A0(new_n18189_), .A1(new_n18170_), .B0(new_n18176_), .Y(new_n18190_));
  OAI21X1  g17998(.A0(new_n18190_), .A1(new_n18171_), .B0(\asqrt[32] ), .Y(new_n18191_));
  NOR3X1   g17999(.A(new_n17514_), .B(new_n17517_), .C(new_n17541_), .Y(new_n18192_));
  AND2X1   g18000(.A(new_n17526_), .B(new_n17508_), .Y(new_n18193_));
  AOI21X1  g18001(.A0(new_n18193_), .A1(\asqrt[11] ), .B0(new_n17513_), .Y(new_n18194_));
  AOI21X1  g18002(.A0(new_n18192_), .A1(\asqrt[11] ), .B0(new_n18194_), .Y(new_n18195_));
  NOR3X1   g18003(.A(new_n18190_), .B(new_n18171_), .C(\asqrt[32] ), .Y(new_n18196_));
  OAI21X1  g18004(.A0(new_n18196_), .A1(new_n18195_), .B0(new_n18191_), .Y(new_n18197_));
  AND2X1   g18005(.A(new_n18197_), .B(\asqrt[33] ), .Y(new_n18198_));
  INVX1    g18006(.A(new_n18195_), .Y(new_n18199_));
  AND2X1   g18007(.A(new_n18188_), .B(\asqrt[30] ), .Y(new_n18200_));
  NAND2X1  g18008(.A(new_n18159_), .B(new_n18158_), .Y(new_n18201_));
  NOR2X1   g18009(.A(new_n18153_), .B(\asqrt[30] ), .Y(new_n18202_));
  AOI21X1  g18010(.A0(new_n18202_), .A1(new_n18201_), .B0(new_n18167_), .Y(new_n18203_));
  OAI21X1  g18011(.A0(new_n18203_), .A1(new_n18200_), .B0(\asqrt[31] ), .Y(new_n18204_));
  INVX1    g18012(.A(new_n18176_), .Y(new_n18205_));
  OAI21X1  g18013(.A0(new_n18160_), .A1(new_n7527_), .B0(new_n7103_), .Y(new_n18206_));
  OAI21X1  g18014(.A0(new_n18206_), .A1(new_n18203_), .B0(new_n18205_), .Y(new_n18207_));
  NAND3X1  g18015(.A(new_n18207_), .B(new_n18204_), .C(new_n6699_), .Y(new_n18208_));
  NAND2X1  g18016(.A(new_n18208_), .B(new_n18199_), .Y(new_n18209_));
  OAI21X1  g18017(.A0(new_n17558_), .A1(new_n17556_), .B0(new_n17532_), .Y(new_n18210_));
  NOR3X1   g18018(.A(new_n18210_), .B(new_n17927_), .C(new_n17516_), .Y(new_n18211_));
  AOI22X1  g18019(.A0(new_n17533_), .A1(new_n17527_), .B0(new_n17515_), .B1(\asqrt[32] ), .Y(new_n18212_));
  AOI21X1  g18020(.A0(new_n18212_), .A1(\asqrt[11] ), .B0(new_n17532_), .Y(new_n18213_));
  NOR2X1   g18021(.A(new_n18213_), .B(new_n18211_), .Y(new_n18214_));
  AND2X1   g18022(.A(new_n18191_), .B(new_n6294_), .Y(new_n18215_));
  AOI21X1  g18023(.A0(new_n18215_), .A1(new_n18209_), .B0(new_n18214_), .Y(new_n18216_));
  OAI21X1  g18024(.A0(new_n18216_), .A1(new_n18198_), .B0(\asqrt[34] ), .Y(new_n18217_));
  AND2X1   g18025(.A(new_n17561_), .B(new_n17559_), .Y(new_n18218_));
  OR4X1    g18026(.A(new_n17927_), .B(new_n18218_), .C(new_n17540_), .D(new_n17560_), .Y(new_n18219_));
  OR2X1    g18027(.A(new_n18218_), .B(new_n17560_), .Y(new_n18220_));
  OAI21X1  g18028(.A0(new_n18220_), .A1(new_n17927_), .B0(new_n17540_), .Y(new_n18221_));
  AND2X1   g18029(.A(new_n18221_), .B(new_n18219_), .Y(new_n18222_));
  INVX1    g18030(.A(new_n18222_), .Y(new_n18223_));
  AOI21X1  g18031(.A0(new_n18207_), .A1(new_n18204_), .B0(new_n6699_), .Y(new_n18224_));
  AOI21X1  g18032(.A0(new_n18208_), .A1(new_n18199_), .B0(new_n18224_), .Y(new_n18225_));
  OAI21X1  g18033(.A0(new_n18225_), .A1(new_n6294_), .B0(new_n5941_), .Y(new_n18226_));
  OAI21X1  g18034(.A0(new_n18226_), .A1(new_n18216_), .B0(new_n18223_), .Y(new_n18227_));
  AOI21X1  g18035(.A0(new_n18227_), .A1(new_n18217_), .B0(new_n5541_), .Y(new_n18228_));
  OR4X1    g18036(.A(new_n17927_), .B(new_n17563_), .C(new_n17551_), .D(new_n17545_), .Y(new_n18229_));
  OR2X1    g18037(.A(new_n17563_), .B(new_n17545_), .Y(new_n18230_));
  OAI21X1  g18038(.A0(new_n18230_), .A1(new_n17927_), .B0(new_n17551_), .Y(new_n18231_));
  AND2X1   g18039(.A(new_n18231_), .B(new_n18229_), .Y(new_n18232_));
  INVX1    g18040(.A(new_n18232_), .Y(new_n18233_));
  NAND3X1  g18041(.A(new_n18227_), .B(new_n18217_), .C(new_n5541_), .Y(new_n18234_));
  AOI21X1  g18042(.A0(new_n18234_), .A1(new_n18233_), .B0(new_n18228_), .Y(new_n18235_));
  OR2X1    g18043(.A(new_n18235_), .B(new_n5176_), .Y(new_n18236_));
  AND2X1   g18044(.A(new_n18234_), .B(new_n18233_), .Y(new_n18237_));
  AND2X1   g18045(.A(new_n17607_), .B(new_n17606_), .Y(new_n18238_));
  NOR4X1   g18046(.A(new_n17927_), .B(new_n18238_), .C(new_n17570_), .D(new_n17605_), .Y(new_n18239_));
  AOI22X1  g18047(.A0(new_n17607_), .A1(new_n17606_), .B0(new_n17579_), .B1(\asqrt[35] ), .Y(new_n18240_));
  AOI21X1  g18048(.A0(new_n18240_), .A1(\asqrt[11] ), .B0(new_n17569_), .Y(new_n18241_));
  NOR2X1   g18049(.A(new_n18241_), .B(new_n18239_), .Y(new_n18242_));
  INVX1    g18050(.A(new_n18242_), .Y(new_n18243_));
  OR2X1    g18051(.A(new_n18228_), .B(\asqrt[36] ), .Y(new_n18244_));
  OAI21X1  g18052(.A0(new_n18244_), .A1(new_n18237_), .B0(new_n18243_), .Y(new_n18245_));
  AOI21X1  g18053(.A0(new_n18245_), .A1(new_n18236_), .B0(new_n4826_), .Y(new_n18246_));
  AND2X1   g18054(.A(new_n17580_), .B(new_n17573_), .Y(new_n18247_));
  OR4X1    g18055(.A(new_n17927_), .B(new_n18247_), .C(new_n17610_), .D(new_n17574_), .Y(new_n18248_));
  OR2X1    g18056(.A(new_n18247_), .B(new_n17574_), .Y(new_n18249_));
  OAI21X1  g18057(.A0(new_n18249_), .A1(new_n17927_), .B0(new_n17610_), .Y(new_n18250_));
  AND2X1   g18058(.A(new_n18250_), .B(new_n18248_), .Y(new_n18251_));
  OR2X1    g18059(.A(new_n18225_), .B(new_n6294_), .Y(new_n18252_));
  AND2X1   g18060(.A(new_n18208_), .B(new_n18199_), .Y(new_n18253_));
  INVX1    g18061(.A(new_n18214_), .Y(new_n18254_));
  NAND2X1  g18062(.A(new_n18191_), .B(new_n6294_), .Y(new_n18255_));
  OAI21X1  g18063(.A0(new_n18255_), .A1(new_n18253_), .B0(new_n18254_), .Y(new_n18256_));
  AOI21X1  g18064(.A0(new_n18256_), .A1(new_n18252_), .B0(new_n5941_), .Y(new_n18257_));
  AOI21X1  g18065(.A0(new_n18197_), .A1(\asqrt[33] ), .B0(\asqrt[34] ), .Y(new_n18258_));
  AOI21X1  g18066(.A0(new_n18258_), .A1(new_n18256_), .B0(new_n18222_), .Y(new_n18259_));
  OAI21X1  g18067(.A0(new_n18259_), .A1(new_n18257_), .B0(\asqrt[35] ), .Y(new_n18260_));
  NOR3X1   g18068(.A(new_n18259_), .B(new_n18257_), .C(\asqrt[35] ), .Y(new_n18261_));
  OAI21X1  g18069(.A0(new_n18261_), .A1(new_n18232_), .B0(new_n18260_), .Y(new_n18262_));
  AOI21X1  g18070(.A0(new_n18262_), .A1(\asqrt[36] ), .B0(\asqrt[37] ), .Y(new_n18263_));
  AOI21X1  g18071(.A0(new_n18263_), .A1(new_n18245_), .B0(new_n18251_), .Y(new_n18264_));
  OAI21X1  g18072(.A0(new_n18264_), .A1(new_n18246_), .B0(\asqrt[38] ), .Y(new_n18265_));
  OR4X1    g18073(.A(new_n17927_), .B(new_n17588_), .C(new_n17614_), .D(new_n17613_), .Y(new_n18266_));
  OR2X1    g18074(.A(new_n17588_), .B(new_n17613_), .Y(new_n18267_));
  OAI21X1  g18075(.A0(new_n18267_), .A1(new_n17927_), .B0(new_n17614_), .Y(new_n18268_));
  AND2X1   g18076(.A(new_n18268_), .B(new_n18266_), .Y(new_n18269_));
  NOR3X1   g18077(.A(new_n18264_), .B(new_n18246_), .C(\asqrt[38] ), .Y(new_n18270_));
  OAI21X1  g18078(.A0(new_n18270_), .A1(new_n18269_), .B0(new_n18265_), .Y(new_n18271_));
  AND2X1   g18079(.A(new_n18271_), .B(\asqrt[39] ), .Y(new_n18272_));
  OR2X1    g18080(.A(new_n18270_), .B(new_n18269_), .Y(new_n18273_));
  OAI21X1  g18081(.A0(new_n17632_), .A1(new_n17630_), .B0(new_n17596_), .Y(new_n18274_));
  NOR3X1   g18082(.A(new_n18274_), .B(new_n17927_), .C(new_n17590_), .Y(new_n18275_));
  AOI22X1  g18083(.A0(new_n17597_), .A1(new_n17591_), .B0(new_n17589_), .B1(\asqrt[38] ), .Y(new_n18276_));
  AOI21X1  g18084(.A0(new_n18276_), .A1(\asqrt[11] ), .B0(new_n17596_), .Y(new_n18277_));
  NOR2X1   g18085(.A(new_n18277_), .B(new_n18275_), .Y(new_n18278_));
  AND2X1   g18086(.A(new_n18265_), .B(new_n4165_), .Y(new_n18279_));
  AOI21X1  g18087(.A0(new_n18279_), .A1(new_n18273_), .B0(new_n18278_), .Y(new_n18280_));
  OAI21X1  g18088(.A0(new_n18280_), .A1(new_n18272_), .B0(\asqrt[40] ), .Y(new_n18281_));
  AND2X1   g18089(.A(new_n17635_), .B(new_n17633_), .Y(new_n18282_));
  OR4X1    g18090(.A(new_n17927_), .B(new_n18282_), .C(new_n17604_), .D(new_n17634_), .Y(new_n18283_));
  OR2X1    g18091(.A(new_n18282_), .B(new_n17634_), .Y(new_n18284_));
  OAI21X1  g18092(.A0(new_n18284_), .A1(new_n17927_), .B0(new_n17604_), .Y(new_n18285_));
  AND2X1   g18093(.A(new_n18285_), .B(new_n18283_), .Y(new_n18286_));
  INVX1    g18094(.A(new_n18286_), .Y(new_n18287_));
  AND2X1   g18095(.A(new_n18262_), .B(\asqrt[36] ), .Y(new_n18288_));
  NAND2X1  g18096(.A(new_n18234_), .B(new_n18233_), .Y(new_n18289_));
  NOR2X1   g18097(.A(new_n18228_), .B(\asqrt[36] ), .Y(new_n18290_));
  AOI21X1  g18098(.A0(new_n18290_), .A1(new_n18289_), .B0(new_n18242_), .Y(new_n18291_));
  OAI21X1  g18099(.A0(new_n18291_), .A1(new_n18288_), .B0(\asqrt[37] ), .Y(new_n18292_));
  INVX1    g18100(.A(new_n18251_), .Y(new_n18293_));
  OAI21X1  g18101(.A0(new_n18235_), .A1(new_n5176_), .B0(new_n4826_), .Y(new_n18294_));
  OAI21X1  g18102(.A0(new_n18294_), .A1(new_n18291_), .B0(new_n18293_), .Y(new_n18295_));
  AOI21X1  g18103(.A0(new_n18295_), .A1(new_n18292_), .B0(new_n4493_), .Y(new_n18296_));
  INVX1    g18104(.A(new_n18269_), .Y(new_n18297_));
  NAND3X1  g18105(.A(new_n18295_), .B(new_n18292_), .C(new_n4493_), .Y(new_n18298_));
  AOI21X1  g18106(.A0(new_n18298_), .A1(new_n18297_), .B0(new_n18296_), .Y(new_n18299_));
  OAI21X1  g18107(.A0(new_n18299_), .A1(new_n4165_), .B0(new_n3863_), .Y(new_n18300_));
  OAI21X1  g18108(.A0(new_n18300_), .A1(new_n18280_), .B0(new_n18287_), .Y(new_n18301_));
  AOI21X1  g18109(.A0(new_n18301_), .A1(new_n18281_), .B0(new_n3564_), .Y(new_n18302_));
  OR4X1    g18110(.A(new_n17927_), .B(new_n17637_), .C(new_n17625_), .D(new_n17619_), .Y(new_n18303_));
  OR2X1    g18111(.A(new_n17637_), .B(new_n17619_), .Y(new_n18304_));
  OAI21X1  g18112(.A0(new_n18304_), .A1(new_n17927_), .B0(new_n17625_), .Y(new_n18305_));
  AND2X1   g18113(.A(new_n18305_), .B(new_n18303_), .Y(new_n18306_));
  INVX1    g18114(.A(new_n18306_), .Y(new_n18307_));
  NAND3X1  g18115(.A(new_n18301_), .B(new_n18281_), .C(new_n3564_), .Y(new_n18308_));
  AOI21X1  g18116(.A0(new_n18308_), .A1(new_n18307_), .B0(new_n18302_), .Y(new_n18309_));
  OR2X1    g18117(.A(new_n18309_), .B(new_n3276_), .Y(new_n18310_));
  OR2X1    g18118(.A(new_n18299_), .B(new_n4165_), .Y(new_n18311_));
  NOR2X1   g18119(.A(new_n18270_), .B(new_n18269_), .Y(new_n18312_));
  INVX1    g18120(.A(new_n18278_), .Y(new_n18313_));
  NAND2X1  g18121(.A(new_n18265_), .B(new_n4165_), .Y(new_n18314_));
  OAI21X1  g18122(.A0(new_n18314_), .A1(new_n18312_), .B0(new_n18313_), .Y(new_n18315_));
  AOI21X1  g18123(.A0(new_n18315_), .A1(new_n18311_), .B0(new_n3863_), .Y(new_n18316_));
  AOI21X1  g18124(.A0(new_n18271_), .A1(\asqrt[39] ), .B0(\asqrt[40] ), .Y(new_n18317_));
  AOI21X1  g18125(.A0(new_n18317_), .A1(new_n18315_), .B0(new_n18286_), .Y(new_n18318_));
  NOR3X1   g18126(.A(new_n18318_), .B(new_n18316_), .C(\asqrt[41] ), .Y(new_n18319_));
  NOR2X1   g18127(.A(new_n18319_), .B(new_n18306_), .Y(new_n18320_));
  AND2X1   g18128(.A(new_n17681_), .B(new_n17680_), .Y(new_n18321_));
  NOR4X1   g18129(.A(new_n17927_), .B(new_n18321_), .C(new_n17644_), .D(new_n17679_), .Y(new_n18322_));
  AOI22X1  g18130(.A0(new_n17681_), .A1(new_n17680_), .B0(new_n17653_), .B1(\asqrt[41] ), .Y(new_n18323_));
  AOI21X1  g18131(.A0(new_n18323_), .A1(\asqrt[11] ), .B0(new_n17643_), .Y(new_n18324_));
  NOR2X1   g18132(.A(new_n18324_), .B(new_n18322_), .Y(new_n18325_));
  INVX1    g18133(.A(new_n18325_), .Y(new_n18326_));
  OAI21X1  g18134(.A0(new_n18318_), .A1(new_n18316_), .B0(\asqrt[41] ), .Y(new_n18327_));
  NAND2X1  g18135(.A(new_n18327_), .B(new_n3276_), .Y(new_n18328_));
  OAI21X1  g18136(.A0(new_n18328_), .A1(new_n18320_), .B0(new_n18326_), .Y(new_n18329_));
  AOI21X1  g18137(.A0(new_n18329_), .A1(new_n18310_), .B0(new_n3008_), .Y(new_n18330_));
  AND2X1   g18138(.A(new_n17654_), .B(new_n17647_), .Y(new_n18331_));
  OR4X1    g18139(.A(new_n17927_), .B(new_n18331_), .C(new_n17684_), .D(new_n17648_), .Y(new_n18332_));
  OR2X1    g18140(.A(new_n18331_), .B(new_n17648_), .Y(new_n18333_));
  OAI21X1  g18141(.A0(new_n18333_), .A1(new_n17927_), .B0(new_n17684_), .Y(new_n18334_));
  AND2X1   g18142(.A(new_n18334_), .B(new_n18332_), .Y(new_n18335_));
  OAI21X1  g18143(.A0(new_n18319_), .A1(new_n18306_), .B0(new_n18327_), .Y(new_n18336_));
  AOI21X1  g18144(.A0(new_n18336_), .A1(\asqrt[42] ), .B0(\asqrt[43] ), .Y(new_n18337_));
  AOI21X1  g18145(.A0(new_n18337_), .A1(new_n18329_), .B0(new_n18335_), .Y(new_n18338_));
  OAI21X1  g18146(.A0(new_n18338_), .A1(new_n18330_), .B0(\asqrt[44] ), .Y(new_n18339_));
  OR4X1    g18147(.A(new_n17927_), .B(new_n17662_), .C(new_n17688_), .D(new_n17687_), .Y(new_n18340_));
  OR2X1    g18148(.A(new_n17662_), .B(new_n17687_), .Y(new_n18341_));
  OAI21X1  g18149(.A0(new_n18341_), .A1(new_n17927_), .B0(new_n17688_), .Y(new_n18342_));
  AND2X1   g18150(.A(new_n18342_), .B(new_n18340_), .Y(new_n18343_));
  NOR3X1   g18151(.A(new_n18338_), .B(new_n18330_), .C(\asqrt[44] ), .Y(new_n18344_));
  OAI21X1  g18152(.A0(new_n18344_), .A1(new_n18343_), .B0(new_n18339_), .Y(new_n18345_));
  AND2X1   g18153(.A(new_n18345_), .B(\asqrt[45] ), .Y(new_n18346_));
  OR2X1    g18154(.A(new_n18344_), .B(new_n18343_), .Y(new_n18347_));
  OAI21X1  g18155(.A0(new_n17706_), .A1(new_n17704_), .B0(new_n17670_), .Y(new_n18348_));
  NOR3X1   g18156(.A(new_n18348_), .B(new_n17927_), .C(new_n17664_), .Y(new_n18349_));
  AOI22X1  g18157(.A0(new_n17671_), .A1(new_n17665_), .B0(new_n17663_), .B1(\asqrt[44] ), .Y(new_n18350_));
  AOI21X1  g18158(.A0(new_n18350_), .A1(\asqrt[11] ), .B0(new_n17670_), .Y(new_n18351_));
  NOR2X1   g18159(.A(new_n18351_), .B(new_n18349_), .Y(new_n18352_));
  AND2X1   g18160(.A(new_n18339_), .B(new_n2570_), .Y(new_n18353_));
  AOI21X1  g18161(.A0(new_n18353_), .A1(new_n18347_), .B0(new_n18352_), .Y(new_n18354_));
  OAI21X1  g18162(.A0(new_n18354_), .A1(new_n18346_), .B0(\asqrt[46] ), .Y(new_n18355_));
  AND2X1   g18163(.A(new_n17709_), .B(new_n17707_), .Y(new_n18356_));
  OR4X1    g18164(.A(new_n17927_), .B(new_n18356_), .C(new_n17678_), .D(new_n17708_), .Y(new_n18357_));
  OR2X1    g18165(.A(new_n18356_), .B(new_n17708_), .Y(new_n18358_));
  OAI21X1  g18166(.A0(new_n18358_), .A1(new_n17927_), .B0(new_n17678_), .Y(new_n18359_));
  AND2X1   g18167(.A(new_n18359_), .B(new_n18357_), .Y(new_n18360_));
  INVX1    g18168(.A(new_n18360_), .Y(new_n18361_));
  AND2X1   g18169(.A(new_n18336_), .B(\asqrt[42] ), .Y(new_n18362_));
  OR2X1    g18170(.A(new_n18319_), .B(new_n18306_), .Y(new_n18363_));
  AND2X1   g18171(.A(new_n18327_), .B(new_n3276_), .Y(new_n18364_));
  AOI21X1  g18172(.A0(new_n18364_), .A1(new_n18363_), .B0(new_n18325_), .Y(new_n18365_));
  OAI21X1  g18173(.A0(new_n18365_), .A1(new_n18362_), .B0(\asqrt[43] ), .Y(new_n18366_));
  INVX1    g18174(.A(new_n18335_), .Y(new_n18367_));
  OAI21X1  g18175(.A0(new_n18309_), .A1(new_n3276_), .B0(new_n3008_), .Y(new_n18368_));
  OAI21X1  g18176(.A0(new_n18368_), .A1(new_n18365_), .B0(new_n18367_), .Y(new_n18369_));
  AOI21X1  g18177(.A0(new_n18369_), .A1(new_n18366_), .B0(new_n2769_), .Y(new_n18370_));
  INVX1    g18178(.A(new_n18343_), .Y(new_n18371_));
  NAND3X1  g18179(.A(new_n18369_), .B(new_n18366_), .C(new_n2769_), .Y(new_n18372_));
  AOI21X1  g18180(.A0(new_n18372_), .A1(new_n18371_), .B0(new_n18370_), .Y(new_n18373_));
  OAI21X1  g18181(.A0(new_n18373_), .A1(new_n2570_), .B0(new_n2263_), .Y(new_n18374_));
  OAI21X1  g18182(.A0(new_n18374_), .A1(new_n18354_), .B0(new_n18361_), .Y(new_n18375_));
  AOI21X1  g18183(.A0(new_n18375_), .A1(new_n18355_), .B0(new_n2040_), .Y(new_n18376_));
  OR4X1    g18184(.A(new_n17927_), .B(new_n17711_), .C(new_n17699_), .D(new_n17693_), .Y(new_n18377_));
  OR2X1    g18185(.A(new_n17711_), .B(new_n17693_), .Y(new_n18378_));
  OAI21X1  g18186(.A0(new_n18378_), .A1(new_n17927_), .B0(new_n17699_), .Y(new_n18379_));
  AND2X1   g18187(.A(new_n18379_), .B(new_n18377_), .Y(new_n18380_));
  INVX1    g18188(.A(new_n18380_), .Y(new_n18381_));
  NAND3X1  g18189(.A(new_n18375_), .B(new_n18355_), .C(new_n2040_), .Y(new_n18382_));
  AOI21X1  g18190(.A0(new_n18382_), .A1(new_n18381_), .B0(new_n18376_), .Y(new_n18383_));
  OR2X1    g18191(.A(new_n18383_), .B(new_n1834_), .Y(new_n18384_));
  OR2X1    g18192(.A(new_n18373_), .B(new_n2570_), .Y(new_n18385_));
  NOR2X1   g18193(.A(new_n18344_), .B(new_n18343_), .Y(new_n18386_));
  INVX1    g18194(.A(new_n18352_), .Y(new_n18387_));
  NAND2X1  g18195(.A(new_n18339_), .B(new_n2570_), .Y(new_n18388_));
  OAI21X1  g18196(.A0(new_n18388_), .A1(new_n18386_), .B0(new_n18387_), .Y(new_n18389_));
  AOI21X1  g18197(.A0(new_n18389_), .A1(new_n18385_), .B0(new_n2263_), .Y(new_n18390_));
  AOI21X1  g18198(.A0(new_n18345_), .A1(\asqrt[45] ), .B0(\asqrt[46] ), .Y(new_n18391_));
  AOI21X1  g18199(.A0(new_n18391_), .A1(new_n18389_), .B0(new_n18360_), .Y(new_n18392_));
  NOR3X1   g18200(.A(new_n18392_), .B(new_n18390_), .C(\asqrt[47] ), .Y(new_n18393_));
  NOR2X1   g18201(.A(new_n18393_), .B(new_n18380_), .Y(new_n18394_));
  AND2X1   g18202(.A(new_n17755_), .B(new_n17754_), .Y(new_n18395_));
  NOR4X1   g18203(.A(new_n17927_), .B(new_n18395_), .C(new_n17718_), .D(new_n17753_), .Y(new_n18396_));
  AOI22X1  g18204(.A0(new_n17755_), .A1(new_n17754_), .B0(new_n17727_), .B1(\asqrt[47] ), .Y(new_n18397_));
  AOI21X1  g18205(.A0(new_n18397_), .A1(\asqrt[11] ), .B0(new_n17717_), .Y(new_n18398_));
  NOR2X1   g18206(.A(new_n18398_), .B(new_n18396_), .Y(new_n18399_));
  INVX1    g18207(.A(new_n18399_), .Y(new_n18400_));
  OAI21X1  g18208(.A0(new_n18392_), .A1(new_n18390_), .B0(\asqrt[47] ), .Y(new_n18401_));
  NAND2X1  g18209(.A(new_n18401_), .B(new_n1834_), .Y(new_n18402_));
  OAI21X1  g18210(.A0(new_n18402_), .A1(new_n18394_), .B0(new_n18400_), .Y(new_n18403_));
  AOI21X1  g18211(.A0(new_n18403_), .A1(new_n18384_), .B0(new_n1632_), .Y(new_n18404_));
  AND2X1   g18212(.A(new_n17728_), .B(new_n17721_), .Y(new_n18405_));
  OR4X1    g18213(.A(new_n17927_), .B(new_n18405_), .C(new_n17758_), .D(new_n17722_), .Y(new_n18406_));
  OR2X1    g18214(.A(new_n18405_), .B(new_n17722_), .Y(new_n18407_));
  OAI21X1  g18215(.A0(new_n18407_), .A1(new_n17927_), .B0(new_n17758_), .Y(new_n18408_));
  AND2X1   g18216(.A(new_n18408_), .B(new_n18406_), .Y(new_n18409_));
  OAI21X1  g18217(.A0(new_n18393_), .A1(new_n18380_), .B0(new_n18401_), .Y(new_n18410_));
  AOI21X1  g18218(.A0(new_n18410_), .A1(\asqrt[48] ), .B0(\asqrt[49] ), .Y(new_n18411_));
  AOI21X1  g18219(.A0(new_n18411_), .A1(new_n18403_), .B0(new_n18409_), .Y(new_n18412_));
  OAI21X1  g18220(.A0(new_n18412_), .A1(new_n18404_), .B0(\asqrt[50] ), .Y(new_n18413_));
  OR4X1    g18221(.A(new_n17927_), .B(new_n17736_), .C(new_n17762_), .D(new_n17761_), .Y(new_n18414_));
  OR2X1    g18222(.A(new_n17736_), .B(new_n17761_), .Y(new_n18415_));
  OAI21X1  g18223(.A0(new_n18415_), .A1(new_n17927_), .B0(new_n17762_), .Y(new_n18416_));
  AND2X1   g18224(.A(new_n18416_), .B(new_n18414_), .Y(new_n18417_));
  NOR3X1   g18225(.A(new_n18412_), .B(new_n18404_), .C(\asqrt[50] ), .Y(new_n18418_));
  OAI21X1  g18226(.A0(new_n18418_), .A1(new_n18417_), .B0(new_n18413_), .Y(new_n18419_));
  AND2X1   g18227(.A(new_n18419_), .B(\asqrt[51] ), .Y(new_n18420_));
  OR2X1    g18228(.A(new_n18418_), .B(new_n18417_), .Y(new_n18421_));
  OAI21X1  g18229(.A0(new_n17780_), .A1(new_n17778_), .B0(new_n17744_), .Y(new_n18422_));
  NOR3X1   g18230(.A(new_n18422_), .B(new_n17927_), .C(new_n17738_), .Y(new_n18423_));
  AOI22X1  g18231(.A0(new_n17745_), .A1(new_n17739_), .B0(new_n17737_), .B1(\asqrt[50] ), .Y(new_n18424_));
  AOI21X1  g18232(.A0(new_n18424_), .A1(\asqrt[11] ), .B0(new_n17744_), .Y(new_n18425_));
  NOR2X1   g18233(.A(new_n18425_), .B(new_n18423_), .Y(new_n18426_));
  AND2X1   g18234(.A(new_n18413_), .B(new_n1277_), .Y(new_n18427_));
  AOI21X1  g18235(.A0(new_n18427_), .A1(new_n18421_), .B0(new_n18426_), .Y(new_n18428_));
  OAI21X1  g18236(.A0(new_n18428_), .A1(new_n18420_), .B0(\asqrt[52] ), .Y(new_n18429_));
  AND2X1   g18237(.A(new_n17783_), .B(new_n17781_), .Y(new_n18430_));
  OR2X1    g18238(.A(new_n17752_), .B(new_n17782_), .Y(new_n18431_));
  OR2X1    g18239(.A(new_n18431_), .B(new_n18430_), .Y(new_n18432_));
  NOR3X1   g18240(.A(new_n17927_), .B(new_n18430_), .C(new_n17782_), .Y(new_n18433_));
  OAI22X1  g18241(.A0(new_n18433_), .A1(new_n17751_), .B0(new_n18432_), .B1(new_n17927_), .Y(new_n18434_));
  AND2X1   g18242(.A(new_n18410_), .B(\asqrt[48] ), .Y(new_n18435_));
  OR2X1    g18243(.A(new_n18393_), .B(new_n18380_), .Y(new_n18436_));
  AND2X1   g18244(.A(new_n18401_), .B(new_n1834_), .Y(new_n18437_));
  AOI21X1  g18245(.A0(new_n18437_), .A1(new_n18436_), .B0(new_n18399_), .Y(new_n18438_));
  OAI21X1  g18246(.A0(new_n18438_), .A1(new_n18435_), .B0(\asqrt[49] ), .Y(new_n18439_));
  INVX1    g18247(.A(new_n18409_), .Y(new_n18440_));
  OAI21X1  g18248(.A0(new_n18383_), .A1(new_n1834_), .B0(new_n1632_), .Y(new_n18441_));
  OAI21X1  g18249(.A0(new_n18441_), .A1(new_n18438_), .B0(new_n18440_), .Y(new_n18442_));
  AOI21X1  g18250(.A0(new_n18442_), .A1(new_n18439_), .B0(new_n1469_), .Y(new_n18443_));
  INVX1    g18251(.A(new_n18417_), .Y(new_n18444_));
  NAND3X1  g18252(.A(new_n18442_), .B(new_n18439_), .C(new_n1469_), .Y(new_n18445_));
  AOI21X1  g18253(.A0(new_n18445_), .A1(new_n18444_), .B0(new_n18443_), .Y(new_n18446_));
  OAI21X1  g18254(.A0(new_n18446_), .A1(new_n1277_), .B0(new_n1111_), .Y(new_n18447_));
  OAI21X1  g18255(.A0(new_n18447_), .A1(new_n18428_), .B0(new_n18434_), .Y(new_n18448_));
  AOI21X1  g18256(.A0(new_n18448_), .A1(new_n18429_), .B0(new_n968_), .Y(new_n18449_));
  OR4X1    g18257(.A(new_n17927_), .B(new_n17785_), .C(new_n17773_), .D(new_n17767_), .Y(new_n18450_));
  OR2X1    g18258(.A(new_n17785_), .B(new_n17767_), .Y(new_n18451_));
  OAI21X1  g18259(.A0(new_n18451_), .A1(new_n17927_), .B0(new_n17773_), .Y(new_n18452_));
  AND2X1   g18260(.A(new_n18452_), .B(new_n18450_), .Y(new_n18453_));
  INVX1    g18261(.A(new_n18453_), .Y(new_n18454_));
  NAND3X1  g18262(.A(new_n18448_), .B(new_n18429_), .C(new_n968_), .Y(new_n18455_));
  AOI21X1  g18263(.A0(new_n18455_), .A1(new_n18454_), .B0(new_n18449_), .Y(new_n18456_));
  OR2X1    g18264(.A(new_n18456_), .B(new_n902_), .Y(new_n18457_));
  OR2X1    g18265(.A(new_n18446_), .B(new_n1277_), .Y(new_n18458_));
  NOR2X1   g18266(.A(new_n18418_), .B(new_n18417_), .Y(new_n18459_));
  INVX1    g18267(.A(new_n18426_), .Y(new_n18460_));
  NAND2X1  g18268(.A(new_n18413_), .B(new_n1277_), .Y(new_n18461_));
  OAI21X1  g18269(.A0(new_n18461_), .A1(new_n18459_), .B0(new_n18460_), .Y(new_n18462_));
  AOI21X1  g18270(.A0(new_n18462_), .A1(new_n18458_), .B0(new_n1111_), .Y(new_n18463_));
  INVX1    g18271(.A(new_n18434_), .Y(new_n18464_));
  AOI21X1  g18272(.A0(new_n18419_), .A1(\asqrt[51] ), .B0(\asqrt[52] ), .Y(new_n18465_));
  AOI21X1  g18273(.A0(new_n18465_), .A1(new_n18462_), .B0(new_n18464_), .Y(new_n18466_));
  NOR3X1   g18274(.A(new_n18466_), .B(new_n18463_), .C(\asqrt[53] ), .Y(new_n18467_));
  NOR2X1   g18275(.A(new_n18467_), .B(new_n18453_), .Y(new_n18468_));
  OAI21X1  g18276(.A0(new_n18466_), .A1(new_n18463_), .B0(\asqrt[53] ), .Y(new_n18469_));
  NAND2X1  g18277(.A(new_n18469_), .B(new_n902_), .Y(new_n18470_));
  AND2X1   g18278(.A(new_n17829_), .B(new_n17828_), .Y(new_n18471_));
  NOR4X1   g18279(.A(new_n17927_), .B(new_n17794_), .C(new_n18471_), .D(new_n17827_), .Y(new_n18472_));
  AOI22X1  g18280(.A0(new_n17829_), .A1(new_n17828_), .B0(new_n17801_), .B1(\asqrt[53] ), .Y(new_n18473_));
  AOI21X1  g18281(.A0(new_n18473_), .A1(\asqrt[11] ), .B0(new_n17793_), .Y(new_n18474_));
  NOR2X1   g18282(.A(new_n18474_), .B(new_n18472_), .Y(new_n18475_));
  INVX1    g18283(.A(new_n18475_), .Y(new_n18476_));
  OAI21X1  g18284(.A0(new_n18470_), .A1(new_n18468_), .B0(new_n18476_), .Y(new_n18477_));
  AOI21X1  g18285(.A0(new_n18477_), .A1(new_n18457_), .B0(new_n697_), .Y(new_n18478_));
  OAI21X1  g18286(.A0(new_n17833_), .A1(new_n17830_), .B0(new_n17800_), .Y(new_n18479_));
  OR2X1    g18287(.A(new_n18479_), .B(new_n17796_), .Y(new_n18480_));
  AND2X1   g18288(.A(new_n17802_), .B(new_n17795_), .Y(new_n18481_));
  NOR3X1   g18289(.A(new_n17927_), .B(new_n18481_), .C(new_n17796_), .Y(new_n18482_));
  OAI22X1  g18290(.A0(new_n18482_), .A1(new_n17800_), .B0(new_n18480_), .B1(new_n17927_), .Y(new_n18483_));
  INVX1    g18291(.A(new_n18483_), .Y(new_n18484_));
  OAI21X1  g18292(.A0(new_n18467_), .A1(new_n18453_), .B0(new_n18469_), .Y(new_n18485_));
  AOI21X1  g18293(.A0(new_n18485_), .A1(\asqrt[54] ), .B0(\asqrt[55] ), .Y(new_n18486_));
  AOI21X1  g18294(.A0(new_n18486_), .A1(new_n18477_), .B0(new_n18484_), .Y(new_n18487_));
  OAI21X1  g18295(.A0(new_n18487_), .A1(new_n18478_), .B0(\asqrt[56] ), .Y(new_n18488_));
  OR4X1    g18296(.A(new_n17927_), .B(new_n17810_), .C(new_n17836_), .D(new_n17835_), .Y(new_n18489_));
  OR2X1    g18297(.A(new_n17810_), .B(new_n17835_), .Y(new_n18490_));
  OAI21X1  g18298(.A0(new_n18490_), .A1(new_n17927_), .B0(new_n17836_), .Y(new_n18491_));
  AND2X1   g18299(.A(new_n18491_), .B(new_n18489_), .Y(new_n18492_));
  NOR3X1   g18300(.A(new_n18487_), .B(new_n18478_), .C(\asqrt[56] ), .Y(new_n18493_));
  OAI21X1  g18301(.A0(new_n18493_), .A1(new_n18492_), .B0(new_n18488_), .Y(new_n18494_));
  AND2X1   g18302(.A(new_n18494_), .B(\asqrt[57] ), .Y(new_n18495_));
  OR2X1    g18303(.A(new_n18493_), .B(new_n18492_), .Y(new_n18496_));
  OAI21X1  g18304(.A0(new_n17854_), .A1(new_n17852_), .B0(new_n17818_), .Y(new_n18497_));
  NOR3X1   g18305(.A(new_n18497_), .B(new_n17927_), .C(new_n17812_), .Y(new_n18498_));
  AOI22X1  g18306(.A0(new_n17819_), .A1(new_n17813_), .B0(new_n17811_), .B1(\asqrt[56] ), .Y(new_n18499_));
  AOI21X1  g18307(.A0(new_n18499_), .A1(\asqrt[11] ), .B0(new_n17818_), .Y(new_n18500_));
  NOR2X1   g18308(.A(new_n18500_), .B(new_n18498_), .Y(new_n18501_));
  AND2X1   g18309(.A(new_n18488_), .B(new_n481_), .Y(new_n18502_));
  AOI21X1  g18310(.A0(new_n18502_), .A1(new_n18496_), .B0(new_n18501_), .Y(new_n18503_));
  OAI21X1  g18311(.A0(new_n18503_), .A1(new_n18495_), .B0(\asqrt[58] ), .Y(new_n18504_));
  AND2X1   g18312(.A(new_n17857_), .B(new_n17855_), .Y(new_n18505_));
  OR4X1    g18313(.A(new_n17927_), .B(new_n18505_), .C(new_n17826_), .D(new_n17856_), .Y(new_n18506_));
  OR2X1    g18314(.A(new_n18505_), .B(new_n17856_), .Y(new_n18507_));
  OAI21X1  g18315(.A0(new_n18507_), .A1(new_n17927_), .B0(new_n17826_), .Y(new_n18508_));
  AND2X1   g18316(.A(new_n18508_), .B(new_n18506_), .Y(new_n18509_));
  INVX1    g18317(.A(new_n18509_), .Y(new_n18510_));
  AND2X1   g18318(.A(new_n18485_), .B(\asqrt[54] ), .Y(new_n18511_));
  OR2X1    g18319(.A(new_n18467_), .B(new_n18453_), .Y(new_n18512_));
  AND2X1   g18320(.A(new_n18469_), .B(new_n902_), .Y(new_n18513_));
  AOI21X1  g18321(.A0(new_n18513_), .A1(new_n18512_), .B0(new_n18475_), .Y(new_n18514_));
  OAI21X1  g18322(.A0(new_n18514_), .A1(new_n18511_), .B0(\asqrt[55] ), .Y(new_n18515_));
  OAI21X1  g18323(.A0(new_n18456_), .A1(new_n902_), .B0(new_n697_), .Y(new_n18516_));
  OAI21X1  g18324(.A0(new_n18516_), .A1(new_n18514_), .B0(new_n18483_), .Y(new_n18517_));
  AOI21X1  g18325(.A0(new_n18517_), .A1(new_n18515_), .B0(new_n582_), .Y(new_n18518_));
  INVX1    g18326(.A(new_n18492_), .Y(new_n18519_));
  NAND3X1  g18327(.A(new_n18517_), .B(new_n18515_), .C(new_n582_), .Y(new_n18520_));
  AOI21X1  g18328(.A0(new_n18520_), .A1(new_n18519_), .B0(new_n18518_), .Y(new_n18521_));
  OAI21X1  g18329(.A0(new_n18521_), .A1(new_n481_), .B0(new_n399_), .Y(new_n18522_));
  OAI21X1  g18330(.A0(new_n18522_), .A1(new_n18503_), .B0(new_n18510_), .Y(new_n18523_));
  AOI21X1  g18331(.A0(new_n18523_), .A1(new_n18504_), .B0(new_n328_), .Y(new_n18524_));
  OR4X1    g18332(.A(new_n17927_), .B(new_n17859_), .C(new_n17847_), .D(new_n17841_), .Y(new_n18525_));
  OR2X1    g18333(.A(new_n17859_), .B(new_n17841_), .Y(new_n18526_));
  OAI21X1  g18334(.A0(new_n18526_), .A1(new_n17927_), .B0(new_n17847_), .Y(new_n18527_));
  AND2X1   g18335(.A(new_n18527_), .B(new_n18525_), .Y(new_n18528_));
  INVX1    g18336(.A(new_n18528_), .Y(new_n18529_));
  NAND3X1  g18337(.A(new_n18523_), .B(new_n18504_), .C(new_n328_), .Y(new_n18530_));
  AOI21X1  g18338(.A0(new_n18530_), .A1(new_n18529_), .B0(new_n18524_), .Y(new_n18531_));
  OR2X1    g18339(.A(new_n18531_), .B(new_n292_), .Y(new_n18532_));
  OR2X1    g18340(.A(new_n18521_), .B(new_n481_), .Y(new_n18533_));
  NOR2X1   g18341(.A(new_n18493_), .B(new_n18492_), .Y(new_n18534_));
  INVX1    g18342(.A(new_n18501_), .Y(new_n18535_));
  NAND2X1  g18343(.A(new_n18488_), .B(new_n481_), .Y(new_n18536_));
  OAI21X1  g18344(.A0(new_n18536_), .A1(new_n18534_), .B0(new_n18535_), .Y(new_n18537_));
  AOI21X1  g18345(.A0(new_n18537_), .A1(new_n18533_), .B0(new_n399_), .Y(new_n18538_));
  AOI21X1  g18346(.A0(new_n18494_), .A1(\asqrt[57] ), .B0(\asqrt[58] ), .Y(new_n18539_));
  AOI21X1  g18347(.A0(new_n18539_), .A1(new_n18537_), .B0(new_n18509_), .Y(new_n18540_));
  NOR3X1   g18348(.A(new_n18540_), .B(new_n18538_), .C(\asqrt[59] ), .Y(new_n18541_));
  NOR2X1   g18349(.A(new_n18541_), .B(new_n18528_), .Y(new_n18542_));
  AND2X1   g18350(.A(new_n17890_), .B(new_n17889_), .Y(new_n18543_));
  NOR4X1   g18351(.A(new_n17927_), .B(new_n18543_), .C(new_n17866_), .D(new_n17888_), .Y(new_n18544_));
  AOI22X1  g18352(.A0(new_n17890_), .A1(new_n17889_), .B0(new_n17875_), .B1(\asqrt[59] ), .Y(new_n18545_));
  AOI21X1  g18353(.A0(new_n18545_), .A1(\asqrt[11] ), .B0(new_n17865_), .Y(new_n18546_));
  NOR2X1   g18354(.A(new_n18546_), .B(new_n18544_), .Y(new_n18547_));
  INVX1    g18355(.A(new_n18547_), .Y(new_n18548_));
  OAI21X1  g18356(.A0(new_n18540_), .A1(new_n18538_), .B0(\asqrt[59] ), .Y(new_n18549_));
  NAND2X1  g18357(.A(new_n18549_), .B(new_n292_), .Y(new_n18550_));
  OAI21X1  g18358(.A0(new_n18550_), .A1(new_n18542_), .B0(new_n18548_), .Y(new_n18551_));
  AOI21X1  g18359(.A0(new_n18551_), .A1(new_n18532_), .B0(new_n217_), .Y(new_n18552_));
  AND2X1   g18360(.A(new_n17876_), .B(new_n17869_), .Y(new_n18553_));
  OR4X1    g18361(.A(new_n17927_), .B(new_n18553_), .C(new_n17893_), .D(new_n17870_), .Y(new_n18554_));
  OR2X1    g18362(.A(new_n18553_), .B(new_n17870_), .Y(new_n18555_));
  OAI21X1  g18363(.A0(new_n18555_), .A1(new_n17927_), .B0(new_n17893_), .Y(new_n18556_));
  AND2X1   g18364(.A(new_n18556_), .B(new_n18554_), .Y(new_n18557_));
  OAI21X1  g18365(.A0(new_n18541_), .A1(new_n18528_), .B0(new_n18549_), .Y(new_n18558_));
  AOI21X1  g18366(.A0(new_n18558_), .A1(\asqrt[60] ), .B0(\asqrt[61] ), .Y(new_n18559_));
  AOI21X1  g18367(.A0(new_n18559_), .A1(new_n18551_), .B0(new_n18557_), .Y(new_n18560_));
  OAI21X1  g18368(.A0(new_n18560_), .A1(new_n18552_), .B0(\asqrt[62] ), .Y(new_n18561_));
  OR4X1    g18369(.A(new_n17927_), .B(new_n17884_), .C(new_n17887_), .D(new_n17903_), .Y(new_n18562_));
  NAND2X1  g18370(.A(new_n17896_), .B(new_n17878_), .Y(new_n18563_));
  OAI21X1  g18371(.A0(new_n18563_), .A1(new_n17927_), .B0(new_n17887_), .Y(new_n18564_));
  AND2X1   g18372(.A(new_n18564_), .B(new_n18562_), .Y(new_n18565_));
  NOR3X1   g18373(.A(new_n18560_), .B(new_n18552_), .C(\asqrt[62] ), .Y(new_n18566_));
  OAI21X1  g18374(.A0(new_n18566_), .A1(new_n18565_), .B0(new_n18561_), .Y(new_n18567_));
  OAI21X1  g18375(.A0(new_n17947_), .A1(new_n17945_), .B0(new_n17902_), .Y(new_n18568_));
  NOR3X1   g18376(.A(new_n18568_), .B(new_n17927_), .C(new_n17886_), .Y(new_n18569_));
  AOI22X1  g18377(.A0(new_n17904_), .A1(new_n17897_), .B0(new_n17885_), .B1(\asqrt[62] ), .Y(new_n18570_));
  AOI21X1  g18378(.A0(new_n18570_), .A1(\asqrt[11] ), .B0(new_n17902_), .Y(new_n18571_));
  NOR2X1   g18379(.A(new_n18571_), .B(new_n18569_), .Y(new_n18572_));
  INVX1    g18380(.A(new_n18572_), .Y(new_n18573_));
  AND2X1   g18381(.A(new_n17951_), .B(new_n17948_), .Y(new_n18574_));
  AOI21X1  g18382(.A0(new_n17948_), .A1(new_n17944_), .B0(new_n17908_), .Y(new_n18575_));
  AOI21X1  g18383(.A0(new_n18575_), .A1(\asqrt[11] ), .B0(new_n18574_), .Y(new_n18576_));
  AND2X1   g18384(.A(new_n18576_), .B(new_n18573_), .Y(new_n18577_));
  AOI21X1  g18385(.A0(new_n18577_), .A1(new_n18567_), .B0(\asqrt[63] ), .Y(new_n18578_));
  NOR2X1   g18386(.A(new_n18566_), .B(new_n18565_), .Y(new_n18579_));
  NAND2X1  g18387(.A(new_n18572_), .B(new_n18561_), .Y(new_n18580_));
  AND2X1   g18388(.A(new_n17948_), .B(new_n17944_), .Y(new_n18581_));
  OAI21X1  g18389(.A0(new_n17927_), .A1(new_n17908_), .B0(new_n18581_), .Y(new_n18582_));
  NOR2X1   g18390(.A(new_n18575_), .B(new_n193_), .Y(new_n18583_));
  AND2X1   g18391(.A(new_n17915_), .B(new_n193_), .Y(new_n18584_));
  OR2X1    g18392(.A(new_n17923_), .B(new_n17906_), .Y(new_n18585_));
  AOI21X1  g18393(.A0(new_n17907_), .A1(new_n17273_), .B0(new_n18585_), .Y(new_n18586_));
  NAND2X1  g18394(.A(new_n18586_), .B(new_n17920_), .Y(new_n18587_));
  NOR3X1   g18395(.A(new_n18587_), .B(new_n18574_), .C(new_n18584_), .Y(new_n18588_));
  AOI21X1  g18396(.A0(new_n18583_), .A1(new_n18582_), .B0(new_n18588_), .Y(new_n18589_));
  OAI21X1  g18397(.A0(new_n18580_), .A1(new_n18579_), .B0(new_n18589_), .Y(new_n18590_));
  NOR2X1   g18398(.A(new_n18590_), .B(new_n18578_), .Y(new_n18591_));
  INVX1    g18399(.A(new_n18591_), .Y(\asqrt[10] ));
  OAI21X1  g18400(.A0(new_n18590_), .A1(new_n18578_), .B0(\a[20] ), .Y(new_n18593_));
  INVX1    g18401(.A(\a[20] ), .Y(new_n18594_));
  NOR2X1   g18402(.A(\a[19] ), .B(\a[18] ), .Y(new_n18595_));
  NAND2X1  g18403(.A(new_n18595_), .B(new_n18594_), .Y(new_n18596_));
  AOI21X1  g18404(.A0(new_n18596_), .A1(new_n18593_), .B0(new_n17927_), .Y(new_n18597_));
  AND2X1   g18405(.A(new_n18558_), .B(\asqrt[60] ), .Y(new_n18598_));
  OR2X1    g18406(.A(new_n18541_), .B(new_n18528_), .Y(new_n18599_));
  AND2X1   g18407(.A(new_n18549_), .B(new_n292_), .Y(new_n18600_));
  AOI21X1  g18408(.A0(new_n18600_), .A1(new_n18599_), .B0(new_n18547_), .Y(new_n18601_));
  OAI21X1  g18409(.A0(new_n18601_), .A1(new_n18598_), .B0(\asqrt[61] ), .Y(new_n18602_));
  INVX1    g18410(.A(new_n18557_), .Y(new_n18603_));
  OAI21X1  g18411(.A0(new_n18531_), .A1(new_n292_), .B0(new_n217_), .Y(new_n18604_));
  OAI21X1  g18412(.A0(new_n18604_), .A1(new_n18601_), .B0(new_n18603_), .Y(new_n18605_));
  AOI21X1  g18413(.A0(new_n18605_), .A1(new_n18602_), .B0(new_n199_), .Y(new_n18606_));
  INVX1    g18414(.A(new_n18565_), .Y(new_n18607_));
  NAND3X1  g18415(.A(new_n18605_), .B(new_n18602_), .C(new_n199_), .Y(new_n18608_));
  AOI21X1  g18416(.A0(new_n18608_), .A1(new_n18607_), .B0(new_n18606_), .Y(new_n18609_));
  INVX1    g18417(.A(new_n18577_), .Y(new_n18610_));
  OAI21X1  g18418(.A0(new_n18610_), .A1(new_n18609_), .B0(new_n193_), .Y(new_n18611_));
  OR2X1    g18419(.A(new_n18566_), .B(new_n18565_), .Y(new_n18612_));
  AND2X1   g18420(.A(new_n18572_), .B(new_n18561_), .Y(new_n18613_));
  INVX1    g18421(.A(new_n18589_), .Y(new_n18614_));
  AOI21X1  g18422(.A0(new_n18613_), .A1(new_n18612_), .B0(new_n18614_), .Y(new_n18615_));
  AOI21X1  g18423(.A0(new_n18615_), .A1(new_n18611_), .B0(new_n18594_), .Y(new_n18616_));
  NAND3X1  g18424(.A(new_n18596_), .B(new_n17924_), .C(new_n17920_), .Y(new_n18617_));
  OR4X1    g18425(.A(new_n18617_), .B(new_n18616_), .C(new_n18574_), .D(new_n18584_), .Y(new_n18618_));
  OAI21X1  g18426(.A0(new_n18590_), .A1(new_n18578_), .B0(new_n18594_), .Y(new_n18619_));
  AOI21X1  g18427(.A0(new_n18615_), .A1(new_n18611_), .B0(new_n17929_), .Y(new_n18620_));
  AOI21X1  g18428(.A0(new_n18619_), .A1(\a[21] ), .B0(new_n18620_), .Y(new_n18621_));
  AOI21X1  g18429(.A0(new_n18621_), .A1(new_n18618_), .B0(new_n18597_), .Y(new_n18622_));
  OR2X1    g18430(.A(new_n18622_), .B(new_n17262_), .Y(new_n18623_));
  AND2X1   g18431(.A(new_n18621_), .B(new_n18618_), .Y(new_n18624_));
  OR2X1    g18432(.A(new_n18597_), .B(\asqrt[12] ), .Y(new_n18625_));
  OAI21X1  g18433(.A0(new_n18590_), .A1(new_n18578_), .B0(new_n17928_), .Y(new_n18626_));
  AND2X1   g18434(.A(new_n18613_), .B(new_n18612_), .Y(new_n18627_));
  AND2X1   g18435(.A(new_n18583_), .B(new_n18582_), .Y(new_n18628_));
  OR2X1    g18436(.A(new_n18588_), .B(new_n17927_), .Y(new_n18629_));
  OR4X1    g18437(.A(new_n18629_), .B(new_n18628_), .C(new_n18627_), .D(new_n18578_), .Y(new_n18630_));
  AOI21X1  g18438(.A0(new_n18630_), .A1(new_n18626_), .B0(new_n17932_), .Y(new_n18631_));
  NOR4X1   g18439(.A(new_n18629_), .B(new_n18628_), .C(new_n18627_), .D(new_n18578_), .Y(new_n18632_));
  NOR3X1   g18440(.A(new_n18632_), .B(new_n18620_), .C(\a[22] ), .Y(new_n18633_));
  OR2X1    g18441(.A(new_n18633_), .B(new_n18631_), .Y(new_n18634_));
  OAI21X1  g18442(.A0(new_n18625_), .A1(new_n18624_), .B0(new_n18634_), .Y(new_n18635_));
  AOI21X1  g18443(.A0(new_n18635_), .A1(new_n18623_), .B0(new_n16617_), .Y(new_n18636_));
  AND2X1   g18444(.A(new_n17941_), .B(new_n17938_), .Y(new_n18637_));
  NOR3X1   g18445(.A(new_n18637_), .B(new_n17978_), .C(new_n17977_), .Y(new_n18638_));
  OAI21X1  g18446(.A0(new_n18590_), .A1(new_n18578_), .B0(new_n18638_), .Y(new_n18639_));
  AOI21X1  g18447(.A0(new_n17955_), .A1(\asqrt[12] ), .B0(new_n17978_), .Y(new_n18640_));
  OAI21X1  g18448(.A0(new_n18590_), .A1(new_n18578_), .B0(new_n18640_), .Y(new_n18641_));
  NAND2X1  g18449(.A(new_n18641_), .B(new_n18637_), .Y(new_n18642_));
  AND2X1   g18450(.A(new_n18596_), .B(new_n18593_), .Y(new_n18643_));
  NOR4X1   g18451(.A(new_n18617_), .B(new_n18616_), .C(new_n18574_), .D(new_n18584_), .Y(new_n18644_));
  INVX1    g18452(.A(\a[21] ), .Y(new_n18645_));
  AOI21X1  g18453(.A0(new_n18615_), .A1(new_n18611_), .B0(\a[20] ), .Y(new_n18646_));
  OAI21X1  g18454(.A0(new_n18646_), .A1(new_n18645_), .B0(new_n18626_), .Y(new_n18647_));
  OAI22X1  g18455(.A0(new_n18647_), .A1(new_n18644_), .B0(new_n18643_), .B1(new_n17927_), .Y(new_n18648_));
  AOI21X1  g18456(.A0(new_n18648_), .A1(\asqrt[12] ), .B0(\asqrt[13] ), .Y(new_n18649_));
  AOI22X1  g18457(.A0(new_n18649_), .A1(new_n18635_), .B0(new_n18642_), .B1(new_n18639_), .Y(new_n18650_));
  OAI21X1  g18458(.A0(new_n18650_), .A1(new_n18636_), .B0(\asqrt[14] ), .Y(new_n18651_));
  AND2X1   g18459(.A(new_n17956_), .B(new_n17942_), .Y(new_n18652_));
  NOR3X1   g18460(.A(new_n17984_), .B(new_n18652_), .C(new_n17943_), .Y(new_n18653_));
  OAI21X1  g18461(.A0(new_n18590_), .A1(new_n18578_), .B0(new_n18653_), .Y(new_n18654_));
  NOR2X1   g18462(.A(new_n18652_), .B(new_n17943_), .Y(new_n18655_));
  OAI21X1  g18463(.A0(new_n18590_), .A1(new_n18578_), .B0(new_n18655_), .Y(new_n18656_));
  NAND2X1  g18464(.A(new_n18656_), .B(new_n17984_), .Y(new_n18657_));
  AND2X1   g18465(.A(new_n18657_), .B(new_n18654_), .Y(new_n18658_));
  NOR3X1   g18466(.A(new_n18650_), .B(new_n18636_), .C(\asqrt[14] ), .Y(new_n18659_));
  OAI21X1  g18467(.A0(new_n18659_), .A1(new_n18658_), .B0(new_n18651_), .Y(new_n18660_));
  AND2X1   g18468(.A(new_n18660_), .B(\asqrt[15] ), .Y(new_n18661_));
  OR2X1    g18469(.A(new_n18659_), .B(new_n18658_), .Y(new_n18662_));
  NOR3X1   g18470(.A(new_n17973_), .B(new_n17976_), .C(new_n17995_), .Y(new_n18663_));
  NAND3X1  g18471(.A(\asqrt[10] ), .B(new_n17986_), .C(new_n17967_), .Y(new_n18664_));
  AOI22X1  g18472(.A0(new_n18664_), .A1(new_n17976_), .B0(new_n18663_), .B1(\asqrt[10] ), .Y(new_n18665_));
  AND2X1   g18473(.A(new_n18648_), .B(\asqrt[12] ), .Y(new_n18666_));
  NAND2X1  g18474(.A(new_n18621_), .B(new_n18618_), .Y(new_n18667_));
  NOR2X1   g18475(.A(new_n18597_), .B(\asqrt[12] ), .Y(new_n18668_));
  NOR2X1   g18476(.A(new_n18633_), .B(new_n18631_), .Y(new_n18669_));
  AOI21X1  g18477(.A0(new_n18668_), .A1(new_n18667_), .B0(new_n18669_), .Y(new_n18670_));
  OAI21X1  g18478(.A0(new_n18670_), .A1(new_n18666_), .B0(\asqrt[13] ), .Y(new_n18671_));
  NAND2X1  g18479(.A(new_n18642_), .B(new_n18639_), .Y(new_n18672_));
  OAI21X1  g18480(.A0(new_n18622_), .A1(new_n17262_), .B0(new_n16617_), .Y(new_n18673_));
  OAI21X1  g18481(.A0(new_n18673_), .A1(new_n18670_), .B0(new_n18672_), .Y(new_n18674_));
  AOI21X1  g18482(.A0(new_n18674_), .A1(new_n18671_), .B0(new_n15990_), .Y(new_n18675_));
  NOR2X1   g18483(.A(new_n18675_), .B(\asqrt[15] ), .Y(new_n18676_));
  AOI21X1  g18484(.A0(new_n18676_), .A1(new_n18662_), .B0(new_n18665_), .Y(new_n18677_));
  OAI21X1  g18485(.A0(new_n18677_), .A1(new_n18661_), .B0(\asqrt[16] ), .Y(new_n18678_));
  AOI21X1  g18486(.A0(new_n17996_), .A1(new_n17987_), .B0(new_n18032_), .Y(new_n18679_));
  AND2X1   g18487(.A(new_n18679_), .B(new_n18030_), .Y(new_n18680_));
  AOI22X1  g18488(.A0(new_n17996_), .A1(new_n17987_), .B0(new_n17974_), .B1(\asqrt[15] ), .Y(new_n18681_));
  AOI21X1  g18489(.A0(new_n18681_), .A1(\asqrt[10] ), .B0(new_n17994_), .Y(new_n18682_));
  AOI21X1  g18490(.A0(new_n18680_), .A1(\asqrt[10] ), .B0(new_n18682_), .Y(new_n18683_));
  INVX1    g18491(.A(new_n18683_), .Y(new_n18684_));
  INVX1    g18492(.A(new_n18658_), .Y(new_n18685_));
  NAND3X1  g18493(.A(new_n18674_), .B(new_n18671_), .C(new_n15990_), .Y(new_n18686_));
  AOI21X1  g18494(.A0(new_n18686_), .A1(new_n18685_), .B0(new_n18675_), .Y(new_n18687_));
  OAI21X1  g18495(.A0(new_n18687_), .A1(new_n15362_), .B0(new_n14754_), .Y(new_n18688_));
  OAI21X1  g18496(.A0(new_n18688_), .A1(new_n18677_), .B0(new_n18684_), .Y(new_n18689_));
  AOI21X1  g18497(.A0(new_n18689_), .A1(new_n18678_), .B0(new_n14165_), .Y(new_n18690_));
  AND2X1   g18498(.A(new_n18036_), .B(new_n18034_), .Y(new_n18691_));
  NOR3X1   g18499(.A(new_n18691_), .B(new_n18004_), .C(new_n18035_), .Y(new_n18692_));
  NOR3X1   g18500(.A(new_n18591_), .B(new_n18691_), .C(new_n18035_), .Y(new_n18693_));
  NOR2X1   g18501(.A(new_n18693_), .B(new_n18003_), .Y(new_n18694_));
  AOI21X1  g18502(.A0(new_n18692_), .A1(\asqrt[10] ), .B0(new_n18694_), .Y(new_n18695_));
  INVX1    g18503(.A(new_n18695_), .Y(new_n18696_));
  NAND3X1  g18504(.A(new_n18689_), .B(new_n18678_), .C(new_n14165_), .Y(new_n18697_));
  AOI21X1  g18505(.A0(new_n18697_), .A1(new_n18696_), .B0(new_n18690_), .Y(new_n18698_));
  OR2X1    g18506(.A(new_n18698_), .B(new_n13571_), .Y(new_n18699_));
  OR2X1    g18507(.A(new_n18687_), .B(new_n15362_), .Y(new_n18700_));
  NOR2X1   g18508(.A(new_n18659_), .B(new_n18658_), .Y(new_n18701_));
  INVX1    g18509(.A(new_n18665_), .Y(new_n18702_));
  OR2X1    g18510(.A(new_n18675_), .B(\asqrt[15] ), .Y(new_n18703_));
  OAI21X1  g18511(.A0(new_n18703_), .A1(new_n18701_), .B0(new_n18702_), .Y(new_n18704_));
  AOI21X1  g18512(.A0(new_n18704_), .A1(new_n18700_), .B0(new_n14754_), .Y(new_n18705_));
  AOI21X1  g18513(.A0(new_n18660_), .A1(\asqrt[15] ), .B0(\asqrt[16] ), .Y(new_n18706_));
  AOI21X1  g18514(.A0(new_n18706_), .A1(new_n18704_), .B0(new_n18683_), .Y(new_n18707_));
  NOR3X1   g18515(.A(new_n18707_), .B(new_n18705_), .C(\asqrt[17] ), .Y(new_n18708_));
  NOR2X1   g18516(.A(new_n18708_), .B(new_n18695_), .Y(new_n18709_));
  NOR3X1   g18517(.A(new_n18040_), .B(new_n18011_), .C(new_n18008_), .Y(new_n18710_));
  NOR3X1   g18518(.A(new_n18591_), .B(new_n18040_), .C(new_n18008_), .Y(new_n18711_));
  NOR2X1   g18519(.A(new_n18711_), .B(new_n18039_), .Y(new_n18712_));
  AOI21X1  g18520(.A0(new_n18710_), .A1(\asqrt[10] ), .B0(new_n18712_), .Y(new_n18713_));
  INVX1    g18521(.A(new_n18713_), .Y(new_n18714_));
  OAI21X1  g18522(.A0(new_n18707_), .A1(new_n18705_), .B0(\asqrt[17] ), .Y(new_n18715_));
  NAND2X1  g18523(.A(new_n18715_), .B(new_n13571_), .Y(new_n18716_));
  OAI21X1  g18524(.A0(new_n18716_), .A1(new_n18709_), .B0(new_n18714_), .Y(new_n18717_));
  AOI21X1  g18525(.A0(new_n18717_), .A1(new_n18699_), .B0(new_n13000_), .Y(new_n18718_));
  AND2X1   g18526(.A(new_n18055_), .B(new_n18054_), .Y(new_n18719_));
  NOR3X1   g18527(.A(new_n18719_), .B(new_n18021_), .C(new_n18053_), .Y(new_n18720_));
  NOR3X1   g18528(.A(new_n18591_), .B(new_n18719_), .C(new_n18053_), .Y(new_n18721_));
  NOR2X1   g18529(.A(new_n18721_), .B(new_n18020_), .Y(new_n18722_));
  AOI21X1  g18530(.A0(new_n18720_), .A1(\asqrt[10] ), .B0(new_n18722_), .Y(new_n18723_));
  OAI21X1  g18531(.A0(new_n18708_), .A1(new_n18695_), .B0(new_n18715_), .Y(new_n18724_));
  AOI21X1  g18532(.A0(new_n18724_), .A1(\asqrt[18] ), .B0(\asqrt[19] ), .Y(new_n18725_));
  AOI21X1  g18533(.A0(new_n18725_), .A1(new_n18717_), .B0(new_n18723_), .Y(new_n18726_));
  OAI21X1  g18534(.A0(new_n18726_), .A1(new_n18718_), .B0(\asqrt[20] ), .Y(new_n18727_));
  AND2X1   g18535(.A(new_n18042_), .B(new_n18023_), .Y(new_n18728_));
  NOR3X1   g18536(.A(new_n18728_), .B(new_n18058_), .C(new_n18024_), .Y(new_n18729_));
  NOR3X1   g18537(.A(new_n18591_), .B(new_n18728_), .C(new_n18024_), .Y(new_n18730_));
  NOR2X1   g18538(.A(new_n18730_), .B(new_n18029_), .Y(new_n18731_));
  AOI21X1  g18539(.A0(new_n18729_), .A1(\asqrt[10] ), .B0(new_n18731_), .Y(new_n18732_));
  NOR3X1   g18540(.A(new_n18726_), .B(new_n18718_), .C(\asqrt[20] ), .Y(new_n18733_));
  OAI21X1  g18541(.A0(new_n18733_), .A1(new_n18732_), .B0(new_n18727_), .Y(new_n18734_));
  AND2X1   g18542(.A(new_n18734_), .B(\asqrt[21] ), .Y(new_n18735_));
  OR2X1    g18543(.A(new_n18733_), .B(new_n18732_), .Y(new_n18736_));
  NAND4X1  g18544(.A(\asqrt[10] ), .B(new_n18061_), .C(new_n18048_), .D(new_n18044_), .Y(new_n18737_));
  NAND2X1  g18545(.A(new_n18061_), .B(new_n18044_), .Y(new_n18738_));
  OAI21X1  g18546(.A0(new_n18738_), .A1(new_n18591_), .B0(new_n18052_), .Y(new_n18739_));
  AND2X1   g18547(.A(new_n18739_), .B(new_n18737_), .Y(new_n18740_));
  AND2X1   g18548(.A(new_n18727_), .B(new_n11896_), .Y(new_n18741_));
  AOI21X1  g18549(.A0(new_n18741_), .A1(new_n18736_), .B0(new_n18740_), .Y(new_n18742_));
  OAI21X1  g18550(.A0(new_n18742_), .A1(new_n18735_), .B0(\asqrt[22] ), .Y(new_n18743_));
  AOI21X1  g18551(.A0(new_n18069_), .A1(new_n18062_), .B0(new_n18106_), .Y(new_n18744_));
  AND2X1   g18552(.A(new_n18744_), .B(new_n18104_), .Y(new_n18745_));
  AOI22X1  g18553(.A0(new_n18069_), .A1(new_n18062_), .B0(new_n18050_), .B1(\asqrt[21] ), .Y(new_n18746_));
  AOI21X1  g18554(.A0(new_n18746_), .A1(\asqrt[10] ), .B0(new_n18067_), .Y(new_n18747_));
  AOI21X1  g18555(.A0(new_n18745_), .A1(\asqrt[10] ), .B0(new_n18747_), .Y(new_n18748_));
  INVX1    g18556(.A(new_n18748_), .Y(new_n18749_));
  AND2X1   g18557(.A(new_n18724_), .B(\asqrt[18] ), .Y(new_n18750_));
  OR2X1    g18558(.A(new_n18708_), .B(new_n18695_), .Y(new_n18751_));
  AND2X1   g18559(.A(new_n18715_), .B(new_n13571_), .Y(new_n18752_));
  AOI21X1  g18560(.A0(new_n18752_), .A1(new_n18751_), .B0(new_n18713_), .Y(new_n18753_));
  OAI21X1  g18561(.A0(new_n18753_), .A1(new_n18750_), .B0(\asqrt[19] ), .Y(new_n18754_));
  INVX1    g18562(.A(new_n18723_), .Y(new_n18755_));
  OAI21X1  g18563(.A0(new_n18698_), .A1(new_n13571_), .B0(new_n13000_), .Y(new_n18756_));
  OAI21X1  g18564(.A0(new_n18756_), .A1(new_n18753_), .B0(new_n18755_), .Y(new_n18757_));
  AOI21X1  g18565(.A0(new_n18757_), .A1(new_n18754_), .B0(new_n12447_), .Y(new_n18758_));
  INVX1    g18566(.A(new_n18732_), .Y(new_n18759_));
  NAND3X1  g18567(.A(new_n18757_), .B(new_n18754_), .C(new_n12447_), .Y(new_n18760_));
  AOI21X1  g18568(.A0(new_n18760_), .A1(new_n18759_), .B0(new_n18758_), .Y(new_n18761_));
  OAI21X1  g18569(.A0(new_n18761_), .A1(new_n11896_), .B0(new_n11362_), .Y(new_n18762_));
  OAI21X1  g18570(.A0(new_n18762_), .A1(new_n18742_), .B0(new_n18749_), .Y(new_n18763_));
  AOI21X1  g18571(.A0(new_n18763_), .A1(new_n18743_), .B0(new_n10849_), .Y(new_n18764_));
  AND2X1   g18572(.A(new_n18110_), .B(new_n18108_), .Y(new_n18765_));
  NOR3X1   g18573(.A(new_n18765_), .B(new_n18077_), .C(new_n18109_), .Y(new_n18766_));
  NOR3X1   g18574(.A(new_n18591_), .B(new_n18765_), .C(new_n18109_), .Y(new_n18767_));
  NOR2X1   g18575(.A(new_n18767_), .B(new_n18076_), .Y(new_n18768_));
  AOI21X1  g18576(.A0(new_n18766_), .A1(\asqrt[10] ), .B0(new_n18768_), .Y(new_n18769_));
  INVX1    g18577(.A(new_n18769_), .Y(new_n18770_));
  NAND3X1  g18578(.A(new_n18763_), .B(new_n18743_), .C(new_n10849_), .Y(new_n18771_));
  AOI21X1  g18579(.A0(new_n18771_), .A1(new_n18770_), .B0(new_n18764_), .Y(new_n18772_));
  OR2X1    g18580(.A(new_n18772_), .B(new_n10332_), .Y(new_n18773_));
  AND2X1   g18581(.A(new_n18771_), .B(new_n18770_), .Y(new_n18774_));
  NAND4X1  g18582(.A(\asqrt[10] ), .B(new_n18085_), .C(new_n18113_), .D(new_n18112_), .Y(new_n18775_));
  NAND2X1  g18583(.A(new_n18085_), .B(new_n18112_), .Y(new_n18776_));
  OAI21X1  g18584(.A0(new_n18776_), .A1(new_n18591_), .B0(new_n18084_), .Y(new_n18777_));
  AND2X1   g18585(.A(new_n18777_), .B(new_n18775_), .Y(new_n18778_));
  INVX1    g18586(.A(new_n18778_), .Y(new_n18779_));
  OR2X1    g18587(.A(new_n18764_), .B(\asqrt[24] ), .Y(new_n18780_));
  OAI21X1  g18588(.A0(new_n18780_), .A1(new_n18774_), .B0(new_n18779_), .Y(new_n18781_));
  AOI21X1  g18589(.A0(new_n18781_), .A1(new_n18773_), .B0(new_n9833_), .Y(new_n18782_));
  AND2X1   g18590(.A(new_n18129_), .B(new_n18128_), .Y(new_n18783_));
  NOR3X1   g18591(.A(new_n18783_), .B(new_n18094_), .C(new_n18127_), .Y(new_n18784_));
  NOR3X1   g18592(.A(new_n18591_), .B(new_n18783_), .C(new_n18127_), .Y(new_n18785_));
  NOR2X1   g18593(.A(new_n18785_), .B(new_n18093_), .Y(new_n18786_));
  AOI21X1  g18594(.A0(new_n18784_), .A1(\asqrt[10] ), .B0(new_n18786_), .Y(new_n18787_));
  OR2X1    g18595(.A(new_n18761_), .B(new_n11896_), .Y(new_n18788_));
  NOR2X1   g18596(.A(new_n18733_), .B(new_n18732_), .Y(new_n18789_));
  INVX1    g18597(.A(new_n18740_), .Y(new_n18790_));
  NAND2X1  g18598(.A(new_n18727_), .B(new_n11896_), .Y(new_n18791_));
  OAI21X1  g18599(.A0(new_n18791_), .A1(new_n18789_), .B0(new_n18790_), .Y(new_n18792_));
  AOI21X1  g18600(.A0(new_n18792_), .A1(new_n18788_), .B0(new_n11362_), .Y(new_n18793_));
  AOI21X1  g18601(.A0(new_n18734_), .A1(\asqrt[21] ), .B0(\asqrt[22] ), .Y(new_n18794_));
  AOI21X1  g18602(.A0(new_n18794_), .A1(new_n18792_), .B0(new_n18748_), .Y(new_n18795_));
  OAI21X1  g18603(.A0(new_n18795_), .A1(new_n18793_), .B0(\asqrt[23] ), .Y(new_n18796_));
  NOR3X1   g18604(.A(new_n18795_), .B(new_n18793_), .C(\asqrt[23] ), .Y(new_n18797_));
  OAI21X1  g18605(.A0(new_n18797_), .A1(new_n18769_), .B0(new_n18796_), .Y(new_n18798_));
  AOI21X1  g18606(.A0(new_n18798_), .A1(\asqrt[24] ), .B0(\asqrt[25] ), .Y(new_n18799_));
  AOI21X1  g18607(.A0(new_n18799_), .A1(new_n18781_), .B0(new_n18787_), .Y(new_n18800_));
  OAI21X1  g18608(.A0(new_n18800_), .A1(new_n18782_), .B0(\asqrt[26] ), .Y(new_n18801_));
  AND2X1   g18609(.A(new_n18116_), .B(new_n18096_), .Y(new_n18802_));
  NOR3X1   g18610(.A(new_n18802_), .B(new_n18102_), .C(new_n18097_), .Y(new_n18803_));
  NOR3X1   g18611(.A(new_n18591_), .B(new_n18802_), .C(new_n18097_), .Y(new_n18804_));
  NOR2X1   g18612(.A(new_n18804_), .B(new_n18103_), .Y(new_n18805_));
  AOI21X1  g18613(.A0(new_n18803_), .A1(\asqrt[10] ), .B0(new_n18805_), .Y(new_n18806_));
  NOR3X1   g18614(.A(new_n18800_), .B(new_n18782_), .C(\asqrt[26] ), .Y(new_n18807_));
  OAI21X1  g18615(.A0(new_n18807_), .A1(new_n18806_), .B0(new_n18801_), .Y(new_n18808_));
  AND2X1   g18616(.A(new_n18808_), .B(\asqrt[27] ), .Y(new_n18809_));
  INVX1    g18617(.A(new_n18806_), .Y(new_n18810_));
  AND2X1   g18618(.A(new_n18798_), .B(\asqrt[24] ), .Y(new_n18811_));
  NAND2X1  g18619(.A(new_n18771_), .B(new_n18770_), .Y(new_n18812_));
  NOR2X1   g18620(.A(new_n18764_), .B(\asqrt[24] ), .Y(new_n18813_));
  AOI21X1  g18621(.A0(new_n18813_), .A1(new_n18812_), .B0(new_n18778_), .Y(new_n18814_));
  OAI21X1  g18622(.A0(new_n18814_), .A1(new_n18811_), .B0(\asqrt[25] ), .Y(new_n18815_));
  INVX1    g18623(.A(new_n18787_), .Y(new_n18816_));
  OAI21X1  g18624(.A0(new_n18772_), .A1(new_n10332_), .B0(new_n9833_), .Y(new_n18817_));
  OAI21X1  g18625(.A0(new_n18817_), .A1(new_n18814_), .B0(new_n18816_), .Y(new_n18818_));
  NAND3X1  g18626(.A(new_n18818_), .B(new_n18815_), .C(new_n9353_), .Y(new_n18819_));
  NAND2X1  g18627(.A(new_n18819_), .B(new_n18810_), .Y(new_n18820_));
  NAND4X1  g18628(.A(\asqrt[10] ), .B(new_n18134_), .C(new_n18122_), .D(new_n18118_), .Y(new_n18821_));
  NAND2X1  g18629(.A(new_n18134_), .B(new_n18118_), .Y(new_n18822_));
  OAI21X1  g18630(.A0(new_n18822_), .A1(new_n18591_), .B0(new_n18126_), .Y(new_n18823_));
  AND2X1   g18631(.A(new_n18823_), .B(new_n18821_), .Y(new_n18824_));
  AOI21X1  g18632(.A0(new_n18818_), .A1(new_n18815_), .B0(new_n9353_), .Y(new_n18825_));
  NOR2X1   g18633(.A(new_n18825_), .B(\asqrt[27] ), .Y(new_n18826_));
  AOI21X1  g18634(.A0(new_n18826_), .A1(new_n18820_), .B0(new_n18824_), .Y(new_n18827_));
  OAI21X1  g18635(.A0(new_n18827_), .A1(new_n18809_), .B0(\asqrt[28] ), .Y(new_n18828_));
  AOI21X1  g18636(.A0(new_n18142_), .A1(new_n18135_), .B0(new_n18179_), .Y(new_n18829_));
  AND2X1   g18637(.A(new_n18829_), .B(new_n18177_), .Y(new_n18830_));
  AOI22X1  g18638(.A0(new_n18142_), .A1(new_n18135_), .B0(new_n18124_), .B1(\asqrt[27] ), .Y(new_n18831_));
  AOI21X1  g18639(.A0(new_n18831_), .A1(\asqrt[10] ), .B0(new_n18140_), .Y(new_n18832_));
  AOI21X1  g18640(.A0(new_n18830_), .A1(\asqrt[10] ), .B0(new_n18832_), .Y(new_n18833_));
  INVX1    g18641(.A(new_n18833_), .Y(new_n18834_));
  AOI21X1  g18642(.A0(new_n18819_), .A1(new_n18810_), .B0(new_n18825_), .Y(new_n18835_));
  OAI21X1  g18643(.A0(new_n18835_), .A1(new_n8874_), .B0(new_n8412_), .Y(new_n18836_));
  OAI21X1  g18644(.A0(new_n18836_), .A1(new_n18827_), .B0(new_n18834_), .Y(new_n18837_));
  AOI21X1  g18645(.A0(new_n18837_), .A1(new_n18828_), .B0(new_n7970_), .Y(new_n18838_));
  AND2X1   g18646(.A(new_n18184_), .B(new_n18181_), .Y(new_n18839_));
  NOR3X1   g18647(.A(new_n18839_), .B(new_n18149_), .C(new_n18182_), .Y(new_n18840_));
  NOR3X1   g18648(.A(new_n18591_), .B(new_n18839_), .C(new_n18182_), .Y(new_n18841_));
  NOR2X1   g18649(.A(new_n18841_), .B(new_n18183_), .Y(new_n18842_));
  AOI21X1  g18650(.A0(new_n18840_), .A1(\asqrt[10] ), .B0(new_n18842_), .Y(new_n18843_));
  INVX1    g18651(.A(new_n18843_), .Y(new_n18844_));
  NAND3X1  g18652(.A(new_n18837_), .B(new_n18828_), .C(new_n7970_), .Y(new_n18845_));
  AOI21X1  g18653(.A0(new_n18845_), .A1(new_n18844_), .B0(new_n18838_), .Y(new_n18846_));
  OR2X1    g18654(.A(new_n18846_), .B(new_n7527_), .Y(new_n18847_));
  OR2X1    g18655(.A(new_n18835_), .B(new_n8874_), .Y(new_n18848_));
  AND2X1   g18656(.A(new_n18819_), .B(new_n18810_), .Y(new_n18849_));
  INVX1    g18657(.A(new_n18824_), .Y(new_n18850_));
  OR2X1    g18658(.A(new_n18825_), .B(\asqrt[27] ), .Y(new_n18851_));
  OAI21X1  g18659(.A0(new_n18851_), .A1(new_n18849_), .B0(new_n18850_), .Y(new_n18852_));
  AOI21X1  g18660(.A0(new_n18852_), .A1(new_n18848_), .B0(new_n8412_), .Y(new_n18853_));
  AOI21X1  g18661(.A0(new_n18808_), .A1(\asqrt[27] ), .B0(\asqrt[28] ), .Y(new_n18854_));
  AOI21X1  g18662(.A0(new_n18854_), .A1(new_n18852_), .B0(new_n18833_), .Y(new_n18855_));
  NOR3X1   g18663(.A(new_n18855_), .B(new_n18853_), .C(\asqrt[29] ), .Y(new_n18856_));
  NOR2X1   g18664(.A(new_n18856_), .B(new_n18843_), .Y(new_n18857_));
  OR4X1    g18665(.A(new_n18591_), .B(new_n18187_), .C(new_n18158_), .D(new_n18153_), .Y(new_n18858_));
  OR2X1    g18666(.A(new_n18187_), .B(new_n18153_), .Y(new_n18859_));
  OAI21X1  g18667(.A0(new_n18859_), .A1(new_n18591_), .B0(new_n18158_), .Y(new_n18860_));
  AND2X1   g18668(.A(new_n18860_), .B(new_n18858_), .Y(new_n18861_));
  INVX1    g18669(.A(new_n18861_), .Y(new_n18862_));
  OAI21X1  g18670(.A0(new_n18855_), .A1(new_n18853_), .B0(\asqrt[29] ), .Y(new_n18863_));
  NAND2X1  g18671(.A(new_n18863_), .B(new_n7527_), .Y(new_n18864_));
  OAI21X1  g18672(.A0(new_n18864_), .A1(new_n18857_), .B0(new_n18862_), .Y(new_n18865_));
  AOI21X1  g18673(.A0(new_n18865_), .A1(new_n18847_), .B0(new_n7103_), .Y(new_n18866_));
  AND2X1   g18674(.A(new_n18202_), .B(new_n18201_), .Y(new_n18867_));
  NOR3X1   g18675(.A(new_n18867_), .B(new_n18168_), .C(new_n18200_), .Y(new_n18868_));
  NOR3X1   g18676(.A(new_n18591_), .B(new_n18867_), .C(new_n18200_), .Y(new_n18869_));
  NOR2X1   g18677(.A(new_n18869_), .B(new_n18167_), .Y(new_n18870_));
  AOI21X1  g18678(.A0(new_n18868_), .A1(\asqrt[10] ), .B0(new_n18870_), .Y(new_n18871_));
  OAI21X1  g18679(.A0(new_n18856_), .A1(new_n18843_), .B0(new_n18863_), .Y(new_n18872_));
  AOI21X1  g18680(.A0(new_n18872_), .A1(\asqrt[30] ), .B0(\asqrt[31] ), .Y(new_n18873_));
  AOI21X1  g18681(.A0(new_n18873_), .A1(new_n18865_), .B0(new_n18871_), .Y(new_n18874_));
  OAI21X1  g18682(.A0(new_n18874_), .A1(new_n18866_), .B0(\asqrt[32] ), .Y(new_n18875_));
  AND2X1   g18683(.A(new_n18189_), .B(new_n18170_), .Y(new_n18876_));
  NOR3X1   g18684(.A(new_n18876_), .B(new_n18205_), .C(new_n18171_), .Y(new_n18877_));
  NOR3X1   g18685(.A(new_n18591_), .B(new_n18876_), .C(new_n18171_), .Y(new_n18878_));
  NOR2X1   g18686(.A(new_n18878_), .B(new_n18176_), .Y(new_n18879_));
  AOI21X1  g18687(.A0(new_n18877_), .A1(\asqrt[10] ), .B0(new_n18879_), .Y(new_n18880_));
  NOR3X1   g18688(.A(new_n18874_), .B(new_n18866_), .C(\asqrt[32] ), .Y(new_n18881_));
  OAI21X1  g18689(.A0(new_n18881_), .A1(new_n18880_), .B0(new_n18875_), .Y(new_n18882_));
  AND2X1   g18690(.A(new_n18882_), .B(\asqrt[33] ), .Y(new_n18883_));
  OR2X1    g18691(.A(new_n18881_), .B(new_n18880_), .Y(new_n18884_));
  OR4X1    g18692(.A(new_n18591_), .B(new_n18196_), .C(new_n18199_), .D(new_n18224_), .Y(new_n18885_));
  OR2X1    g18693(.A(new_n18196_), .B(new_n18224_), .Y(new_n18886_));
  OAI21X1  g18694(.A0(new_n18886_), .A1(new_n18591_), .B0(new_n18199_), .Y(new_n18887_));
  AND2X1   g18695(.A(new_n18887_), .B(new_n18885_), .Y(new_n18888_));
  AND2X1   g18696(.A(new_n18875_), .B(new_n6294_), .Y(new_n18889_));
  AOI21X1  g18697(.A0(new_n18889_), .A1(new_n18884_), .B0(new_n18888_), .Y(new_n18890_));
  OAI21X1  g18698(.A0(new_n18890_), .A1(new_n18883_), .B0(\asqrt[34] ), .Y(new_n18891_));
  AOI21X1  g18699(.A0(new_n18215_), .A1(new_n18209_), .B0(new_n18254_), .Y(new_n18892_));
  AND2X1   g18700(.A(new_n18892_), .B(new_n18252_), .Y(new_n18893_));
  AOI22X1  g18701(.A0(new_n18215_), .A1(new_n18209_), .B0(new_n18197_), .B1(\asqrt[33] ), .Y(new_n18894_));
  AOI21X1  g18702(.A0(new_n18894_), .A1(\asqrt[10] ), .B0(new_n18214_), .Y(new_n18895_));
  AOI21X1  g18703(.A0(new_n18893_), .A1(\asqrt[10] ), .B0(new_n18895_), .Y(new_n18896_));
  INVX1    g18704(.A(new_n18896_), .Y(new_n18897_));
  AND2X1   g18705(.A(new_n18872_), .B(\asqrt[30] ), .Y(new_n18898_));
  OR2X1    g18706(.A(new_n18856_), .B(new_n18843_), .Y(new_n18899_));
  AND2X1   g18707(.A(new_n18863_), .B(new_n7527_), .Y(new_n18900_));
  AOI21X1  g18708(.A0(new_n18900_), .A1(new_n18899_), .B0(new_n18861_), .Y(new_n18901_));
  OAI21X1  g18709(.A0(new_n18901_), .A1(new_n18898_), .B0(\asqrt[31] ), .Y(new_n18902_));
  INVX1    g18710(.A(new_n18871_), .Y(new_n18903_));
  OAI21X1  g18711(.A0(new_n18846_), .A1(new_n7527_), .B0(new_n7103_), .Y(new_n18904_));
  OAI21X1  g18712(.A0(new_n18904_), .A1(new_n18901_), .B0(new_n18903_), .Y(new_n18905_));
  AOI21X1  g18713(.A0(new_n18905_), .A1(new_n18902_), .B0(new_n6699_), .Y(new_n18906_));
  INVX1    g18714(.A(new_n18880_), .Y(new_n18907_));
  NAND3X1  g18715(.A(new_n18905_), .B(new_n18902_), .C(new_n6699_), .Y(new_n18908_));
  AOI21X1  g18716(.A0(new_n18908_), .A1(new_n18907_), .B0(new_n18906_), .Y(new_n18909_));
  OAI21X1  g18717(.A0(new_n18909_), .A1(new_n6294_), .B0(new_n5941_), .Y(new_n18910_));
  OAI21X1  g18718(.A0(new_n18910_), .A1(new_n18890_), .B0(new_n18897_), .Y(new_n18911_));
  AOI21X1  g18719(.A0(new_n18911_), .A1(new_n18891_), .B0(new_n5541_), .Y(new_n18912_));
  AND2X1   g18720(.A(new_n18258_), .B(new_n18256_), .Y(new_n18913_));
  NOR3X1   g18721(.A(new_n18913_), .B(new_n18223_), .C(new_n18257_), .Y(new_n18914_));
  NOR3X1   g18722(.A(new_n18591_), .B(new_n18913_), .C(new_n18257_), .Y(new_n18915_));
  NOR2X1   g18723(.A(new_n18915_), .B(new_n18222_), .Y(new_n18916_));
  AOI21X1  g18724(.A0(new_n18914_), .A1(\asqrt[10] ), .B0(new_n18916_), .Y(new_n18917_));
  INVX1    g18725(.A(new_n18917_), .Y(new_n18918_));
  NAND3X1  g18726(.A(new_n18911_), .B(new_n18891_), .C(new_n5541_), .Y(new_n18919_));
  AOI21X1  g18727(.A0(new_n18919_), .A1(new_n18918_), .B0(new_n18912_), .Y(new_n18920_));
  OR2X1    g18728(.A(new_n18920_), .B(new_n5176_), .Y(new_n18921_));
  AND2X1   g18729(.A(new_n18919_), .B(new_n18918_), .Y(new_n18922_));
  NAND4X1  g18730(.A(\asqrt[10] ), .B(new_n18234_), .C(new_n18232_), .D(new_n18260_), .Y(new_n18923_));
  NAND2X1  g18731(.A(new_n18234_), .B(new_n18260_), .Y(new_n18924_));
  OAI21X1  g18732(.A0(new_n18924_), .A1(new_n18591_), .B0(new_n18233_), .Y(new_n18925_));
  AND2X1   g18733(.A(new_n18925_), .B(new_n18923_), .Y(new_n18926_));
  INVX1    g18734(.A(new_n18926_), .Y(new_n18927_));
  OR2X1    g18735(.A(new_n18912_), .B(\asqrt[36] ), .Y(new_n18928_));
  OAI21X1  g18736(.A0(new_n18928_), .A1(new_n18922_), .B0(new_n18927_), .Y(new_n18929_));
  AOI21X1  g18737(.A0(new_n18929_), .A1(new_n18921_), .B0(new_n4826_), .Y(new_n18930_));
  AND2X1   g18738(.A(new_n18290_), .B(new_n18289_), .Y(new_n18931_));
  NOR3X1   g18739(.A(new_n18931_), .B(new_n18243_), .C(new_n18288_), .Y(new_n18932_));
  NOR3X1   g18740(.A(new_n18591_), .B(new_n18931_), .C(new_n18288_), .Y(new_n18933_));
  NOR2X1   g18741(.A(new_n18933_), .B(new_n18242_), .Y(new_n18934_));
  AOI21X1  g18742(.A0(new_n18932_), .A1(\asqrt[10] ), .B0(new_n18934_), .Y(new_n18935_));
  OR2X1    g18743(.A(new_n18909_), .B(new_n6294_), .Y(new_n18936_));
  NOR2X1   g18744(.A(new_n18881_), .B(new_n18880_), .Y(new_n18937_));
  INVX1    g18745(.A(new_n18888_), .Y(new_n18938_));
  NAND2X1  g18746(.A(new_n18875_), .B(new_n6294_), .Y(new_n18939_));
  OAI21X1  g18747(.A0(new_n18939_), .A1(new_n18937_), .B0(new_n18938_), .Y(new_n18940_));
  AOI21X1  g18748(.A0(new_n18940_), .A1(new_n18936_), .B0(new_n5941_), .Y(new_n18941_));
  AOI21X1  g18749(.A0(new_n18882_), .A1(\asqrt[33] ), .B0(\asqrt[34] ), .Y(new_n18942_));
  AOI21X1  g18750(.A0(new_n18942_), .A1(new_n18940_), .B0(new_n18896_), .Y(new_n18943_));
  OAI21X1  g18751(.A0(new_n18943_), .A1(new_n18941_), .B0(\asqrt[35] ), .Y(new_n18944_));
  NOR3X1   g18752(.A(new_n18943_), .B(new_n18941_), .C(\asqrt[35] ), .Y(new_n18945_));
  OAI21X1  g18753(.A0(new_n18945_), .A1(new_n18917_), .B0(new_n18944_), .Y(new_n18946_));
  AOI21X1  g18754(.A0(new_n18946_), .A1(\asqrt[36] ), .B0(\asqrt[37] ), .Y(new_n18947_));
  AOI21X1  g18755(.A0(new_n18947_), .A1(new_n18929_), .B0(new_n18935_), .Y(new_n18948_));
  OAI21X1  g18756(.A0(new_n18948_), .A1(new_n18930_), .B0(\asqrt[38] ), .Y(new_n18949_));
  AND2X1   g18757(.A(new_n18263_), .B(new_n18245_), .Y(new_n18950_));
  NOR3X1   g18758(.A(new_n18950_), .B(new_n18293_), .C(new_n18246_), .Y(new_n18951_));
  NOR3X1   g18759(.A(new_n18591_), .B(new_n18950_), .C(new_n18246_), .Y(new_n18952_));
  NOR2X1   g18760(.A(new_n18952_), .B(new_n18251_), .Y(new_n18953_));
  AOI21X1  g18761(.A0(new_n18951_), .A1(\asqrt[10] ), .B0(new_n18953_), .Y(new_n18954_));
  NOR3X1   g18762(.A(new_n18948_), .B(new_n18930_), .C(\asqrt[38] ), .Y(new_n18955_));
  OAI21X1  g18763(.A0(new_n18955_), .A1(new_n18954_), .B0(new_n18949_), .Y(new_n18956_));
  AND2X1   g18764(.A(new_n18956_), .B(\asqrt[39] ), .Y(new_n18957_));
  OR2X1    g18765(.A(new_n18955_), .B(new_n18954_), .Y(new_n18958_));
  OR4X1    g18766(.A(new_n18591_), .B(new_n18270_), .C(new_n18297_), .D(new_n18296_), .Y(new_n18959_));
  OR2X1    g18767(.A(new_n18270_), .B(new_n18296_), .Y(new_n18960_));
  OAI21X1  g18768(.A0(new_n18960_), .A1(new_n18591_), .B0(new_n18297_), .Y(new_n18961_));
  AND2X1   g18769(.A(new_n18961_), .B(new_n18959_), .Y(new_n18962_));
  AND2X1   g18770(.A(new_n18949_), .B(new_n4165_), .Y(new_n18963_));
  AOI21X1  g18771(.A0(new_n18963_), .A1(new_n18958_), .B0(new_n18962_), .Y(new_n18964_));
  OAI21X1  g18772(.A0(new_n18964_), .A1(new_n18957_), .B0(\asqrt[40] ), .Y(new_n18965_));
  AOI21X1  g18773(.A0(new_n18279_), .A1(new_n18273_), .B0(new_n18313_), .Y(new_n18966_));
  AND2X1   g18774(.A(new_n18966_), .B(new_n18311_), .Y(new_n18967_));
  AOI22X1  g18775(.A0(new_n18279_), .A1(new_n18273_), .B0(new_n18271_), .B1(\asqrt[39] ), .Y(new_n18968_));
  AOI21X1  g18776(.A0(new_n18968_), .A1(\asqrt[10] ), .B0(new_n18278_), .Y(new_n18969_));
  AOI21X1  g18777(.A0(new_n18967_), .A1(\asqrt[10] ), .B0(new_n18969_), .Y(new_n18970_));
  INVX1    g18778(.A(new_n18970_), .Y(new_n18971_));
  AND2X1   g18779(.A(new_n18946_), .B(\asqrt[36] ), .Y(new_n18972_));
  NAND2X1  g18780(.A(new_n18919_), .B(new_n18918_), .Y(new_n18973_));
  NOR2X1   g18781(.A(new_n18912_), .B(\asqrt[36] ), .Y(new_n18974_));
  AOI21X1  g18782(.A0(new_n18974_), .A1(new_n18973_), .B0(new_n18926_), .Y(new_n18975_));
  OAI21X1  g18783(.A0(new_n18975_), .A1(new_n18972_), .B0(\asqrt[37] ), .Y(new_n18976_));
  INVX1    g18784(.A(new_n18935_), .Y(new_n18977_));
  OAI21X1  g18785(.A0(new_n18920_), .A1(new_n5176_), .B0(new_n4826_), .Y(new_n18978_));
  OAI21X1  g18786(.A0(new_n18978_), .A1(new_n18975_), .B0(new_n18977_), .Y(new_n18979_));
  AOI21X1  g18787(.A0(new_n18979_), .A1(new_n18976_), .B0(new_n4493_), .Y(new_n18980_));
  INVX1    g18788(.A(new_n18954_), .Y(new_n18981_));
  NAND3X1  g18789(.A(new_n18979_), .B(new_n18976_), .C(new_n4493_), .Y(new_n18982_));
  AOI21X1  g18790(.A0(new_n18982_), .A1(new_n18981_), .B0(new_n18980_), .Y(new_n18983_));
  OAI21X1  g18791(.A0(new_n18983_), .A1(new_n4165_), .B0(new_n3863_), .Y(new_n18984_));
  OAI21X1  g18792(.A0(new_n18984_), .A1(new_n18964_), .B0(new_n18971_), .Y(new_n18985_));
  AOI21X1  g18793(.A0(new_n18985_), .A1(new_n18965_), .B0(new_n3564_), .Y(new_n18986_));
  AND2X1   g18794(.A(new_n18317_), .B(new_n18315_), .Y(new_n18987_));
  NOR3X1   g18795(.A(new_n18987_), .B(new_n18287_), .C(new_n18316_), .Y(new_n18988_));
  NOR3X1   g18796(.A(new_n18591_), .B(new_n18987_), .C(new_n18316_), .Y(new_n18989_));
  NOR2X1   g18797(.A(new_n18989_), .B(new_n18286_), .Y(new_n18990_));
  AOI21X1  g18798(.A0(new_n18988_), .A1(\asqrt[10] ), .B0(new_n18990_), .Y(new_n18991_));
  INVX1    g18799(.A(new_n18991_), .Y(new_n18992_));
  NAND3X1  g18800(.A(new_n18985_), .B(new_n18965_), .C(new_n3564_), .Y(new_n18993_));
  AOI21X1  g18801(.A0(new_n18993_), .A1(new_n18992_), .B0(new_n18986_), .Y(new_n18994_));
  OR2X1    g18802(.A(new_n18994_), .B(new_n3276_), .Y(new_n18995_));
  OR2X1    g18803(.A(new_n18983_), .B(new_n4165_), .Y(new_n18996_));
  NOR2X1   g18804(.A(new_n18955_), .B(new_n18954_), .Y(new_n18997_));
  INVX1    g18805(.A(new_n18962_), .Y(new_n18998_));
  NAND2X1  g18806(.A(new_n18949_), .B(new_n4165_), .Y(new_n18999_));
  OAI21X1  g18807(.A0(new_n18999_), .A1(new_n18997_), .B0(new_n18998_), .Y(new_n19000_));
  AOI21X1  g18808(.A0(new_n19000_), .A1(new_n18996_), .B0(new_n3863_), .Y(new_n19001_));
  AOI21X1  g18809(.A0(new_n18956_), .A1(\asqrt[39] ), .B0(\asqrt[40] ), .Y(new_n19002_));
  AOI21X1  g18810(.A0(new_n19002_), .A1(new_n19000_), .B0(new_n18970_), .Y(new_n19003_));
  NOR3X1   g18811(.A(new_n19003_), .B(new_n19001_), .C(\asqrt[41] ), .Y(new_n19004_));
  NOR2X1   g18812(.A(new_n19004_), .B(new_n18991_), .Y(new_n19005_));
  OR4X1    g18813(.A(new_n18591_), .B(new_n18319_), .C(new_n18307_), .D(new_n18302_), .Y(new_n19006_));
  OR2X1    g18814(.A(new_n18319_), .B(new_n18302_), .Y(new_n19007_));
  OAI21X1  g18815(.A0(new_n19007_), .A1(new_n18591_), .B0(new_n18307_), .Y(new_n19008_));
  AND2X1   g18816(.A(new_n19008_), .B(new_n19006_), .Y(new_n19009_));
  INVX1    g18817(.A(new_n19009_), .Y(new_n19010_));
  OAI21X1  g18818(.A0(new_n19003_), .A1(new_n19001_), .B0(\asqrt[41] ), .Y(new_n19011_));
  NAND2X1  g18819(.A(new_n19011_), .B(new_n3276_), .Y(new_n19012_));
  OAI21X1  g18820(.A0(new_n19012_), .A1(new_n19005_), .B0(new_n19010_), .Y(new_n19013_));
  AOI21X1  g18821(.A0(new_n19013_), .A1(new_n18995_), .B0(new_n3008_), .Y(new_n19014_));
  AND2X1   g18822(.A(new_n18364_), .B(new_n18363_), .Y(new_n19015_));
  NOR3X1   g18823(.A(new_n19015_), .B(new_n18326_), .C(new_n18362_), .Y(new_n19016_));
  NOR3X1   g18824(.A(new_n18591_), .B(new_n19015_), .C(new_n18362_), .Y(new_n19017_));
  NOR2X1   g18825(.A(new_n19017_), .B(new_n18325_), .Y(new_n19018_));
  AOI21X1  g18826(.A0(new_n19016_), .A1(\asqrt[10] ), .B0(new_n19018_), .Y(new_n19019_));
  OAI21X1  g18827(.A0(new_n19004_), .A1(new_n18991_), .B0(new_n19011_), .Y(new_n19020_));
  AOI21X1  g18828(.A0(new_n19020_), .A1(\asqrt[42] ), .B0(\asqrt[43] ), .Y(new_n19021_));
  AOI21X1  g18829(.A0(new_n19021_), .A1(new_n19013_), .B0(new_n19019_), .Y(new_n19022_));
  OAI21X1  g18830(.A0(new_n19022_), .A1(new_n19014_), .B0(\asqrt[44] ), .Y(new_n19023_));
  AND2X1   g18831(.A(new_n18337_), .B(new_n18329_), .Y(new_n19024_));
  NOR3X1   g18832(.A(new_n19024_), .B(new_n18367_), .C(new_n18330_), .Y(new_n19025_));
  NOR3X1   g18833(.A(new_n18591_), .B(new_n19024_), .C(new_n18330_), .Y(new_n19026_));
  NOR2X1   g18834(.A(new_n19026_), .B(new_n18335_), .Y(new_n19027_));
  AOI21X1  g18835(.A0(new_n19025_), .A1(\asqrt[10] ), .B0(new_n19027_), .Y(new_n19028_));
  NOR3X1   g18836(.A(new_n19022_), .B(new_n19014_), .C(\asqrt[44] ), .Y(new_n19029_));
  OAI21X1  g18837(.A0(new_n19029_), .A1(new_n19028_), .B0(new_n19023_), .Y(new_n19030_));
  AND2X1   g18838(.A(new_n19030_), .B(\asqrt[45] ), .Y(new_n19031_));
  OR2X1    g18839(.A(new_n19029_), .B(new_n19028_), .Y(new_n19032_));
  OR4X1    g18840(.A(new_n18591_), .B(new_n18344_), .C(new_n18371_), .D(new_n18370_), .Y(new_n19033_));
  OR2X1    g18841(.A(new_n18344_), .B(new_n18370_), .Y(new_n19034_));
  OAI21X1  g18842(.A0(new_n19034_), .A1(new_n18591_), .B0(new_n18371_), .Y(new_n19035_));
  AND2X1   g18843(.A(new_n19035_), .B(new_n19033_), .Y(new_n19036_));
  AND2X1   g18844(.A(new_n19023_), .B(new_n2570_), .Y(new_n19037_));
  AOI21X1  g18845(.A0(new_n19037_), .A1(new_n19032_), .B0(new_n19036_), .Y(new_n19038_));
  OAI21X1  g18846(.A0(new_n19038_), .A1(new_n19031_), .B0(\asqrt[46] ), .Y(new_n19039_));
  AOI21X1  g18847(.A0(new_n18353_), .A1(new_n18347_), .B0(new_n18387_), .Y(new_n19040_));
  AND2X1   g18848(.A(new_n19040_), .B(new_n18385_), .Y(new_n19041_));
  AOI22X1  g18849(.A0(new_n18353_), .A1(new_n18347_), .B0(new_n18345_), .B1(\asqrt[45] ), .Y(new_n19042_));
  AOI21X1  g18850(.A0(new_n19042_), .A1(\asqrt[10] ), .B0(new_n18352_), .Y(new_n19043_));
  AOI21X1  g18851(.A0(new_n19041_), .A1(\asqrt[10] ), .B0(new_n19043_), .Y(new_n19044_));
  INVX1    g18852(.A(new_n19044_), .Y(new_n19045_));
  AND2X1   g18853(.A(new_n19020_), .B(\asqrt[42] ), .Y(new_n19046_));
  OR2X1    g18854(.A(new_n19004_), .B(new_n18991_), .Y(new_n19047_));
  AND2X1   g18855(.A(new_n19011_), .B(new_n3276_), .Y(new_n19048_));
  AOI21X1  g18856(.A0(new_n19048_), .A1(new_n19047_), .B0(new_n19009_), .Y(new_n19049_));
  OAI21X1  g18857(.A0(new_n19049_), .A1(new_n19046_), .B0(\asqrt[43] ), .Y(new_n19050_));
  INVX1    g18858(.A(new_n19019_), .Y(new_n19051_));
  OAI21X1  g18859(.A0(new_n18994_), .A1(new_n3276_), .B0(new_n3008_), .Y(new_n19052_));
  OAI21X1  g18860(.A0(new_n19052_), .A1(new_n19049_), .B0(new_n19051_), .Y(new_n19053_));
  AOI21X1  g18861(.A0(new_n19053_), .A1(new_n19050_), .B0(new_n2769_), .Y(new_n19054_));
  INVX1    g18862(.A(new_n19028_), .Y(new_n19055_));
  NAND3X1  g18863(.A(new_n19053_), .B(new_n19050_), .C(new_n2769_), .Y(new_n19056_));
  AOI21X1  g18864(.A0(new_n19056_), .A1(new_n19055_), .B0(new_n19054_), .Y(new_n19057_));
  OAI21X1  g18865(.A0(new_n19057_), .A1(new_n2570_), .B0(new_n2263_), .Y(new_n19058_));
  OAI21X1  g18866(.A0(new_n19058_), .A1(new_n19038_), .B0(new_n19045_), .Y(new_n19059_));
  AOI21X1  g18867(.A0(new_n19059_), .A1(new_n19039_), .B0(new_n2040_), .Y(new_n19060_));
  AND2X1   g18868(.A(new_n18391_), .B(new_n18389_), .Y(new_n19061_));
  NOR3X1   g18869(.A(new_n19061_), .B(new_n18361_), .C(new_n18390_), .Y(new_n19062_));
  NOR3X1   g18870(.A(new_n18591_), .B(new_n19061_), .C(new_n18390_), .Y(new_n19063_));
  NOR2X1   g18871(.A(new_n19063_), .B(new_n18360_), .Y(new_n19064_));
  AOI21X1  g18872(.A0(new_n19062_), .A1(\asqrt[10] ), .B0(new_n19064_), .Y(new_n19065_));
  INVX1    g18873(.A(new_n19065_), .Y(new_n19066_));
  NAND3X1  g18874(.A(new_n19059_), .B(new_n19039_), .C(new_n2040_), .Y(new_n19067_));
  AOI21X1  g18875(.A0(new_n19067_), .A1(new_n19066_), .B0(new_n19060_), .Y(new_n19068_));
  OR2X1    g18876(.A(new_n19068_), .B(new_n1834_), .Y(new_n19069_));
  OR2X1    g18877(.A(new_n19057_), .B(new_n2570_), .Y(new_n19070_));
  NOR2X1   g18878(.A(new_n19029_), .B(new_n19028_), .Y(new_n19071_));
  INVX1    g18879(.A(new_n19036_), .Y(new_n19072_));
  NAND2X1  g18880(.A(new_n19023_), .B(new_n2570_), .Y(new_n19073_));
  OAI21X1  g18881(.A0(new_n19073_), .A1(new_n19071_), .B0(new_n19072_), .Y(new_n19074_));
  AOI21X1  g18882(.A0(new_n19074_), .A1(new_n19070_), .B0(new_n2263_), .Y(new_n19075_));
  AOI21X1  g18883(.A0(new_n19030_), .A1(\asqrt[45] ), .B0(\asqrt[46] ), .Y(new_n19076_));
  AOI21X1  g18884(.A0(new_n19076_), .A1(new_n19074_), .B0(new_n19044_), .Y(new_n19077_));
  NOR3X1   g18885(.A(new_n19077_), .B(new_n19075_), .C(\asqrt[47] ), .Y(new_n19078_));
  NOR2X1   g18886(.A(new_n19078_), .B(new_n19065_), .Y(new_n19079_));
  OR4X1    g18887(.A(new_n18591_), .B(new_n18393_), .C(new_n18381_), .D(new_n18376_), .Y(new_n19080_));
  OR2X1    g18888(.A(new_n18393_), .B(new_n18376_), .Y(new_n19081_));
  OAI21X1  g18889(.A0(new_n19081_), .A1(new_n18591_), .B0(new_n18381_), .Y(new_n19082_));
  AND2X1   g18890(.A(new_n19082_), .B(new_n19080_), .Y(new_n19083_));
  INVX1    g18891(.A(new_n19083_), .Y(new_n19084_));
  OAI21X1  g18892(.A0(new_n19077_), .A1(new_n19075_), .B0(\asqrt[47] ), .Y(new_n19085_));
  NAND2X1  g18893(.A(new_n19085_), .B(new_n1834_), .Y(new_n19086_));
  OAI21X1  g18894(.A0(new_n19086_), .A1(new_n19079_), .B0(new_n19084_), .Y(new_n19087_));
  AOI21X1  g18895(.A0(new_n19087_), .A1(new_n19069_), .B0(new_n1632_), .Y(new_n19088_));
  AND2X1   g18896(.A(new_n18437_), .B(new_n18436_), .Y(new_n19089_));
  NOR3X1   g18897(.A(new_n19089_), .B(new_n18400_), .C(new_n18435_), .Y(new_n19090_));
  NOR3X1   g18898(.A(new_n18591_), .B(new_n19089_), .C(new_n18435_), .Y(new_n19091_));
  NOR2X1   g18899(.A(new_n19091_), .B(new_n18399_), .Y(new_n19092_));
  AOI21X1  g18900(.A0(new_n19090_), .A1(\asqrt[10] ), .B0(new_n19092_), .Y(new_n19093_));
  OAI21X1  g18901(.A0(new_n19078_), .A1(new_n19065_), .B0(new_n19085_), .Y(new_n19094_));
  AOI21X1  g18902(.A0(new_n19094_), .A1(\asqrt[48] ), .B0(\asqrt[49] ), .Y(new_n19095_));
  AOI21X1  g18903(.A0(new_n19095_), .A1(new_n19087_), .B0(new_n19093_), .Y(new_n19096_));
  OAI21X1  g18904(.A0(new_n19096_), .A1(new_n19088_), .B0(\asqrt[50] ), .Y(new_n19097_));
  AND2X1   g18905(.A(new_n18411_), .B(new_n18403_), .Y(new_n19098_));
  NOR3X1   g18906(.A(new_n19098_), .B(new_n18440_), .C(new_n18404_), .Y(new_n19099_));
  NOR3X1   g18907(.A(new_n18591_), .B(new_n19098_), .C(new_n18404_), .Y(new_n19100_));
  NOR2X1   g18908(.A(new_n19100_), .B(new_n18409_), .Y(new_n19101_));
  AOI21X1  g18909(.A0(new_n19099_), .A1(\asqrt[10] ), .B0(new_n19101_), .Y(new_n19102_));
  NOR3X1   g18910(.A(new_n19096_), .B(new_n19088_), .C(\asqrt[50] ), .Y(new_n19103_));
  OAI21X1  g18911(.A0(new_n19103_), .A1(new_n19102_), .B0(new_n19097_), .Y(new_n19104_));
  AND2X1   g18912(.A(new_n19104_), .B(\asqrt[51] ), .Y(new_n19105_));
  OR2X1    g18913(.A(new_n19103_), .B(new_n19102_), .Y(new_n19106_));
  OR4X1    g18914(.A(new_n18591_), .B(new_n18418_), .C(new_n18444_), .D(new_n18443_), .Y(new_n19107_));
  OR2X1    g18915(.A(new_n18418_), .B(new_n18443_), .Y(new_n19108_));
  OAI21X1  g18916(.A0(new_n19108_), .A1(new_n18591_), .B0(new_n18444_), .Y(new_n19109_));
  AND2X1   g18917(.A(new_n19109_), .B(new_n19107_), .Y(new_n19110_));
  AND2X1   g18918(.A(new_n19097_), .B(new_n1277_), .Y(new_n19111_));
  AOI21X1  g18919(.A0(new_n19111_), .A1(new_n19106_), .B0(new_n19110_), .Y(new_n19112_));
  OAI21X1  g18920(.A0(new_n19112_), .A1(new_n19105_), .B0(\asqrt[52] ), .Y(new_n19113_));
  AOI21X1  g18921(.A0(new_n18427_), .A1(new_n18421_), .B0(new_n18460_), .Y(new_n19114_));
  AND2X1   g18922(.A(new_n19114_), .B(new_n18458_), .Y(new_n19115_));
  AOI22X1  g18923(.A0(new_n18427_), .A1(new_n18421_), .B0(new_n18419_), .B1(\asqrt[51] ), .Y(new_n19116_));
  AOI21X1  g18924(.A0(new_n19116_), .A1(\asqrt[10] ), .B0(new_n18426_), .Y(new_n19117_));
  AOI21X1  g18925(.A0(new_n19115_), .A1(\asqrt[10] ), .B0(new_n19117_), .Y(new_n19118_));
  INVX1    g18926(.A(new_n19118_), .Y(new_n19119_));
  AND2X1   g18927(.A(new_n19094_), .B(\asqrt[48] ), .Y(new_n19120_));
  OR2X1    g18928(.A(new_n19078_), .B(new_n19065_), .Y(new_n19121_));
  AND2X1   g18929(.A(new_n19085_), .B(new_n1834_), .Y(new_n19122_));
  AOI21X1  g18930(.A0(new_n19122_), .A1(new_n19121_), .B0(new_n19083_), .Y(new_n19123_));
  OAI21X1  g18931(.A0(new_n19123_), .A1(new_n19120_), .B0(\asqrt[49] ), .Y(new_n19124_));
  INVX1    g18932(.A(new_n19093_), .Y(new_n19125_));
  OAI21X1  g18933(.A0(new_n19068_), .A1(new_n1834_), .B0(new_n1632_), .Y(new_n19126_));
  OAI21X1  g18934(.A0(new_n19126_), .A1(new_n19123_), .B0(new_n19125_), .Y(new_n19127_));
  AOI21X1  g18935(.A0(new_n19127_), .A1(new_n19124_), .B0(new_n1469_), .Y(new_n19128_));
  INVX1    g18936(.A(new_n19102_), .Y(new_n19129_));
  NAND3X1  g18937(.A(new_n19127_), .B(new_n19124_), .C(new_n1469_), .Y(new_n19130_));
  AOI21X1  g18938(.A0(new_n19130_), .A1(new_n19129_), .B0(new_n19128_), .Y(new_n19131_));
  OAI21X1  g18939(.A0(new_n19131_), .A1(new_n1277_), .B0(new_n1111_), .Y(new_n19132_));
  OAI21X1  g18940(.A0(new_n19132_), .A1(new_n19112_), .B0(new_n19119_), .Y(new_n19133_));
  AOI21X1  g18941(.A0(new_n19133_), .A1(new_n19113_), .B0(new_n968_), .Y(new_n19134_));
  AND2X1   g18942(.A(new_n18465_), .B(new_n18462_), .Y(new_n19135_));
  NOR3X1   g18943(.A(new_n19135_), .B(new_n18434_), .C(new_n18463_), .Y(new_n19136_));
  NOR3X1   g18944(.A(new_n18591_), .B(new_n19135_), .C(new_n18463_), .Y(new_n19137_));
  NOR2X1   g18945(.A(new_n19137_), .B(new_n18464_), .Y(new_n19138_));
  AOI21X1  g18946(.A0(new_n19136_), .A1(\asqrt[10] ), .B0(new_n19138_), .Y(new_n19139_));
  INVX1    g18947(.A(new_n19139_), .Y(new_n19140_));
  NAND3X1  g18948(.A(new_n19133_), .B(new_n19113_), .C(new_n968_), .Y(new_n19141_));
  AOI21X1  g18949(.A0(new_n19141_), .A1(new_n19140_), .B0(new_n19134_), .Y(new_n19142_));
  OR2X1    g18950(.A(new_n19142_), .B(new_n902_), .Y(new_n19143_));
  OR2X1    g18951(.A(new_n19131_), .B(new_n1277_), .Y(new_n19144_));
  NOR2X1   g18952(.A(new_n19103_), .B(new_n19102_), .Y(new_n19145_));
  INVX1    g18953(.A(new_n19110_), .Y(new_n19146_));
  NAND2X1  g18954(.A(new_n19097_), .B(new_n1277_), .Y(new_n19147_));
  OAI21X1  g18955(.A0(new_n19147_), .A1(new_n19145_), .B0(new_n19146_), .Y(new_n19148_));
  AOI21X1  g18956(.A0(new_n19148_), .A1(new_n19144_), .B0(new_n1111_), .Y(new_n19149_));
  AOI21X1  g18957(.A0(new_n19104_), .A1(\asqrt[51] ), .B0(\asqrt[52] ), .Y(new_n19150_));
  AOI21X1  g18958(.A0(new_n19150_), .A1(new_n19148_), .B0(new_n19118_), .Y(new_n19151_));
  NOR3X1   g18959(.A(new_n19151_), .B(new_n19149_), .C(\asqrt[53] ), .Y(new_n19152_));
  NOR2X1   g18960(.A(new_n19152_), .B(new_n19139_), .Y(new_n19153_));
  OR4X1    g18961(.A(new_n18591_), .B(new_n18467_), .C(new_n18454_), .D(new_n18449_), .Y(new_n19154_));
  OR2X1    g18962(.A(new_n18467_), .B(new_n18449_), .Y(new_n19155_));
  OAI21X1  g18963(.A0(new_n19155_), .A1(new_n18591_), .B0(new_n18454_), .Y(new_n19156_));
  AND2X1   g18964(.A(new_n19156_), .B(new_n19154_), .Y(new_n19157_));
  INVX1    g18965(.A(new_n19157_), .Y(new_n19158_));
  OAI21X1  g18966(.A0(new_n19151_), .A1(new_n19149_), .B0(\asqrt[53] ), .Y(new_n19159_));
  NAND2X1  g18967(.A(new_n19159_), .B(new_n902_), .Y(new_n19160_));
  OAI21X1  g18968(.A0(new_n19160_), .A1(new_n19153_), .B0(new_n19158_), .Y(new_n19161_));
  AOI21X1  g18969(.A0(new_n19161_), .A1(new_n19143_), .B0(new_n697_), .Y(new_n19162_));
  OAI21X1  g18970(.A0(new_n19152_), .A1(new_n19139_), .B0(new_n19159_), .Y(new_n19163_));
  AOI21X1  g18971(.A0(new_n19163_), .A1(\asqrt[54] ), .B0(\asqrt[55] ), .Y(new_n19164_));
  AND2X1   g18972(.A(new_n18513_), .B(new_n18512_), .Y(new_n19165_));
  NOR3X1   g18973(.A(new_n18476_), .B(new_n19165_), .C(new_n18511_), .Y(new_n19166_));
  NOR3X1   g18974(.A(new_n18591_), .B(new_n19165_), .C(new_n18511_), .Y(new_n19167_));
  NOR2X1   g18975(.A(new_n19167_), .B(new_n18475_), .Y(new_n19168_));
  AOI21X1  g18976(.A0(new_n19166_), .A1(\asqrt[10] ), .B0(new_n19168_), .Y(new_n19169_));
  AOI21X1  g18977(.A0(new_n19164_), .A1(new_n19161_), .B0(new_n19169_), .Y(new_n19170_));
  OAI21X1  g18978(.A0(new_n19170_), .A1(new_n19162_), .B0(\asqrt[56] ), .Y(new_n19171_));
  AND2X1   g18979(.A(new_n18486_), .B(new_n18477_), .Y(new_n19172_));
  NOR3X1   g18980(.A(new_n19172_), .B(new_n18483_), .C(new_n18478_), .Y(new_n19173_));
  NOR3X1   g18981(.A(new_n18591_), .B(new_n19172_), .C(new_n18478_), .Y(new_n19174_));
  NOR2X1   g18982(.A(new_n19174_), .B(new_n18484_), .Y(new_n19175_));
  AOI21X1  g18983(.A0(new_n19173_), .A1(\asqrt[10] ), .B0(new_n19175_), .Y(new_n19176_));
  NOR3X1   g18984(.A(new_n19170_), .B(new_n19162_), .C(\asqrt[56] ), .Y(new_n19177_));
  OAI21X1  g18985(.A0(new_n19177_), .A1(new_n19176_), .B0(new_n19171_), .Y(new_n19178_));
  AND2X1   g18986(.A(new_n19178_), .B(\asqrt[57] ), .Y(new_n19179_));
  OR2X1    g18987(.A(new_n19177_), .B(new_n19176_), .Y(new_n19180_));
  OR4X1    g18988(.A(new_n18591_), .B(new_n18493_), .C(new_n18519_), .D(new_n18518_), .Y(new_n19181_));
  OR2X1    g18989(.A(new_n18493_), .B(new_n18518_), .Y(new_n19182_));
  OAI21X1  g18990(.A0(new_n19182_), .A1(new_n18591_), .B0(new_n18519_), .Y(new_n19183_));
  AND2X1   g18991(.A(new_n19183_), .B(new_n19181_), .Y(new_n19184_));
  AND2X1   g18992(.A(new_n19171_), .B(new_n481_), .Y(new_n19185_));
  AOI21X1  g18993(.A0(new_n19185_), .A1(new_n19180_), .B0(new_n19184_), .Y(new_n19186_));
  OAI21X1  g18994(.A0(new_n19186_), .A1(new_n19179_), .B0(\asqrt[58] ), .Y(new_n19187_));
  AOI21X1  g18995(.A0(new_n18502_), .A1(new_n18496_), .B0(new_n18535_), .Y(new_n19188_));
  AND2X1   g18996(.A(new_n19188_), .B(new_n18533_), .Y(new_n19189_));
  AOI22X1  g18997(.A0(new_n18502_), .A1(new_n18496_), .B0(new_n18494_), .B1(\asqrt[57] ), .Y(new_n19190_));
  AOI21X1  g18998(.A0(new_n19190_), .A1(\asqrt[10] ), .B0(new_n18501_), .Y(new_n19191_));
  AOI21X1  g18999(.A0(new_n19189_), .A1(\asqrt[10] ), .B0(new_n19191_), .Y(new_n19192_));
  INVX1    g19000(.A(new_n19192_), .Y(new_n19193_));
  AND2X1   g19001(.A(new_n19163_), .B(\asqrt[54] ), .Y(new_n19194_));
  OR2X1    g19002(.A(new_n19152_), .B(new_n19139_), .Y(new_n19195_));
  AND2X1   g19003(.A(new_n19159_), .B(new_n902_), .Y(new_n19196_));
  AOI21X1  g19004(.A0(new_n19196_), .A1(new_n19195_), .B0(new_n19157_), .Y(new_n19197_));
  OAI21X1  g19005(.A0(new_n19197_), .A1(new_n19194_), .B0(\asqrt[55] ), .Y(new_n19198_));
  OAI21X1  g19006(.A0(new_n19142_), .A1(new_n902_), .B0(new_n697_), .Y(new_n19199_));
  INVX1    g19007(.A(new_n19169_), .Y(new_n19200_));
  OAI21X1  g19008(.A0(new_n19199_), .A1(new_n19197_), .B0(new_n19200_), .Y(new_n19201_));
  AOI21X1  g19009(.A0(new_n19201_), .A1(new_n19198_), .B0(new_n582_), .Y(new_n19202_));
  INVX1    g19010(.A(new_n19176_), .Y(new_n19203_));
  NAND3X1  g19011(.A(new_n19201_), .B(new_n19198_), .C(new_n582_), .Y(new_n19204_));
  AOI21X1  g19012(.A0(new_n19204_), .A1(new_n19203_), .B0(new_n19202_), .Y(new_n19205_));
  OAI21X1  g19013(.A0(new_n19205_), .A1(new_n481_), .B0(new_n399_), .Y(new_n19206_));
  OAI21X1  g19014(.A0(new_n19206_), .A1(new_n19186_), .B0(new_n19193_), .Y(new_n19207_));
  AOI21X1  g19015(.A0(new_n19207_), .A1(new_n19187_), .B0(new_n328_), .Y(new_n19208_));
  AND2X1   g19016(.A(new_n18539_), .B(new_n18537_), .Y(new_n19209_));
  NOR3X1   g19017(.A(new_n19209_), .B(new_n18510_), .C(new_n18538_), .Y(new_n19210_));
  NOR3X1   g19018(.A(new_n18591_), .B(new_n19209_), .C(new_n18538_), .Y(new_n19211_));
  NOR2X1   g19019(.A(new_n19211_), .B(new_n18509_), .Y(new_n19212_));
  AOI21X1  g19020(.A0(new_n19210_), .A1(\asqrt[10] ), .B0(new_n19212_), .Y(new_n19213_));
  INVX1    g19021(.A(new_n19213_), .Y(new_n19214_));
  NAND3X1  g19022(.A(new_n19207_), .B(new_n19187_), .C(new_n328_), .Y(new_n19215_));
  AOI21X1  g19023(.A0(new_n19215_), .A1(new_n19214_), .B0(new_n19208_), .Y(new_n19216_));
  OR2X1    g19024(.A(new_n19216_), .B(new_n292_), .Y(new_n19217_));
  OR2X1    g19025(.A(new_n19205_), .B(new_n481_), .Y(new_n19218_));
  NOR2X1   g19026(.A(new_n19177_), .B(new_n19176_), .Y(new_n19219_));
  INVX1    g19027(.A(new_n19184_), .Y(new_n19220_));
  NAND2X1  g19028(.A(new_n19171_), .B(new_n481_), .Y(new_n19221_));
  OAI21X1  g19029(.A0(new_n19221_), .A1(new_n19219_), .B0(new_n19220_), .Y(new_n19222_));
  AOI21X1  g19030(.A0(new_n19222_), .A1(new_n19218_), .B0(new_n399_), .Y(new_n19223_));
  AOI21X1  g19031(.A0(new_n19178_), .A1(\asqrt[57] ), .B0(\asqrt[58] ), .Y(new_n19224_));
  AOI21X1  g19032(.A0(new_n19224_), .A1(new_n19222_), .B0(new_n19192_), .Y(new_n19225_));
  NOR3X1   g19033(.A(new_n19225_), .B(new_n19223_), .C(\asqrt[59] ), .Y(new_n19226_));
  NOR2X1   g19034(.A(new_n19226_), .B(new_n19213_), .Y(new_n19227_));
  OR4X1    g19035(.A(new_n18591_), .B(new_n18541_), .C(new_n18529_), .D(new_n18524_), .Y(new_n19228_));
  OR2X1    g19036(.A(new_n18541_), .B(new_n18524_), .Y(new_n19229_));
  OAI21X1  g19037(.A0(new_n19229_), .A1(new_n18591_), .B0(new_n18529_), .Y(new_n19230_));
  AND2X1   g19038(.A(new_n19230_), .B(new_n19228_), .Y(new_n19231_));
  INVX1    g19039(.A(new_n19231_), .Y(new_n19232_));
  OAI21X1  g19040(.A0(new_n19225_), .A1(new_n19223_), .B0(\asqrt[59] ), .Y(new_n19233_));
  NAND2X1  g19041(.A(new_n19233_), .B(new_n292_), .Y(new_n19234_));
  OAI21X1  g19042(.A0(new_n19234_), .A1(new_n19227_), .B0(new_n19232_), .Y(new_n19235_));
  AOI21X1  g19043(.A0(new_n19235_), .A1(new_n19217_), .B0(new_n217_), .Y(new_n19236_));
  AND2X1   g19044(.A(new_n18600_), .B(new_n18599_), .Y(new_n19237_));
  NOR3X1   g19045(.A(new_n19237_), .B(new_n18548_), .C(new_n18598_), .Y(new_n19238_));
  NOR3X1   g19046(.A(new_n18591_), .B(new_n19237_), .C(new_n18598_), .Y(new_n19239_));
  NOR2X1   g19047(.A(new_n19239_), .B(new_n18547_), .Y(new_n19240_));
  AOI21X1  g19048(.A0(new_n19238_), .A1(\asqrt[10] ), .B0(new_n19240_), .Y(new_n19241_));
  OAI21X1  g19049(.A0(new_n19226_), .A1(new_n19213_), .B0(new_n19233_), .Y(new_n19242_));
  AOI21X1  g19050(.A0(new_n19242_), .A1(\asqrt[60] ), .B0(\asqrt[61] ), .Y(new_n19243_));
  AOI21X1  g19051(.A0(new_n19243_), .A1(new_n19235_), .B0(new_n19241_), .Y(new_n19244_));
  OAI21X1  g19052(.A0(new_n19244_), .A1(new_n19236_), .B0(\asqrt[62] ), .Y(new_n19245_));
  AND2X1   g19053(.A(new_n18559_), .B(new_n18551_), .Y(new_n19246_));
  NOR3X1   g19054(.A(new_n19246_), .B(new_n18603_), .C(new_n18552_), .Y(new_n19247_));
  NOR3X1   g19055(.A(new_n18591_), .B(new_n19246_), .C(new_n18552_), .Y(new_n19248_));
  NOR2X1   g19056(.A(new_n19248_), .B(new_n18557_), .Y(new_n19249_));
  AOI21X1  g19057(.A0(new_n19247_), .A1(\asqrt[10] ), .B0(new_n19249_), .Y(new_n19250_));
  NOR3X1   g19058(.A(new_n19244_), .B(new_n19236_), .C(\asqrt[62] ), .Y(new_n19251_));
  OAI21X1  g19059(.A0(new_n19251_), .A1(new_n19250_), .B0(new_n19245_), .Y(new_n19252_));
  NOR4X1   g19060(.A(new_n18591_), .B(new_n18566_), .C(new_n18607_), .D(new_n18606_), .Y(new_n19253_));
  NOR3X1   g19061(.A(new_n18591_), .B(new_n18566_), .C(new_n18606_), .Y(new_n19254_));
  NOR2X1   g19062(.A(new_n19254_), .B(new_n18565_), .Y(new_n19255_));
  NOR2X1   g19063(.A(new_n19255_), .B(new_n19253_), .Y(new_n19256_));
  INVX1    g19064(.A(new_n19256_), .Y(new_n19257_));
  AND2X1   g19065(.A(new_n18573_), .B(new_n18567_), .Y(new_n19258_));
  AOI21X1  g19066(.A0(new_n19258_), .A1(\asqrt[10] ), .B0(new_n18627_), .Y(new_n19259_));
  AND2X1   g19067(.A(new_n19259_), .B(new_n19257_), .Y(new_n19260_));
  AOI21X1  g19068(.A0(new_n19260_), .A1(new_n19252_), .B0(\asqrt[63] ), .Y(new_n19261_));
  NOR2X1   g19069(.A(new_n19251_), .B(new_n19250_), .Y(new_n19262_));
  NAND2X1  g19070(.A(new_n19256_), .B(new_n19245_), .Y(new_n19263_));
  AOI21X1  g19071(.A0(new_n18615_), .A1(new_n18611_), .B0(new_n18572_), .Y(new_n19264_));
  AOI21X1  g19072(.A0(new_n18573_), .A1(new_n18567_), .B0(new_n193_), .Y(new_n19265_));
  OAI21X1  g19073(.A0(new_n19264_), .A1(new_n18567_), .B0(new_n19265_), .Y(new_n19266_));
  NOR4X1   g19074(.A(new_n18588_), .B(new_n18628_), .C(new_n18571_), .D(new_n18569_), .Y(new_n19267_));
  OAI21X1  g19075(.A0(new_n18580_), .A1(new_n18579_), .B0(new_n19267_), .Y(new_n19268_));
  NOR2X1   g19076(.A(new_n19268_), .B(new_n18578_), .Y(new_n19269_));
  INVX1    g19077(.A(new_n19269_), .Y(new_n19270_));
  AND2X1   g19078(.A(new_n19270_), .B(new_n19266_), .Y(new_n19271_));
  OAI21X1  g19079(.A0(new_n19263_), .A1(new_n19262_), .B0(new_n19271_), .Y(new_n19272_));
  NOR2X1   g19080(.A(new_n19272_), .B(new_n19261_), .Y(new_n19273_));
  OAI21X1  g19081(.A0(new_n19272_), .A1(new_n19261_), .B0(\a[18] ), .Y(new_n19274_));
  NOR3X1   g19082(.A(\a[18] ), .B(\a[17] ), .C(\a[16] ), .Y(new_n19275_));
  INVX1    g19083(.A(new_n19275_), .Y(new_n19276_));
  AOI21X1  g19084(.A0(new_n19276_), .A1(new_n19274_), .B0(new_n18591_), .Y(new_n19277_));
  OR2X1    g19085(.A(new_n19275_), .B(new_n18588_), .Y(new_n19278_));
  NOR4X1   g19086(.A(new_n19278_), .B(new_n18628_), .C(new_n18627_), .D(new_n18578_), .Y(new_n19279_));
  NAND2X1  g19087(.A(new_n19279_), .B(new_n19274_), .Y(new_n19280_));
  INVX1    g19088(.A(\a[18] ), .Y(new_n19281_));
  OAI21X1  g19089(.A0(new_n19272_), .A1(new_n19261_), .B0(new_n19281_), .Y(new_n19282_));
  INVX1    g19090(.A(new_n18595_), .Y(new_n19283_));
  AND2X1   g19091(.A(new_n19242_), .B(\asqrt[60] ), .Y(new_n19284_));
  OR2X1    g19092(.A(new_n19226_), .B(new_n19213_), .Y(new_n19285_));
  AND2X1   g19093(.A(new_n19233_), .B(new_n292_), .Y(new_n19286_));
  AOI21X1  g19094(.A0(new_n19286_), .A1(new_n19285_), .B0(new_n19231_), .Y(new_n19287_));
  OAI21X1  g19095(.A0(new_n19287_), .A1(new_n19284_), .B0(\asqrt[61] ), .Y(new_n19288_));
  INVX1    g19096(.A(new_n19241_), .Y(new_n19289_));
  OAI21X1  g19097(.A0(new_n19216_), .A1(new_n292_), .B0(new_n217_), .Y(new_n19290_));
  OAI21X1  g19098(.A0(new_n19290_), .A1(new_n19287_), .B0(new_n19289_), .Y(new_n19291_));
  AOI21X1  g19099(.A0(new_n19291_), .A1(new_n19288_), .B0(new_n199_), .Y(new_n19292_));
  INVX1    g19100(.A(new_n19250_), .Y(new_n19293_));
  NAND3X1  g19101(.A(new_n19291_), .B(new_n19288_), .C(new_n199_), .Y(new_n19294_));
  AOI21X1  g19102(.A0(new_n19294_), .A1(new_n19293_), .B0(new_n19292_), .Y(new_n19295_));
  INVX1    g19103(.A(new_n19260_), .Y(new_n19296_));
  OAI21X1  g19104(.A0(new_n19296_), .A1(new_n19295_), .B0(new_n193_), .Y(new_n19297_));
  OR2X1    g19105(.A(new_n19251_), .B(new_n19250_), .Y(new_n19298_));
  AND2X1   g19106(.A(new_n19256_), .B(new_n19245_), .Y(new_n19299_));
  INVX1    g19107(.A(new_n19271_), .Y(new_n19300_));
  AOI21X1  g19108(.A0(new_n19299_), .A1(new_n19298_), .B0(new_n19300_), .Y(new_n19301_));
  AOI21X1  g19109(.A0(new_n19301_), .A1(new_n19297_), .B0(new_n19283_), .Y(new_n19302_));
  AOI21X1  g19110(.A0(new_n19282_), .A1(\a[19] ), .B0(new_n19302_), .Y(new_n19303_));
  AOI21X1  g19111(.A0(new_n19303_), .A1(new_n19280_), .B0(new_n19277_), .Y(new_n19304_));
  OR2X1    g19112(.A(new_n19304_), .B(new_n17927_), .Y(new_n19305_));
  AND2X1   g19113(.A(new_n19303_), .B(new_n19280_), .Y(new_n19306_));
  OR2X1    g19114(.A(new_n19277_), .B(\asqrt[11] ), .Y(new_n19307_));
  OAI21X1  g19115(.A0(new_n19272_), .A1(new_n19261_), .B0(new_n18595_), .Y(new_n19308_));
  INVX1    g19116(.A(new_n19266_), .Y(new_n19309_));
  NOR3X1   g19117(.A(new_n19269_), .B(new_n19309_), .C(new_n18591_), .Y(new_n19310_));
  OAI21X1  g19118(.A0(new_n19263_), .A1(new_n19262_), .B0(new_n19310_), .Y(new_n19311_));
  OR2X1    g19119(.A(new_n19311_), .B(new_n19261_), .Y(new_n19312_));
  AOI21X1  g19120(.A0(new_n19312_), .A1(new_n19308_), .B0(new_n18594_), .Y(new_n19313_));
  OAI21X1  g19121(.A0(new_n19311_), .A1(new_n19261_), .B0(new_n18594_), .Y(new_n19314_));
  NOR2X1   g19122(.A(new_n19314_), .B(new_n19302_), .Y(new_n19315_));
  OR2X1    g19123(.A(new_n19315_), .B(new_n19313_), .Y(new_n19316_));
  OAI21X1  g19124(.A0(new_n19307_), .A1(new_n19306_), .B0(new_n19316_), .Y(new_n19317_));
  AOI21X1  g19125(.A0(new_n19317_), .A1(new_n19305_), .B0(new_n17262_), .Y(new_n19318_));
  NOR3X1   g19126(.A(new_n18621_), .B(new_n18644_), .C(new_n18597_), .Y(new_n19319_));
  OAI21X1  g19127(.A0(new_n19272_), .A1(new_n19261_), .B0(new_n19319_), .Y(new_n19320_));
  NOR2X1   g19128(.A(new_n18644_), .B(new_n18597_), .Y(new_n19321_));
  OAI21X1  g19129(.A0(new_n19272_), .A1(new_n19261_), .B0(new_n19321_), .Y(new_n19322_));
  NAND2X1  g19130(.A(new_n19322_), .B(new_n18621_), .Y(new_n19323_));
  AND2X1   g19131(.A(new_n19323_), .B(new_n19320_), .Y(new_n19324_));
  AOI21X1  g19132(.A0(new_n19301_), .A1(new_n19297_), .B0(new_n19281_), .Y(new_n19325_));
  OAI21X1  g19133(.A0(new_n19275_), .A1(new_n19325_), .B0(\asqrt[10] ), .Y(new_n19326_));
  AND2X1   g19134(.A(new_n19279_), .B(new_n19274_), .Y(new_n19327_));
  INVX1    g19135(.A(\a[19] ), .Y(new_n19328_));
  AOI21X1  g19136(.A0(new_n19301_), .A1(new_n19297_), .B0(\a[18] ), .Y(new_n19329_));
  OAI21X1  g19137(.A0(new_n19329_), .A1(new_n19328_), .B0(new_n19308_), .Y(new_n19330_));
  OAI21X1  g19138(.A0(new_n19330_), .A1(new_n19327_), .B0(new_n19326_), .Y(new_n19331_));
  AOI21X1  g19139(.A0(new_n19331_), .A1(\asqrt[11] ), .B0(\asqrt[12] ), .Y(new_n19332_));
  AOI21X1  g19140(.A0(new_n19332_), .A1(new_n19317_), .B0(new_n19324_), .Y(new_n19333_));
  OAI21X1  g19141(.A0(new_n19333_), .A1(new_n19318_), .B0(\asqrt[13] ), .Y(new_n19334_));
  AOI21X1  g19142(.A0(new_n18668_), .A1(new_n18667_), .B0(new_n18634_), .Y(new_n19335_));
  AND2X1   g19143(.A(new_n19335_), .B(new_n18623_), .Y(new_n19336_));
  OAI21X1  g19144(.A0(new_n19272_), .A1(new_n19261_), .B0(new_n19336_), .Y(new_n19337_));
  AOI22X1  g19145(.A0(new_n18668_), .A1(new_n18667_), .B0(new_n18648_), .B1(\asqrt[12] ), .Y(new_n19338_));
  OAI21X1  g19146(.A0(new_n19272_), .A1(new_n19261_), .B0(new_n19338_), .Y(new_n19339_));
  NAND2X1  g19147(.A(new_n19339_), .B(new_n18634_), .Y(new_n19340_));
  AND2X1   g19148(.A(new_n19340_), .B(new_n19337_), .Y(new_n19341_));
  NOR3X1   g19149(.A(new_n19333_), .B(new_n19318_), .C(\asqrt[13] ), .Y(new_n19342_));
  OAI21X1  g19150(.A0(new_n19342_), .A1(new_n19341_), .B0(new_n19334_), .Y(new_n19343_));
  AND2X1   g19151(.A(new_n19343_), .B(\asqrt[14] ), .Y(new_n19344_));
  OR2X1    g19152(.A(new_n19342_), .B(new_n19341_), .Y(new_n19345_));
  INVX1    g19153(.A(new_n19273_), .Y(\asqrt[9] ));
  AND2X1   g19154(.A(new_n18649_), .B(new_n18635_), .Y(new_n19347_));
  NOR3X1   g19155(.A(new_n19347_), .B(new_n18672_), .C(new_n18636_), .Y(new_n19348_));
  NOR2X1   g19156(.A(new_n19347_), .B(new_n18636_), .Y(new_n19349_));
  OAI21X1  g19157(.A0(new_n19272_), .A1(new_n19261_), .B0(new_n19349_), .Y(new_n19350_));
  AOI22X1  g19158(.A0(new_n19350_), .A1(new_n18672_), .B0(new_n19348_), .B1(\asqrt[9] ), .Y(new_n19351_));
  AND2X1   g19159(.A(new_n19334_), .B(new_n15990_), .Y(new_n19352_));
  AOI21X1  g19160(.A0(new_n19352_), .A1(new_n19345_), .B0(new_n19351_), .Y(new_n19353_));
  OAI21X1  g19161(.A0(new_n19353_), .A1(new_n19344_), .B0(\asqrt[15] ), .Y(new_n19354_));
  NAND4X1  g19162(.A(\asqrt[9] ), .B(new_n18686_), .C(new_n18658_), .D(new_n18651_), .Y(new_n19355_));
  NOR3X1   g19163(.A(new_n19273_), .B(new_n18659_), .C(new_n18675_), .Y(new_n19356_));
  OAI21X1  g19164(.A0(new_n19356_), .A1(new_n18658_), .B0(new_n19355_), .Y(new_n19357_));
  AND2X1   g19165(.A(new_n19331_), .B(\asqrt[11] ), .Y(new_n19358_));
  NAND2X1  g19166(.A(new_n19303_), .B(new_n19280_), .Y(new_n19359_));
  AND2X1   g19167(.A(new_n19326_), .B(new_n17927_), .Y(new_n19360_));
  NOR2X1   g19168(.A(new_n19315_), .B(new_n19313_), .Y(new_n19361_));
  AOI21X1  g19169(.A0(new_n19360_), .A1(new_n19359_), .B0(new_n19361_), .Y(new_n19362_));
  OAI21X1  g19170(.A0(new_n19362_), .A1(new_n19358_), .B0(\asqrt[12] ), .Y(new_n19363_));
  NAND2X1  g19171(.A(new_n19323_), .B(new_n19320_), .Y(new_n19364_));
  OAI21X1  g19172(.A0(new_n19304_), .A1(new_n17927_), .B0(new_n17262_), .Y(new_n19365_));
  OAI21X1  g19173(.A0(new_n19365_), .A1(new_n19362_), .B0(new_n19364_), .Y(new_n19366_));
  AOI21X1  g19174(.A0(new_n19366_), .A1(new_n19363_), .B0(new_n16617_), .Y(new_n19367_));
  INVX1    g19175(.A(new_n19341_), .Y(new_n19368_));
  NAND3X1  g19176(.A(new_n19366_), .B(new_n19363_), .C(new_n16617_), .Y(new_n19369_));
  AOI21X1  g19177(.A0(new_n19369_), .A1(new_n19368_), .B0(new_n19367_), .Y(new_n19370_));
  OAI21X1  g19178(.A0(new_n19370_), .A1(new_n15990_), .B0(new_n15362_), .Y(new_n19371_));
  OAI21X1  g19179(.A0(new_n19371_), .A1(new_n19353_), .B0(new_n19357_), .Y(new_n19372_));
  AOI21X1  g19180(.A0(new_n19372_), .A1(new_n19354_), .B0(new_n14754_), .Y(new_n19373_));
  AND2X1   g19181(.A(new_n18676_), .B(new_n18662_), .Y(new_n19374_));
  NOR3X1   g19182(.A(new_n19374_), .B(new_n18702_), .C(new_n18661_), .Y(new_n19375_));
  NOR3X1   g19183(.A(new_n19273_), .B(new_n19374_), .C(new_n18661_), .Y(new_n19376_));
  NOR2X1   g19184(.A(new_n19376_), .B(new_n18665_), .Y(new_n19377_));
  AOI21X1  g19185(.A0(new_n19375_), .A1(\asqrt[9] ), .B0(new_n19377_), .Y(new_n19378_));
  INVX1    g19186(.A(new_n19378_), .Y(new_n19379_));
  NAND3X1  g19187(.A(new_n19372_), .B(new_n19354_), .C(new_n14754_), .Y(new_n19380_));
  AOI21X1  g19188(.A0(new_n19380_), .A1(new_n19379_), .B0(new_n19373_), .Y(new_n19381_));
  OR2X1    g19189(.A(new_n19381_), .B(new_n14165_), .Y(new_n19382_));
  AND2X1   g19190(.A(new_n19380_), .B(new_n19379_), .Y(new_n19383_));
  AND2X1   g19191(.A(new_n18706_), .B(new_n18704_), .Y(new_n19384_));
  NOR3X1   g19192(.A(new_n19384_), .B(new_n18684_), .C(new_n18705_), .Y(new_n19385_));
  NOR3X1   g19193(.A(new_n19273_), .B(new_n19384_), .C(new_n18705_), .Y(new_n19386_));
  NOR2X1   g19194(.A(new_n19386_), .B(new_n18683_), .Y(new_n19387_));
  AOI21X1  g19195(.A0(new_n19385_), .A1(\asqrt[9] ), .B0(new_n19387_), .Y(new_n19388_));
  INVX1    g19196(.A(new_n19388_), .Y(new_n19389_));
  OR2X1    g19197(.A(new_n19370_), .B(new_n15990_), .Y(new_n19390_));
  NOR2X1   g19198(.A(new_n19342_), .B(new_n19341_), .Y(new_n19391_));
  INVX1    g19199(.A(new_n19351_), .Y(new_n19392_));
  NAND2X1  g19200(.A(new_n19334_), .B(new_n15990_), .Y(new_n19393_));
  OAI21X1  g19201(.A0(new_n19393_), .A1(new_n19391_), .B0(new_n19392_), .Y(new_n19394_));
  AOI21X1  g19202(.A0(new_n19394_), .A1(new_n19390_), .B0(new_n15362_), .Y(new_n19395_));
  INVX1    g19203(.A(new_n19357_), .Y(new_n19396_));
  AOI21X1  g19204(.A0(new_n19343_), .A1(\asqrt[14] ), .B0(\asqrt[15] ), .Y(new_n19397_));
  AOI21X1  g19205(.A0(new_n19397_), .A1(new_n19394_), .B0(new_n19396_), .Y(new_n19398_));
  OAI21X1  g19206(.A0(new_n19398_), .A1(new_n19395_), .B0(\asqrt[16] ), .Y(new_n19399_));
  NAND2X1  g19207(.A(new_n19399_), .B(new_n14165_), .Y(new_n19400_));
  OAI21X1  g19208(.A0(new_n19400_), .A1(new_n19383_), .B0(new_n19389_), .Y(new_n19401_));
  AOI21X1  g19209(.A0(new_n19401_), .A1(new_n19382_), .B0(new_n13571_), .Y(new_n19402_));
  OR4X1    g19210(.A(new_n19273_), .B(new_n18708_), .C(new_n18696_), .D(new_n18690_), .Y(new_n19403_));
  OR2X1    g19211(.A(new_n18708_), .B(new_n18690_), .Y(new_n19404_));
  OAI21X1  g19212(.A0(new_n19404_), .A1(new_n19273_), .B0(new_n18696_), .Y(new_n19405_));
  AND2X1   g19213(.A(new_n19405_), .B(new_n19403_), .Y(new_n19406_));
  NOR3X1   g19214(.A(new_n19398_), .B(new_n19395_), .C(\asqrt[16] ), .Y(new_n19407_));
  OAI21X1  g19215(.A0(new_n19407_), .A1(new_n19378_), .B0(new_n19399_), .Y(new_n19408_));
  AOI21X1  g19216(.A0(new_n19408_), .A1(\asqrt[17] ), .B0(\asqrt[18] ), .Y(new_n19409_));
  AOI21X1  g19217(.A0(new_n19409_), .A1(new_n19401_), .B0(new_n19406_), .Y(new_n19410_));
  OAI21X1  g19218(.A0(new_n19410_), .A1(new_n19402_), .B0(\asqrt[19] ), .Y(new_n19411_));
  OAI21X1  g19219(.A0(new_n18716_), .A1(new_n18709_), .B0(new_n18713_), .Y(new_n19412_));
  NOR2X1   g19220(.A(new_n19412_), .B(new_n18750_), .Y(new_n19413_));
  AOI22X1  g19221(.A0(new_n18752_), .A1(new_n18751_), .B0(new_n18724_), .B1(\asqrt[18] ), .Y(new_n19414_));
  AOI21X1  g19222(.A0(new_n19414_), .A1(\asqrt[9] ), .B0(new_n18713_), .Y(new_n19415_));
  AOI21X1  g19223(.A0(new_n19413_), .A1(\asqrt[9] ), .B0(new_n19415_), .Y(new_n19416_));
  NOR3X1   g19224(.A(new_n19410_), .B(new_n19402_), .C(\asqrt[19] ), .Y(new_n19417_));
  OAI21X1  g19225(.A0(new_n19417_), .A1(new_n19416_), .B0(new_n19411_), .Y(new_n19418_));
  AND2X1   g19226(.A(new_n19418_), .B(\asqrt[20] ), .Y(new_n19419_));
  INVX1    g19227(.A(new_n19416_), .Y(new_n19420_));
  AND2X1   g19228(.A(new_n19408_), .B(\asqrt[17] ), .Y(new_n19421_));
  NAND2X1  g19229(.A(new_n19380_), .B(new_n19379_), .Y(new_n19422_));
  AND2X1   g19230(.A(new_n19399_), .B(new_n14165_), .Y(new_n19423_));
  AOI21X1  g19231(.A0(new_n19423_), .A1(new_n19422_), .B0(new_n19388_), .Y(new_n19424_));
  OAI21X1  g19232(.A0(new_n19424_), .A1(new_n19421_), .B0(\asqrt[18] ), .Y(new_n19425_));
  INVX1    g19233(.A(new_n19406_), .Y(new_n19426_));
  OAI21X1  g19234(.A0(new_n19381_), .A1(new_n14165_), .B0(new_n13571_), .Y(new_n19427_));
  OAI21X1  g19235(.A0(new_n19427_), .A1(new_n19424_), .B0(new_n19426_), .Y(new_n19428_));
  NAND3X1  g19236(.A(new_n19428_), .B(new_n19425_), .C(new_n13000_), .Y(new_n19429_));
  NAND2X1  g19237(.A(new_n19429_), .B(new_n19420_), .Y(new_n19430_));
  AND2X1   g19238(.A(new_n18725_), .B(new_n18717_), .Y(new_n19431_));
  NOR3X1   g19239(.A(new_n19431_), .B(new_n18755_), .C(new_n18718_), .Y(new_n19432_));
  NOR3X1   g19240(.A(new_n19273_), .B(new_n19431_), .C(new_n18718_), .Y(new_n19433_));
  NOR2X1   g19241(.A(new_n19433_), .B(new_n18723_), .Y(new_n19434_));
  AOI21X1  g19242(.A0(new_n19432_), .A1(\asqrt[9] ), .B0(new_n19434_), .Y(new_n19435_));
  AND2X1   g19243(.A(new_n19411_), .B(new_n12447_), .Y(new_n19436_));
  AOI21X1  g19244(.A0(new_n19436_), .A1(new_n19430_), .B0(new_n19435_), .Y(new_n19437_));
  OAI21X1  g19245(.A0(new_n19437_), .A1(new_n19419_), .B0(\asqrt[21] ), .Y(new_n19438_));
  OR4X1    g19246(.A(new_n19273_), .B(new_n18733_), .C(new_n18759_), .D(new_n18758_), .Y(new_n19439_));
  OR2X1    g19247(.A(new_n18733_), .B(new_n18758_), .Y(new_n19440_));
  OAI21X1  g19248(.A0(new_n19440_), .A1(new_n19273_), .B0(new_n18759_), .Y(new_n19441_));
  AND2X1   g19249(.A(new_n19441_), .B(new_n19439_), .Y(new_n19442_));
  INVX1    g19250(.A(new_n19442_), .Y(new_n19443_));
  AOI21X1  g19251(.A0(new_n19428_), .A1(new_n19425_), .B0(new_n13000_), .Y(new_n19444_));
  AOI21X1  g19252(.A0(new_n19429_), .A1(new_n19420_), .B0(new_n19444_), .Y(new_n19445_));
  OAI21X1  g19253(.A0(new_n19445_), .A1(new_n12447_), .B0(new_n11896_), .Y(new_n19446_));
  OAI21X1  g19254(.A0(new_n19446_), .A1(new_n19437_), .B0(new_n19443_), .Y(new_n19447_));
  AOI21X1  g19255(.A0(new_n19447_), .A1(new_n19438_), .B0(new_n11362_), .Y(new_n19448_));
  AND2X1   g19256(.A(new_n18741_), .B(new_n18736_), .Y(new_n19449_));
  NOR3X1   g19257(.A(new_n19449_), .B(new_n18790_), .C(new_n18735_), .Y(new_n19450_));
  NOR3X1   g19258(.A(new_n19273_), .B(new_n19449_), .C(new_n18735_), .Y(new_n19451_));
  NOR2X1   g19259(.A(new_n19451_), .B(new_n18740_), .Y(new_n19452_));
  AOI21X1  g19260(.A0(new_n19450_), .A1(\asqrt[9] ), .B0(new_n19452_), .Y(new_n19453_));
  INVX1    g19261(.A(new_n19453_), .Y(new_n19454_));
  NAND3X1  g19262(.A(new_n19447_), .B(new_n19438_), .C(new_n11362_), .Y(new_n19455_));
  AOI21X1  g19263(.A0(new_n19455_), .A1(new_n19454_), .B0(new_n19448_), .Y(new_n19456_));
  OR2X1    g19264(.A(new_n19456_), .B(new_n10849_), .Y(new_n19457_));
  AND2X1   g19265(.A(new_n19455_), .B(new_n19454_), .Y(new_n19458_));
  AND2X1   g19266(.A(new_n18794_), .B(new_n18792_), .Y(new_n19459_));
  NOR3X1   g19267(.A(new_n19459_), .B(new_n18749_), .C(new_n18793_), .Y(new_n19460_));
  NOR3X1   g19268(.A(new_n19273_), .B(new_n19459_), .C(new_n18793_), .Y(new_n19461_));
  NOR2X1   g19269(.A(new_n19461_), .B(new_n18748_), .Y(new_n19462_));
  AOI21X1  g19270(.A0(new_n19460_), .A1(\asqrt[9] ), .B0(new_n19462_), .Y(new_n19463_));
  INVX1    g19271(.A(new_n19463_), .Y(new_n19464_));
  OR2X1    g19272(.A(new_n19445_), .B(new_n12447_), .Y(new_n19465_));
  AND2X1   g19273(.A(new_n19429_), .B(new_n19420_), .Y(new_n19466_));
  INVX1    g19274(.A(new_n19435_), .Y(new_n19467_));
  NAND2X1  g19275(.A(new_n19411_), .B(new_n12447_), .Y(new_n19468_));
  OAI21X1  g19276(.A0(new_n19468_), .A1(new_n19466_), .B0(new_n19467_), .Y(new_n19469_));
  AOI21X1  g19277(.A0(new_n19469_), .A1(new_n19465_), .B0(new_n11896_), .Y(new_n19470_));
  AOI21X1  g19278(.A0(new_n19418_), .A1(\asqrt[20] ), .B0(\asqrt[21] ), .Y(new_n19471_));
  AOI21X1  g19279(.A0(new_n19471_), .A1(new_n19469_), .B0(new_n19442_), .Y(new_n19472_));
  OAI21X1  g19280(.A0(new_n19472_), .A1(new_n19470_), .B0(\asqrt[22] ), .Y(new_n19473_));
  NAND2X1  g19281(.A(new_n19473_), .B(new_n10849_), .Y(new_n19474_));
  OAI21X1  g19282(.A0(new_n19474_), .A1(new_n19458_), .B0(new_n19464_), .Y(new_n19475_));
  AOI21X1  g19283(.A0(new_n19475_), .A1(new_n19457_), .B0(new_n10332_), .Y(new_n19476_));
  NAND4X1  g19284(.A(\asqrt[9] ), .B(new_n18771_), .C(new_n18769_), .D(new_n18796_), .Y(new_n19477_));
  NAND2X1  g19285(.A(new_n18771_), .B(new_n18796_), .Y(new_n19478_));
  OAI21X1  g19286(.A0(new_n19478_), .A1(new_n19273_), .B0(new_n18770_), .Y(new_n19479_));
  AND2X1   g19287(.A(new_n19479_), .B(new_n19477_), .Y(new_n19480_));
  NOR3X1   g19288(.A(new_n19472_), .B(new_n19470_), .C(\asqrt[22] ), .Y(new_n19481_));
  OAI21X1  g19289(.A0(new_n19481_), .A1(new_n19453_), .B0(new_n19473_), .Y(new_n19482_));
  AOI21X1  g19290(.A0(new_n19482_), .A1(\asqrt[23] ), .B0(\asqrt[24] ), .Y(new_n19483_));
  AOI21X1  g19291(.A0(new_n19483_), .A1(new_n19475_), .B0(new_n19480_), .Y(new_n19484_));
  OAI21X1  g19292(.A0(new_n19484_), .A1(new_n19476_), .B0(\asqrt[25] ), .Y(new_n19485_));
  AOI21X1  g19293(.A0(new_n18813_), .A1(new_n18812_), .B0(new_n18779_), .Y(new_n19486_));
  AND2X1   g19294(.A(new_n19486_), .B(new_n18773_), .Y(new_n19487_));
  AOI22X1  g19295(.A0(new_n18813_), .A1(new_n18812_), .B0(new_n18798_), .B1(\asqrt[24] ), .Y(new_n19488_));
  AOI21X1  g19296(.A0(new_n19488_), .A1(\asqrt[9] ), .B0(new_n18778_), .Y(new_n19489_));
  AOI21X1  g19297(.A0(new_n19487_), .A1(\asqrt[9] ), .B0(new_n19489_), .Y(new_n19490_));
  NOR3X1   g19298(.A(new_n19484_), .B(new_n19476_), .C(\asqrt[25] ), .Y(new_n19491_));
  OAI21X1  g19299(.A0(new_n19491_), .A1(new_n19490_), .B0(new_n19485_), .Y(new_n19492_));
  AND2X1   g19300(.A(new_n19492_), .B(\asqrt[26] ), .Y(new_n19493_));
  INVX1    g19301(.A(new_n19490_), .Y(new_n19494_));
  AND2X1   g19302(.A(new_n19482_), .B(\asqrt[23] ), .Y(new_n19495_));
  NAND2X1  g19303(.A(new_n19455_), .B(new_n19454_), .Y(new_n19496_));
  AND2X1   g19304(.A(new_n19473_), .B(new_n10849_), .Y(new_n19497_));
  AOI21X1  g19305(.A0(new_n19497_), .A1(new_n19496_), .B0(new_n19463_), .Y(new_n19498_));
  OAI21X1  g19306(.A0(new_n19498_), .A1(new_n19495_), .B0(\asqrt[24] ), .Y(new_n19499_));
  INVX1    g19307(.A(new_n19480_), .Y(new_n19500_));
  OAI21X1  g19308(.A0(new_n19456_), .A1(new_n10849_), .B0(new_n10332_), .Y(new_n19501_));
  OAI21X1  g19309(.A0(new_n19501_), .A1(new_n19498_), .B0(new_n19500_), .Y(new_n19502_));
  NAND3X1  g19310(.A(new_n19502_), .B(new_n19499_), .C(new_n9833_), .Y(new_n19503_));
  NAND2X1  g19311(.A(new_n19503_), .B(new_n19494_), .Y(new_n19504_));
  AND2X1   g19312(.A(new_n18799_), .B(new_n18781_), .Y(new_n19505_));
  NOR3X1   g19313(.A(new_n19505_), .B(new_n18816_), .C(new_n18782_), .Y(new_n19506_));
  NOR3X1   g19314(.A(new_n19273_), .B(new_n19505_), .C(new_n18782_), .Y(new_n19507_));
  NOR2X1   g19315(.A(new_n19507_), .B(new_n18787_), .Y(new_n19508_));
  AOI21X1  g19316(.A0(new_n19506_), .A1(\asqrt[9] ), .B0(new_n19508_), .Y(new_n19509_));
  AND2X1   g19317(.A(new_n19485_), .B(new_n9353_), .Y(new_n19510_));
  AOI21X1  g19318(.A0(new_n19510_), .A1(new_n19504_), .B0(new_n19509_), .Y(new_n19511_));
  OAI21X1  g19319(.A0(new_n19511_), .A1(new_n19493_), .B0(\asqrt[27] ), .Y(new_n19512_));
  NAND4X1  g19320(.A(\asqrt[9] ), .B(new_n18819_), .C(new_n18806_), .D(new_n18801_), .Y(new_n19513_));
  NAND2X1  g19321(.A(new_n18819_), .B(new_n18801_), .Y(new_n19514_));
  OAI21X1  g19322(.A0(new_n19514_), .A1(new_n19273_), .B0(new_n18810_), .Y(new_n19515_));
  AND2X1   g19323(.A(new_n19515_), .B(new_n19513_), .Y(new_n19516_));
  INVX1    g19324(.A(new_n19516_), .Y(new_n19517_));
  AOI21X1  g19325(.A0(new_n19502_), .A1(new_n19499_), .B0(new_n9833_), .Y(new_n19518_));
  AOI21X1  g19326(.A0(new_n19503_), .A1(new_n19494_), .B0(new_n19518_), .Y(new_n19519_));
  OAI21X1  g19327(.A0(new_n19519_), .A1(new_n9353_), .B0(new_n8874_), .Y(new_n19520_));
  OAI21X1  g19328(.A0(new_n19520_), .A1(new_n19511_), .B0(new_n19517_), .Y(new_n19521_));
  AOI21X1  g19329(.A0(new_n19521_), .A1(new_n19512_), .B0(new_n8412_), .Y(new_n19522_));
  AND2X1   g19330(.A(new_n18826_), .B(new_n18820_), .Y(new_n19523_));
  NOR3X1   g19331(.A(new_n19523_), .B(new_n18850_), .C(new_n18809_), .Y(new_n19524_));
  NOR3X1   g19332(.A(new_n19273_), .B(new_n19523_), .C(new_n18809_), .Y(new_n19525_));
  NOR2X1   g19333(.A(new_n19525_), .B(new_n18824_), .Y(new_n19526_));
  AOI21X1  g19334(.A0(new_n19524_), .A1(\asqrt[9] ), .B0(new_n19526_), .Y(new_n19527_));
  INVX1    g19335(.A(new_n19527_), .Y(new_n19528_));
  NAND3X1  g19336(.A(new_n19521_), .B(new_n19512_), .C(new_n8412_), .Y(new_n19529_));
  AOI21X1  g19337(.A0(new_n19529_), .A1(new_n19528_), .B0(new_n19522_), .Y(new_n19530_));
  OR2X1    g19338(.A(new_n19530_), .B(new_n7970_), .Y(new_n19531_));
  AND2X1   g19339(.A(new_n19529_), .B(new_n19528_), .Y(new_n19532_));
  AND2X1   g19340(.A(new_n18854_), .B(new_n18852_), .Y(new_n19533_));
  NOR3X1   g19341(.A(new_n19533_), .B(new_n18834_), .C(new_n18853_), .Y(new_n19534_));
  NOR3X1   g19342(.A(new_n19273_), .B(new_n19533_), .C(new_n18853_), .Y(new_n19535_));
  NOR2X1   g19343(.A(new_n19535_), .B(new_n18833_), .Y(new_n19536_));
  AOI21X1  g19344(.A0(new_n19534_), .A1(\asqrt[9] ), .B0(new_n19536_), .Y(new_n19537_));
  INVX1    g19345(.A(new_n19537_), .Y(new_n19538_));
  OR2X1    g19346(.A(new_n19519_), .B(new_n9353_), .Y(new_n19539_));
  AND2X1   g19347(.A(new_n19503_), .B(new_n19494_), .Y(new_n19540_));
  INVX1    g19348(.A(new_n19509_), .Y(new_n19541_));
  NAND2X1  g19349(.A(new_n19485_), .B(new_n9353_), .Y(new_n19542_));
  OAI21X1  g19350(.A0(new_n19542_), .A1(new_n19540_), .B0(new_n19541_), .Y(new_n19543_));
  AOI21X1  g19351(.A0(new_n19543_), .A1(new_n19539_), .B0(new_n8874_), .Y(new_n19544_));
  AOI21X1  g19352(.A0(new_n19492_), .A1(\asqrt[26] ), .B0(\asqrt[27] ), .Y(new_n19545_));
  AOI21X1  g19353(.A0(new_n19545_), .A1(new_n19543_), .B0(new_n19516_), .Y(new_n19546_));
  OAI21X1  g19354(.A0(new_n19546_), .A1(new_n19544_), .B0(\asqrt[28] ), .Y(new_n19547_));
  NAND2X1  g19355(.A(new_n19547_), .B(new_n7970_), .Y(new_n19548_));
  OAI21X1  g19356(.A0(new_n19548_), .A1(new_n19532_), .B0(new_n19538_), .Y(new_n19549_));
  AOI21X1  g19357(.A0(new_n19549_), .A1(new_n19531_), .B0(new_n7527_), .Y(new_n19550_));
  NAND4X1  g19358(.A(\asqrt[9] ), .B(new_n18845_), .C(new_n18843_), .D(new_n18863_), .Y(new_n19551_));
  OR2X1    g19359(.A(new_n18856_), .B(new_n18838_), .Y(new_n19552_));
  OAI21X1  g19360(.A0(new_n19552_), .A1(new_n19273_), .B0(new_n18844_), .Y(new_n19553_));
  AND2X1   g19361(.A(new_n19553_), .B(new_n19551_), .Y(new_n19554_));
  NOR3X1   g19362(.A(new_n19546_), .B(new_n19544_), .C(\asqrt[28] ), .Y(new_n19555_));
  OAI21X1  g19363(.A0(new_n19555_), .A1(new_n19527_), .B0(new_n19547_), .Y(new_n19556_));
  AOI21X1  g19364(.A0(new_n19556_), .A1(\asqrt[29] ), .B0(\asqrt[30] ), .Y(new_n19557_));
  AOI21X1  g19365(.A0(new_n19557_), .A1(new_n19549_), .B0(new_n19554_), .Y(new_n19558_));
  OAI21X1  g19366(.A0(new_n19558_), .A1(new_n19550_), .B0(\asqrt[31] ), .Y(new_n19559_));
  AOI21X1  g19367(.A0(new_n18900_), .A1(new_n18899_), .B0(new_n18862_), .Y(new_n19560_));
  AND2X1   g19368(.A(new_n19560_), .B(new_n18847_), .Y(new_n19561_));
  AOI22X1  g19369(.A0(new_n18900_), .A1(new_n18899_), .B0(new_n18872_), .B1(\asqrt[30] ), .Y(new_n19562_));
  AOI21X1  g19370(.A0(new_n19562_), .A1(\asqrt[9] ), .B0(new_n18861_), .Y(new_n19563_));
  AOI21X1  g19371(.A0(new_n19561_), .A1(\asqrt[9] ), .B0(new_n19563_), .Y(new_n19564_));
  NOR3X1   g19372(.A(new_n19558_), .B(new_n19550_), .C(\asqrt[31] ), .Y(new_n19565_));
  OAI21X1  g19373(.A0(new_n19565_), .A1(new_n19564_), .B0(new_n19559_), .Y(new_n19566_));
  AND2X1   g19374(.A(new_n19566_), .B(\asqrt[32] ), .Y(new_n19567_));
  INVX1    g19375(.A(new_n19564_), .Y(new_n19568_));
  AND2X1   g19376(.A(new_n19556_), .B(\asqrt[29] ), .Y(new_n19569_));
  NAND2X1  g19377(.A(new_n19529_), .B(new_n19528_), .Y(new_n19570_));
  AND2X1   g19378(.A(new_n19547_), .B(new_n7970_), .Y(new_n19571_));
  AOI21X1  g19379(.A0(new_n19571_), .A1(new_n19570_), .B0(new_n19537_), .Y(new_n19572_));
  OAI21X1  g19380(.A0(new_n19572_), .A1(new_n19569_), .B0(\asqrt[30] ), .Y(new_n19573_));
  INVX1    g19381(.A(new_n19554_), .Y(new_n19574_));
  OAI21X1  g19382(.A0(new_n19530_), .A1(new_n7970_), .B0(new_n7527_), .Y(new_n19575_));
  OAI21X1  g19383(.A0(new_n19575_), .A1(new_n19572_), .B0(new_n19574_), .Y(new_n19576_));
  NAND3X1  g19384(.A(new_n19576_), .B(new_n19573_), .C(new_n7103_), .Y(new_n19577_));
  NAND2X1  g19385(.A(new_n19577_), .B(new_n19568_), .Y(new_n19578_));
  AND2X1   g19386(.A(new_n18873_), .B(new_n18865_), .Y(new_n19579_));
  NOR3X1   g19387(.A(new_n19579_), .B(new_n18903_), .C(new_n18866_), .Y(new_n19580_));
  NOR3X1   g19388(.A(new_n19273_), .B(new_n19579_), .C(new_n18866_), .Y(new_n19581_));
  NOR2X1   g19389(.A(new_n19581_), .B(new_n18871_), .Y(new_n19582_));
  AOI21X1  g19390(.A0(new_n19580_), .A1(\asqrt[9] ), .B0(new_n19582_), .Y(new_n19583_));
  AND2X1   g19391(.A(new_n19559_), .B(new_n6699_), .Y(new_n19584_));
  AOI21X1  g19392(.A0(new_n19584_), .A1(new_n19578_), .B0(new_n19583_), .Y(new_n19585_));
  OAI21X1  g19393(.A0(new_n19585_), .A1(new_n19567_), .B0(\asqrt[33] ), .Y(new_n19586_));
  OR4X1    g19394(.A(new_n19273_), .B(new_n18881_), .C(new_n18907_), .D(new_n18906_), .Y(new_n19587_));
  OR2X1    g19395(.A(new_n18881_), .B(new_n18906_), .Y(new_n19588_));
  OAI21X1  g19396(.A0(new_n19588_), .A1(new_n19273_), .B0(new_n18907_), .Y(new_n19589_));
  AND2X1   g19397(.A(new_n19589_), .B(new_n19587_), .Y(new_n19590_));
  INVX1    g19398(.A(new_n19590_), .Y(new_n19591_));
  AOI21X1  g19399(.A0(new_n19576_), .A1(new_n19573_), .B0(new_n7103_), .Y(new_n19592_));
  AOI21X1  g19400(.A0(new_n19577_), .A1(new_n19568_), .B0(new_n19592_), .Y(new_n19593_));
  OAI21X1  g19401(.A0(new_n19593_), .A1(new_n6699_), .B0(new_n6294_), .Y(new_n19594_));
  OAI21X1  g19402(.A0(new_n19594_), .A1(new_n19585_), .B0(new_n19591_), .Y(new_n19595_));
  AOI21X1  g19403(.A0(new_n19595_), .A1(new_n19586_), .B0(new_n5941_), .Y(new_n19596_));
  AND2X1   g19404(.A(new_n18889_), .B(new_n18884_), .Y(new_n19597_));
  NOR3X1   g19405(.A(new_n19597_), .B(new_n18938_), .C(new_n18883_), .Y(new_n19598_));
  NOR3X1   g19406(.A(new_n19273_), .B(new_n19597_), .C(new_n18883_), .Y(new_n19599_));
  NOR2X1   g19407(.A(new_n19599_), .B(new_n18888_), .Y(new_n19600_));
  AOI21X1  g19408(.A0(new_n19598_), .A1(\asqrt[9] ), .B0(new_n19600_), .Y(new_n19601_));
  INVX1    g19409(.A(new_n19601_), .Y(new_n19602_));
  NAND3X1  g19410(.A(new_n19595_), .B(new_n19586_), .C(new_n5941_), .Y(new_n19603_));
  AOI21X1  g19411(.A0(new_n19603_), .A1(new_n19602_), .B0(new_n19596_), .Y(new_n19604_));
  OR2X1    g19412(.A(new_n19604_), .B(new_n5541_), .Y(new_n19605_));
  AND2X1   g19413(.A(new_n19603_), .B(new_n19602_), .Y(new_n19606_));
  AND2X1   g19414(.A(new_n18942_), .B(new_n18940_), .Y(new_n19607_));
  NOR3X1   g19415(.A(new_n19607_), .B(new_n18897_), .C(new_n18941_), .Y(new_n19608_));
  NOR3X1   g19416(.A(new_n19273_), .B(new_n19607_), .C(new_n18941_), .Y(new_n19609_));
  NOR2X1   g19417(.A(new_n19609_), .B(new_n18896_), .Y(new_n19610_));
  AOI21X1  g19418(.A0(new_n19608_), .A1(\asqrt[9] ), .B0(new_n19610_), .Y(new_n19611_));
  INVX1    g19419(.A(new_n19611_), .Y(new_n19612_));
  OR2X1    g19420(.A(new_n19593_), .B(new_n6699_), .Y(new_n19613_));
  AND2X1   g19421(.A(new_n19577_), .B(new_n19568_), .Y(new_n19614_));
  INVX1    g19422(.A(new_n19583_), .Y(new_n19615_));
  NAND2X1  g19423(.A(new_n19559_), .B(new_n6699_), .Y(new_n19616_));
  OAI21X1  g19424(.A0(new_n19616_), .A1(new_n19614_), .B0(new_n19615_), .Y(new_n19617_));
  AOI21X1  g19425(.A0(new_n19617_), .A1(new_n19613_), .B0(new_n6294_), .Y(new_n19618_));
  AOI21X1  g19426(.A0(new_n19566_), .A1(\asqrt[32] ), .B0(\asqrt[33] ), .Y(new_n19619_));
  AOI21X1  g19427(.A0(new_n19619_), .A1(new_n19617_), .B0(new_n19590_), .Y(new_n19620_));
  OAI21X1  g19428(.A0(new_n19620_), .A1(new_n19618_), .B0(\asqrt[34] ), .Y(new_n19621_));
  NAND2X1  g19429(.A(new_n19621_), .B(new_n5541_), .Y(new_n19622_));
  OAI21X1  g19430(.A0(new_n19622_), .A1(new_n19606_), .B0(new_n19612_), .Y(new_n19623_));
  AOI21X1  g19431(.A0(new_n19623_), .A1(new_n19605_), .B0(new_n5176_), .Y(new_n19624_));
  NAND4X1  g19432(.A(\asqrt[9] ), .B(new_n18919_), .C(new_n18917_), .D(new_n18944_), .Y(new_n19625_));
  NAND2X1  g19433(.A(new_n18919_), .B(new_n18944_), .Y(new_n19626_));
  OAI21X1  g19434(.A0(new_n19626_), .A1(new_n19273_), .B0(new_n18918_), .Y(new_n19627_));
  AND2X1   g19435(.A(new_n19627_), .B(new_n19625_), .Y(new_n19628_));
  NOR3X1   g19436(.A(new_n19620_), .B(new_n19618_), .C(\asqrt[34] ), .Y(new_n19629_));
  OAI21X1  g19437(.A0(new_n19629_), .A1(new_n19601_), .B0(new_n19621_), .Y(new_n19630_));
  AOI21X1  g19438(.A0(new_n19630_), .A1(\asqrt[35] ), .B0(\asqrt[36] ), .Y(new_n19631_));
  AOI21X1  g19439(.A0(new_n19631_), .A1(new_n19623_), .B0(new_n19628_), .Y(new_n19632_));
  OAI21X1  g19440(.A0(new_n19632_), .A1(new_n19624_), .B0(\asqrt[37] ), .Y(new_n19633_));
  AOI21X1  g19441(.A0(new_n18974_), .A1(new_n18973_), .B0(new_n18927_), .Y(new_n19634_));
  AND2X1   g19442(.A(new_n19634_), .B(new_n18921_), .Y(new_n19635_));
  AOI22X1  g19443(.A0(new_n18974_), .A1(new_n18973_), .B0(new_n18946_), .B1(\asqrt[36] ), .Y(new_n19636_));
  AOI21X1  g19444(.A0(new_n19636_), .A1(\asqrt[9] ), .B0(new_n18926_), .Y(new_n19637_));
  AOI21X1  g19445(.A0(new_n19635_), .A1(\asqrt[9] ), .B0(new_n19637_), .Y(new_n19638_));
  NOR3X1   g19446(.A(new_n19632_), .B(new_n19624_), .C(\asqrt[37] ), .Y(new_n19639_));
  OAI21X1  g19447(.A0(new_n19639_), .A1(new_n19638_), .B0(new_n19633_), .Y(new_n19640_));
  AND2X1   g19448(.A(new_n19640_), .B(\asqrt[38] ), .Y(new_n19641_));
  INVX1    g19449(.A(new_n19638_), .Y(new_n19642_));
  AND2X1   g19450(.A(new_n19630_), .B(\asqrt[35] ), .Y(new_n19643_));
  NAND2X1  g19451(.A(new_n19603_), .B(new_n19602_), .Y(new_n19644_));
  AND2X1   g19452(.A(new_n19621_), .B(new_n5541_), .Y(new_n19645_));
  AOI21X1  g19453(.A0(new_n19645_), .A1(new_n19644_), .B0(new_n19611_), .Y(new_n19646_));
  OAI21X1  g19454(.A0(new_n19646_), .A1(new_n19643_), .B0(\asqrt[36] ), .Y(new_n19647_));
  INVX1    g19455(.A(new_n19628_), .Y(new_n19648_));
  OAI21X1  g19456(.A0(new_n19604_), .A1(new_n5541_), .B0(new_n5176_), .Y(new_n19649_));
  OAI21X1  g19457(.A0(new_n19649_), .A1(new_n19646_), .B0(new_n19648_), .Y(new_n19650_));
  NAND3X1  g19458(.A(new_n19650_), .B(new_n19647_), .C(new_n4826_), .Y(new_n19651_));
  NAND2X1  g19459(.A(new_n19651_), .B(new_n19642_), .Y(new_n19652_));
  AND2X1   g19460(.A(new_n18947_), .B(new_n18929_), .Y(new_n19653_));
  NOR3X1   g19461(.A(new_n19653_), .B(new_n18977_), .C(new_n18930_), .Y(new_n19654_));
  NOR3X1   g19462(.A(new_n19273_), .B(new_n19653_), .C(new_n18930_), .Y(new_n19655_));
  NOR2X1   g19463(.A(new_n19655_), .B(new_n18935_), .Y(new_n19656_));
  AOI21X1  g19464(.A0(new_n19654_), .A1(\asqrt[9] ), .B0(new_n19656_), .Y(new_n19657_));
  AND2X1   g19465(.A(new_n19633_), .B(new_n4493_), .Y(new_n19658_));
  AOI21X1  g19466(.A0(new_n19658_), .A1(new_n19652_), .B0(new_n19657_), .Y(new_n19659_));
  OAI21X1  g19467(.A0(new_n19659_), .A1(new_n19641_), .B0(\asqrt[39] ), .Y(new_n19660_));
  OR4X1    g19468(.A(new_n19273_), .B(new_n18955_), .C(new_n18981_), .D(new_n18980_), .Y(new_n19661_));
  OR2X1    g19469(.A(new_n18955_), .B(new_n18980_), .Y(new_n19662_));
  OAI21X1  g19470(.A0(new_n19662_), .A1(new_n19273_), .B0(new_n18981_), .Y(new_n19663_));
  AND2X1   g19471(.A(new_n19663_), .B(new_n19661_), .Y(new_n19664_));
  INVX1    g19472(.A(new_n19664_), .Y(new_n19665_));
  AOI21X1  g19473(.A0(new_n19650_), .A1(new_n19647_), .B0(new_n4826_), .Y(new_n19666_));
  AOI21X1  g19474(.A0(new_n19651_), .A1(new_n19642_), .B0(new_n19666_), .Y(new_n19667_));
  OAI21X1  g19475(.A0(new_n19667_), .A1(new_n4493_), .B0(new_n4165_), .Y(new_n19668_));
  OAI21X1  g19476(.A0(new_n19668_), .A1(new_n19659_), .B0(new_n19665_), .Y(new_n19669_));
  AOI21X1  g19477(.A0(new_n19669_), .A1(new_n19660_), .B0(new_n3863_), .Y(new_n19670_));
  AND2X1   g19478(.A(new_n18963_), .B(new_n18958_), .Y(new_n19671_));
  NOR3X1   g19479(.A(new_n19671_), .B(new_n18998_), .C(new_n18957_), .Y(new_n19672_));
  NOR3X1   g19480(.A(new_n19273_), .B(new_n19671_), .C(new_n18957_), .Y(new_n19673_));
  NOR2X1   g19481(.A(new_n19673_), .B(new_n18962_), .Y(new_n19674_));
  AOI21X1  g19482(.A0(new_n19672_), .A1(\asqrt[9] ), .B0(new_n19674_), .Y(new_n19675_));
  INVX1    g19483(.A(new_n19675_), .Y(new_n19676_));
  NAND3X1  g19484(.A(new_n19669_), .B(new_n19660_), .C(new_n3863_), .Y(new_n19677_));
  AOI21X1  g19485(.A0(new_n19677_), .A1(new_n19676_), .B0(new_n19670_), .Y(new_n19678_));
  OR2X1    g19486(.A(new_n19678_), .B(new_n3564_), .Y(new_n19679_));
  OR2X1    g19487(.A(new_n19667_), .B(new_n4493_), .Y(new_n19680_));
  AND2X1   g19488(.A(new_n19651_), .B(new_n19642_), .Y(new_n19681_));
  INVX1    g19489(.A(new_n19657_), .Y(new_n19682_));
  NAND2X1  g19490(.A(new_n19633_), .B(new_n4493_), .Y(new_n19683_));
  OAI21X1  g19491(.A0(new_n19683_), .A1(new_n19681_), .B0(new_n19682_), .Y(new_n19684_));
  AOI21X1  g19492(.A0(new_n19684_), .A1(new_n19680_), .B0(new_n4165_), .Y(new_n19685_));
  AOI21X1  g19493(.A0(new_n19640_), .A1(\asqrt[38] ), .B0(\asqrt[39] ), .Y(new_n19686_));
  AOI21X1  g19494(.A0(new_n19686_), .A1(new_n19684_), .B0(new_n19664_), .Y(new_n19687_));
  NOR3X1   g19495(.A(new_n19687_), .B(new_n19685_), .C(\asqrt[40] ), .Y(new_n19688_));
  NOR2X1   g19496(.A(new_n19688_), .B(new_n19675_), .Y(new_n19689_));
  AND2X1   g19497(.A(new_n19002_), .B(new_n19000_), .Y(new_n19690_));
  NOR3X1   g19498(.A(new_n19690_), .B(new_n18971_), .C(new_n19001_), .Y(new_n19691_));
  NOR3X1   g19499(.A(new_n19273_), .B(new_n19690_), .C(new_n19001_), .Y(new_n19692_));
  NOR2X1   g19500(.A(new_n19692_), .B(new_n18970_), .Y(new_n19693_));
  AOI21X1  g19501(.A0(new_n19691_), .A1(\asqrt[9] ), .B0(new_n19693_), .Y(new_n19694_));
  INVX1    g19502(.A(new_n19694_), .Y(new_n19695_));
  OAI21X1  g19503(.A0(new_n19687_), .A1(new_n19685_), .B0(\asqrt[40] ), .Y(new_n19696_));
  NAND2X1  g19504(.A(new_n19696_), .B(new_n3564_), .Y(new_n19697_));
  OAI21X1  g19505(.A0(new_n19697_), .A1(new_n19689_), .B0(new_n19695_), .Y(new_n19698_));
  AOI21X1  g19506(.A0(new_n19698_), .A1(new_n19679_), .B0(new_n3276_), .Y(new_n19699_));
  OR4X1    g19507(.A(new_n19273_), .B(new_n19004_), .C(new_n18992_), .D(new_n18986_), .Y(new_n19700_));
  OR2X1    g19508(.A(new_n19004_), .B(new_n18986_), .Y(new_n19701_));
  OAI21X1  g19509(.A0(new_n19701_), .A1(new_n19273_), .B0(new_n18992_), .Y(new_n19702_));
  AND2X1   g19510(.A(new_n19702_), .B(new_n19700_), .Y(new_n19703_));
  OAI21X1  g19511(.A0(new_n19688_), .A1(new_n19675_), .B0(new_n19696_), .Y(new_n19704_));
  AOI21X1  g19512(.A0(new_n19704_), .A1(\asqrt[41] ), .B0(\asqrt[42] ), .Y(new_n19705_));
  AOI21X1  g19513(.A0(new_n19705_), .A1(new_n19698_), .B0(new_n19703_), .Y(new_n19706_));
  OAI21X1  g19514(.A0(new_n19706_), .A1(new_n19699_), .B0(\asqrt[43] ), .Y(new_n19707_));
  AOI21X1  g19515(.A0(new_n19048_), .A1(new_n19047_), .B0(new_n19010_), .Y(new_n19708_));
  AND2X1   g19516(.A(new_n19708_), .B(new_n18995_), .Y(new_n19709_));
  AOI22X1  g19517(.A0(new_n19048_), .A1(new_n19047_), .B0(new_n19020_), .B1(\asqrt[42] ), .Y(new_n19710_));
  AOI21X1  g19518(.A0(new_n19710_), .A1(\asqrt[9] ), .B0(new_n19009_), .Y(new_n19711_));
  AOI21X1  g19519(.A0(new_n19709_), .A1(\asqrt[9] ), .B0(new_n19711_), .Y(new_n19712_));
  NOR3X1   g19520(.A(new_n19706_), .B(new_n19699_), .C(\asqrt[43] ), .Y(new_n19713_));
  OAI21X1  g19521(.A0(new_n19713_), .A1(new_n19712_), .B0(new_n19707_), .Y(new_n19714_));
  AND2X1   g19522(.A(new_n19714_), .B(\asqrt[44] ), .Y(new_n19715_));
  OR2X1    g19523(.A(new_n19713_), .B(new_n19712_), .Y(new_n19716_));
  AND2X1   g19524(.A(new_n19021_), .B(new_n19013_), .Y(new_n19717_));
  NOR3X1   g19525(.A(new_n19717_), .B(new_n19051_), .C(new_n19014_), .Y(new_n19718_));
  NOR3X1   g19526(.A(new_n19273_), .B(new_n19717_), .C(new_n19014_), .Y(new_n19719_));
  NOR2X1   g19527(.A(new_n19719_), .B(new_n19019_), .Y(new_n19720_));
  AOI21X1  g19528(.A0(new_n19718_), .A1(\asqrt[9] ), .B0(new_n19720_), .Y(new_n19721_));
  AND2X1   g19529(.A(new_n19707_), .B(new_n2769_), .Y(new_n19722_));
  AOI21X1  g19530(.A0(new_n19722_), .A1(new_n19716_), .B0(new_n19721_), .Y(new_n19723_));
  OAI21X1  g19531(.A0(new_n19723_), .A1(new_n19715_), .B0(\asqrt[45] ), .Y(new_n19724_));
  OR4X1    g19532(.A(new_n19273_), .B(new_n19029_), .C(new_n19055_), .D(new_n19054_), .Y(new_n19725_));
  OR2X1    g19533(.A(new_n19029_), .B(new_n19054_), .Y(new_n19726_));
  OAI21X1  g19534(.A0(new_n19726_), .A1(new_n19273_), .B0(new_n19055_), .Y(new_n19727_));
  AND2X1   g19535(.A(new_n19727_), .B(new_n19725_), .Y(new_n19728_));
  INVX1    g19536(.A(new_n19728_), .Y(new_n19729_));
  AND2X1   g19537(.A(new_n19704_), .B(\asqrt[41] ), .Y(new_n19730_));
  OR2X1    g19538(.A(new_n19688_), .B(new_n19675_), .Y(new_n19731_));
  AND2X1   g19539(.A(new_n19696_), .B(new_n3564_), .Y(new_n19732_));
  AOI21X1  g19540(.A0(new_n19732_), .A1(new_n19731_), .B0(new_n19694_), .Y(new_n19733_));
  OAI21X1  g19541(.A0(new_n19733_), .A1(new_n19730_), .B0(\asqrt[42] ), .Y(new_n19734_));
  INVX1    g19542(.A(new_n19703_), .Y(new_n19735_));
  OAI21X1  g19543(.A0(new_n19678_), .A1(new_n3564_), .B0(new_n3276_), .Y(new_n19736_));
  OAI21X1  g19544(.A0(new_n19736_), .A1(new_n19733_), .B0(new_n19735_), .Y(new_n19737_));
  AOI21X1  g19545(.A0(new_n19737_), .A1(new_n19734_), .B0(new_n3008_), .Y(new_n19738_));
  INVX1    g19546(.A(new_n19712_), .Y(new_n19739_));
  NAND3X1  g19547(.A(new_n19737_), .B(new_n19734_), .C(new_n3008_), .Y(new_n19740_));
  AOI21X1  g19548(.A0(new_n19740_), .A1(new_n19739_), .B0(new_n19738_), .Y(new_n19741_));
  OAI21X1  g19549(.A0(new_n19741_), .A1(new_n2769_), .B0(new_n2570_), .Y(new_n19742_));
  OAI21X1  g19550(.A0(new_n19742_), .A1(new_n19723_), .B0(new_n19729_), .Y(new_n19743_));
  AOI21X1  g19551(.A0(new_n19743_), .A1(new_n19724_), .B0(new_n2263_), .Y(new_n19744_));
  AND2X1   g19552(.A(new_n19037_), .B(new_n19032_), .Y(new_n19745_));
  NOR3X1   g19553(.A(new_n19745_), .B(new_n19072_), .C(new_n19031_), .Y(new_n19746_));
  NOR3X1   g19554(.A(new_n19273_), .B(new_n19745_), .C(new_n19031_), .Y(new_n19747_));
  NOR2X1   g19555(.A(new_n19747_), .B(new_n19036_), .Y(new_n19748_));
  AOI21X1  g19556(.A0(new_n19746_), .A1(\asqrt[9] ), .B0(new_n19748_), .Y(new_n19749_));
  INVX1    g19557(.A(new_n19749_), .Y(new_n19750_));
  NAND3X1  g19558(.A(new_n19743_), .B(new_n19724_), .C(new_n2263_), .Y(new_n19751_));
  AOI21X1  g19559(.A0(new_n19751_), .A1(new_n19750_), .B0(new_n19744_), .Y(new_n19752_));
  OR2X1    g19560(.A(new_n19752_), .B(new_n2040_), .Y(new_n19753_));
  OR2X1    g19561(.A(new_n19741_), .B(new_n2769_), .Y(new_n19754_));
  NOR2X1   g19562(.A(new_n19713_), .B(new_n19712_), .Y(new_n19755_));
  INVX1    g19563(.A(new_n19721_), .Y(new_n19756_));
  NAND2X1  g19564(.A(new_n19707_), .B(new_n2769_), .Y(new_n19757_));
  OAI21X1  g19565(.A0(new_n19757_), .A1(new_n19755_), .B0(new_n19756_), .Y(new_n19758_));
  AOI21X1  g19566(.A0(new_n19758_), .A1(new_n19754_), .B0(new_n2570_), .Y(new_n19759_));
  AOI21X1  g19567(.A0(new_n19714_), .A1(\asqrt[44] ), .B0(\asqrt[45] ), .Y(new_n19760_));
  AOI21X1  g19568(.A0(new_n19760_), .A1(new_n19758_), .B0(new_n19728_), .Y(new_n19761_));
  NOR3X1   g19569(.A(new_n19761_), .B(new_n19759_), .C(\asqrt[46] ), .Y(new_n19762_));
  NOR2X1   g19570(.A(new_n19762_), .B(new_n19749_), .Y(new_n19763_));
  AND2X1   g19571(.A(new_n19076_), .B(new_n19074_), .Y(new_n19764_));
  NOR3X1   g19572(.A(new_n19764_), .B(new_n19045_), .C(new_n19075_), .Y(new_n19765_));
  NOR3X1   g19573(.A(new_n19273_), .B(new_n19764_), .C(new_n19075_), .Y(new_n19766_));
  NOR2X1   g19574(.A(new_n19766_), .B(new_n19044_), .Y(new_n19767_));
  AOI21X1  g19575(.A0(new_n19765_), .A1(\asqrt[9] ), .B0(new_n19767_), .Y(new_n19768_));
  INVX1    g19576(.A(new_n19768_), .Y(new_n19769_));
  OAI21X1  g19577(.A0(new_n19761_), .A1(new_n19759_), .B0(\asqrt[46] ), .Y(new_n19770_));
  NAND2X1  g19578(.A(new_n19770_), .B(new_n2040_), .Y(new_n19771_));
  OAI21X1  g19579(.A0(new_n19771_), .A1(new_n19763_), .B0(new_n19769_), .Y(new_n19772_));
  AOI21X1  g19580(.A0(new_n19772_), .A1(new_n19753_), .B0(new_n1834_), .Y(new_n19773_));
  OR4X1    g19581(.A(new_n19273_), .B(new_n19078_), .C(new_n19066_), .D(new_n19060_), .Y(new_n19774_));
  OR2X1    g19582(.A(new_n19078_), .B(new_n19060_), .Y(new_n19775_));
  OAI21X1  g19583(.A0(new_n19775_), .A1(new_n19273_), .B0(new_n19066_), .Y(new_n19776_));
  AND2X1   g19584(.A(new_n19776_), .B(new_n19774_), .Y(new_n19777_));
  OAI21X1  g19585(.A0(new_n19762_), .A1(new_n19749_), .B0(new_n19770_), .Y(new_n19778_));
  AOI21X1  g19586(.A0(new_n19778_), .A1(\asqrt[47] ), .B0(\asqrt[48] ), .Y(new_n19779_));
  AOI21X1  g19587(.A0(new_n19779_), .A1(new_n19772_), .B0(new_n19777_), .Y(new_n19780_));
  OAI21X1  g19588(.A0(new_n19780_), .A1(new_n19773_), .B0(\asqrt[49] ), .Y(new_n19781_));
  AOI21X1  g19589(.A0(new_n19122_), .A1(new_n19121_), .B0(new_n19084_), .Y(new_n19782_));
  AND2X1   g19590(.A(new_n19782_), .B(new_n19069_), .Y(new_n19783_));
  AOI22X1  g19591(.A0(new_n19122_), .A1(new_n19121_), .B0(new_n19094_), .B1(\asqrt[48] ), .Y(new_n19784_));
  AOI21X1  g19592(.A0(new_n19784_), .A1(\asqrt[9] ), .B0(new_n19083_), .Y(new_n19785_));
  AOI21X1  g19593(.A0(new_n19783_), .A1(\asqrt[9] ), .B0(new_n19785_), .Y(new_n19786_));
  NOR3X1   g19594(.A(new_n19780_), .B(new_n19773_), .C(\asqrt[49] ), .Y(new_n19787_));
  OAI21X1  g19595(.A0(new_n19787_), .A1(new_n19786_), .B0(new_n19781_), .Y(new_n19788_));
  AND2X1   g19596(.A(new_n19788_), .B(\asqrt[50] ), .Y(new_n19789_));
  OR2X1    g19597(.A(new_n19787_), .B(new_n19786_), .Y(new_n19790_));
  AND2X1   g19598(.A(new_n19095_), .B(new_n19087_), .Y(new_n19791_));
  NOR3X1   g19599(.A(new_n19791_), .B(new_n19125_), .C(new_n19088_), .Y(new_n19792_));
  NOR3X1   g19600(.A(new_n19273_), .B(new_n19791_), .C(new_n19088_), .Y(new_n19793_));
  NOR2X1   g19601(.A(new_n19793_), .B(new_n19093_), .Y(new_n19794_));
  AOI21X1  g19602(.A0(new_n19792_), .A1(\asqrt[9] ), .B0(new_n19794_), .Y(new_n19795_));
  AND2X1   g19603(.A(new_n19781_), .B(new_n1469_), .Y(new_n19796_));
  AOI21X1  g19604(.A0(new_n19796_), .A1(new_n19790_), .B0(new_n19795_), .Y(new_n19797_));
  OAI21X1  g19605(.A0(new_n19797_), .A1(new_n19789_), .B0(\asqrt[51] ), .Y(new_n19798_));
  OR4X1    g19606(.A(new_n19273_), .B(new_n19103_), .C(new_n19129_), .D(new_n19128_), .Y(new_n19799_));
  OR2X1    g19607(.A(new_n19103_), .B(new_n19128_), .Y(new_n19800_));
  OAI21X1  g19608(.A0(new_n19800_), .A1(new_n19273_), .B0(new_n19129_), .Y(new_n19801_));
  AND2X1   g19609(.A(new_n19801_), .B(new_n19799_), .Y(new_n19802_));
  INVX1    g19610(.A(new_n19802_), .Y(new_n19803_));
  AND2X1   g19611(.A(new_n19778_), .B(\asqrt[47] ), .Y(new_n19804_));
  OR2X1    g19612(.A(new_n19762_), .B(new_n19749_), .Y(new_n19805_));
  AND2X1   g19613(.A(new_n19770_), .B(new_n2040_), .Y(new_n19806_));
  AOI21X1  g19614(.A0(new_n19806_), .A1(new_n19805_), .B0(new_n19768_), .Y(new_n19807_));
  OAI21X1  g19615(.A0(new_n19807_), .A1(new_n19804_), .B0(\asqrt[48] ), .Y(new_n19808_));
  INVX1    g19616(.A(new_n19777_), .Y(new_n19809_));
  OAI21X1  g19617(.A0(new_n19752_), .A1(new_n2040_), .B0(new_n1834_), .Y(new_n19810_));
  OAI21X1  g19618(.A0(new_n19810_), .A1(new_n19807_), .B0(new_n19809_), .Y(new_n19811_));
  AOI21X1  g19619(.A0(new_n19811_), .A1(new_n19808_), .B0(new_n1632_), .Y(new_n19812_));
  INVX1    g19620(.A(new_n19786_), .Y(new_n19813_));
  NAND3X1  g19621(.A(new_n19811_), .B(new_n19808_), .C(new_n1632_), .Y(new_n19814_));
  AOI21X1  g19622(.A0(new_n19814_), .A1(new_n19813_), .B0(new_n19812_), .Y(new_n19815_));
  OAI21X1  g19623(.A0(new_n19815_), .A1(new_n1469_), .B0(new_n1277_), .Y(new_n19816_));
  OAI21X1  g19624(.A0(new_n19816_), .A1(new_n19797_), .B0(new_n19803_), .Y(new_n19817_));
  AOI21X1  g19625(.A0(new_n19817_), .A1(new_n19798_), .B0(new_n1111_), .Y(new_n19818_));
  AND2X1   g19626(.A(new_n19111_), .B(new_n19106_), .Y(new_n19819_));
  NOR3X1   g19627(.A(new_n19819_), .B(new_n19146_), .C(new_n19105_), .Y(new_n19820_));
  NOR3X1   g19628(.A(new_n19273_), .B(new_n19819_), .C(new_n19105_), .Y(new_n19821_));
  NOR2X1   g19629(.A(new_n19821_), .B(new_n19110_), .Y(new_n19822_));
  AOI21X1  g19630(.A0(new_n19820_), .A1(\asqrt[9] ), .B0(new_n19822_), .Y(new_n19823_));
  INVX1    g19631(.A(new_n19823_), .Y(new_n19824_));
  NAND3X1  g19632(.A(new_n19817_), .B(new_n19798_), .C(new_n1111_), .Y(new_n19825_));
  AOI21X1  g19633(.A0(new_n19825_), .A1(new_n19824_), .B0(new_n19818_), .Y(new_n19826_));
  OR2X1    g19634(.A(new_n19826_), .B(new_n968_), .Y(new_n19827_));
  OR2X1    g19635(.A(new_n19815_), .B(new_n1469_), .Y(new_n19828_));
  NOR2X1   g19636(.A(new_n19787_), .B(new_n19786_), .Y(new_n19829_));
  INVX1    g19637(.A(new_n19795_), .Y(new_n19830_));
  NAND2X1  g19638(.A(new_n19781_), .B(new_n1469_), .Y(new_n19831_));
  OAI21X1  g19639(.A0(new_n19831_), .A1(new_n19829_), .B0(new_n19830_), .Y(new_n19832_));
  AOI21X1  g19640(.A0(new_n19832_), .A1(new_n19828_), .B0(new_n1277_), .Y(new_n19833_));
  AOI21X1  g19641(.A0(new_n19788_), .A1(\asqrt[50] ), .B0(\asqrt[51] ), .Y(new_n19834_));
  AOI21X1  g19642(.A0(new_n19834_), .A1(new_n19832_), .B0(new_n19802_), .Y(new_n19835_));
  NOR3X1   g19643(.A(new_n19835_), .B(new_n19833_), .C(\asqrt[52] ), .Y(new_n19836_));
  NOR2X1   g19644(.A(new_n19836_), .B(new_n19823_), .Y(new_n19837_));
  AND2X1   g19645(.A(new_n19150_), .B(new_n19148_), .Y(new_n19838_));
  NOR3X1   g19646(.A(new_n19838_), .B(new_n19119_), .C(new_n19149_), .Y(new_n19839_));
  NOR3X1   g19647(.A(new_n19273_), .B(new_n19838_), .C(new_n19149_), .Y(new_n19840_));
  NOR2X1   g19648(.A(new_n19840_), .B(new_n19118_), .Y(new_n19841_));
  AOI21X1  g19649(.A0(new_n19839_), .A1(\asqrt[9] ), .B0(new_n19841_), .Y(new_n19842_));
  INVX1    g19650(.A(new_n19842_), .Y(new_n19843_));
  OAI21X1  g19651(.A0(new_n19835_), .A1(new_n19833_), .B0(\asqrt[52] ), .Y(new_n19844_));
  NAND2X1  g19652(.A(new_n19844_), .B(new_n968_), .Y(new_n19845_));
  OAI21X1  g19653(.A0(new_n19845_), .A1(new_n19837_), .B0(new_n19843_), .Y(new_n19846_));
  AOI21X1  g19654(.A0(new_n19846_), .A1(new_n19827_), .B0(new_n902_), .Y(new_n19847_));
  NAND4X1  g19655(.A(\asqrt[9] ), .B(new_n19141_), .C(new_n19139_), .D(new_n19159_), .Y(new_n19848_));
  OR2X1    g19656(.A(new_n19152_), .B(new_n19134_), .Y(new_n19849_));
  OAI21X1  g19657(.A0(new_n19849_), .A1(new_n19273_), .B0(new_n19140_), .Y(new_n19850_));
  AND2X1   g19658(.A(new_n19850_), .B(new_n19848_), .Y(new_n19851_));
  OAI21X1  g19659(.A0(new_n19836_), .A1(new_n19823_), .B0(new_n19844_), .Y(new_n19852_));
  AOI21X1  g19660(.A0(new_n19852_), .A1(\asqrt[53] ), .B0(\asqrt[54] ), .Y(new_n19853_));
  AOI21X1  g19661(.A0(new_n19853_), .A1(new_n19846_), .B0(new_n19851_), .Y(new_n19854_));
  OAI21X1  g19662(.A0(new_n19854_), .A1(new_n19847_), .B0(\asqrt[55] ), .Y(new_n19855_));
  AOI21X1  g19663(.A0(new_n19196_), .A1(new_n19195_), .B0(new_n19158_), .Y(new_n19856_));
  AND2X1   g19664(.A(new_n19856_), .B(new_n19143_), .Y(new_n19857_));
  AOI22X1  g19665(.A0(new_n19196_), .A1(new_n19195_), .B0(new_n19163_), .B1(\asqrt[54] ), .Y(new_n19858_));
  AOI21X1  g19666(.A0(new_n19858_), .A1(\asqrt[9] ), .B0(new_n19157_), .Y(new_n19859_));
  AOI21X1  g19667(.A0(new_n19857_), .A1(\asqrt[9] ), .B0(new_n19859_), .Y(new_n19860_));
  NOR3X1   g19668(.A(new_n19854_), .B(new_n19847_), .C(\asqrt[55] ), .Y(new_n19861_));
  OAI21X1  g19669(.A0(new_n19861_), .A1(new_n19860_), .B0(new_n19855_), .Y(new_n19862_));
  AND2X1   g19670(.A(new_n19862_), .B(\asqrt[56] ), .Y(new_n19863_));
  OR2X1    g19671(.A(new_n19861_), .B(new_n19860_), .Y(new_n19864_));
  AND2X1   g19672(.A(new_n19855_), .B(new_n582_), .Y(new_n19865_));
  AND2X1   g19673(.A(new_n19164_), .B(new_n19161_), .Y(new_n19866_));
  NOR3X1   g19674(.A(new_n19200_), .B(new_n19866_), .C(new_n19162_), .Y(new_n19867_));
  NOR3X1   g19675(.A(new_n19273_), .B(new_n19866_), .C(new_n19162_), .Y(new_n19868_));
  NOR2X1   g19676(.A(new_n19868_), .B(new_n19169_), .Y(new_n19869_));
  AOI21X1  g19677(.A0(new_n19867_), .A1(\asqrt[9] ), .B0(new_n19869_), .Y(new_n19870_));
  AOI21X1  g19678(.A0(new_n19865_), .A1(new_n19864_), .B0(new_n19870_), .Y(new_n19871_));
  OAI21X1  g19679(.A0(new_n19871_), .A1(new_n19863_), .B0(\asqrt[57] ), .Y(new_n19872_));
  NAND4X1  g19680(.A(\asqrt[9] ), .B(new_n19204_), .C(new_n19176_), .D(new_n19171_), .Y(new_n19873_));
  OR2X1    g19681(.A(new_n19177_), .B(new_n19202_), .Y(new_n19874_));
  OAI21X1  g19682(.A0(new_n19874_), .A1(new_n19273_), .B0(new_n19203_), .Y(new_n19875_));
  AND2X1   g19683(.A(new_n19875_), .B(new_n19873_), .Y(new_n19876_));
  INVX1    g19684(.A(new_n19876_), .Y(new_n19877_));
  AND2X1   g19685(.A(new_n19852_), .B(\asqrt[53] ), .Y(new_n19878_));
  OR2X1    g19686(.A(new_n19836_), .B(new_n19823_), .Y(new_n19879_));
  AND2X1   g19687(.A(new_n19844_), .B(new_n968_), .Y(new_n19880_));
  AOI21X1  g19688(.A0(new_n19880_), .A1(new_n19879_), .B0(new_n19842_), .Y(new_n19881_));
  OAI21X1  g19689(.A0(new_n19881_), .A1(new_n19878_), .B0(\asqrt[54] ), .Y(new_n19882_));
  INVX1    g19690(.A(new_n19851_), .Y(new_n19883_));
  OAI21X1  g19691(.A0(new_n19826_), .A1(new_n968_), .B0(new_n902_), .Y(new_n19884_));
  OAI21X1  g19692(.A0(new_n19884_), .A1(new_n19881_), .B0(new_n19883_), .Y(new_n19885_));
  AOI21X1  g19693(.A0(new_n19885_), .A1(new_n19882_), .B0(new_n697_), .Y(new_n19886_));
  INVX1    g19694(.A(new_n19860_), .Y(new_n19887_));
  NAND3X1  g19695(.A(new_n19885_), .B(new_n19882_), .C(new_n697_), .Y(new_n19888_));
  AOI21X1  g19696(.A0(new_n19888_), .A1(new_n19887_), .B0(new_n19886_), .Y(new_n19889_));
  OAI21X1  g19697(.A0(new_n19889_), .A1(new_n582_), .B0(new_n481_), .Y(new_n19890_));
  OAI21X1  g19698(.A0(new_n19890_), .A1(new_n19871_), .B0(new_n19877_), .Y(new_n19891_));
  AOI21X1  g19699(.A0(new_n19891_), .A1(new_n19872_), .B0(new_n399_), .Y(new_n19892_));
  AND2X1   g19700(.A(new_n19185_), .B(new_n19180_), .Y(new_n19893_));
  NOR3X1   g19701(.A(new_n19893_), .B(new_n19220_), .C(new_n19179_), .Y(new_n19894_));
  NOR3X1   g19702(.A(new_n19273_), .B(new_n19893_), .C(new_n19179_), .Y(new_n19895_));
  NOR2X1   g19703(.A(new_n19895_), .B(new_n19184_), .Y(new_n19896_));
  AOI21X1  g19704(.A0(new_n19894_), .A1(\asqrt[9] ), .B0(new_n19896_), .Y(new_n19897_));
  INVX1    g19705(.A(new_n19897_), .Y(new_n19898_));
  NAND3X1  g19706(.A(new_n19891_), .B(new_n19872_), .C(new_n399_), .Y(new_n19899_));
  AOI21X1  g19707(.A0(new_n19899_), .A1(new_n19898_), .B0(new_n19892_), .Y(new_n19900_));
  OR2X1    g19708(.A(new_n19900_), .B(new_n328_), .Y(new_n19901_));
  OR2X1    g19709(.A(new_n19889_), .B(new_n582_), .Y(new_n19902_));
  NOR2X1   g19710(.A(new_n19861_), .B(new_n19860_), .Y(new_n19903_));
  NAND2X1  g19711(.A(new_n19855_), .B(new_n582_), .Y(new_n19904_));
  INVX1    g19712(.A(new_n19870_), .Y(new_n19905_));
  OAI21X1  g19713(.A0(new_n19904_), .A1(new_n19903_), .B0(new_n19905_), .Y(new_n19906_));
  AOI21X1  g19714(.A0(new_n19906_), .A1(new_n19902_), .B0(new_n481_), .Y(new_n19907_));
  AOI21X1  g19715(.A0(new_n19862_), .A1(\asqrt[56] ), .B0(\asqrt[57] ), .Y(new_n19908_));
  AOI21X1  g19716(.A0(new_n19908_), .A1(new_n19906_), .B0(new_n19876_), .Y(new_n19909_));
  NOR3X1   g19717(.A(new_n19909_), .B(new_n19907_), .C(\asqrt[58] ), .Y(new_n19910_));
  NOR2X1   g19718(.A(new_n19910_), .B(new_n19897_), .Y(new_n19911_));
  AND2X1   g19719(.A(new_n19224_), .B(new_n19222_), .Y(new_n19912_));
  NOR3X1   g19720(.A(new_n19912_), .B(new_n19193_), .C(new_n19223_), .Y(new_n19913_));
  NOR3X1   g19721(.A(new_n19273_), .B(new_n19912_), .C(new_n19223_), .Y(new_n19914_));
  NOR2X1   g19722(.A(new_n19914_), .B(new_n19192_), .Y(new_n19915_));
  AOI21X1  g19723(.A0(new_n19913_), .A1(\asqrt[9] ), .B0(new_n19915_), .Y(new_n19916_));
  INVX1    g19724(.A(new_n19916_), .Y(new_n19917_));
  OAI21X1  g19725(.A0(new_n19909_), .A1(new_n19907_), .B0(\asqrt[58] ), .Y(new_n19918_));
  NAND2X1  g19726(.A(new_n19918_), .B(new_n328_), .Y(new_n19919_));
  OAI21X1  g19727(.A0(new_n19919_), .A1(new_n19911_), .B0(new_n19917_), .Y(new_n19920_));
  AOI21X1  g19728(.A0(new_n19920_), .A1(new_n19901_), .B0(new_n292_), .Y(new_n19921_));
  OR4X1    g19729(.A(new_n19273_), .B(new_n19226_), .C(new_n19214_), .D(new_n19208_), .Y(new_n19922_));
  OR2X1    g19730(.A(new_n19226_), .B(new_n19208_), .Y(new_n19923_));
  OAI21X1  g19731(.A0(new_n19923_), .A1(new_n19273_), .B0(new_n19214_), .Y(new_n19924_));
  AND2X1   g19732(.A(new_n19924_), .B(new_n19922_), .Y(new_n19925_));
  OAI21X1  g19733(.A0(new_n19910_), .A1(new_n19897_), .B0(new_n19918_), .Y(new_n19926_));
  AOI21X1  g19734(.A0(new_n19926_), .A1(\asqrt[59] ), .B0(\asqrt[60] ), .Y(new_n19927_));
  AOI21X1  g19735(.A0(new_n19927_), .A1(new_n19920_), .B0(new_n19925_), .Y(new_n19928_));
  OAI21X1  g19736(.A0(new_n19928_), .A1(new_n19921_), .B0(\asqrt[61] ), .Y(new_n19929_));
  AOI21X1  g19737(.A0(new_n19286_), .A1(new_n19285_), .B0(new_n19232_), .Y(new_n19930_));
  AND2X1   g19738(.A(new_n19930_), .B(new_n19217_), .Y(new_n19931_));
  AOI22X1  g19739(.A0(new_n19286_), .A1(new_n19285_), .B0(new_n19242_), .B1(\asqrt[60] ), .Y(new_n19932_));
  AOI21X1  g19740(.A0(new_n19932_), .A1(\asqrt[9] ), .B0(new_n19231_), .Y(new_n19933_));
  AOI21X1  g19741(.A0(new_n19931_), .A1(\asqrt[9] ), .B0(new_n19933_), .Y(new_n19934_));
  NOR3X1   g19742(.A(new_n19928_), .B(new_n19921_), .C(\asqrt[61] ), .Y(new_n19935_));
  OAI21X1  g19743(.A0(new_n19935_), .A1(new_n19934_), .B0(new_n19929_), .Y(new_n19936_));
  AND2X1   g19744(.A(new_n19936_), .B(\asqrt[62] ), .Y(new_n19937_));
  OR2X1    g19745(.A(new_n19935_), .B(new_n19934_), .Y(new_n19938_));
  AND2X1   g19746(.A(new_n19243_), .B(new_n19235_), .Y(new_n19939_));
  NOR3X1   g19747(.A(new_n19939_), .B(new_n19289_), .C(new_n19236_), .Y(new_n19940_));
  NOR3X1   g19748(.A(new_n19273_), .B(new_n19939_), .C(new_n19236_), .Y(new_n19941_));
  NOR2X1   g19749(.A(new_n19941_), .B(new_n19241_), .Y(new_n19942_));
  AOI21X1  g19750(.A0(new_n19940_), .A1(\asqrt[9] ), .B0(new_n19942_), .Y(new_n19943_));
  AND2X1   g19751(.A(new_n19929_), .B(new_n199_), .Y(new_n19944_));
  AOI21X1  g19752(.A0(new_n19944_), .A1(new_n19938_), .B0(new_n19943_), .Y(new_n19945_));
  NAND3X1  g19753(.A(new_n19294_), .B(new_n19250_), .C(new_n19245_), .Y(new_n19946_));
  AOI21X1  g19754(.A0(new_n19301_), .A1(new_n19297_), .B0(new_n19946_), .Y(new_n19947_));
  NAND3X1  g19755(.A(\asqrt[9] ), .B(new_n19294_), .C(new_n19245_), .Y(new_n19948_));
  AOI21X1  g19756(.A0(new_n19948_), .A1(new_n19293_), .B0(new_n19947_), .Y(new_n19949_));
  INVX1    g19757(.A(new_n19949_), .Y(new_n19950_));
  NOR3X1   g19758(.A(new_n19273_), .B(new_n19256_), .C(new_n19295_), .Y(new_n19951_));
  AOI21X1  g19759(.A0(new_n19299_), .A1(new_n19298_), .B0(new_n19951_), .Y(new_n19952_));
  AND2X1   g19760(.A(new_n19952_), .B(new_n19950_), .Y(new_n19953_));
  OAI21X1  g19761(.A0(new_n19945_), .A1(new_n19937_), .B0(new_n19953_), .Y(new_n19954_));
  AND2X1   g19762(.A(new_n19926_), .B(\asqrt[59] ), .Y(new_n19955_));
  OR2X1    g19763(.A(new_n19910_), .B(new_n19897_), .Y(new_n19956_));
  AND2X1   g19764(.A(new_n19918_), .B(new_n328_), .Y(new_n19957_));
  AOI21X1  g19765(.A0(new_n19957_), .A1(new_n19956_), .B0(new_n19916_), .Y(new_n19958_));
  OAI21X1  g19766(.A0(new_n19958_), .A1(new_n19955_), .B0(\asqrt[60] ), .Y(new_n19959_));
  INVX1    g19767(.A(new_n19925_), .Y(new_n19960_));
  OAI21X1  g19768(.A0(new_n19900_), .A1(new_n328_), .B0(new_n292_), .Y(new_n19961_));
  OAI21X1  g19769(.A0(new_n19961_), .A1(new_n19958_), .B0(new_n19960_), .Y(new_n19962_));
  AOI21X1  g19770(.A0(new_n19962_), .A1(new_n19959_), .B0(new_n217_), .Y(new_n19963_));
  INVX1    g19771(.A(new_n19934_), .Y(new_n19964_));
  NAND3X1  g19772(.A(new_n19962_), .B(new_n19959_), .C(new_n217_), .Y(new_n19965_));
  AOI21X1  g19773(.A0(new_n19965_), .A1(new_n19964_), .B0(new_n19963_), .Y(new_n19966_));
  OAI21X1  g19774(.A0(new_n19966_), .A1(new_n199_), .B0(new_n19949_), .Y(new_n19967_));
  AOI21X1  g19775(.A0(new_n19301_), .A1(new_n19297_), .B0(new_n19256_), .Y(new_n19968_));
  AOI21X1  g19776(.A0(new_n19257_), .A1(new_n19252_), .B0(new_n193_), .Y(new_n19969_));
  OAI21X1  g19777(.A0(new_n19968_), .A1(new_n19252_), .B0(new_n19969_), .Y(new_n19970_));
  OR2X1    g19778(.A(new_n19263_), .B(new_n19262_), .Y(new_n19971_));
  NOR4X1   g19779(.A(new_n19269_), .B(new_n19309_), .C(new_n19255_), .D(new_n19253_), .Y(new_n19972_));
  NAND3X1  g19780(.A(new_n19972_), .B(new_n19971_), .C(new_n19297_), .Y(new_n19973_));
  AND2X1   g19781(.A(new_n19973_), .B(new_n19970_), .Y(new_n19974_));
  OAI21X1  g19782(.A0(new_n19967_), .A1(new_n19945_), .B0(new_n19974_), .Y(new_n19975_));
  AOI21X1  g19783(.A0(new_n19954_), .A1(new_n193_), .B0(new_n19975_), .Y(new_n19976_));
  OR2X1    g19784(.A(new_n19966_), .B(new_n199_), .Y(new_n19977_));
  NOR2X1   g19785(.A(new_n19935_), .B(new_n19934_), .Y(new_n19978_));
  INVX1    g19786(.A(new_n19943_), .Y(new_n19979_));
  NAND2X1  g19787(.A(new_n19929_), .B(new_n199_), .Y(new_n19980_));
  OAI21X1  g19788(.A0(new_n19980_), .A1(new_n19978_), .B0(new_n19979_), .Y(new_n19981_));
  INVX1    g19789(.A(new_n19953_), .Y(new_n19982_));
  AOI21X1  g19790(.A0(new_n19981_), .A1(new_n19977_), .B0(new_n19982_), .Y(new_n19983_));
  AOI21X1  g19791(.A0(new_n19936_), .A1(\asqrt[62] ), .B0(new_n19950_), .Y(new_n19984_));
  INVX1    g19792(.A(new_n19974_), .Y(new_n19985_));
  AOI21X1  g19793(.A0(new_n19984_), .A1(new_n19981_), .B0(new_n19985_), .Y(new_n19986_));
  OAI21X1  g19794(.A0(new_n19983_), .A1(\asqrt[63] ), .B0(new_n19986_), .Y(\asqrt[8] ));
  NOR2X1   g19795(.A(\a[15] ), .B(\a[14] ), .Y(new_n19988_));
  MX2X1    g19796(.A(new_n19988_), .B(\asqrt[8] ), .S0(\a[16] ), .Y(new_n19989_));
  AND2X1   g19797(.A(new_n19989_), .B(\asqrt[9] ), .Y(new_n19990_));
  NOR3X1   g19798(.A(\a[16] ), .B(\a[15] ), .C(\a[14] ), .Y(new_n19991_));
  NOR3X1   g19799(.A(new_n19991_), .B(new_n19269_), .C(new_n19309_), .Y(new_n19992_));
  NAND3X1  g19800(.A(new_n19992_), .B(new_n19971_), .C(new_n19297_), .Y(new_n19993_));
  AOI21X1  g19801(.A0(\asqrt[8] ), .A1(\a[16] ), .B0(new_n19993_), .Y(new_n19994_));
  INVX1    g19802(.A(\a[16] ), .Y(new_n19995_));
  INVX1    g19803(.A(\a[17] ), .Y(new_n19996_));
  AOI21X1  g19804(.A0(\asqrt[8] ), .A1(new_n19995_), .B0(new_n19996_), .Y(new_n19997_));
  NOR2X1   g19805(.A(\a[17] ), .B(\a[16] ), .Y(new_n19998_));
  AND2X1   g19806(.A(\asqrt[8] ), .B(new_n19998_), .Y(new_n19999_));
  NOR3X1   g19807(.A(new_n19999_), .B(new_n19997_), .C(new_n19994_), .Y(new_n20000_));
  OAI21X1  g19808(.A0(new_n20000_), .A1(new_n19990_), .B0(\asqrt[10] ), .Y(new_n20001_));
  INVX1    g19809(.A(new_n19988_), .Y(new_n20002_));
  MX2X1    g19810(.A(new_n20002_), .B(new_n19976_), .S0(\a[16] ), .Y(new_n20003_));
  OAI21X1  g19811(.A0(new_n20003_), .A1(new_n19273_), .B0(new_n18591_), .Y(new_n20004_));
  NAND3X1  g19812(.A(new_n19973_), .B(new_n19970_), .C(\asqrt[9] ), .Y(new_n20005_));
  INVX1    g19813(.A(new_n20005_), .Y(new_n20006_));
  OAI21X1  g19814(.A0(new_n19967_), .A1(new_n19945_), .B0(new_n20006_), .Y(new_n20007_));
  AOI21X1  g19815(.A0(new_n19954_), .A1(new_n193_), .B0(new_n20007_), .Y(new_n20008_));
  AOI21X1  g19816(.A0(\asqrt[8] ), .A1(new_n19998_), .B0(new_n20008_), .Y(new_n20009_));
  OR2X1    g19817(.A(new_n20008_), .B(\a[18] ), .Y(new_n20010_));
  OAI22X1  g19818(.A0(new_n20010_), .A1(new_n19999_), .B0(new_n20009_), .B1(new_n19281_), .Y(new_n20011_));
  OAI21X1  g19819(.A0(new_n20004_), .A1(new_n20000_), .B0(new_n20011_), .Y(new_n20012_));
  AOI21X1  g19820(.A0(new_n20012_), .A1(new_n20001_), .B0(new_n17927_), .Y(new_n20013_));
  NOR4X1   g19821(.A(new_n19976_), .B(new_n19303_), .C(new_n19327_), .D(new_n19277_), .Y(new_n20014_));
  AND2X1   g19822(.A(new_n19280_), .B(new_n19326_), .Y(new_n20015_));
  AOI21X1  g19823(.A0(new_n20015_), .A1(\asqrt[8] ), .B0(new_n19330_), .Y(new_n20016_));
  NOR2X1   g19824(.A(new_n20016_), .B(new_n20014_), .Y(new_n20017_));
  INVX1    g19825(.A(new_n20017_), .Y(new_n20018_));
  NAND3X1  g19826(.A(new_n20012_), .B(new_n20001_), .C(new_n17927_), .Y(new_n20019_));
  AOI21X1  g19827(.A0(new_n20019_), .A1(new_n20018_), .B0(new_n20013_), .Y(new_n20020_));
  OR2X1    g19828(.A(new_n20020_), .B(new_n17262_), .Y(new_n20021_));
  AND2X1   g19829(.A(new_n20019_), .B(new_n20018_), .Y(new_n20022_));
  AOI21X1  g19830(.A0(new_n19360_), .A1(new_n19359_), .B0(new_n19316_), .Y(new_n20023_));
  NAND3X1  g19831(.A(new_n20023_), .B(\asqrt[8] ), .C(new_n19305_), .Y(new_n20024_));
  OAI22X1  g19832(.A0(new_n19307_), .A1(new_n19306_), .B0(new_n19304_), .B1(new_n17927_), .Y(new_n20025_));
  OAI21X1  g19833(.A0(new_n20025_), .A1(new_n19976_), .B0(new_n19316_), .Y(new_n20026_));
  AND2X1   g19834(.A(new_n20026_), .B(new_n20024_), .Y(new_n20027_));
  INVX1    g19835(.A(new_n20027_), .Y(new_n20028_));
  OR2X1    g19836(.A(new_n20013_), .B(\asqrt[12] ), .Y(new_n20029_));
  OAI21X1  g19837(.A0(new_n20029_), .A1(new_n20022_), .B0(new_n20028_), .Y(new_n20030_));
  AOI21X1  g19838(.A0(new_n20030_), .A1(new_n20021_), .B0(new_n16617_), .Y(new_n20031_));
  AND2X1   g19839(.A(new_n19332_), .B(new_n19317_), .Y(new_n20032_));
  INVX1    g19840(.A(new_n20032_), .Y(new_n20033_));
  NAND3X1  g19841(.A(new_n20033_), .B(new_n19324_), .C(new_n19363_), .Y(new_n20034_));
  NOR3X1   g19842(.A(new_n19976_), .B(new_n20032_), .C(new_n19318_), .Y(new_n20035_));
  OAI22X1  g19843(.A0(new_n20035_), .A1(new_n19324_), .B0(new_n20034_), .B1(new_n19976_), .Y(new_n20036_));
  INVX1    g19844(.A(new_n20036_), .Y(new_n20037_));
  OR2X1    g19845(.A(new_n20003_), .B(new_n19273_), .Y(new_n20038_));
  INVX1    g19846(.A(new_n19993_), .Y(new_n20039_));
  OAI21X1  g19847(.A0(new_n19976_), .A1(new_n19995_), .B0(new_n20039_), .Y(new_n20040_));
  OAI21X1  g19848(.A0(new_n19976_), .A1(\a[16] ), .B0(\a[17] ), .Y(new_n20041_));
  INVX1    g19849(.A(new_n19998_), .Y(new_n20042_));
  OR2X1    g19850(.A(new_n19976_), .B(new_n20042_), .Y(new_n20043_));
  NAND3X1  g19851(.A(new_n20043_), .B(new_n20041_), .C(new_n20040_), .Y(new_n20044_));
  AOI21X1  g19852(.A0(new_n20044_), .A1(new_n20038_), .B0(new_n18591_), .Y(new_n20045_));
  AOI21X1  g19853(.A0(new_n19989_), .A1(\asqrt[9] ), .B0(\asqrt[10] ), .Y(new_n20046_));
  OR2X1    g19854(.A(new_n20009_), .B(new_n19281_), .Y(new_n20047_));
  OR2X1    g19855(.A(new_n20010_), .B(new_n19999_), .Y(new_n20048_));
  AOI22X1  g19856(.A0(new_n20048_), .A1(new_n20047_), .B0(new_n20046_), .B1(new_n20044_), .Y(new_n20049_));
  OAI21X1  g19857(.A0(new_n20049_), .A1(new_n20045_), .B0(\asqrt[11] ), .Y(new_n20050_));
  NOR3X1   g19858(.A(new_n20049_), .B(new_n20045_), .C(\asqrt[11] ), .Y(new_n20051_));
  OAI21X1  g19859(.A0(new_n20051_), .A1(new_n20017_), .B0(new_n20050_), .Y(new_n20052_));
  AOI21X1  g19860(.A0(new_n20052_), .A1(\asqrt[12] ), .B0(\asqrt[13] ), .Y(new_n20053_));
  AOI21X1  g19861(.A0(new_n20053_), .A1(new_n20030_), .B0(new_n20037_), .Y(new_n20054_));
  OAI21X1  g19862(.A0(new_n20054_), .A1(new_n20031_), .B0(\asqrt[14] ), .Y(new_n20055_));
  OR4X1    g19863(.A(new_n19976_), .B(new_n19342_), .C(new_n19368_), .D(new_n19367_), .Y(new_n20056_));
  NAND2X1  g19864(.A(new_n19369_), .B(new_n19334_), .Y(new_n20057_));
  OAI21X1  g19865(.A0(new_n20057_), .A1(new_n19976_), .B0(new_n19368_), .Y(new_n20058_));
  AND2X1   g19866(.A(new_n20058_), .B(new_n20056_), .Y(new_n20059_));
  NOR3X1   g19867(.A(new_n20054_), .B(new_n20031_), .C(\asqrt[14] ), .Y(new_n20060_));
  OAI21X1  g19868(.A0(new_n20060_), .A1(new_n20059_), .B0(new_n20055_), .Y(new_n20061_));
  AND2X1   g19869(.A(new_n20061_), .B(\asqrt[15] ), .Y(new_n20062_));
  INVX1    g19870(.A(new_n20059_), .Y(new_n20063_));
  AND2X1   g19871(.A(new_n20052_), .B(\asqrt[12] ), .Y(new_n20064_));
  NAND2X1  g19872(.A(new_n20019_), .B(new_n20018_), .Y(new_n20065_));
  NOR2X1   g19873(.A(new_n20013_), .B(\asqrt[12] ), .Y(new_n20066_));
  AOI21X1  g19874(.A0(new_n20066_), .A1(new_n20065_), .B0(new_n20027_), .Y(new_n20067_));
  OAI21X1  g19875(.A0(new_n20067_), .A1(new_n20064_), .B0(\asqrt[13] ), .Y(new_n20068_));
  OAI21X1  g19876(.A0(new_n20020_), .A1(new_n17262_), .B0(new_n16617_), .Y(new_n20069_));
  OAI21X1  g19877(.A0(new_n20069_), .A1(new_n20067_), .B0(new_n20036_), .Y(new_n20070_));
  NAND3X1  g19878(.A(new_n20070_), .B(new_n20068_), .C(new_n15990_), .Y(new_n20071_));
  NAND2X1  g19879(.A(new_n20071_), .B(new_n20063_), .Y(new_n20072_));
  AND2X1   g19880(.A(new_n19352_), .B(new_n19345_), .Y(new_n20073_));
  NOR4X1   g19881(.A(new_n19976_), .B(new_n20073_), .C(new_n19392_), .D(new_n19344_), .Y(new_n20074_));
  AOI22X1  g19882(.A0(new_n19352_), .A1(new_n19345_), .B0(new_n19343_), .B1(\asqrt[14] ), .Y(new_n20075_));
  AOI21X1  g19883(.A0(new_n20075_), .A1(\asqrt[8] ), .B0(new_n19351_), .Y(new_n20076_));
  NOR2X1   g19884(.A(new_n20076_), .B(new_n20074_), .Y(new_n20077_));
  AOI21X1  g19885(.A0(new_n20070_), .A1(new_n20068_), .B0(new_n15990_), .Y(new_n20078_));
  NOR2X1   g19886(.A(new_n20078_), .B(\asqrt[15] ), .Y(new_n20079_));
  AOI21X1  g19887(.A0(new_n20079_), .A1(new_n20072_), .B0(new_n20077_), .Y(new_n20080_));
  OAI21X1  g19888(.A0(new_n20080_), .A1(new_n20062_), .B0(\asqrt[16] ), .Y(new_n20081_));
  AND2X1   g19889(.A(new_n19397_), .B(new_n19394_), .Y(new_n20082_));
  OR4X1    g19890(.A(new_n19976_), .B(new_n20082_), .C(new_n19357_), .D(new_n19395_), .Y(new_n20083_));
  OR2X1    g19891(.A(new_n20082_), .B(new_n19395_), .Y(new_n20084_));
  OAI21X1  g19892(.A0(new_n20084_), .A1(new_n19976_), .B0(new_n19357_), .Y(new_n20085_));
  AND2X1   g19893(.A(new_n20085_), .B(new_n20083_), .Y(new_n20086_));
  INVX1    g19894(.A(new_n20086_), .Y(new_n20087_));
  AOI21X1  g19895(.A0(new_n20071_), .A1(new_n20063_), .B0(new_n20078_), .Y(new_n20088_));
  OAI21X1  g19896(.A0(new_n20088_), .A1(new_n15362_), .B0(new_n14754_), .Y(new_n20089_));
  OAI21X1  g19897(.A0(new_n20089_), .A1(new_n20080_), .B0(new_n20087_), .Y(new_n20090_));
  AOI21X1  g19898(.A0(new_n20090_), .A1(new_n20081_), .B0(new_n14165_), .Y(new_n20091_));
  OR4X1    g19899(.A(new_n19976_), .B(new_n19407_), .C(new_n19379_), .D(new_n19373_), .Y(new_n20092_));
  NAND2X1  g19900(.A(new_n19380_), .B(new_n19399_), .Y(new_n20093_));
  OAI21X1  g19901(.A0(new_n20093_), .A1(new_n19976_), .B0(new_n19379_), .Y(new_n20094_));
  AND2X1   g19902(.A(new_n20094_), .B(new_n20092_), .Y(new_n20095_));
  INVX1    g19903(.A(new_n20095_), .Y(new_n20096_));
  NAND3X1  g19904(.A(new_n20090_), .B(new_n20081_), .C(new_n14165_), .Y(new_n20097_));
  AOI21X1  g19905(.A0(new_n20097_), .A1(new_n20096_), .B0(new_n20091_), .Y(new_n20098_));
  OR2X1    g19906(.A(new_n20098_), .B(new_n13571_), .Y(new_n20099_));
  AND2X1   g19907(.A(new_n20097_), .B(new_n20096_), .Y(new_n20100_));
  OAI21X1  g19908(.A0(new_n19400_), .A1(new_n19383_), .B0(new_n19388_), .Y(new_n20101_));
  NOR3X1   g19909(.A(new_n20101_), .B(new_n19976_), .C(new_n19421_), .Y(new_n20102_));
  AOI22X1  g19910(.A0(new_n19423_), .A1(new_n19422_), .B0(new_n19408_), .B1(\asqrt[17] ), .Y(new_n20103_));
  AOI21X1  g19911(.A0(new_n20103_), .A1(\asqrt[8] ), .B0(new_n19388_), .Y(new_n20104_));
  NOR2X1   g19912(.A(new_n20104_), .B(new_n20102_), .Y(new_n20105_));
  INVX1    g19913(.A(new_n20105_), .Y(new_n20106_));
  OR2X1    g19914(.A(new_n20091_), .B(\asqrt[18] ), .Y(new_n20107_));
  OAI21X1  g19915(.A0(new_n20107_), .A1(new_n20100_), .B0(new_n20106_), .Y(new_n20108_));
  AOI21X1  g19916(.A0(new_n20108_), .A1(new_n20099_), .B0(new_n13000_), .Y(new_n20109_));
  AND2X1   g19917(.A(new_n19409_), .B(new_n19401_), .Y(new_n20110_));
  OR4X1    g19918(.A(new_n19976_), .B(new_n20110_), .C(new_n19426_), .D(new_n19402_), .Y(new_n20111_));
  OR2X1    g19919(.A(new_n20110_), .B(new_n19402_), .Y(new_n20112_));
  OAI21X1  g19920(.A0(new_n20112_), .A1(new_n19976_), .B0(new_n19426_), .Y(new_n20113_));
  AND2X1   g19921(.A(new_n20113_), .B(new_n20111_), .Y(new_n20114_));
  OR2X1    g19922(.A(new_n20088_), .B(new_n15362_), .Y(new_n20115_));
  AND2X1   g19923(.A(new_n20071_), .B(new_n20063_), .Y(new_n20116_));
  INVX1    g19924(.A(new_n20077_), .Y(new_n20117_));
  OR2X1    g19925(.A(new_n20078_), .B(\asqrt[15] ), .Y(new_n20118_));
  OAI21X1  g19926(.A0(new_n20118_), .A1(new_n20116_), .B0(new_n20117_), .Y(new_n20119_));
  AOI21X1  g19927(.A0(new_n20119_), .A1(new_n20115_), .B0(new_n14754_), .Y(new_n20120_));
  AOI21X1  g19928(.A0(new_n20061_), .A1(\asqrt[15] ), .B0(\asqrt[16] ), .Y(new_n20121_));
  AOI21X1  g19929(.A0(new_n20121_), .A1(new_n20119_), .B0(new_n20086_), .Y(new_n20122_));
  OAI21X1  g19930(.A0(new_n20122_), .A1(new_n20120_), .B0(\asqrt[17] ), .Y(new_n20123_));
  NOR3X1   g19931(.A(new_n20122_), .B(new_n20120_), .C(\asqrt[17] ), .Y(new_n20124_));
  OAI21X1  g19932(.A0(new_n20124_), .A1(new_n20095_), .B0(new_n20123_), .Y(new_n20125_));
  AOI21X1  g19933(.A0(new_n20125_), .A1(\asqrt[18] ), .B0(\asqrt[19] ), .Y(new_n20126_));
  AOI21X1  g19934(.A0(new_n20126_), .A1(new_n20108_), .B0(new_n20114_), .Y(new_n20127_));
  OAI21X1  g19935(.A0(new_n20127_), .A1(new_n20109_), .B0(\asqrt[20] ), .Y(new_n20128_));
  OR4X1    g19936(.A(new_n19976_), .B(new_n19417_), .C(new_n19420_), .D(new_n19444_), .Y(new_n20129_));
  NAND2X1  g19937(.A(new_n19429_), .B(new_n19411_), .Y(new_n20130_));
  OAI21X1  g19938(.A0(new_n20130_), .A1(new_n19976_), .B0(new_n19420_), .Y(new_n20131_));
  AND2X1   g19939(.A(new_n20131_), .B(new_n20129_), .Y(new_n20132_));
  NOR3X1   g19940(.A(new_n20127_), .B(new_n20109_), .C(\asqrt[20] ), .Y(new_n20133_));
  OAI21X1  g19941(.A0(new_n20133_), .A1(new_n20132_), .B0(new_n20128_), .Y(new_n20134_));
  AND2X1   g19942(.A(new_n20134_), .B(\asqrt[21] ), .Y(new_n20135_));
  INVX1    g19943(.A(new_n20132_), .Y(new_n20136_));
  AND2X1   g19944(.A(new_n20125_), .B(\asqrt[18] ), .Y(new_n20137_));
  NAND2X1  g19945(.A(new_n20097_), .B(new_n20096_), .Y(new_n20138_));
  NOR2X1   g19946(.A(new_n20091_), .B(\asqrt[18] ), .Y(new_n20139_));
  AOI21X1  g19947(.A0(new_n20139_), .A1(new_n20138_), .B0(new_n20105_), .Y(new_n20140_));
  OAI21X1  g19948(.A0(new_n20140_), .A1(new_n20137_), .B0(\asqrt[19] ), .Y(new_n20141_));
  INVX1    g19949(.A(new_n20114_), .Y(new_n20142_));
  OAI21X1  g19950(.A0(new_n20098_), .A1(new_n13571_), .B0(new_n13000_), .Y(new_n20143_));
  OAI21X1  g19951(.A0(new_n20143_), .A1(new_n20140_), .B0(new_n20142_), .Y(new_n20144_));
  NAND3X1  g19952(.A(new_n20144_), .B(new_n20141_), .C(new_n12447_), .Y(new_n20145_));
  NAND2X1  g19953(.A(new_n20145_), .B(new_n20136_), .Y(new_n20146_));
  AND2X1   g19954(.A(new_n19436_), .B(new_n19430_), .Y(new_n20147_));
  NOR4X1   g19955(.A(new_n19976_), .B(new_n20147_), .C(new_n19467_), .D(new_n19419_), .Y(new_n20148_));
  AOI22X1  g19956(.A0(new_n19436_), .A1(new_n19430_), .B0(new_n19418_), .B1(\asqrt[20] ), .Y(new_n20149_));
  AOI21X1  g19957(.A0(new_n20149_), .A1(\asqrt[8] ), .B0(new_n19435_), .Y(new_n20150_));
  NOR2X1   g19958(.A(new_n20150_), .B(new_n20148_), .Y(new_n20151_));
  AOI21X1  g19959(.A0(new_n20144_), .A1(new_n20141_), .B0(new_n12447_), .Y(new_n20152_));
  NOR2X1   g19960(.A(new_n20152_), .B(\asqrt[21] ), .Y(new_n20153_));
  AOI21X1  g19961(.A0(new_n20153_), .A1(new_n20146_), .B0(new_n20151_), .Y(new_n20154_));
  OAI21X1  g19962(.A0(new_n20154_), .A1(new_n20135_), .B0(\asqrt[22] ), .Y(new_n20155_));
  AND2X1   g19963(.A(new_n19471_), .B(new_n19469_), .Y(new_n20156_));
  OR4X1    g19964(.A(new_n19976_), .B(new_n20156_), .C(new_n19443_), .D(new_n19470_), .Y(new_n20157_));
  OR2X1    g19965(.A(new_n20156_), .B(new_n19470_), .Y(new_n20158_));
  OAI21X1  g19966(.A0(new_n20158_), .A1(new_n19976_), .B0(new_n19443_), .Y(new_n20159_));
  AND2X1   g19967(.A(new_n20159_), .B(new_n20157_), .Y(new_n20160_));
  INVX1    g19968(.A(new_n20160_), .Y(new_n20161_));
  AOI21X1  g19969(.A0(new_n20145_), .A1(new_n20136_), .B0(new_n20152_), .Y(new_n20162_));
  OAI21X1  g19970(.A0(new_n20162_), .A1(new_n11896_), .B0(new_n11362_), .Y(new_n20163_));
  OAI21X1  g19971(.A0(new_n20163_), .A1(new_n20154_), .B0(new_n20161_), .Y(new_n20164_));
  AOI21X1  g19972(.A0(new_n20164_), .A1(new_n20155_), .B0(new_n10849_), .Y(new_n20165_));
  OR4X1    g19973(.A(new_n19976_), .B(new_n19481_), .C(new_n19454_), .D(new_n19448_), .Y(new_n20166_));
  NAND2X1  g19974(.A(new_n19455_), .B(new_n19473_), .Y(new_n20167_));
  OAI21X1  g19975(.A0(new_n20167_), .A1(new_n19976_), .B0(new_n19454_), .Y(new_n20168_));
  AND2X1   g19976(.A(new_n20168_), .B(new_n20166_), .Y(new_n20169_));
  INVX1    g19977(.A(new_n20169_), .Y(new_n20170_));
  NAND3X1  g19978(.A(new_n20164_), .B(new_n20155_), .C(new_n10849_), .Y(new_n20171_));
  AOI21X1  g19979(.A0(new_n20171_), .A1(new_n20170_), .B0(new_n20165_), .Y(new_n20172_));
  OR2X1    g19980(.A(new_n20172_), .B(new_n10332_), .Y(new_n20173_));
  AND2X1   g19981(.A(new_n20171_), .B(new_n20170_), .Y(new_n20174_));
  OAI21X1  g19982(.A0(new_n19474_), .A1(new_n19458_), .B0(new_n19463_), .Y(new_n20175_));
  NOR3X1   g19983(.A(new_n20175_), .B(new_n19976_), .C(new_n19495_), .Y(new_n20176_));
  AOI22X1  g19984(.A0(new_n19497_), .A1(new_n19496_), .B0(new_n19482_), .B1(\asqrt[23] ), .Y(new_n20177_));
  AOI21X1  g19985(.A0(new_n20177_), .A1(\asqrt[8] ), .B0(new_n19463_), .Y(new_n20178_));
  NOR2X1   g19986(.A(new_n20178_), .B(new_n20176_), .Y(new_n20179_));
  INVX1    g19987(.A(new_n20179_), .Y(new_n20180_));
  OR2X1    g19988(.A(new_n20165_), .B(\asqrt[24] ), .Y(new_n20181_));
  OAI21X1  g19989(.A0(new_n20181_), .A1(new_n20174_), .B0(new_n20180_), .Y(new_n20182_));
  AOI21X1  g19990(.A0(new_n20182_), .A1(new_n20173_), .B0(new_n9833_), .Y(new_n20183_));
  AND2X1   g19991(.A(new_n19483_), .B(new_n19475_), .Y(new_n20184_));
  OR4X1    g19992(.A(new_n19976_), .B(new_n20184_), .C(new_n19500_), .D(new_n19476_), .Y(new_n20185_));
  OR2X1    g19993(.A(new_n20184_), .B(new_n19476_), .Y(new_n20186_));
  OAI21X1  g19994(.A0(new_n20186_), .A1(new_n19976_), .B0(new_n19500_), .Y(new_n20187_));
  AND2X1   g19995(.A(new_n20187_), .B(new_n20185_), .Y(new_n20188_));
  OR2X1    g19996(.A(new_n20162_), .B(new_n11896_), .Y(new_n20189_));
  AND2X1   g19997(.A(new_n20145_), .B(new_n20136_), .Y(new_n20190_));
  INVX1    g19998(.A(new_n20151_), .Y(new_n20191_));
  OR2X1    g19999(.A(new_n20152_), .B(\asqrt[21] ), .Y(new_n20192_));
  OAI21X1  g20000(.A0(new_n20192_), .A1(new_n20190_), .B0(new_n20191_), .Y(new_n20193_));
  AOI21X1  g20001(.A0(new_n20193_), .A1(new_n20189_), .B0(new_n11362_), .Y(new_n20194_));
  AOI21X1  g20002(.A0(new_n20134_), .A1(\asqrt[21] ), .B0(\asqrt[22] ), .Y(new_n20195_));
  AOI21X1  g20003(.A0(new_n20195_), .A1(new_n20193_), .B0(new_n20160_), .Y(new_n20196_));
  OAI21X1  g20004(.A0(new_n20196_), .A1(new_n20194_), .B0(\asqrt[23] ), .Y(new_n20197_));
  NOR3X1   g20005(.A(new_n20196_), .B(new_n20194_), .C(\asqrt[23] ), .Y(new_n20198_));
  OAI21X1  g20006(.A0(new_n20198_), .A1(new_n20169_), .B0(new_n20197_), .Y(new_n20199_));
  AOI21X1  g20007(.A0(new_n20199_), .A1(\asqrt[24] ), .B0(\asqrt[25] ), .Y(new_n20200_));
  AOI21X1  g20008(.A0(new_n20200_), .A1(new_n20182_), .B0(new_n20188_), .Y(new_n20201_));
  OAI21X1  g20009(.A0(new_n20201_), .A1(new_n20183_), .B0(\asqrt[26] ), .Y(new_n20202_));
  OR4X1    g20010(.A(new_n19976_), .B(new_n19491_), .C(new_n19494_), .D(new_n19518_), .Y(new_n20203_));
  NAND2X1  g20011(.A(new_n19503_), .B(new_n19485_), .Y(new_n20204_));
  OAI21X1  g20012(.A0(new_n20204_), .A1(new_n19976_), .B0(new_n19494_), .Y(new_n20205_));
  AND2X1   g20013(.A(new_n20205_), .B(new_n20203_), .Y(new_n20206_));
  NOR3X1   g20014(.A(new_n20201_), .B(new_n20183_), .C(\asqrt[26] ), .Y(new_n20207_));
  OAI21X1  g20015(.A0(new_n20207_), .A1(new_n20206_), .B0(new_n20202_), .Y(new_n20208_));
  AND2X1   g20016(.A(new_n20208_), .B(\asqrt[27] ), .Y(new_n20209_));
  OR2X1    g20017(.A(new_n20207_), .B(new_n20206_), .Y(new_n20210_));
  AND2X1   g20018(.A(new_n19510_), .B(new_n19504_), .Y(new_n20211_));
  NOR4X1   g20019(.A(new_n19976_), .B(new_n20211_), .C(new_n19541_), .D(new_n19493_), .Y(new_n20212_));
  AOI22X1  g20020(.A0(new_n19510_), .A1(new_n19504_), .B0(new_n19492_), .B1(\asqrt[26] ), .Y(new_n20213_));
  AOI21X1  g20021(.A0(new_n20213_), .A1(\asqrt[8] ), .B0(new_n19509_), .Y(new_n20214_));
  NOR2X1   g20022(.A(new_n20214_), .B(new_n20212_), .Y(new_n20215_));
  AND2X1   g20023(.A(new_n20202_), .B(new_n8874_), .Y(new_n20216_));
  AOI21X1  g20024(.A0(new_n20216_), .A1(new_n20210_), .B0(new_n20215_), .Y(new_n20217_));
  OAI21X1  g20025(.A0(new_n20217_), .A1(new_n20209_), .B0(\asqrt[28] ), .Y(new_n20218_));
  AND2X1   g20026(.A(new_n19545_), .B(new_n19543_), .Y(new_n20219_));
  OR4X1    g20027(.A(new_n19976_), .B(new_n20219_), .C(new_n19517_), .D(new_n19544_), .Y(new_n20220_));
  OR2X1    g20028(.A(new_n20219_), .B(new_n19544_), .Y(new_n20221_));
  OAI21X1  g20029(.A0(new_n20221_), .A1(new_n19976_), .B0(new_n19517_), .Y(new_n20222_));
  AND2X1   g20030(.A(new_n20222_), .B(new_n20220_), .Y(new_n20223_));
  INVX1    g20031(.A(new_n20223_), .Y(new_n20224_));
  AND2X1   g20032(.A(new_n20199_), .B(\asqrt[24] ), .Y(new_n20225_));
  NAND2X1  g20033(.A(new_n20171_), .B(new_n20170_), .Y(new_n20226_));
  NOR2X1   g20034(.A(new_n20165_), .B(\asqrt[24] ), .Y(new_n20227_));
  AOI21X1  g20035(.A0(new_n20227_), .A1(new_n20226_), .B0(new_n20179_), .Y(new_n20228_));
  OAI21X1  g20036(.A0(new_n20228_), .A1(new_n20225_), .B0(\asqrt[25] ), .Y(new_n20229_));
  INVX1    g20037(.A(new_n20188_), .Y(new_n20230_));
  OAI21X1  g20038(.A0(new_n20172_), .A1(new_n10332_), .B0(new_n9833_), .Y(new_n20231_));
  OAI21X1  g20039(.A0(new_n20231_), .A1(new_n20228_), .B0(new_n20230_), .Y(new_n20232_));
  AOI21X1  g20040(.A0(new_n20232_), .A1(new_n20229_), .B0(new_n9353_), .Y(new_n20233_));
  INVX1    g20041(.A(new_n20206_), .Y(new_n20234_));
  NAND3X1  g20042(.A(new_n20232_), .B(new_n20229_), .C(new_n9353_), .Y(new_n20235_));
  AOI21X1  g20043(.A0(new_n20235_), .A1(new_n20234_), .B0(new_n20233_), .Y(new_n20236_));
  OAI21X1  g20044(.A0(new_n20236_), .A1(new_n8874_), .B0(new_n8412_), .Y(new_n20237_));
  OAI21X1  g20045(.A0(new_n20237_), .A1(new_n20217_), .B0(new_n20224_), .Y(new_n20238_));
  AOI21X1  g20046(.A0(new_n20238_), .A1(new_n20218_), .B0(new_n7970_), .Y(new_n20239_));
  OR4X1    g20047(.A(new_n19976_), .B(new_n19555_), .C(new_n19528_), .D(new_n19522_), .Y(new_n20240_));
  NAND2X1  g20048(.A(new_n19529_), .B(new_n19547_), .Y(new_n20241_));
  OAI21X1  g20049(.A0(new_n20241_), .A1(new_n19976_), .B0(new_n19528_), .Y(new_n20242_));
  AND2X1   g20050(.A(new_n20242_), .B(new_n20240_), .Y(new_n20243_));
  INVX1    g20051(.A(new_n20243_), .Y(new_n20244_));
  NAND3X1  g20052(.A(new_n20238_), .B(new_n20218_), .C(new_n7970_), .Y(new_n20245_));
  AOI21X1  g20053(.A0(new_n20245_), .A1(new_n20244_), .B0(new_n20239_), .Y(new_n20246_));
  OR2X1    g20054(.A(new_n20246_), .B(new_n7527_), .Y(new_n20247_));
  OR2X1    g20055(.A(new_n20236_), .B(new_n8874_), .Y(new_n20248_));
  NOR2X1   g20056(.A(new_n20207_), .B(new_n20206_), .Y(new_n20249_));
  INVX1    g20057(.A(new_n20215_), .Y(new_n20250_));
  NAND2X1  g20058(.A(new_n20202_), .B(new_n8874_), .Y(new_n20251_));
  OAI21X1  g20059(.A0(new_n20251_), .A1(new_n20249_), .B0(new_n20250_), .Y(new_n20252_));
  AOI21X1  g20060(.A0(new_n20252_), .A1(new_n20248_), .B0(new_n8412_), .Y(new_n20253_));
  AOI21X1  g20061(.A0(new_n20208_), .A1(\asqrt[27] ), .B0(\asqrt[28] ), .Y(new_n20254_));
  AOI21X1  g20062(.A0(new_n20254_), .A1(new_n20252_), .B0(new_n20223_), .Y(new_n20255_));
  NOR3X1   g20063(.A(new_n20255_), .B(new_n20253_), .C(\asqrt[29] ), .Y(new_n20256_));
  NOR2X1   g20064(.A(new_n20256_), .B(new_n20243_), .Y(new_n20257_));
  OAI21X1  g20065(.A0(new_n19548_), .A1(new_n19532_), .B0(new_n19537_), .Y(new_n20258_));
  NOR3X1   g20066(.A(new_n20258_), .B(new_n19976_), .C(new_n19569_), .Y(new_n20259_));
  AOI22X1  g20067(.A0(new_n19571_), .A1(new_n19570_), .B0(new_n19556_), .B1(\asqrt[29] ), .Y(new_n20260_));
  AOI21X1  g20068(.A0(new_n20260_), .A1(\asqrt[8] ), .B0(new_n19537_), .Y(new_n20261_));
  NOR2X1   g20069(.A(new_n20261_), .B(new_n20259_), .Y(new_n20262_));
  INVX1    g20070(.A(new_n20262_), .Y(new_n20263_));
  OAI21X1  g20071(.A0(new_n20255_), .A1(new_n20253_), .B0(\asqrt[29] ), .Y(new_n20264_));
  NAND2X1  g20072(.A(new_n20264_), .B(new_n7527_), .Y(new_n20265_));
  OAI21X1  g20073(.A0(new_n20265_), .A1(new_n20257_), .B0(new_n20263_), .Y(new_n20266_));
  AOI21X1  g20074(.A0(new_n20266_), .A1(new_n20247_), .B0(new_n7103_), .Y(new_n20267_));
  AND2X1   g20075(.A(new_n19557_), .B(new_n19549_), .Y(new_n20268_));
  OR4X1    g20076(.A(new_n19976_), .B(new_n20268_), .C(new_n19574_), .D(new_n19550_), .Y(new_n20269_));
  OR2X1    g20077(.A(new_n20268_), .B(new_n19550_), .Y(new_n20270_));
  OAI21X1  g20078(.A0(new_n20270_), .A1(new_n19976_), .B0(new_n19574_), .Y(new_n20271_));
  AND2X1   g20079(.A(new_n20271_), .B(new_n20269_), .Y(new_n20272_));
  OAI21X1  g20080(.A0(new_n20256_), .A1(new_n20243_), .B0(new_n20264_), .Y(new_n20273_));
  AOI21X1  g20081(.A0(new_n20273_), .A1(\asqrt[30] ), .B0(\asqrt[31] ), .Y(new_n20274_));
  AOI21X1  g20082(.A0(new_n20274_), .A1(new_n20266_), .B0(new_n20272_), .Y(new_n20275_));
  OAI21X1  g20083(.A0(new_n20275_), .A1(new_n20267_), .B0(\asqrt[32] ), .Y(new_n20276_));
  OR4X1    g20084(.A(new_n19976_), .B(new_n19565_), .C(new_n19568_), .D(new_n19592_), .Y(new_n20277_));
  NAND2X1  g20085(.A(new_n19577_), .B(new_n19559_), .Y(new_n20278_));
  OAI21X1  g20086(.A0(new_n20278_), .A1(new_n19976_), .B0(new_n19568_), .Y(new_n20279_));
  AND2X1   g20087(.A(new_n20279_), .B(new_n20277_), .Y(new_n20280_));
  NOR3X1   g20088(.A(new_n20275_), .B(new_n20267_), .C(\asqrt[32] ), .Y(new_n20281_));
  OAI21X1  g20089(.A0(new_n20281_), .A1(new_n20280_), .B0(new_n20276_), .Y(new_n20282_));
  AND2X1   g20090(.A(new_n20282_), .B(\asqrt[33] ), .Y(new_n20283_));
  OR2X1    g20091(.A(new_n20281_), .B(new_n20280_), .Y(new_n20284_));
  AND2X1   g20092(.A(new_n19584_), .B(new_n19578_), .Y(new_n20285_));
  NOR4X1   g20093(.A(new_n19976_), .B(new_n20285_), .C(new_n19615_), .D(new_n19567_), .Y(new_n20286_));
  AOI22X1  g20094(.A0(new_n19584_), .A1(new_n19578_), .B0(new_n19566_), .B1(\asqrt[32] ), .Y(new_n20287_));
  AOI21X1  g20095(.A0(new_n20287_), .A1(\asqrt[8] ), .B0(new_n19583_), .Y(new_n20288_));
  NOR2X1   g20096(.A(new_n20288_), .B(new_n20286_), .Y(new_n20289_));
  AND2X1   g20097(.A(new_n20276_), .B(new_n6294_), .Y(new_n20290_));
  AOI21X1  g20098(.A0(new_n20290_), .A1(new_n20284_), .B0(new_n20289_), .Y(new_n20291_));
  OAI21X1  g20099(.A0(new_n20291_), .A1(new_n20283_), .B0(\asqrt[34] ), .Y(new_n20292_));
  AND2X1   g20100(.A(new_n19619_), .B(new_n19617_), .Y(new_n20293_));
  OR4X1    g20101(.A(new_n19976_), .B(new_n20293_), .C(new_n19591_), .D(new_n19618_), .Y(new_n20294_));
  OR2X1    g20102(.A(new_n20293_), .B(new_n19618_), .Y(new_n20295_));
  OAI21X1  g20103(.A0(new_n20295_), .A1(new_n19976_), .B0(new_n19591_), .Y(new_n20296_));
  AND2X1   g20104(.A(new_n20296_), .B(new_n20294_), .Y(new_n20297_));
  INVX1    g20105(.A(new_n20297_), .Y(new_n20298_));
  AND2X1   g20106(.A(new_n20273_), .B(\asqrt[30] ), .Y(new_n20299_));
  OR2X1    g20107(.A(new_n20256_), .B(new_n20243_), .Y(new_n20300_));
  AND2X1   g20108(.A(new_n20264_), .B(new_n7527_), .Y(new_n20301_));
  AOI21X1  g20109(.A0(new_n20301_), .A1(new_n20300_), .B0(new_n20262_), .Y(new_n20302_));
  OAI21X1  g20110(.A0(new_n20302_), .A1(new_n20299_), .B0(\asqrt[31] ), .Y(new_n20303_));
  INVX1    g20111(.A(new_n20272_), .Y(new_n20304_));
  OAI21X1  g20112(.A0(new_n20246_), .A1(new_n7527_), .B0(new_n7103_), .Y(new_n20305_));
  OAI21X1  g20113(.A0(new_n20305_), .A1(new_n20302_), .B0(new_n20304_), .Y(new_n20306_));
  AOI21X1  g20114(.A0(new_n20306_), .A1(new_n20303_), .B0(new_n6699_), .Y(new_n20307_));
  INVX1    g20115(.A(new_n20280_), .Y(new_n20308_));
  NAND3X1  g20116(.A(new_n20306_), .B(new_n20303_), .C(new_n6699_), .Y(new_n20309_));
  AOI21X1  g20117(.A0(new_n20309_), .A1(new_n20308_), .B0(new_n20307_), .Y(new_n20310_));
  OAI21X1  g20118(.A0(new_n20310_), .A1(new_n6294_), .B0(new_n5941_), .Y(new_n20311_));
  OAI21X1  g20119(.A0(new_n20311_), .A1(new_n20291_), .B0(new_n20298_), .Y(new_n20312_));
  AOI21X1  g20120(.A0(new_n20312_), .A1(new_n20292_), .B0(new_n5541_), .Y(new_n20313_));
  OR4X1    g20121(.A(new_n19976_), .B(new_n19629_), .C(new_n19602_), .D(new_n19596_), .Y(new_n20314_));
  OR2X1    g20122(.A(new_n19629_), .B(new_n19596_), .Y(new_n20315_));
  OAI21X1  g20123(.A0(new_n20315_), .A1(new_n19976_), .B0(new_n19602_), .Y(new_n20316_));
  AND2X1   g20124(.A(new_n20316_), .B(new_n20314_), .Y(new_n20317_));
  INVX1    g20125(.A(new_n20317_), .Y(new_n20318_));
  NAND3X1  g20126(.A(new_n20312_), .B(new_n20292_), .C(new_n5541_), .Y(new_n20319_));
  AOI21X1  g20127(.A0(new_n20319_), .A1(new_n20318_), .B0(new_n20313_), .Y(new_n20320_));
  OR2X1    g20128(.A(new_n20320_), .B(new_n5176_), .Y(new_n20321_));
  OR2X1    g20129(.A(new_n20310_), .B(new_n6294_), .Y(new_n20322_));
  NOR2X1   g20130(.A(new_n20281_), .B(new_n20280_), .Y(new_n20323_));
  INVX1    g20131(.A(new_n20289_), .Y(new_n20324_));
  NAND2X1  g20132(.A(new_n20276_), .B(new_n6294_), .Y(new_n20325_));
  OAI21X1  g20133(.A0(new_n20325_), .A1(new_n20323_), .B0(new_n20324_), .Y(new_n20326_));
  AOI21X1  g20134(.A0(new_n20326_), .A1(new_n20322_), .B0(new_n5941_), .Y(new_n20327_));
  AOI21X1  g20135(.A0(new_n20282_), .A1(\asqrt[33] ), .B0(\asqrt[34] ), .Y(new_n20328_));
  AOI21X1  g20136(.A0(new_n20328_), .A1(new_n20326_), .B0(new_n20297_), .Y(new_n20329_));
  NOR3X1   g20137(.A(new_n20329_), .B(new_n20327_), .C(\asqrt[35] ), .Y(new_n20330_));
  NOR2X1   g20138(.A(new_n20330_), .B(new_n20317_), .Y(new_n20331_));
  OAI21X1  g20139(.A0(new_n19622_), .A1(new_n19606_), .B0(new_n19611_), .Y(new_n20332_));
  NOR3X1   g20140(.A(new_n20332_), .B(new_n19976_), .C(new_n19643_), .Y(new_n20333_));
  AOI22X1  g20141(.A0(new_n19645_), .A1(new_n19644_), .B0(new_n19630_), .B1(\asqrt[35] ), .Y(new_n20334_));
  AOI21X1  g20142(.A0(new_n20334_), .A1(\asqrt[8] ), .B0(new_n19611_), .Y(new_n20335_));
  NOR2X1   g20143(.A(new_n20335_), .B(new_n20333_), .Y(new_n20336_));
  INVX1    g20144(.A(new_n20336_), .Y(new_n20337_));
  OAI21X1  g20145(.A0(new_n20329_), .A1(new_n20327_), .B0(\asqrt[35] ), .Y(new_n20338_));
  NAND2X1  g20146(.A(new_n20338_), .B(new_n5176_), .Y(new_n20339_));
  OAI21X1  g20147(.A0(new_n20339_), .A1(new_n20331_), .B0(new_n20337_), .Y(new_n20340_));
  AOI21X1  g20148(.A0(new_n20340_), .A1(new_n20321_), .B0(new_n4826_), .Y(new_n20341_));
  AND2X1   g20149(.A(new_n19631_), .B(new_n19623_), .Y(new_n20342_));
  OR4X1    g20150(.A(new_n19976_), .B(new_n20342_), .C(new_n19648_), .D(new_n19624_), .Y(new_n20343_));
  OR2X1    g20151(.A(new_n20342_), .B(new_n19624_), .Y(new_n20344_));
  OAI21X1  g20152(.A0(new_n20344_), .A1(new_n19976_), .B0(new_n19648_), .Y(new_n20345_));
  AND2X1   g20153(.A(new_n20345_), .B(new_n20343_), .Y(new_n20346_));
  OAI21X1  g20154(.A0(new_n20330_), .A1(new_n20317_), .B0(new_n20338_), .Y(new_n20347_));
  AOI21X1  g20155(.A0(new_n20347_), .A1(\asqrt[36] ), .B0(\asqrt[37] ), .Y(new_n20348_));
  AOI21X1  g20156(.A0(new_n20348_), .A1(new_n20340_), .B0(new_n20346_), .Y(new_n20349_));
  OAI21X1  g20157(.A0(new_n20349_), .A1(new_n20341_), .B0(\asqrt[38] ), .Y(new_n20350_));
  OR4X1    g20158(.A(new_n19976_), .B(new_n19639_), .C(new_n19642_), .D(new_n19666_), .Y(new_n20351_));
  NAND2X1  g20159(.A(new_n19651_), .B(new_n19633_), .Y(new_n20352_));
  OAI21X1  g20160(.A0(new_n20352_), .A1(new_n19976_), .B0(new_n19642_), .Y(new_n20353_));
  AND2X1   g20161(.A(new_n20353_), .B(new_n20351_), .Y(new_n20354_));
  NOR3X1   g20162(.A(new_n20349_), .B(new_n20341_), .C(\asqrt[38] ), .Y(new_n20355_));
  OAI21X1  g20163(.A0(new_n20355_), .A1(new_n20354_), .B0(new_n20350_), .Y(new_n20356_));
  AND2X1   g20164(.A(new_n20356_), .B(\asqrt[39] ), .Y(new_n20357_));
  OR2X1    g20165(.A(new_n20355_), .B(new_n20354_), .Y(new_n20358_));
  AND2X1   g20166(.A(new_n19658_), .B(new_n19652_), .Y(new_n20359_));
  NOR4X1   g20167(.A(new_n19976_), .B(new_n20359_), .C(new_n19682_), .D(new_n19641_), .Y(new_n20360_));
  AOI22X1  g20168(.A0(new_n19658_), .A1(new_n19652_), .B0(new_n19640_), .B1(\asqrt[38] ), .Y(new_n20361_));
  AOI21X1  g20169(.A0(new_n20361_), .A1(\asqrt[8] ), .B0(new_n19657_), .Y(new_n20362_));
  NOR2X1   g20170(.A(new_n20362_), .B(new_n20360_), .Y(new_n20363_));
  AND2X1   g20171(.A(new_n20350_), .B(new_n4165_), .Y(new_n20364_));
  AOI21X1  g20172(.A0(new_n20364_), .A1(new_n20358_), .B0(new_n20363_), .Y(new_n20365_));
  OAI21X1  g20173(.A0(new_n20365_), .A1(new_n20357_), .B0(\asqrt[40] ), .Y(new_n20366_));
  AND2X1   g20174(.A(new_n19686_), .B(new_n19684_), .Y(new_n20367_));
  OR4X1    g20175(.A(new_n19976_), .B(new_n20367_), .C(new_n19665_), .D(new_n19685_), .Y(new_n20368_));
  OR2X1    g20176(.A(new_n20367_), .B(new_n19685_), .Y(new_n20369_));
  OAI21X1  g20177(.A0(new_n20369_), .A1(new_n19976_), .B0(new_n19665_), .Y(new_n20370_));
  AND2X1   g20178(.A(new_n20370_), .B(new_n20368_), .Y(new_n20371_));
  INVX1    g20179(.A(new_n20371_), .Y(new_n20372_));
  AND2X1   g20180(.A(new_n20347_), .B(\asqrt[36] ), .Y(new_n20373_));
  OR2X1    g20181(.A(new_n20330_), .B(new_n20317_), .Y(new_n20374_));
  AND2X1   g20182(.A(new_n20338_), .B(new_n5176_), .Y(new_n20375_));
  AOI21X1  g20183(.A0(new_n20375_), .A1(new_n20374_), .B0(new_n20336_), .Y(new_n20376_));
  OAI21X1  g20184(.A0(new_n20376_), .A1(new_n20373_), .B0(\asqrt[37] ), .Y(new_n20377_));
  INVX1    g20185(.A(new_n20346_), .Y(new_n20378_));
  OAI21X1  g20186(.A0(new_n20320_), .A1(new_n5176_), .B0(new_n4826_), .Y(new_n20379_));
  OAI21X1  g20187(.A0(new_n20379_), .A1(new_n20376_), .B0(new_n20378_), .Y(new_n20380_));
  AOI21X1  g20188(.A0(new_n20380_), .A1(new_n20377_), .B0(new_n4493_), .Y(new_n20381_));
  INVX1    g20189(.A(new_n20354_), .Y(new_n20382_));
  NAND3X1  g20190(.A(new_n20380_), .B(new_n20377_), .C(new_n4493_), .Y(new_n20383_));
  AOI21X1  g20191(.A0(new_n20383_), .A1(new_n20382_), .B0(new_n20381_), .Y(new_n20384_));
  OAI21X1  g20192(.A0(new_n20384_), .A1(new_n4165_), .B0(new_n3863_), .Y(new_n20385_));
  OAI21X1  g20193(.A0(new_n20385_), .A1(new_n20365_), .B0(new_n20372_), .Y(new_n20386_));
  AOI21X1  g20194(.A0(new_n20386_), .A1(new_n20366_), .B0(new_n3564_), .Y(new_n20387_));
  OR4X1    g20195(.A(new_n19976_), .B(new_n19688_), .C(new_n19676_), .D(new_n19670_), .Y(new_n20388_));
  OR2X1    g20196(.A(new_n19688_), .B(new_n19670_), .Y(new_n20389_));
  OAI21X1  g20197(.A0(new_n20389_), .A1(new_n19976_), .B0(new_n19676_), .Y(new_n20390_));
  AND2X1   g20198(.A(new_n20390_), .B(new_n20388_), .Y(new_n20391_));
  INVX1    g20199(.A(new_n20391_), .Y(new_n20392_));
  NAND3X1  g20200(.A(new_n20386_), .B(new_n20366_), .C(new_n3564_), .Y(new_n20393_));
  AOI21X1  g20201(.A0(new_n20393_), .A1(new_n20392_), .B0(new_n20387_), .Y(new_n20394_));
  OR2X1    g20202(.A(new_n20394_), .B(new_n3276_), .Y(new_n20395_));
  OR2X1    g20203(.A(new_n20384_), .B(new_n4165_), .Y(new_n20396_));
  NOR2X1   g20204(.A(new_n20355_), .B(new_n20354_), .Y(new_n20397_));
  INVX1    g20205(.A(new_n20363_), .Y(new_n20398_));
  NAND2X1  g20206(.A(new_n20350_), .B(new_n4165_), .Y(new_n20399_));
  OAI21X1  g20207(.A0(new_n20399_), .A1(new_n20397_), .B0(new_n20398_), .Y(new_n20400_));
  AOI21X1  g20208(.A0(new_n20400_), .A1(new_n20396_), .B0(new_n3863_), .Y(new_n20401_));
  AOI21X1  g20209(.A0(new_n20356_), .A1(\asqrt[39] ), .B0(\asqrt[40] ), .Y(new_n20402_));
  AOI21X1  g20210(.A0(new_n20402_), .A1(new_n20400_), .B0(new_n20371_), .Y(new_n20403_));
  NOR3X1   g20211(.A(new_n20403_), .B(new_n20401_), .C(\asqrt[41] ), .Y(new_n20404_));
  NOR2X1   g20212(.A(new_n20404_), .B(new_n20391_), .Y(new_n20405_));
  OAI21X1  g20213(.A0(new_n19697_), .A1(new_n19689_), .B0(new_n19694_), .Y(new_n20406_));
  NOR3X1   g20214(.A(new_n20406_), .B(new_n19976_), .C(new_n19730_), .Y(new_n20407_));
  AOI22X1  g20215(.A0(new_n19732_), .A1(new_n19731_), .B0(new_n19704_), .B1(\asqrt[41] ), .Y(new_n20408_));
  AOI21X1  g20216(.A0(new_n20408_), .A1(\asqrt[8] ), .B0(new_n19694_), .Y(new_n20409_));
  NOR2X1   g20217(.A(new_n20409_), .B(new_n20407_), .Y(new_n20410_));
  INVX1    g20218(.A(new_n20410_), .Y(new_n20411_));
  OAI21X1  g20219(.A0(new_n20403_), .A1(new_n20401_), .B0(\asqrt[41] ), .Y(new_n20412_));
  NAND2X1  g20220(.A(new_n20412_), .B(new_n3276_), .Y(new_n20413_));
  OAI21X1  g20221(.A0(new_n20413_), .A1(new_n20405_), .B0(new_n20411_), .Y(new_n20414_));
  AOI21X1  g20222(.A0(new_n20414_), .A1(new_n20395_), .B0(new_n3008_), .Y(new_n20415_));
  AND2X1   g20223(.A(new_n19705_), .B(new_n19698_), .Y(new_n20416_));
  OR4X1    g20224(.A(new_n19976_), .B(new_n20416_), .C(new_n19735_), .D(new_n19699_), .Y(new_n20417_));
  OR2X1    g20225(.A(new_n20416_), .B(new_n19699_), .Y(new_n20418_));
  OAI21X1  g20226(.A0(new_n20418_), .A1(new_n19976_), .B0(new_n19735_), .Y(new_n20419_));
  AND2X1   g20227(.A(new_n20419_), .B(new_n20417_), .Y(new_n20420_));
  OAI21X1  g20228(.A0(new_n20404_), .A1(new_n20391_), .B0(new_n20412_), .Y(new_n20421_));
  AOI21X1  g20229(.A0(new_n20421_), .A1(\asqrt[42] ), .B0(\asqrt[43] ), .Y(new_n20422_));
  AOI21X1  g20230(.A0(new_n20422_), .A1(new_n20414_), .B0(new_n20420_), .Y(new_n20423_));
  OAI21X1  g20231(.A0(new_n20423_), .A1(new_n20415_), .B0(\asqrt[44] ), .Y(new_n20424_));
  OR4X1    g20232(.A(new_n19976_), .B(new_n19713_), .C(new_n19739_), .D(new_n19738_), .Y(new_n20425_));
  OR2X1    g20233(.A(new_n19713_), .B(new_n19738_), .Y(new_n20426_));
  OAI21X1  g20234(.A0(new_n20426_), .A1(new_n19976_), .B0(new_n19739_), .Y(new_n20427_));
  AND2X1   g20235(.A(new_n20427_), .B(new_n20425_), .Y(new_n20428_));
  NOR3X1   g20236(.A(new_n20423_), .B(new_n20415_), .C(\asqrt[44] ), .Y(new_n20429_));
  OAI21X1  g20237(.A0(new_n20429_), .A1(new_n20428_), .B0(new_n20424_), .Y(new_n20430_));
  AND2X1   g20238(.A(new_n20430_), .B(\asqrt[45] ), .Y(new_n20431_));
  OR2X1    g20239(.A(new_n20429_), .B(new_n20428_), .Y(new_n20432_));
  AND2X1   g20240(.A(new_n19722_), .B(new_n19716_), .Y(new_n20433_));
  NOR4X1   g20241(.A(new_n19976_), .B(new_n20433_), .C(new_n19756_), .D(new_n19715_), .Y(new_n20434_));
  AOI22X1  g20242(.A0(new_n19722_), .A1(new_n19716_), .B0(new_n19714_), .B1(\asqrt[44] ), .Y(new_n20435_));
  AOI21X1  g20243(.A0(new_n20435_), .A1(\asqrt[8] ), .B0(new_n19721_), .Y(new_n20436_));
  NOR2X1   g20244(.A(new_n20436_), .B(new_n20434_), .Y(new_n20437_));
  AND2X1   g20245(.A(new_n20424_), .B(new_n2570_), .Y(new_n20438_));
  AOI21X1  g20246(.A0(new_n20438_), .A1(new_n20432_), .B0(new_n20437_), .Y(new_n20439_));
  OAI21X1  g20247(.A0(new_n20439_), .A1(new_n20431_), .B0(\asqrt[46] ), .Y(new_n20440_));
  AND2X1   g20248(.A(new_n19760_), .B(new_n19758_), .Y(new_n20441_));
  OR4X1    g20249(.A(new_n19976_), .B(new_n20441_), .C(new_n19729_), .D(new_n19759_), .Y(new_n20442_));
  OR2X1    g20250(.A(new_n20441_), .B(new_n19759_), .Y(new_n20443_));
  OAI21X1  g20251(.A0(new_n20443_), .A1(new_n19976_), .B0(new_n19729_), .Y(new_n20444_));
  AND2X1   g20252(.A(new_n20444_), .B(new_n20442_), .Y(new_n20445_));
  INVX1    g20253(.A(new_n20445_), .Y(new_n20446_));
  AND2X1   g20254(.A(new_n20421_), .B(\asqrt[42] ), .Y(new_n20447_));
  OR2X1    g20255(.A(new_n20404_), .B(new_n20391_), .Y(new_n20448_));
  AND2X1   g20256(.A(new_n20412_), .B(new_n3276_), .Y(new_n20449_));
  AOI21X1  g20257(.A0(new_n20449_), .A1(new_n20448_), .B0(new_n20410_), .Y(new_n20450_));
  OAI21X1  g20258(.A0(new_n20450_), .A1(new_n20447_), .B0(\asqrt[43] ), .Y(new_n20451_));
  INVX1    g20259(.A(new_n20420_), .Y(new_n20452_));
  OAI21X1  g20260(.A0(new_n20394_), .A1(new_n3276_), .B0(new_n3008_), .Y(new_n20453_));
  OAI21X1  g20261(.A0(new_n20453_), .A1(new_n20450_), .B0(new_n20452_), .Y(new_n20454_));
  AOI21X1  g20262(.A0(new_n20454_), .A1(new_n20451_), .B0(new_n2769_), .Y(new_n20455_));
  INVX1    g20263(.A(new_n20428_), .Y(new_n20456_));
  NAND3X1  g20264(.A(new_n20454_), .B(new_n20451_), .C(new_n2769_), .Y(new_n20457_));
  AOI21X1  g20265(.A0(new_n20457_), .A1(new_n20456_), .B0(new_n20455_), .Y(new_n20458_));
  OAI21X1  g20266(.A0(new_n20458_), .A1(new_n2570_), .B0(new_n2263_), .Y(new_n20459_));
  OAI21X1  g20267(.A0(new_n20459_), .A1(new_n20439_), .B0(new_n20446_), .Y(new_n20460_));
  AOI21X1  g20268(.A0(new_n20460_), .A1(new_n20440_), .B0(new_n2040_), .Y(new_n20461_));
  OR4X1    g20269(.A(new_n19976_), .B(new_n19762_), .C(new_n19750_), .D(new_n19744_), .Y(new_n20462_));
  OR2X1    g20270(.A(new_n19762_), .B(new_n19744_), .Y(new_n20463_));
  OAI21X1  g20271(.A0(new_n20463_), .A1(new_n19976_), .B0(new_n19750_), .Y(new_n20464_));
  AND2X1   g20272(.A(new_n20464_), .B(new_n20462_), .Y(new_n20465_));
  INVX1    g20273(.A(new_n20465_), .Y(new_n20466_));
  NAND3X1  g20274(.A(new_n20460_), .B(new_n20440_), .C(new_n2040_), .Y(new_n20467_));
  AOI21X1  g20275(.A0(new_n20467_), .A1(new_n20466_), .B0(new_n20461_), .Y(new_n20468_));
  OR2X1    g20276(.A(new_n20468_), .B(new_n1834_), .Y(new_n20469_));
  OR2X1    g20277(.A(new_n20458_), .B(new_n2570_), .Y(new_n20470_));
  NOR2X1   g20278(.A(new_n20429_), .B(new_n20428_), .Y(new_n20471_));
  INVX1    g20279(.A(new_n20437_), .Y(new_n20472_));
  NAND2X1  g20280(.A(new_n20424_), .B(new_n2570_), .Y(new_n20473_));
  OAI21X1  g20281(.A0(new_n20473_), .A1(new_n20471_), .B0(new_n20472_), .Y(new_n20474_));
  AOI21X1  g20282(.A0(new_n20474_), .A1(new_n20470_), .B0(new_n2263_), .Y(new_n20475_));
  AOI21X1  g20283(.A0(new_n20430_), .A1(\asqrt[45] ), .B0(\asqrt[46] ), .Y(new_n20476_));
  AOI21X1  g20284(.A0(new_n20476_), .A1(new_n20474_), .B0(new_n20445_), .Y(new_n20477_));
  NOR3X1   g20285(.A(new_n20477_), .B(new_n20475_), .C(\asqrt[47] ), .Y(new_n20478_));
  NOR2X1   g20286(.A(new_n20478_), .B(new_n20465_), .Y(new_n20479_));
  OAI21X1  g20287(.A0(new_n19771_), .A1(new_n19763_), .B0(new_n19768_), .Y(new_n20480_));
  NOR3X1   g20288(.A(new_n20480_), .B(new_n19976_), .C(new_n19804_), .Y(new_n20481_));
  AOI22X1  g20289(.A0(new_n19806_), .A1(new_n19805_), .B0(new_n19778_), .B1(\asqrt[47] ), .Y(new_n20482_));
  AOI21X1  g20290(.A0(new_n20482_), .A1(\asqrt[8] ), .B0(new_n19768_), .Y(new_n20483_));
  NOR2X1   g20291(.A(new_n20483_), .B(new_n20481_), .Y(new_n20484_));
  INVX1    g20292(.A(new_n20484_), .Y(new_n20485_));
  OAI21X1  g20293(.A0(new_n20477_), .A1(new_n20475_), .B0(\asqrt[47] ), .Y(new_n20486_));
  NAND2X1  g20294(.A(new_n20486_), .B(new_n1834_), .Y(new_n20487_));
  OAI21X1  g20295(.A0(new_n20487_), .A1(new_n20479_), .B0(new_n20485_), .Y(new_n20488_));
  AOI21X1  g20296(.A0(new_n20488_), .A1(new_n20469_), .B0(new_n1632_), .Y(new_n20489_));
  AND2X1   g20297(.A(new_n19779_), .B(new_n19772_), .Y(new_n20490_));
  OR2X1    g20298(.A(new_n19809_), .B(new_n19773_), .Y(new_n20491_));
  OR2X1    g20299(.A(new_n20491_), .B(new_n20490_), .Y(new_n20492_));
  NOR3X1   g20300(.A(new_n19976_), .B(new_n20490_), .C(new_n19773_), .Y(new_n20493_));
  OAI22X1  g20301(.A0(new_n20493_), .A1(new_n19777_), .B0(new_n20492_), .B1(new_n19976_), .Y(new_n20494_));
  INVX1    g20302(.A(new_n20494_), .Y(new_n20495_));
  OAI21X1  g20303(.A0(new_n20478_), .A1(new_n20465_), .B0(new_n20486_), .Y(new_n20496_));
  AOI21X1  g20304(.A0(new_n20496_), .A1(\asqrt[48] ), .B0(\asqrt[49] ), .Y(new_n20497_));
  AOI21X1  g20305(.A0(new_n20497_), .A1(new_n20488_), .B0(new_n20495_), .Y(new_n20498_));
  OAI21X1  g20306(.A0(new_n20498_), .A1(new_n20489_), .B0(\asqrt[50] ), .Y(new_n20499_));
  OR4X1    g20307(.A(new_n19976_), .B(new_n19787_), .C(new_n19813_), .D(new_n19812_), .Y(new_n20500_));
  OR2X1    g20308(.A(new_n19787_), .B(new_n19812_), .Y(new_n20501_));
  OAI21X1  g20309(.A0(new_n20501_), .A1(new_n19976_), .B0(new_n19813_), .Y(new_n20502_));
  AND2X1   g20310(.A(new_n20502_), .B(new_n20500_), .Y(new_n20503_));
  NOR3X1   g20311(.A(new_n20498_), .B(new_n20489_), .C(\asqrt[50] ), .Y(new_n20504_));
  OAI21X1  g20312(.A0(new_n20504_), .A1(new_n20503_), .B0(new_n20499_), .Y(new_n20505_));
  AND2X1   g20313(.A(new_n20505_), .B(\asqrt[51] ), .Y(new_n20506_));
  OR2X1    g20314(.A(new_n20504_), .B(new_n20503_), .Y(new_n20507_));
  AND2X1   g20315(.A(new_n19796_), .B(new_n19790_), .Y(new_n20508_));
  NOR4X1   g20316(.A(new_n19976_), .B(new_n20508_), .C(new_n19830_), .D(new_n19789_), .Y(new_n20509_));
  AOI22X1  g20317(.A0(new_n19796_), .A1(new_n19790_), .B0(new_n19788_), .B1(\asqrt[50] ), .Y(new_n20510_));
  AOI21X1  g20318(.A0(new_n20510_), .A1(\asqrt[8] ), .B0(new_n19795_), .Y(new_n20511_));
  NOR2X1   g20319(.A(new_n20511_), .B(new_n20509_), .Y(new_n20512_));
  AND2X1   g20320(.A(new_n20499_), .B(new_n1277_), .Y(new_n20513_));
  AOI21X1  g20321(.A0(new_n20513_), .A1(new_n20507_), .B0(new_n20512_), .Y(new_n20514_));
  OAI21X1  g20322(.A0(new_n20514_), .A1(new_n20506_), .B0(\asqrt[52] ), .Y(new_n20515_));
  AND2X1   g20323(.A(new_n19834_), .B(new_n19832_), .Y(new_n20516_));
  OR4X1    g20324(.A(new_n19976_), .B(new_n20516_), .C(new_n19803_), .D(new_n19833_), .Y(new_n20517_));
  OR2X1    g20325(.A(new_n20516_), .B(new_n19833_), .Y(new_n20518_));
  OAI21X1  g20326(.A0(new_n20518_), .A1(new_n19976_), .B0(new_n19803_), .Y(new_n20519_));
  AND2X1   g20327(.A(new_n20519_), .B(new_n20517_), .Y(new_n20520_));
  INVX1    g20328(.A(new_n20520_), .Y(new_n20521_));
  AND2X1   g20329(.A(new_n20496_), .B(\asqrt[48] ), .Y(new_n20522_));
  OR2X1    g20330(.A(new_n20478_), .B(new_n20465_), .Y(new_n20523_));
  AND2X1   g20331(.A(new_n20486_), .B(new_n1834_), .Y(new_n20524_));
  AOI21X1  g20332(.A0(new_n20524_), .A1(new_n20523_), .B0(new_n20484_), .Y(new_n20525_));
  OAI21X1  g20333(.A0(new_n20525_), .A1(new_n20522_), .B0(\asqrt[49] ), .Y(new_n20526_));
  OAI21X1  g20334(.A0(new_n20468_), .A1(new_n1834_), .B0(new_n1632_), .Y(new_n20527_));
  OAI21X1  g20335(.A0(new_n20527_), .A1(new_n20525_), .B0(new_n20494_), .Y(new_n20528_));
  AOI21X1  g20336(.A0(new_n20528_), .A1(new_n20526_), .B0(new_n1469_), .Y(new_n20529_));
  INVX1    g20337(.A(new_n20503_), .Y(new_n20530_));
  NAND3X1  g20338(.A(new_n20528_), .B(new_n20526_), .C(new_n1469_), .Y(new_n20531_));
  AOI21X1  g20339(.A0(new_n20531_), .A1(new_n20530_), .B0(new_n20529_), .Y(new_n20532_));
  OAI21X1  g20340(.A0(new_n20532_), .A1(new_n1277_), .B0(new_n1111_), .Y(new_n20533_));
  OAI21X1  g20341(.A0(new_n20533_), .A1(new_n20514_), .B0(new_n20521_), .Y(new_n20534_));
  AOI21X1  g20342(.A0(new_n20534_), .A1(new_n20515_), .B0(new_n968_), .Y(new_n20535_));
  OR4X1    g20343(.A(new_n19976_), .B(new_n19836_), .C(new_n19824_), .D(new_n19818_), .Y(new_n20536_));
  OR2X1    g20344(.A(new_n19836_), .B(new_n19818_), .Y(new_n20537_));
  OAI21X1  g20345(.A0(new_n20537_), .A1(new_n19976_), .B0(new_n19824_), .Y(new_n20538_));
  AND2X1   g20346(.A(new_n20538_), .B(new_n20536_), .Y(new_n20539_));
  INVX1    g20347(.A(new_n20539_), .Y(new_n20540_));
  NAND3X1  g20348(.A(new_n20534_), .B(new_n20515_), .C(new_n968_), .Y(new_n20541_));
  AOI21X1  g20349(.A0(new_n20541_), .A1(new_n20540_), .B0(new_n20535_), .Y(new_n20542_));
  OR2X1    g20350(.A(new_n20542_), .B(new_n902_), .Y(new_n20543_));
  OR2X1    g20351(.A(new_n20532_), .B(new_n1277_), .Y(new_n20544_));
  NOR2X1   g20352(.A(new_n20504_), .B(new_n20503_), .Y(new_n20545_));
  INVX1    g20353(.A(new_n20512_), .Y(new_n20546_));
  NAND2X1  g20354(.A(new_n20499_), .B(new_n1277_), .Y(new_n20547_));
  OAI21X1  g20355(.A0(new_n20547_), .A1(new_n20545_), .B0(new_n20546_), .Y(new_n20548_));
  AOI21X1  g20356(.A0(new_n20548_), .A1(new_n20544_), .B0(new_n1111_), .Y(new_n20549_));
  AOI21X1  g20357(.A0(new_n20505_), .A1(\asqrt[51] ), .B0(\asqrt[52] ), .Y(new_n20550_));
  AOI21X1  g20358(.A0(new_n20550_), .A1(new_n20548_), .B0(new_n20520_), .Y(new_n20551_));
  NOR3X1   g20359(.A(new_n20551_), .B(new_n20549_), .C(\asqrt[53] ), .Y(new_n20552_));
  NOR2X1   g20360(.A(new_n20552_), .B(new_n20539_), .Y(new_n20553_));
  OAI21X1  g20361(.A0(new_n19845_), .A1(new_n19837_), .B0(new_n19842_), .Y(new_n20554_));
  NOR3X1   g20362(.A(new_n20554_), .B(new_n19976_), .C(new_n19878_), .Y(new_n20555_));
  AOI22X1  g20363(.A0(new_n19880_), .A1(new_n19879_), .B0(new_n19852_), .B1(\asqrt[53] ), .Y(new_n20556_));
  AOI21X1  g20364(.A0(new_n20556_), .A1(\asqrt[8] ), .B0(new_n19842_), .Y(new_n20557_));
  NOR2X1   g20365(.A(new_n20557_), .B(new_n20555_), .Y(new_n20558_));
  INVX1    g20366(.A(new_n20558_), .Y(new_n20559_));
  OAI21X1  g20367(.A0(new_n20551_), .A1(new_n20549_), .B0(\asqrt[53] ), .Y(new_n20560_));
  NAND2X1  g20368(.A(new_n20560_), .B(new_n902_), .Y(new_n20561_));
  OAI21X1  g20369(.A0(new_n20561_), .A1(new_n20553_), .B0(new_n20559_), .Y(new_n20562_));
  AOI21X1  g20370(.A0(new_n20562_), .A1(new_n20543_), .B0(new_n697_), .Y(new_n20563_));
  AND2X1   g20371(.A(new_n19853_), .B(new_n19846_), .Y(new_n20564_));
  OR4X1    g20372(.A(new_n19976_), .B(new_n20564_), .C(new_n19883_), .D(new_n19847_), .Y(new_n20565_));
  OR2X1    g20373(.A(new_n20564_), .B(new_n19847_), .Y(new_n20566_));
  OAI21X1  g20374(.A0(new_n20566_), .A1(new_n19976_), .B0(new_n19883_), .Y(new_n20567_));
  AND2X1   g20375(.A(new_n20567_), .B(new_n20565_), .Y(new_n20568_));
  OAI21X1  g20376(.A0(new_n20552_), .A1(new_n20539_), .B0(new_n20560_), .Y(new_n20569_));
  AOI21X1  g20377(.A0(new_n20569_), .A1(\asqrt[54] ), .B0(\asqrt[55] ), .Y(new_n20570_));
  AOI21X1  g20378(.A0(new_n20570_), .A1(new_n20562_), .B0(new_n20568_), .Y(new_n20571_));
  OAI21X1  g20379(.A0(new_n20571_), .A1(new_n20563_), .B0(\asqrt[56] ), .Y(new_n20572_));
  OR4X1    g20380(.A(new_n19976_), .B(new_n19861_), .C(new_n19887_), .D(new_n19886_), .Y(new_n20573_));
  OR2X1    g20381(.A(new_n19861_), .B(new_n19886_), .Y(new_n20574_));
  OAI21X1  g20382(.A0(new_n20574_), .A1(new_n19976_), .B0(new_n19887_), .Y(new_n20575_));
  AND2X1   g20383(.A(new_n20575_), .B(new_n20573_), .Y(new_n20576_));
  NOR3X1   g20384(.A(new_n20571_), .B(new_n20563_), .C(\asqrt[56] ), .Y(new_n20577_));
  OAI21X1  g20385(.A0(new_n20577_), .A1(new_n20576_), .B0(new_n20572_), .Y(new_n20578_));
  AND2X1   g20386(.A(new_n20578_), .B(\asqrt[57] ), .Y(new_n20579_));
  OR2X1    g20387(.A(new_n20577_), .B(new_n20576_), .Y(new_n20580_));
  AND2X1   g20388(.A(new_n20572_), .B(new_n481_), .Y(new_n20581_));
  AND2X1   g20389(.A(new_n19865_), .B(new_n19864_), .Y(new_n20582_));
  NOR4X1   g20390(.A(new_n19976_), .B(new_n19905_), .C(new_n20582_), .D(new_n19863_), .Y(new_n20583_));
  AOI22X1  g20391(.A0(new_n19865_), .A1(new_n19864_), .B0(new_n19862_), .B1(\asqrt[56] ), .Y(new_n20584_));
  AOI21X1  g20392(.A0(new_n20584_), .A1(\asqrt[8] ), .B0(new_n19870_), .Y(new_n20585_));
  NOR2X1   g20393(.A(new_n20585_), .B(new_n20583_), .Y(new_n20586_));
  AOI21X1  g20394(.A0(new_n20581_), .A1(new_n20580_), .B0(new_n20586_), .Y(new_n20587_));
  OAI21X1  g20395(.A0(new_n20587_), .A1(new_n20579_), .B0(\asqrt[58] ), .Y(new_n20588_));
  AND2X1   g20396(.A(new_n19908_), .B(new_n19906_), .Y(new_n20589_));
  OR4X1    g20397(.A(new_n19976_), .B(new_n20589_), .C(new_n19877_), .D(new_n19907_), .Y(new_n20590_));
  OR2X1    g20398(.A(new_n20589_), .B(new_n19907_), .Y(new_n20591_));
  OAI21X1  g20399(.A0(new_n20591_), .A1(new_n19976_), .B0(new_n19877_), .Y(new_n20592_));
  AND2X1   g20400(.A(new_n20592_), .B(new_n20590_), .Y(new_n20593_));
  INVX1    g20401(.A(new_n20593_), .Y(new_n20594_));
  AND2X1   g20402(.A(new_n20569_), .B(\asqrt[54] ), .Y(new_n20595_));
  OR2X1    g20403(.A(new_n20552_), .B(new_n20539_), .Y(new_n20596_));
  AND2X1   g20404(.A(new_n20560_), .B(new_n902_), .Y(new_n20597_));
  AOI21X1  g20405(.A0(new_n20597_), .A1(new_n20596_), .B0(new_n20558_), .Y(new_n20598_));
  OAI21X1  g20406(.A0(new_n20598_), .A1(new_n20595_), .B0(\asqrt[55] ), .Y(new_n20599_));
  INVX1    g20407(.A(new_n20568_), .Y(new_n20600_));
  OAI21X1  g20408(.A0(new_n20542_), .A1(new_n902_), .B0(new_n697_), .Y(new_n20601_));
  OAI21X1  g20409(.A0(new_n20601_), .A1(new_n20598_), .B0(new_n20600_), .Y(new_n20602_));
  AOI21X1  g20410(.A0(new_n20602_), .A1(new_n20599_), .B0(new_n582_), .Y(new_n20603_));
  INVX1    g20411(.A(new_n20576_), .Y(new_n20604_));
  NAND3X1  g20412(.A(new_n20602_), .B(new_n20599_), .C(new_n582_), .Y(new_n20605_));
  AOI21X1  g20413(.A0(new_n20605_), .A1(new_n20604_), .B0(new_n20603_), .Y(new_n20606_));
  OAI21X1  g20414(.A0(new_n20606_), .A1(new_n481_), .B0(new_n399_), .Y(new_n20607_));
  OAI21X1  g20415(.A0(new_n20607_), .A1(new_n20587_), .B0(new_n20594_), .Y(new_n20608_));
  AOI21X1  g20416(.A0(new_n20608_), .A1(new_n20588_), .B0(new_n328_), .Y(new_n20609_));
  NAND3X1  g20417(.A(new_n19899_), .B(new_n19897_), .C(new_n19918_), .Y(new_n20610_));
  NOR3X1   g20418(.A(new_n19976_), .B(new_n19910_), .C(new_n19892_), .Y(new_n20611_));
  OAI22X1  g20419(.A0(new_n20611_), .A1(new_n19897_), .B0(new_n20610_), .B1(new_n19976_), .Y(new_n20612_));
  NAND3X1  g20420(.A(new_n20608_), .B(new_n20588_), .C(new_n328_), .Y(new_n20613_));
  AOI21X1  g20421(.A0(new_n20613_), .A1(new_n20612_), .B0(new_n20609_), .Y(new_n20614_));
  OR2X1    g20422(.A(new_n20614_), .B(new_n292_), .Y(new_n20615_));
  INVX1    g20423(.A(new_n20612_), .Y(new_n20616_));
  OR2X1    g20424(.A(new_n20606_), .B(new_n481_), .Y(new_n20617_));
  NOR2X1   g20425(.A(new_n20577_), .B(new_n20576_), .Y(new_n20618_));
  NAND2X1  g20426(.A(new_n20572_), .B(new_n481_), .Y(new_n20619_));
  INVX1    g20427(.A(new_n20586_), .Y(new_n20620_));
  OAI21X1  g20428(.A0(new_n20619_), .A1(new_n20618_), .B0(new_n20620_), .Y(new_n20621_));
  AOI21X1  g20429(.A0(new_n20621_), .A1(new_n20617_), .B0(new_n399_), .Y(new_n20622_));
  AOI21X1  g20430(.A0(new_n20578_), .A1(\asqrt[57] ), .B0(\asqrt[58] ), .Y(new_n20623_));
  AOI21X1  g20431(.A0(new_n20623_), .A1(new_n20621_), .B0(new_n20593_), .Y(new_n20624_));
  NOR3X1   g20432(.A(new_n20624_), .B(new_n20622_), .C(\asqrt[59] ), .Y(new_n20625_));
  NOR2X1   g20433(.A(new_n20625_), .B(new_n20616_), .Y(new_n20626_));
  OAI21X1  g20434(.A0(new_n19919_), .A1(new_n19911_), .B0(new_n19916_), .Y(new_n20627_));
  NOR3X1   g20435(.A(new_n20627_), .B(new_n19976_), .C(new_n19955_), .Y(new_n20628_));
  AOI22X1  g20436(.A0(new_n19957_), .A1(new_n19956_), .B0(new_n19926_), .B1(\asqrt[59] ), .Y(new_n20629_));
  AOI21X1  g20437(.A0(new_n20629_), .A1(\asqrt[8] ), .B0(new_n19916_), .Y(new_n20630_));
  NOR2X1   g20438(.A(new_n20630_), .B(new_n20628_), .Y(new_n20631_));
  INVX1    g20439(.A(new_n20631_), .Y(new_n20632_));
  OAI21X1  g20440(.A0(new_n20624_), .A1(new_n20622_), .B0(\asqrt[59] ), .Y(new_n20633_));
  NAND2X1  g20441(.A(new_n20633_), .B(new_n292_), .Y(new_n20634_));
  OAI21X1  g20442(.A0(new_n20634_), .A1(new_n20626_), .B0(new_n20632_), .Y(new_n20635_));
  AOI21X1  g20443(.A0(new_n20635_), .A1(new_n20615_), .B0(new_n217_), .Y(new_n20636_));
  AND2X1   g20444(.A(new_n19927_), .B(new_n19920_), .Y(new_n20637_));
  OR4X1    g20445(.A(new_n19976_), .B(new_n20637_), .C(new_n19960_), .D(new_n19921_), .Y(new_n20638_));
  OR2X1    g20446(.A(new_n20637_), .B(new_n19921_), .Y(new_n20639_));
  OAI21X1  g20447(.A0(new_n20639_), .A1(new_n19976_), .B0(new_n19960_), .Y(new_n20640_));
  AND2X1   g20448(.A(new_n20640_), .B(new_n20638_), .Y(new_n20641_));
  OAI21X1  g20449(.A0(new_n20625_), .A1(new_n20616_), .B0(new_n20633_), .Y(new_n20642_));
  AOI21X1  g20450(.A0(new_n20642_), .A1(\asqrt[60] ), .B0(\asqrt[61] ), .Y(new_n20643_));
  AOI21X1  g20451(.A0(new_n20643_), .A1(new_n20635_), .B0(new_n20641_), .Y(new_n20644_));
  OAI21X1  g20452(.A0(new_n20644_), .A1(new_n20636_), .B0(\asqrt[62] ), .Y(new_n20645_));
  OR4X1    g20453(.A(new_n19976_), .B(new_n19935_), .C(new_n19964_), .D(new_n19963_), .Y(new_n20646_));
  OR2X1    g20454(.A(new_n19935_), .B(new_n19963_), .Y(new_n20647_));
  OAI21X1  g20455(.A0(new_n20647_), .A1(new_n19976_), .B0(new_n19964_), .Y(new_n20648_));
  AND2X1   g20456(.A(new_n20648_), .B(new_n20646_), .Y(new_n20649_));
  NOR3X1   g20457(.A(new_n20644_), .B(new_n20636_), .C(\asqrt[62] ), .Y(new_n20650_));
  OAI21X1  g20458(.A0(new_n20650_), .A1(new_n20649_), .B0(new_n20645_), .Y(new_n20651_));
  AND2X1   g20459(.A(new_n19944_), .B(new_n19938_), .Y(new_n20652_));
  NOR4X1   g20460(.A(new_n19976_), .B(new_n20652_), .C(new_n19979_), .D(new_n19937_), .Y(new_n20653_));
  AOI22X1  g20461(.A0(new_n19944_), .A1(new_n19938_), .B0(new_n19936_), .B1(\asqrt[62] ), .Y(new_n20654_));
  AOI21X1  g20462(.A0(new_n20654_), .A1(\asqrt[8] ), .B0(new_n19943_), .Y(new_n20655_));
  NOR2X1   g20463(.A(new_n20655_), .B(new_n20653_), .Y(new_n20656_));
  INVX1    g20464(.A(new_n20656_), .Y(new_n20657_));
  AND2X1   g20465(.A(new_n19984_), .B(new_n19981_), .Y(new_n20658_));
  AOI21X1  g20466(.A0(new_n19981_), .A1(new_n19977_), .B0(new_n19949_), .Y(new_n20659_));
  AOI21X1  g20467(.A0(new_n20659_), .A1(\asqrt[8] ), .B0(new_n20658_), .Y(new_n20660_));
  AND2X1   g20468(.A(new_n20660_), .B(new_n20657_), .Y(new_n20661_));
  AOI21X1  g20469(.A0(new_n20661_), .A1(new_n20651_), .B0(\asqrt[63] ), .Y(new_n20662_));
  NOR2X1   g20470(.A(new_n20650_), .B(new_n20649_), .Y(new_n20663_));
  NAND2X1  g20471(.A(new_n20656_), .B(new_n20645_), .Y(new_n20664_));
  AND2X1   g20472(.A(new_n19981_), .B(new_n19977_), .Y(new_n20665_));
  OAI21X1  g20473(.A0(new_n19976_), .A1(new_n19949_), .B0(new_n20665_), .Y(new_n20666_));
  NOR2X1   g20474(.A(new_n20659_), .B(new_n193_), .Y(new_n20667_));
  AND2X1   g20475(.A(new_n19954_), .B(new_n193_), .Y(new_n20668_));
  OAI21X1  g20476(.A0(new_n19946_), .A1(new_n19273_), .B0(new_n19973_), .Y(new_n20669_));
  AOI21X1  g20477(.A0(new_n19948_), .A1(new_n19293_), .B0(new_n20669_), .Y(new_n20670_));
  NAND2X1  g20478(.A(new_n20670_), .B(new_n19970_), .Y(new_n20671_));
  OR2X1    g20479(.A(new_n20671_), .B(new_n20658_), .Y(new_n20672_));
  NOR2X1   g20480(.A(new_n20672_), .B(new_n20668_), .Y(new_n20673_));
  AOI21X1  g20481(.A0(new_n20667_), .A1(new_n20666_), .B0(new_n20673_), .Y(new_n20674_));
  OAI21X1  g20482(.A0(new_n20664_), .A1(new_n20663_), .B0(new_n20674_), .Y(new_n20675_));
  NOR2X1   g20483(.A(new_n20675_), .B(new_n20662_), .Y(new_n20676_));
  INVX1    g20484(.A(new_n20676_), .Y(\asqrt[7] ));
  OAI21X1  g20485(.A0(new_n20675_), .A1(new_n20662_), .B0(\a[14] ), .Y(new_n20678_));
  INVX1    g20486(.A(\a[14] ), .Y(new_n20679_));
  NOR2X1   g20487(.A(\a[13] ), .B(\a[12] ), .Y(new_n20680_));
  NAND2X1  g20488(.A(new_n20680_), .B(new_n20679_), .Y(new_n20681_));
  AND2X1   g20489(.A(new_n20681_), .B(new_n20678_), .Y(new_n20682_));
  AND2X1   g20490(.A(new_n20642_), .B(\asqrt[60] ), .Y(new_n20683_));
  OR2X1    g20491(.A(new_n20625_), .B(new_n20616_), .Y(new_n20684_));
  AND2X1   g20492(.A(new_n20633_), .B(new_n292_), .Y(new_n20685_));
  AOI21X1  g20493(.A0(new_n20685_), .A1(new_n20684_), .B0(new_n20631_), .Y(new_n20686_));
  OAI21X1  g20494(.A0(new_n20686_), .A1(new_n20683_), .B0(\asqrt[61] ), .Y(new_n20687_));
  INVX1    g20495(.A(new_n20641_), .Y(new_n20688_));
  OAI21X1  g20496(.A0(new_n20614_), .A1(new_n292_), .B0(new_n217_), .Y(new_n20689_));
  OAI21X1  g20497(.A0(new_n20689_), .A1(new_n20686_), .B0(new_n20688_), .Y(new_n20690_));
  AOI21X1  g20498(.A0(new_n20690_), .A1(new_n20687_), .B0(new_n199_), .Y(new_n20691_));
  INVX1    g20499(.A(new_n20649_), .Y(new_n20692_));
  NAND3X1  g20500(.A(new_n20690_), .B(new_n20687_), .C(new_n199_), .Y(new_n20693_));
  AOI21X1  g20501(.A0(new_n20693_), .A1(new_n20692_), .B0(new_n20691_), .Y(new_n20694_));
  INVX1    g20502(.A(new_n20661_), .Y(new_n20695_));
  OAI21X1  g20503(.A0(new_n20695_), .A1(new_n20694_), .B0(new_n193_), .Y(new_n20696_));
  OR2X1    g20504(.A(new_n20650_), .B(new_n20649_), .Y(new_n20697_));
  AND2X1   g20505(.A(new_n20656_), .B(new_n20645_), .Y(new_n20698_));
  INVX1    g20506(.A(new_n20674_), .Y(new_n20699_));
  AOI21X1  g20507(.A0(new_n20698_), .A1(new_n20697_), .B0(new_n20699_), .Y(new_n20700_));
  AOI21X1  g20508(.A0(new_n20700_), .A1(new_n20696_), .B0(new_n20679_), .Y(new_n20701_));
  NAND3X1  g20509(.A(new_n20681_), .B(new_n19973_), .C(new_n19970_), .Y(new_n20702_));
  NOR4X1   g20510(.A(new_n20702_), .B(new_n20701_), .C(new_n20658_), .D(new_n20668_), .Y(new_n20703_));
  INVX1    g20511(.A(\a[15] ), .Y(new_n20704_));
  AOI21X1  g20512(.A0(new_n20700_), .A1(new_n20696_), .B0(\a[14] ), .Y(new_n20705_));
  OAI21X1  g20513(.A0(new_n20675_), .A1(new_n20662_), .B0(new_n19988_), .Y(new_n20706_));
  OAI21X1  g20514(.A0(new_n20705_), .A1(new_n20704_), .B0(new_n20706_), .Y(new_n20707_));
  OAI22X1  g20515(.A0(new_n20707_), .A1(new_n20703_), .B0(new_n20682_), .B1(new_n19976_), .Y(new_n20708_));
  AND2X1   g20516(.A(new_n20708_), .B(\asqrt[9] ), .Y(new_n20709_));
  OR4X1    g20517(.A(new_n20702_), .B(new_n20701_), .C(new_n20658_), .D(new_n20668_), .Y(new_n20710_));
  OAI21X1  g20518(.A0(new_n20675_), .A1(new_n20662_), .B0(new_n20679_), .Y(new_n20711_));
  AOI21X1  g20519(.A0(new_n20700_), .A1(new_n20696_), .B0(new_n20002_), .Y(new_n20712_));
  AOI21X1  g20520(.A0(new_n20711_), .A1(\a[15] ), .B0(new_n20712_), .Y(new_n20713_));
  NAND2X1  g20521(.A(new_n20713_), .B(new_n20710_), .Y(new_n20714_));
  AOI21X1  g20522(.A0(new_n20681_), .A1(new_n20678_), .B0(new_n19976_), .Y(new_n20715_));
  NOR2X1   g20523(.A(new_n20715_), .B(\asqrt[9] ), .Y(new_n20716_));
  AND2X1   g20524(.A(new_n20698_), .B(new_n20697_), .Y(new_n20717_));
  AND2X1   g20525(.A(new_n20667_), .B(new_n20666_), .Y(new_n20718_));
  OAI21X1  g20526(.A0(new_n20672_), .A1(new_n20668_), .B0(\asqrt[8] ), .Y(new_n20719_));
  OR4X1    g20527(.A(new_n20719_), .B(new_n20718_), .C(new_n20717_), .D(new_n20662_), .Y(new_n20720_));
  AOI21X1  g20528(.A0(new_n20720_), .A1(new_n20706_), .B0(new_n19995_), .Y(new_n20721_));
  NOR4X1   g20529(.A(new_n20719_), .B(new_n20718_), .C(new_n20717_), .D(new_n20662_), .Y(new_n20722_));
  NOR3X1   g20530(.A(new_n20722_), .B(new_n20712_), .C(\a[16] ), .Y(new_n20723_));
  NOR2X1   g20531(.A(new_n20723_), .B(new_n20721_), .Y(new_n20724_));
  AOI21X1  g20532(.A0(new_n20716_), .A1(new_n20714_), .B0(new_n20724_), .Y(new_n20725_));
  OAI21X1  g20533(.A0(new_n20725_), .A1(new_n20709_), .B0(\asqrt[10] ), .Y(new_n20726_));
  AND2X1   g20534(.A(new_n20043_), .B(new_n20041_), .Y(new_n20727_));
  NOR3X1   g20535(.A(new_n20727_), .B(new_n19994_), .C(new_n19990_), .Y(new_n20728_));
  OAI21X1  g20536(.A0(new_n20675_), .A1(new_n20662_), .B0(new_n20728_), .Y(new_n20729_));
  AOI21X1  g20537(.A0(new_n19989_), .A1(\asqrt[9] ), .B0(new_n19994_), .Y(new_n20730_));
  OAI21X1  g20538(.A0(new_n20675_), .A1(new_n20662_), .B0(new_n20730_), .Y(new_n20731_));
  NAND2X1  g20539(.A(new_n20731_), .B(new_n20727_), .Y(new_n20732_));
  NAND2X1  g20540(.A(new_n20732_), .B(new_n20729_), .Y(new_n20733_));
  AOI21X1  g20541(.A0(new_n20713_), .A1(new_n20710_), .B0(new_n20715_), .Y(new_n20734_));
  OAI21X1  g20542(.A0(new_n20734_), .A1(new_n19273_), .B0(new_n18591_), .Y(new_n20735_));
  OAI21X1  g20543(.A0(new_n20735_), .A1(new_n20725_), .B0(new_n20733_), .Y(new_n20736_));
  AOI21X1  g20544(.A0(new_n20736_), .A1(new_n20726_), .B0(new_n17927_), .Y(new_n20737_));
  AND2X1   g20545(.A(new_n20046_), .B(new_n20044_), .Y(new_n20738_));
  NOR3X1   g20546(.A(new_n20011_), .B(new_n20738_), .C(new_n20045_), .Y(new_n20739_));
  OAI21X1  g20547(.A0(new_n20675_), .A1(new_n20662_), .B0(new_n20739_), .Y(new_n20740_));
  NOR2X1   g20548(.A(new_n20738_), .B(new_n20045_), .Y(new_n20741_));
  OAI21X1  g20549(.A0(new_n20675_), .A1(new_n20662_), .B0(new_n20741_), .Y(new_n20742_));
  NAND2X1  g20550(.A(new_n20742_), .B(new_n20011_), .Y(new_n20743_));
  AND2X1   g20551(.A(new_n20743_), .B(new_n20740_), .Y(new_n20744_));
  INVX1    g20552(.A(new_n20744_), .Y(new_n20745_));
  NAND3X1  g20553(.A(new_n20736_), .B(new_n20726_), .C(new_n17927_), .Y(new_n20746_));
  AOI21X1  g20554(.A0(new_n20746_), .A1(new_n20745_), .B0(new_n20737_), .Y(new_n20747_));
  OR2X1    g20555(.A(new_n20747_), .B(new_n17262_), .Y(new_n20748_));
  OR2X1    g20556(.A(new_n20734_), .B(new_n19273_), .Y(new_n20749_));
  AND2X1   g20557(.A(new_n20713_), .B(new_n20710_), .Y(new_n20750_));
  OR2X1    g20558(.A(new_n20715_), .B(\asqrt[9] ), .Y(new_n20751_));
  OR2X1    g20559(.A(new_n20723_), .B(new_n20721_), .Y(new_n20752_));
  OAI21X1  g20560(.A0(new_n20751_), .A1(new_n20750_), .B0(new_n20752_), .Y(new_n20753_));
  AOI21X1  g20561(.A0(new_n20753_), .A1(new_n20749_), .B0(new_n18591_), .Y(new_n20754_));
  AOI21X1  g20562(.A0(new_n20708_), .A1(\asqrt[9] ), .B0(\asqrt[10] ), .Y(new_n20755_));
  AOI22X1  g20563(.A0(new_n20755_), .A1(new_n20753_), .B0(new_n20732_), .B1(new_n20729_), .Y(new_n20756_));
  NOR3X1   g20564(.A(new_n20756_), .B(new_n20754_), .C(\asqrt[11] ), .Y(new_n20757_));
  NOR2X1   g20565(.A(new_n20757_), .B(new_n20744_), .Y(new_n20758_));
  NOR3X1   g20566(.A(new_n20051_), .B(new_n20018_), .C(new_n20013_), .Y(new_n20759_));
  NAND3X1  g20567(.A(\asqrt[7] ), .B(new_n20019_), .C(new_n20050_), .Y(new_n20760_));
  AOI22X1  g20568(.A0(new_n20760_), .A1(new_n20018_), .B0(new_n20759_), .B1(\asqrt[7] ), .Y(new_n20761_));
  INVX1    g20569(.A(new_n20761_), .Y(new_n20762_));
  OR2X1    g20570(.A(new_n20737_), .B(\asqrt[12] ), .Y(new_n20763_));
  OAI21X1  g20571(.A0(new_n20763_), .A1(new_n20758_), .B0(new_n20762_), .Y(new_n20764_));
  AOI21X1  g20572(.A0(new_n20764_), .A1(new_n20748_), .B0(new_n16617_), .Y(new_n20765_));
  AOI21X1  g20573(.A0(new_n20066_), .A1(new_n20065_), .B0(new_n20028_), .Y(new_n20766_));
  AND2X1   g20574(.A(new_n20766_), .B(new_n20021_), .Y(new_n20767_));
  AOI22X1  g20575(.A0(new_n20066_), .A1(new_n20065_), .B0(new_n20052_), .B1(\asqrt[12] ), .Y(new_n20768_));
  AOI21X1  g20576(.A0(new_n20768_), .A1(\asqrt[7] ), .B0(new_n20027_), .Y(new_n20769_));
  AOI21X1  g20577(.A0(new_n20767_), .A1(\asqrt[7] ), .B0(new_n20769_), .Y(new_n20770_));
  OAI21X1  g20578(.A0(new_n20756_), .A1(new_n20754_), .B0(\asqrt[11] ), .Y(new_n20771_));
  OAI21X1  g20579(.A0(new_n20757_), .A1(new_n20744_), .B0(new_n20771_), .Y(new_n20772_));
  AOI21X1  g20580(.A0(new_n20772_), .A1(\asqrt[12] ), .B0(\asqrt[13] ), .Y(new_n20773_));
  AOI21X1  g20581(.A0(new_n20773_), .A1(new_n20764_), .B0(new_n20770_), .Y(new_n20774_));
  OAI21X1  g20582(.A0(new_n20774_), .A1(new_n20765_), .B0(\asqrt[14] ), .Y(new_n20775_));
  AND2X1   g20583(.A(new_n20053_), .B(new_n20030_), .Y(new_n20776_));
  NOR3X1   g20584(.A(new_n20776_), .B(new_n20036_), .C(new_n20031_), .Y(new_n20777_));
  NOR3X1   g20585(.A(new_n20676_), .B(new_n20776_), .C(new_n20031_), .Y(new_n20778_));
  NOR2X1   g20586(.A(new_n20778_), .B(new_n20037_), .Y(new_n20779_));
  AOI21X1  g20587(.A0(new_n20777_), .A1(\asqrt[7] ), .B0(new_n20779_), .Y(new_n20780_));
  NOR3X1   g20588(.A(new_n20774_), .B(new_n20765_), .C(\asqrt[14] ), .Y(new_n20781_));
  OAI21X1  g20589(.A0(new_n20781_), .A1(new_n20780_), .B0(new_n20775_), .Y(new_n20782_));
  AND2X1   g20590(.A(new_n20782_), .B(\asqrt[15] ), .Y(new_n20783_));
  OR2X1    g20591(.A(new_n20781_), .B(new_n20780_), .Y(new_n20784_));
  NOR3X1   g20592(.A(new_n20060_), .B(new_n20063_), .C(new_n20078_), .Y(new_n20785_));
  NOR3X1   g20593(.A(new_n20676_), .B(new_n20060_), .C(new_n20078_), .Y(new_n20786_));
  NOR2X1   g20594(.A(new_n20786_), .B(new_n20059_), .Y(new_n20787_));
  AOI21X1  g20595(.A0(new_n20785_), .A1(\asqrt[7] ), .B0(new_n20787_), .Y(new_n20788_));
  AND2X1   g20596(.A(new_n20775_), .B(new_n15362_), .Y(new_n20789_));
  AOI21X1  g20597(.A0(new_n20789_), .A1(new_n20784_), .B0(new_n20788_), .Y(new_n20790_));
  OAI21X1  g20598(.A0(new_n20790_), .A1(new_n20783_), .B0(\asqrt[16] ), .Y(new_n20791_));
  AND2X1   g20599(.A(new_n20079_), .B(new_n20072_), .Y(new_n20792_));
  NOR3X1   g20600(.A(new_n20792_), .B(new_n20117_), .C(new_n20062_), .Y(new_n20793_));
  NOR3X1   g20601(.A(new_n20676_), .B(new_n20792_), .C(new_n20062_), .Y(new_n20794_));
  NOR2X1   g20602(.A(new_n20794_), .B(new_n20077_), .Y(new_n20795_));
  AOI21X1  g20603(.A0(new_n20793_), .A1(\asqrt[7] ), .B0(new_n20795_), .Y(new_n20796_));
  INVX1    g20604(.A(new_n20796_), .Y(new_n20797_));
  AND2X1   g20605(.A(new_n20772_), .B(\asqrt[12] ), .Y(new_n20798_));
  OR2X1    g20606(.A(new_n20757_), .B(new_n20744_), .Y(new_n20799_));
  NOR2X1   g20607(.A(new_n20737_), .B(\asqrt[12] ), .Y(new_n20800_));
  AOI21X1  g20608(.A0(new_n20800_), .A1(new_n20799_), .B0(new_n20761_), .Y(new_n20801_));
  OAI21X1  g20609(.A0(new_n20801_), .A1(new_n20798_), .B0(\asqrt[13] ), .Y(new_n20802_));
  INVX1    g20610(.A(new_n20770_), .Y(new_n20803_));
  OAI21X1  g20611(.A0(new_n20747_), .A1(new_n17262_), .B0(new_n16617_), .Y(new_n20804_));
  OAI21X1  g20612(.A0(new_n20804_), .A1(new_n20801_), .B0(new_n20803_), .Y(new_n20805_));
  AOI21X1  g20613(.A0(new_n20805_), .A1(new_n20802_), .B0(new_n15990_), .Y(new_n20806_));
  INVX1    g20614(.A(new_n20780_), .Y(new_n20807_));
  NAND3X1  g20615(.A(new_n20805_), .B(new_n20802_), .C(new_n15990_), .Y(new_n20808_));
  AOI21X1  g20616(.A0(new_n20808_), .A1(new_n20807_), .B0(new_n20806_), .Y(new_n20809_));
  OAI21X1  g20617(.A0(new_n20809_), .A1(new_n15362_), .B0(new_n14754_), .Y(new_n20810_));
  OAI21X1  g20618(.A0(new_n20810_), .A1(new_n20790_), .B0(new_n20797_), .Y(new_n20811_));
  AOI21X1  g20619(.A0(new_n20811_), .A1(new_n20791_), .B0(new_n14165_), .Y(new_n20812_));
  AND2X1   g20620(.A(new_n20121_), .B(new_n20119_), .Y(new_n20813_));
  NOR3X1   g20621(.A(new_n20813_), .B(new_n20087_), .C(new_n20120_), .Y(new_n20814_));
  NOR3X1   g20622(.A(new_n20676_), .B(new_n20813_), .C(new_n20120_), .Y(new_n20815_));
  NOR2X1   g20623(.A(new_n20815_), .B(new_n20086_), .Y(new_n20816_));
  AOI21X1  g20624(.A0(new_n20814_), .A1(\asqrt[7] ), .B0(new_n20816_), .Y(new_n20817_));
  INVX1    g20625(.A(new_n20817_), .Y(new_n20818_));
  NAND3X1  g20626(.A(new_n20811_), .B(new_n20791_), .C(new_n14165_), .Y(new_n20819_));
  AOI21X1  g20627(.A0(new_n20819_), .A1(new_n20818_), .B0(new_n20812_), .Y(new_n20820_));
  OR2X1    g20628(.A(new_n20820_), .B(new_n13571_), .Y(new_n20821_));
  OR2X1    g20629(.A(new_n20809_), .B(new_n15362_), .Y(new_n20822_));
  NOR2X1   g20630(.A(new_n20781_), .B(new_n20780_), .Y(new_n20823_));
  INVX1    g20631(.A(new_n20788_), .Y(new_n20824_));
  NAND2X1  g20632(.A(new_n20775_), .B(new_n15362_), .Y(new_n20825_));
  OAI21X1  g20633(.A0(new_n20825_), .A1(new_n20823_), .B0(new_n20824_), .Y(new_n20826_));
  AOI21X1  g20634(.A0(new_n20826_), .A1(new_n20822_), .B0(new_n14754_), .Y(new_n20827_));
  AOI21X1  g20635(.A0(new_n20782_), .A1(\asqrt[15] ), .B0(\asqrt[16] ), .Y(new_n20828_));
  AOI21X1  g20636(.A0(new_n20828_), .A1(new_n20826_), .B0(new_n20796_), .Y(new_n20829_));
  NOR3X1   g20637(.A(new_n20829_), .B(new_n20827_), .C(\asqrt[17] ), .Y(new_n20830_));
  NOR2X1   g20638(.A(new_n20830_), .B(new_n20817_), .Y(new_n20831_));
  NAND4X1  g20639(.A(\asqrt[7] ), .B(new_n20097_), .C(new_n20095_), .D(new_n20123_), .Y(new_n20832_));
  NAND2X1  g20640(.A(new_n20097_), .B(new_n20123_), .Y(new_n20833_));
  OAI21X1  g20641(.A0(new_n20833_), .A1(new_n20676_), .B0(new_n20096_), .Y(new_n20834_));
  AND2X1   g20642(.A(new_n20834_), .B(new_n20832_), .Y(new_n20835_));
  INVX1    g20643(.A(new_n20835_), .Y(new_n20836_));
  OAI21X1  g20644(.A0(new_n20829_), .A1(new_n20827_), .B0(\asqrt[17] ), .Y(new_n20837_));
  NAND2X1  g20645(.A(new_n20837_), .B(new_n13571_), .Y(new_n20838_));
  OAI21X1  g20646(.A0(new_n20838_), .A1(new_n20831_), .B0(new_n20836_), .Y(new_n20839_));
  AOI21X1  g20647(.A0(new_n20839_), .A1(new_n20821_), .B0(new_n13000_), .Y(new_n20840_));
  AOI21X1  g20648(.A0(new_n20139_), .A1(new_n20138_), .B0(new_n20106_), .Y(new_n20841_));
  AND2X1   g20649(.A(new_n20841_), .B(new_n20099_), .Y(new_n20842_));
  AOI22X1  g20650(.A0(new_n20139_), .A1(new_n20138_), .B0(new_n20125_), .B1(\asqrt[18] ), .Y(new_n20843_));
  AOI21X1  g20651(.A0(new_n20843_), .A1(\asqrt[7] ), .B0(new_n20105_), .Y(new_n20844_));
  AOI21X1  g20652(.A0(new_n20842_), .A1(\asqrt[7] ), .B0(new_n20844_), .Y(new_n20845_));
  OAI21X1  g20653(.A0(new_n20830_), .A1(new_n20817_), .B0(new_n20837_), .Y(new_n20846_));
  AOI21X1  g20654(.A0(new_n20846_), .A1(\asqrt[18] ), .B0(\asqrt[19] ), .Y(new_n20847_));
  AOI21X1  g20655(.A0(new_n20847_), .A1(new_n20839_), .B0(new_n20845_), .Y(new_n20848_));
  OAI21X1  g20656(.A0(new_n20848_), .A1(new_n20840_), .B0(\asqrt[20] ), .Y(new_n20849_));
  AND2X1   g20657(.A(new_n20126_), .B(new_n20108_), .Y(new_n20850_));
  NOR3X1   g20658(.A(new_n20850_), .B(new_n20142_), .C(new_n20109_), .Y(new_n20851_));
  NOR3X1   g20659(.A(new_n20676_), .B(new_n20850_), .C(new_n20109_), .Y(new_n20852_));
  NOR2X1   g20660(.A(new_n20852_), .B(new_n20114_), .Y(new_n20853_));
  AOI21X1  g20661(.A0(new_n20851_), .A1(\asqrt[7] ), .B0(new_n20853_), .Y(new_n20854_));
  NOR3X1   g20662(.A(new_n20848_), .B(new_n20840_), .C(\asqrt[20] ), .Y(new_n20855_));
  OAI21X1  g20663(.A0(new_n20855_), .A1(new_n20854_), .B0(new_n20849_), .Y(new_n20856_));
  AND2X1   g20664(.A(new_n20856_), .B(\asqrt[21] ), .Y(new_n20857_));
  INVX1    g20665(.A(new_n20854_), .Y(new_n20858_));
  AND2X1   g20666(.A(new_n20846_), .B(\asqrt[18] ), .Y(new_n20859_));
  OR2X1    g20667(.A(new_n20830_), .B(new_n20817_), .Y(new_n20860_));
  AND2X1   g20668(.A(new_n20837_), .B(new_n13571_), .Y(new_n20861_));
  AOI21X1  g20669(.A0(new_n20861_), .A1(new_n20860_), .B0(new_n20835_), .Y(new_n20862_));
  OAI21X1  g20670(.A0(new_n20862_), .A1(new_n20859_), .B0(\asqrt[19] ), .Y(new_n20863_));
  INVX1    g20671(.A(new_n20845_), .Y(new_n20864_));
  OAI21X1  g20672(.A0(new_n20820_), .A1(new_n13571_), .B0(new_n13000_), .Y(new_n20865_));
  OAI21X1  g20673(.A0(new_n20865_), .A1(new_n20862_), .B0(new_n20864_), .Y(new_n20866_));
  NAND3X1  g20674(.A(new_n20866_), .B(new_n20863_), .C(new_n12447_), .Y(new_n20867_));
  NAND2X1  g20675(.A(new_n20867_), .B(new_n20858_), .Y(new_n20868_));
  NAND4X1  g20676(.A(\asqrt[7] ), .B(new_n20145_), .C(new_n20132_), .D(new_n20128_), .Y(new_n20869_));
  NAND2X1  g20677(.A(new_n20145_), .B(new_n20128_), .Y(new_n20870_));
  OAI21X1  g20678(.A0(new_n20870_), .A1(new_n20676_), .B0(new_n20136_), .Y(new_n20871_));
  AND2X1   g20679(.A(new_n20871_), .B(new_n20869_), .Y(new_n20872_));
  AOI21X1  g20680(.A0(new_n20866_), .A1(new_n20863_), .B0(new_n12447_), .Y(new_n20873_));
  NOR2X1   g20681(.A(new_n20873_), .B(\asqrt[21] ), .Y(new_n20874_));
  AOI21X1  g20682(.A0(new_n20874_), .A1(new_n20868_), .B0(new_n20872_), .Y(new_n20875_));
  OAI21X1  g20683(.A0(new_n20875_), .A1(new_n20857_), .B0(\asqrt[22] ), .Y(new_n20876_));
  AND2X1   g20684(.A(new_n20153_), .B(new_n20146_), .Y(new_n20877_));
  NOR3X1   g20685(.A(new_n20877_), .B(new_n20191_), .C(new_n20135_), .Y(new_n20878_));
  NOR3X1   g20686(.A(new_n20676_), .B(new_n20877_), .C(new_n20135_), .Y(new_n20879_));
  NOR2X1   g20687(.A(new_n20879_), .B(new_n20151_), .Y(new_n20880_));
  AOI21X1  g20688(.A0(new_n20878_), .A1(\asqrt[7] ), .B0(new_n20880_), .Y(new_n20881_));
  INVX1    g20689(.A(new_n20881_), .Y(new_n20882_));
  AOI21X1  g20690(.A0(new_n20867_), .A1(new_n20858_), .B0(new_n20873_), .Y(new_n20883_));
  OAI21X1  g20691(.A0(new_n20883_), .A1(new_n11896_), .B0(new_n11362_), .Y(new_n20884_));
  OAI21X1  g20692(.A0(new_n20884_), .A1(new_n20875_), .B0(new_n20882_), .Y(new_n20885_));
  AOI21X1  g20693(.A0(new_n20885_), .A1(new_n20876_), .B0(new_n10849_), .Y(new_n20886_));
  AND2X1   g20694(.A(new_n20195_), .B(new_n20193_), .Y(new_n20887_));
  NOR3X1   g20695(.A(new_n20887_), .B(new_n20161_), .C(new_n20194_), .Y(new_n20888_));
  NOR3X1   g20696(.A(new_n20676_), .B(new_n20887_), .C(new_n20194_), .Y(new_n20889_));
  NOR2X1   g20697(.A(new_n20889_), .B(new_n20160_), .Y(new_n20890_));
  AOI21X1  g20698(.A0(new_n20888_), .A1(\asqrt[7] ), .B0(new_n20890_), .Y(new_n20891_));
  INVX1    g20699(.A(new_n20891_), .Y(new_n20892_));
  NAND3X1  g20700(.A(new_n20885_), .B(new_n20876_), .C(new_n10849_), .Y(new_n20893_));
  AOI21X1  g20701(.A0(new_n20893_), .A1(new_n20892_), .B0(new_n20886_), .Y(new_n20894_));
  OR2X1    g20702(.A(new_n20894_), .B(new_n10332_), .Y(new_n20895_));
  AND2X1   g20703(.A(new_n20893_), .B(new_n20892_), .Y(new_n20896_));
  NAND4X1  g20704(.A(\asqrt[7] ), .B(new_n20171_), .C(new_n20169_), .D(new_n20197_), .Y(new_n20897_));
  NAND2X1  g20705(.A(new_n20171_), .B(new_n20197_), .Y(new_n20898_));
  OAI21X1  g20706(.A0(new_n20898_), .A1(new_n20676_), .B0(new_n20170_), .Y(new_n20899_));
  AND2X1   g20707(.A(new_n20899_), .B(new_n20897_), .Y(new_n20900_));
  INVX1    g20708(.A(new_n20900_), .Y(new_n20901_));
  OR2X1    g20709(.A(new_n20886_), .B(\asqrt[24] ), .Y(new_n20902_));
  OAI21X1  g20710(.A0(new_n20902_), .A1(new_n20896_), .B0(new_n20901_), .Y(new_n20903_));
  AOI21X1  g20711(.A0(new_n20903_), .A1(new_n20895_), .B0(new_n9833_), .Y(new_n20904_));
  AOI21X1  g20712(.A0(new_n20227_), .A1(new_n20226_), .B0(new_n20180_), .Y(new_n20905_));
  AND2X1   g20713(.A(new_n20905_), .B(new_n20173_), .Y(new_n20906_));
  AOI22X1  g20714(.A0(new_n20227_), .A1(new_n20226_), .B0(new_n20199_), .B1(\asqrt[24] ), .Y(new_n20907_));
  AOI21X1  g20715(.A0(new_n20907_), .A1(\asqrt[7] ), .B0(new_n20179_), .Y(new_n20908_));
  AOI21X1  g20716(.A0(new_n20906_), .A1(\asqrt[7] ), .B0(new_n20908_), .Y(new_n20909_));
  OR2X1    g20717(.A(new_n20883_), .B(new_n11896_), .Y(new_n20910_));
  AND2X1   g20718(.A(new_n20867_), .B(new_n20858_), .Y(new_n20911_));
  INVX1    g20719(.A(new_n20872_), .Y(new_n20912_));
  OR2X1    g20720(.A(new_n20873_), .B(\asqrt[21] ), .Y(new_n20913_));
  OAI21X1  g20721(.A0(new_n20913_), .A1(new_n20911_), .B0(new_n20912_), .Y(new_n20914_));
  AOI21X1  g20722(.A0(new_n20914_), .A1(new_n20910_), .B0(new_n11362_), .Y(new_n20915_));
  AOI21X1  g20723(.A0(new_n20856_), .A1(\asqrt[21] ), .B0(\asqrt[22] ), .Y(new_n20916_));
  AOI21X1  g20724(.A0(new_n20916_), .A1(new_n20914_), .B0(new_n20881_), .Y(new_n20917_));
  OAI21X1  g20725(.A0(new_n20917_), .A1(new_n20915_), .B0(\asqrt[23] ), .Y(new_n20918_));
  NOR3X1   g20726(.A(new_n20917_), .B(new_n20915_), .C(\asqrt[23] ), .Y(new_n20919_));
  OAI21X1  g20727(.A0(new_n20919_), .A1(new_n20891_), .B0(new_n20918_), .Y(new_n20920_));
  AOI21X1  g20728(.A0(new_n20920_), .A1(\asqrt[24] ), .B0(\asqrt[25] ), .Y(new_n20921_));
  AOI21X1  g20729(.A0(new_n20921_), .A1(new_n20903_), .B0(new_n20909_), .Y(new_n20922_));
  OAI21X1  g20730(.A0(new_n20922_), .A1(new_n20904_), .B0(\asqrt[26] ), .Y(new_n20923_));
  AND2X1   g20731(.A(new_n20200_), .B(new_n20182_), .Y(new_n20924_));
  NOR3X1   g20732(.A(new_n20924_), .B(new_n20230_), .C(new_n20183_), .Y(new_n20925_));
  NOR3X1   g20733(.A(new_n20676_), .B(new_n20924_), .C(new_n20183_), .Y(new_n20926_));
  NOR2X1   g20734(.A(new_n20926_), .B(new_n20188_), .Y(new_n20927_));
  AOI21X1  g20735(.A0(new_n20925_), .A1(\asqrt[7] ), .B0(new_n20927_), .Y(new_n20928_));
  NOR3X1   g20736(.A(new_n20922_), .B(new_n20904_), .C(\asqrt[26] ), .Y(new_n20929_));
  OAI21X1  g20737(.A0(new_n20929_), .A1(new_n20928_), .B0(new_n20923_), .Y(new_n20930_));
  AND2X1   g20738(.A(new_n20930_), .B(\asqrt[27] ), .Y(new_n20931_));
  OR2X1    g20739(.A(new_n20929_), .B(new_n20928_), .Y(new_n20932_));
  OR4X1    g20740(.A(new_n20676_), .B(new_n20207_), .C(new_n20234_), .D(new_n20233_), .Y(new_n20933_));
  OR2X1    g20741(.A(new_n20207_), .B(new_n20233_), .Y(new_n20934_));
  OAI21X1  g20742(.A0(new_n20934_), .A1(new_n20676_), .B0(new_n20234_), .Y(new_n20935_));
  AND2X1   g20743(.A(new_n20935_), .B(new_n20933_), .Y(new_n20936_));
  AND2X1   g20744(.A(new_n20923_), .B(new_n8874_), .Y(new_n20937_));
  AOI21X1  g20745(.A0(new_n20937_), .A1(new_n20932_), .B0(new_n20936_), .Y(new_n20938_));
  OAI21X1  g20746(.A0(new_n20938_), .A1(new_n20931_), .B0(\asqrt[28] ), .Y(new_n20939_));
  AND2X1   g20747(.A(new_n20216_), .B(new_n20210_), .Y(new_n20940_));
  NOR3X1   g20748(.A(new_n20940_), .B(new_n20250_), .C(new_n20209_), .Y(new_n20941_));
  NOR3X1   g20749(.A(new_n20676_), .B(new_n20940_), .C(new_n20209_), .Y(new_n20942_));
  NOR2X1   g20750(.A(new_n20942_), .B(new_n20215_), .Y(new_n20943_));
  AOI21X1  g20751(.A0(new_n20941_), .A1(\asqrt[7] ), .B0(new_n20943_), .Y(new_n20944_));
  INVX1    g20752(.A(new_n20944_), .Y(new_n20945_));
  AND2X1   g20753(.A(new_n20920_), .B(\asqrt[24] ), .Y(new_n20946_));
  NAND2X1  g20754(.A(new_n20893_), .B(new_n20892_), .Y(new_n20947_));
  NOR2X1   g20755(.A(new_n20886_), .B(\asqrt[24] ), .Y(new_n20948_));
  AOI21X1  g20756(.A0(new_n20948_), .A1(new_n20947_), .B0(new_n20900_), .Y(new_n20949_));
  OAI21X1  g20757(.A0(new_n20949_), .A1(new_n20946_), .B0(\asqrt[25] ), .Y(new_n20950_));
  INVX1    g20758(.A(new_n20909_), .Y(new_n20951_));
  OAI21X1  g20759(.A0(new_n20894_), .A1(new_n10332_), .B0(new_n9833_), .Y(new_n20952_));
  OAI21X1  g20760(.A0(new_n20952_), .A1(new_n20949_), .B0(new_n20951_), .Y(new_n20953_));
  AOI21X1  g20761(.A0(new_n20953_), .A1(new_n20950_), .B0(new_n9353_), .Y(new_n20954_));
  INVX1    g20762(.A(new_n20928_), .Y(new_n20955_));
  NAND3X1  g20763(.A(new_n20953_), .B(new_n20950_), .C(new_n9353_), .Y(new_n20956_));
  AOI21X1  g20764(.A0(new_n20956_), .A1(new_n20955_), .B0(new_n20954_), .Y(new_n20957_));
  OAI21X1  g20765(.A0(new_n20957_), .A1(new_n8874_), .B0(new_n8412_), .Y(new_n20958_));
  OAI21X1  g20766(.A0(new_n20958_), .A1(new_n20938_), .B0(new_n20945_), .Y(new_n20959_));
  AOI21X1  g20767(.A0(new_n20959_), .A1(new_n20939_), .B0(new_n7970_), .Y(new_n20960_));
  AND2X1   g20768(.A(new_n20254_), .B(new_n20252_), .Y(new_n20961_));
  NOR3X1   g20769(.A(new_n20961_), .B(new_n20224_), .C(new_n20253_), .Y(new_n20962_));
  NOR3X1   g20770(.A(new_n20676_), .B(new_n20961_), .C(new_n20253_), .Y(new_n20963_));
  NOR2X1   g20771(.A(new_n20963_), .B(new_n20223_), .Y(new_n20964_));
  AOI21X1  g20772(.A0(new_n20962_), .A1(\asqrt[7] ), .B0(new_n20964_), .Y(new_n20965_));
  INVX1    g20773(.A(new_n20965_), .Y(new_n20966_));
  NAND3X1  g20774(.A(new_n20959_), .B(new_n20939_), .C(new_n7970_), .Y(new_n20967_));
  AOI21X1  g20775(.A0(new_n20967_), .A1(new_n20966_), .B0(new_n20960_), .Y(new_n20968_));
  OR2X1    g20776(.A(new_n20968_), .B(new_n7527_), .Y(new_n20969_));
  OR2X1    g20777(.A(new_n20957_), .B(new_n8874_), .Y(new_n20970_));
  NOR2X1   g20778(.A(new_n20929_), .B(new_n20928_), .Y(new_n20971_));
  INVX1    g20779(.A(new_n20936_), .Y(new_n20972_));
  NAND2X1  g20780(.A(new_n20923_), .B(new_n8874_), .Y(new_n20973_));
  OAI21X1  g20781(.A0(new_n20973_), .A1(new_n20971_), .B0(new_n20972_), .Y(new_n20974_));
  AOI21X1  g20782(.A0(new_n20974_), .A1(new_n20970_), .B0(new_n8412_), .Y(new_n20975_));
  AOI21X1  g20783(.A0(new_n20930_), .A1(\asqrt[27] ), .B0(\asqrt[28] ), .Y(new_n20976_));
  AOI21X1  g20784(.A0(new_n20976_), .A1(new_n20974_), .B0(new_n20944_), .Y(new_n20977_));
  NOR3X1   g20785(.A(new_n20977_), .B(new_n20975_), .C(\asqrt[29] ), .Y(new_n20978_));
  NOR2X1   g20786(.A(new_n20978_), .B(new_n20965_), .Y(new_n20979_));
  OR4X1    g20787(.A(new_n20676_), .B(new_n20256_), .C(new_n20244_), .D(new_n20239_), .Y(new_n20980_));
  OR2X1    g20788(.A(new_n20256_), .B(new_n20239_), .Y(new_n20981_));
  OAI21X1  g20789(.A0(new_n20981_), .A1(new_n20676_), .B0(new_n20244_), .Y(new_n20982_));
  AND2X1   g20790(.A(new_n20982_), .B(new_n20980_), .Y(new_n20983_));
  INVX1    g20791(.A(new_n20983_), .Y(new_n20984_));
  OAI21X1  g20792(.A0(new_n20977_), .A1(new_n20975_), .B0(\asqrt[29] ), .Y(new_n20985_));
  NAND2X1  g20793(.A(new_n20985_), .B(new_n7527_), .Y(new_n20986_));
  OAI21X1  g20794(.A0(new_n20986_), .A1(new_n20979_), .B0(new_n20984_), .Y(new_n20987_));
  AOI21X1  g20795(.A0(new_n20987_), .A1(new_n20969_), .B0(new_n7103_), .Y(new_n20988_));
  AOI21X1  g20796(.A0(new_n20301_), .A1(new_n20300_), .B0(new_n20263_), .Y(new_n20989_));
  AND2X1   g20797(.A(new_n20989_), .B(new_n20247_), .Y(new_n20990_));
  AOI22X1  g20798(.A0(new_n20301_), .A1(new_n20300_), .B0(new_n20273_), .B1(\asqrt[30] ), .Y(new_n20991_));
  AOI21X1  g20799(.A0(new_n20991_), .A1(\asqrt[7] ), .B0(new_n20262_), .Y(new_n20992_));
  AOI21X1  g20800(.A0(new_n20990_), .A1(\asqrt[7] ), .B0(new_n20992_), .Y(new_n20993_));
  OAI21X1  g20801(.A0(new_n20978_), .A1(new_n20965_), .B0(new_n20985_), .Y(new_n20994_));
  AOI21X1  g20802(.A0(new_n20994_), .A1(\asqrt[30] ), .B0(\asqrt[31] ), .Y(new_n20995_));
  AOI21X1  g20803(.A0(new_n20995_), .A1(new_n20987_), .B0(new_n20993_), .Y(new_n20996_));
  OAI21X1  g20804(.A0(new_n20996_), .A1(new_n20988_), .B0(\asqrt[32] ), .Y(new_n20997_));
  AND2X1   g20805(.A(new_n20274_), .B(new_n20266_), .Y(new_n20998_));
  NOR3X1   g20806(.A(new_n20998_), .B(new_n20304_), .C(new_n20267_), .Y(new_n20999_));
  NOR3X1   g20807(.A(new_n20676_), .B(new_n20998_), .C(new_n20267_), .Y(new_n21000_));
  NOR2X1   g20808(.A(new_n21000_), .B(new_n20272_), .Y(new_n21001_));
  AOI21X1  g20809(.A0(new_n20999_), .A1(\asqrt[7] ), .B0(new_n21001_), .Y(new_n21002_));
  NOR3X1   g20810(.A(new_n20996_), .B(new_n20988_), .C(\asqrt[32] ), .Y(new_n21003_));
  OAI21X1  g20811(.A0(new_n21003_), .A1(new_n21002_), .B0(new_n20997_), .Y(new_n21004_));
  AND2X1   g20812(.A(new_n21004_), .B(\asqrt[33] ), .Y(new_n21005_));
  OR2X1    g20813(.A(new_n21003_), .B(new_n21002_), .Y(new_n21006_));
  OR4X1    g20814(.A(new_n20676_), .B(new_n20281_), .C(new_n20308_), .D(new_n20307_), .Y(new_n21007_));
  OR2X1    g20815(.A(new_n20281_), .B(new_n20307_), .Y(new_n21008_));
  OAI21X1  g20816(.A0(new_n21008_), .A1(new_n20676_), .B0(new_n20308_), .Y(new_n21009_));
  AND2X1   g20817(.A(new_n21009_), .B(new_n21007_), .Y(new_n21010_));
  AND2X1   g20818(.A(new_n20997_), .B(new_n6294_), .Y(new_n21011_));
  AOI21X1  g20819(.A0(new_n21011_), .A1(new_n21006_), .B0(new_n21010_), .Y(new_n21012_));
  OAI21X1  g20820(.A0(new_n21012_), .A1(new_n21005_), .B0(\asqrt[34] ), .Y(new_n21013_));
  AND2X1   g20821(.A(new_n20290_), .B(new_n20284_), .Y(new_n21014_));
  NOR3X1   g20822(.A(new_n21014_), .B(new_n20324_), .C(new_n20283_), .Y(new_n21015_));
  NOR3X1   g20823(.A(new_n20676_), .B(new_n21014_), .C(new_n20283_), .Y(new_n21016_));
  NOR2X1   g20824(.A(new_n21016_), .B(new_n20289_), .Y(new_n21017_));
  AOI21X1  g20825(.A0(new_n21015_), .A1(\asqrt[7] ), .B0(new_n21017_), .Y(new_n21018_));
  INVX1    g20826(.A(new_n21018_), .Y(new_n21019_));
  AND2X1   g20827(.A(new_n20994_), .B(\asqrt[30] ), .Y(new_n21020_));
  OR2X1    g20828(.A(new_n20978_), .B(new_n20965_), .Y(new_n21021_));
  AND2X1   g20829(.A(new_n20985_), .B(new_n7527_), .Y(new_n21022_));
  AOI21X1  g20830(.A0(new_n21022_), .A1(new_n21021_), .B0(new_n20983_), .Y(new_n21023_));
  OAI21X1  g20831(.A0(new_n21023_), .A1(new_n21020_), .B0(\asqrt[31] ), .Y(new_n21024_));
  INVX1    g20832(.A(new_n20993_), .Y(new_n21025_));
  OAI21X1  g20833(.A0(new_n20968_), .A1(new_n7527_), .B0(new_n7103_), .Y(new_n21026_));
  OAI21X1  g20834(.A0(new_n21026_), .A1(new_n21023_), .B0(new_n21025_), .Y(new_n21027_));
  AOI21X1  g20835(.A0(new_n21027_), .A1(new_n21024_), .B0(new_n6699_), .Y(new_n21028_));
  INVX1    g20836(.A(new_n21002_), .Y(new_n21029_));
  NAND3X1  g20837(.A(new_n21027_), .B(new_n21024_), .C(new_n6699_), .Y(new_n21030_));
  AOI21X1  g20838(.A0(new_n21030_), .A1(new_n21029_), .B0(new_n21028_), .Y(new_n21031_));
  OAI21X1  g20839(.A0(new_n21031_), .A1(new_n6294_), .B0(new_n5941_), .Y(new_n21032_));
  OAI21X1  g20840(.A0(new_n21032_), .A1(new_n21012_), .B0(new_n21019_), .Y(new_n21033_));
  AOI21X1  g20841(.A0(new_n21033_), .A1(new_n21013_), .B0(new_n5541_), .Y(new_n21034_));
  AND2X1   g20842(.A(new_n20328_), .B(new_n20326_), .Y(new_n21035_));
  NOR3X1   g20843(.A(new_n21035_), .B(new_n20298_), .C(new_n20327_), .Y(new_n21036_));
  NOR3X1   g20844(.A(new_n20676_), .B(new_n21035_), .C(new_n20327_), .Y(new_n21037_));
  NOR2X1   g20845(.A(new_n21037_), .B(new_n20297_), .Y(new_n21038_));
  AOI21X1  g20846(.A0(new_n21036_), .A1(\asqrt[7] ), .B0(new_n21038_), .Y(new_n21039_));
  INVX1    g20847(.A(new_n21039_), .Y(new_n21040_));
  NAND3X1  g20848(.A(new_n21033_), .B(new_n21013_), .C(new_n5541_), .Y(new_n21041_));
  AOI21X1  g20849(.A0(new_n21041_), .A1(new_n21040_), .B0(new_n21034_), .Y(new_n21042_));
  OR2X1    g20850(.A(new_n21042_), .B(new_n5176_), .Y(new_n21043_));
  OR2X1    g20851(.A(new_n21031_), .B(new_n6294_), .Y(new_n21044_));
  NOR2X1   g20852(.A(new_n21003_), .B(new_n21002_), .Y(new_n21045_));
  INVX1    g20853(.A(new_n21010_), .Y(new_n21046_));
  NAND2X1  g20854(.A(new_n20997_), .B(new_n6294_), .Y(new_n21047_));
  OAI21X1  g20855(.A0(new_n21047_), .A1(new_n21045_), .B0(new_n21046_), .Y(new_n21048_));
  AOI21X1  g20856(.A0(new_n21048_), .A1(new_n21044_), .B0(new_n5941_), .Y(new_n21049_));
  AOI21X1  g20857(.A0(new_n21004_), .A1(\asqrt[33] ), .B0(\asqrt[34] ), .Y(new_n21050_));
  AOI21X1  g20858(.A0(new_n21050_), .A1(new_n21048_), .B0(new_n21018_), .Y(new_n21051_));
  NOR3X1   g20859(.A(new_n21051_), .B(new_n21049_), .C(\asqrt[35] ), .Y(new_n21052_));
  NOR2X1   g20860(.A(new_n21052_), .B(new_n21039_), .Y(new_n21053_));
  OR4X1    g20861(.A(new_n20676_), .B(new_n20330_), .C(new_n20318_), .D(new_n20313_), .Y(new_n21054_));
  OR2X1    g20862(.A(new_n20330_), .B(new_n20313_), .Y(new_n21055_));
  OAI21X1  g20863(.A0(new_n21055_), .A1(new_n20676_), .B0(new_n20318_), .Y(new_n21056_));
  AND2X1   g20864(.A(new_n21056_), .B(new_n21054_), .Y(new_n21057_));
  INVX1    g20865(.A(new_n21057_), .Y(new_n21058_));
  OAI21X1  g20866(.A0(new_n21051_), .A1(new_n21049_), .B0(\asqrt[35] ), .Y(new_n21059_));
  NAND2X1  g20867(.A(new_n21059_), .B(new_n5176_), .Y(new_n21060_));
  OAI21X1  g20868(.A0(new_n21060_), .A1(new_n21053_), .B0(new_n21058_), .Y(new_n21061_));
  AOI21X1  g20869(.A0(new_n21061_), .A1(new_n21043_), .B0(new_n4826_), .Y(new_n21062_));
  AOI21X1  g20870(.A0(new_n20375_), .A1(new_n20374_), .B0(new_n20337_), .Y(new_n21063_));
  AND2X1   g20871(.A(new_n21063_), .B(new_n20321_), .Y(new_n21064_));
  AOI22X1  g20872(.A0(new_n20375_), .A1(new_n20374_), .B0(new_n20347_), .B1(\asqrt[36] ), .Y(new_n21065_));
  AOI21X1  g20873(.A0(new_n21065_), .A1(\asqrt[7] ), .B0(new_n20336_), .Y(new_n21066_));
  AOI21X1  g20874(.A0(new_n21064_), .A1(\asqrt[7] ), .B0(new_n21066_), .Y(new_n21067_));
  OAI21X1  g20875(.A0(new_n21052_), .A1(new_n21039_), .B0(new_n21059_), .Y(new_n21068_));
  AOI21X1  g20876(.A0(new_n21068_), .A1(\asqrt[36] ), .B0(\asqrt[37] ), .Y(new_n21069_));
  AOI21X1  g20877(.A0(new_n21069_), .A1(new_n21061_), .B0(new_n21067_), .Y(new_n21070_));
  OAI21X1  g20878(.A0(new_n21070_), .A1(new_n21062_), .B0(\asqrt[38] ), .Y(new_n21071_));
  AND2X1   g20879(.A(new_n20348_), .B(new_n20340_), .Y(new_n21072_));
  NOR3X1   g20880(.A(new_n21072_), .B(new_n20378_), .C(new_n20341_), .Y(new_n21073_));
  NOR3X1   g20881(.A(new_n20676_), .B(new_n21072_), .C(new_n20341_), .Y(new_n21074_));
  NOR2X1   g20882(.A(new_n21074_), .B(new_n20346_), .Y(new_n21075_));
  AOI21X1  g20883(.A0(new_n21073_), .A1(\asqrt[7] ), .B0(new_n21075_), .Y(new_n21076_));
  NOR3X1   g20884(.A(new_n21070_), .B(new_n21062_), .C(\asqrt[38] ), .Y(new_n21077_));
  OAI21X1  g20885(.A0(new_n21077_), .A1(new_n21076_), .B0(new_n21071_), .Y(new_n21078_));
  AND2X1   g20886(.A(new_n21078_), .B(\asqrt[39] ), .Y(new_n21079_));
  OR2X1    g20887(.A(new_n21077_), .B(new_n21076_), .Y(new_n21080_));
  OR4X1    g20888(.A(new_n20676_), .B(new_n20355_), .C(new_n20382_), .D(new_n20381_), .Y(new_n21081_));
  OR2X1    g20889(.A(new_n20355_), .B(new_n20381_), .Y(new_n21082_));
  OAI21X1  g20890(.A0(new_n21082_), .A1(new_n20676_), .B0(new_n20382_), .Y(new_n21083_));
  AND2X1   g20891(.A(new_n21083_), .B(new_n21081_), .Y(new_n21084_));
  AND2X1   g20892(.A(new_n21071_), .B(new_n4165_), .Y(new_n21085_));
  AOI21X1  g20893(.A0(new_n21085_), .A1(new_n21080_), .B0(new_n21084_), .Y(new_n21086_));
  OAI21X1  g20894(.A0(new_n21086_), .A1(new_n21079_), .B0(\asqrt[40] ), .Y(new_n21087_));
  AND2X1   g20895(.A(new_n20364_), .B(new_n20358_), .Y(new_n21088_));
  NOR3X1   g20896(.A(new_n21088_), .B(new_n20398_), .C(new_n20357_), .Y(new_n21089_));
  NOR3X1   g20897(.A(new_n20676_), .B(new_n21088_), .C(new_n20357_), .Y(new_n21090_));
  NOR2X1   g20898(.A(new_n21090_), .B(new_n20363_), .Y(new_n21091_));
  AOI21X1  g20899(.A0(new_n21089_), .A1(\asqrt[7] ), .B0(new_n21091_), .Y(new_n21092_));
  INVX1    g20900(.A(new_n21092_), .Y(new_n21093_));
  AND2X1   g20901(.A(new_n21068_), .B(\asqrt[36] ), .Y(new_n21094_));
  OR2X1    g20902(.A(new_n21052_), .B(new_n21039_), .Y(new_n21095_));
  AND2X1   g20903(.A(new_n21059_), .B(new_n5176_), .Y(new_n21096_));
  AOI21X1  g20904(.A0(new_n21096_), .A1(new_n21095_), .B0(new_n21057_), .Y(new_n21097_));
  OAI21X1  g20905(.A0(new_n21097_), .A1(new_n21094_), .B0(\asqrt[37] ), .Y(new_n21098_));
  INVX1    g20906(.A(new_n21067_), .Y(new_n21099_));
  OAI21X1  g20907(.A0(new_n21042_), .A1(new_n5176_), .B0(new_n4826_), .Y(new_n21100_));
  OAI21X1  g20908(.A0(new_n21100_), .A1(new_n21097_), .B0(new_n21099_), .Y(new_n21101_));
  AOI21X1  g20909(.A0(new_n21101_), .A1(new_n21098_), .B0(new_n4493_), .Y(new_n21102_));
  INVX1    g20910(.A(new_n21076_), .Y(new_n21103_));
  NAND3X1  g20911(.A(new_n21101_), .B(new_n21098_), .C(new_n4493_), .Y(new_n21104_));
  AOI21X1  g20912(.A0(new_n21104_), .A1(new_n21103_), .B0(new_n21102_), .Y(new_n21105_));
  OAI21X1  g20913(.A0(new_n21105_), .A1(new_n4165_), .B0(new_n3863_), .Y(new_n21106_));
  OAI21X1  g20914(.A0(new_n21106_), .A1(new_n21086_), .B0(new_n21093_), .Y(new_n21107_));
  AOI21X1  g20915(.A0(new_n21107_), .A1(new_n21087_), .B0(new_n3564_), .Y(new_n21108_));
  AND2X1   g20916(.A(new_n20402_), .B(new_n20400_), .Y(new_n21109_));
  NOR3X1   g20917(.A(new_n21109_), .B(new_n20372_), .C(new_n20401_), .Y(new_n21110_));
  NOR3X1   g20918(.A(new_n20676_), .B(new_n21109_), .C(new_n20401_), .Y(new_n21111_));
  NOR2X1   g20919(.A(new_n21111_), .B(new_n20371_), .Y(new_n21112_));
  AOI21X1  g20920(.A0(new_n21110_), .A1(\asqrt[7] ), .B0(new_n21112_), .Y(new_n21113_));
  INVX1    g20921(.A(new_n21113_), .Y(new_n21114_));
  NAND3X1  g20922(.A(new_n21107_), .B(new_n21087_), .C(new_n3564_), .Y(new_n21115_));
  AOI21X1  g20923(.A0(new_n21115_), .A1(new_n21114_), .B0(new_n21108_), .Y(new_n21116_));
  OR2X1    g20924(.A(new_n21116_), .B(new_n3276_), .Y(new_n21117_));
  OR2X1    g20925(.A(new_n21105_), .B(new_n4165_), .Y(new_n21118_));
  NOR2X1   g20926(.A(new_n21077_), .B(new_n21076_), .Y(new_n21119_));
  INVX1    g20927(.A(new_n21084_), .Y(new_n21120_));
  NAND2X1  g20928(.A(new_n21071_), .B(new_n4165_), .Y(new_n21121_));
  OAI21X1  g20929(.A0(new_n21121_), .A1(new_n21119_), .B0(new_n21120_), .Y(new_n21122_));
  AOI21X1  g20930(.A0(new_n21122_), .A1(new_n21118_), .B0(new_n3863_), .Y(new_n21123_));
  AOI21X1  g20931(.A0(new_n21078_), .A1(\asqrt[39] ), .B0(\asqrt[40] ), .Y(new_n21124_));
  AOI21X1  g20932(.A0(new_n21124_), .A1(new_n21122_), .B0(new_n21092_), .Y(new_n21125_));
  NOR3X1   g20933(.A(new_n21125_), .B(new_n21123_), .C(\asqrt[41] ), .Y(new_n21126_));
  NOR2X1   g20934(.A(new_n21126_), .B(new_n21113_), .Y(new_n21127_));
  OR4X1    g20935(.A(new_n20676_), .B(new_n20404_), .C(new_n20392_), .D(new_n20387_), .Y(new_n21128_));
  OR2X1    g20936(.A(new_n20404_), .B(new_n20387_), .Y(new_n21129_));
  OAI21X1  g20937(.A0(new_n21129_), .A1(new_n20676_), .B0(new_n20392_), .Y(new_n21130_));
  AND2X1   g20938(.A(new_n21130_), .B(new_n21128_), .Y(new_n21131_));
  INVX1    g20939(.A(new_n21131_), .Y(new_n21132_));
  OAI21X1  g20940(.A0(new_n21125_), .A1(new_n21123_), .B0(\asqrt[41] ), .Y(new_n21133_));
  NAND2X1  g20941(.A(new_n21133_), .B(new_n3276_), .Y(new_n21134_));
  OAI21X1  g20942(.A0(new_n21134_), .A1(new_n21127_), .B0(new_n21132_), .Y(new_n21135_));
  AOI21X1  g20943(.A0(new_n21135_), .A1(new_n21117_), .B0(new_n3008_), .Y(new_n21136_));
  AOI21X1  g20944(.A0(new_n20449_), .A1(new_n20448_), .B0(new_n20411_), .Y(new_n21137_));
  AND2X1   g20945(.A(new_n21137_), .B(new_n20395_), .Y(new_n21138_));
  AOI22X1  g20946(.A0(new_n20449_), .A1(new_n20448_), .B0(new_n20421_), .B1(\asqrt[42] ), .Y(new_n21139_));
  AOI21X1  g20947(.A0(new_n21139_), .A1(\asqrt[7] ), .B0(new_n20410_), .Y(new_n21140_));
  AOI21X1  g20948(.A0(new_n21138_), .A1(\asqrt[7] ), .B0(new_n21140_), .Y(new_n21141_));
  OAI21X1  g20949(.A0(new_n21126_), .A1(new_n21113_), .B0(new_n21133_), .Y(new_n21142_));
  AOI21X1  g20950(.A0(new_n21142_), .A1(\asqrt[42] ), .B0(\asqrt[43] ), .Y(new_n21143_));
  AOI21X1  g20951(.A0(new_n21143_), .A1(new_n21135_), .B0(new_n21141_), .Y(new_n21144_));
  OAI21X1  g20952(.A0(new_n21144_), .A1(new_n21136_), .B0(\asqrt[44] ), .Y(new_n21145_));
  AND2X1   g20953(.A(new_n20422_), .B(new_n20414_), .Y(new_n21146_));
  NOR3X1   g20954(.A(new_n21146_), .B(new_n20452_), .C(new_n20415_), .Y(new_n21147_));
  NOR3X1   g20955(.A(new_n20676_), .B(new_n21146_), .C(new_n20415_), .Y(new_n21148_));
  NOR2X1   g20956(.A(new_n21148_), .B(new_n20420_), .Y(new_n21149_));
  AOI21X1  g20957(.A0(new_n21147_), .A1(\asqrt[7] ), .B0(new_n21149_), .Y(new_n21150_));
  NOR3X1   g20958(.A(new_n21144_), .B(new_n21136_), .C(\asqrt[44] ), .Y(new_n21151_));
  OAI21X1  g20959(.A0(new_n21151_), .A1(new_n21150_), .B0(new_n21145_), .Y(new_n21152_));
  AND2X1   g20960(.A(new_n21152_), .B(\asqrt[45] ), .Y(new_n21153_));
  OR2X1    g20961(.A(new_n21151_), .B(new_n21150_), .Y(new_n21154_));
  OR4X1    g20962(.A(new_n20676_), .B(new_n20429_), .C(new_n20456_), .D(new_n20455_), .Y(new_n21155_));
  OR2X1    g20963(.A(new_n20429_), .B(new_n20455_), .Y(new_n21156_));
  OAI21X1  g20964(.A0(new_n21156_), .A1(new_n20676_), .B0(new_n20456_), .Y(new_n21157_));
  AND2X1   g20965(.A(new_n21157_), .B(new_n21155_), .Y(new_n21158_));
  AND2X1   g20966(.A(new_n21145_), .B(new_n2570_), .Y(new_n21159_));
  AOI21X1  g20967(.A0(new_n21159_), .A1(new_n21154_), .B0(new_n21158_), .Y(new_n21160_));
  OAI21X1  g20968(.A0(new_n21160_), .A1(new_n21153_), .B0(\asqrt[46] ), .Y(new_n21161_));
  AND2X1   g20969(.A(new_n20438_), .B(new_n20432_), .Y(new_n21162_));
  NOR3X1   g20970(.A(new_n21162_), .B(new_n20472_), .C(new_n20431_), .Y(new_n21163_));
  NOR3X1   g20971(.A(new_n20676_), .B(new_n21162_), .C(new_n20431_), .Y(new_n21164_));
  NOR2X1   g20972(.A(new_n21164_), .B(new_n20437_), .Y(new_n21165_));
  AOI21X1  g20973(.A0(new_n21163_), .A1(\asqrt[7] ), .B0(new_n21165_), .Y(new_n21166_));
  INVX1    g20974(.A(new_n21166_), .Y(new_n21167_));
  AND2X1   g20975(.A(new_n21142_), .B(\asqrt[42] ), .Y(new_n21168_));
  OR2X1    g20976(.A(new_n21126_), .B(new_n21113_), .Y(new_n21169_));
  AND2X1   g20977(.A(new_n21133_), .B(new_n3276_), .Y(new_n21170_));
  AOI21X1  g20978(.A0(new_n21170_), .A1(new_n21169_), .B0(new_n21131_), .Y(new_n21171_));
  OAI21X1  g20979(.A0(new_n21171_), .A1(new_n21168_), .B0(\asqrt[43] ), .Y(new_n21172_));
  INVX1    g20980(.A(new_n21141_), .Y(new_n21173_));
  OAI21X1  g20981(.A0(new_n21116_), .A1(new_n3276_), .B0(new_n3008_), .Y(new_n21174_));
  OAI21X1  g20982(.A0(new_n21174_), .A1(new_n21171_), .B0(new_n21173_), .Y(new_n21175_));
  AOI21X1  g20983(.A0(new_n21175_), .A1(new_n21172_), .B0(new_n2769_), .Y(new_n21176_));
  INVX1    g20984(.A(new_n21150_), .Y(new_n21177_));
  NAND3X1  g20985(.A(new_n21175_), .B(new_n21172_), .C(new_n2769_), .Y(new_n21178_));
  AOI21X1  g20986(.A0(new_n21178_), .A1(new_n21177_), .B0(new_n21176_), .Y(new_n21179_));
  OAI21X1  g20987(.A0(new_n21179_), .A1(new_n2570_), .B0(new_n2263_), .Y(new_n21180_));
  OAI21X1  g20988(.A0(new_n21180_), .A1(new_n21160_), .B0(new_n21167_), .Y(new_n21181_));
  AOI21X1  g20989(.A0(new_n21181_), .A1(new_n21161_), .B0(new_n2040_), .Y(new_n21182_));
  AND2X1   g20990(.A(new_n20476_), .B(new_n20474_), .Y(new_n21183_));
  NOR3X1   g20991(.A(new_n21183_), .B(new_n20446_), .C(new_n20475_), .Y(new_n21184_));
  NOR3X1   g20992(.A(new_n20676_), .B(new_n21183_), .C(new_n20475_), .Y(new_n21185_));
  NOR2X1   g20993(.A(new_n21185_), .B(new_n20445_), .Y(new_n21186_));
  AOI21X1  g20994(.A0(new_n21184_), .A1(\asqrt[7] ), .B0(new_n21186_), .Y(new_n21187_));
  INVX1    g20995(.A(new_n21187_), .Y(new_n21188_));
  NAND3X1  g20996(.A(new_n21181_), .B(new_n21161_), .C(new_n2040_), .Y(new_n21189_));
  AOI21X1  g20997(.A0(new_n21189_), .A1(new_n21188_), .B0(new_n21182_), .Y(new_n21190_));
  OR2X1    g20998(.A(new_n21190_), .B(new_n1834_), .Y(new_n21191_));
  OR2X1    g20999(.A(new_n21179_), .B(new_n2570_), .Y(new_n21192_));
  NOR2X1   g21000(.A(new_n21151_), .B(new_n21150_), .Y(new_n21193_));
  INVX1    g21001(.A(new_n21158_), .Y(new_n21194_));
  NAND2X1  g21002(.A(new_n21145_), .B(new_n2570_), .Y(new_n21195_));
  OAI21X1  g21003(.A0(new_n21195_), .A1(new_n21193_), .B0(new_n21194_), .Y(new_n21196_));
  AOI21X1  g21004(.A0(new_n21196_), .A1(new_n21192_), .B0(new_n2263_), .Y(new_n21197_));
  AOI21X1  g21005(.A0(new_n21152_), .A1(\asqrt[45] ), .B0(\asqrt[46] ), .Y(new_n21198_));
  AOI21X1  g21006(.A0(new_n21198_), .A1(new_n21196_), .B0(new_n21166_), .Y(new_n21199_));
  NOR3X1   g21007(.A(new_n21199_), .B(new_n21197_), .C(\asqrt[47] ), .Y(new_n21200_));
  NOR2X1   g21008(.A(new_n21200_), .B(new_n21187_), .Y(new_n21201_));
  OR4X1    g21009(.A(new_n20676_), .B(new_n20478_), .C(new_n20466_), .D(new_n20461_), .Y(new_n21202_));
  OR2X1    g21010(.A(new_n20478_), .B(new_n20461_), .Y(new_n21203_));
  OAI21X1  g21011(.A0(new_n21203_), .A1(new_n20676_), .B0(new_n20466_), .Y(new_n21204_));
  AND2X1   g21012(.A(new_n21204_), .B(new_n21202_), .Y(new_n21205_));
  INVX1    g21013(.A(new_n21205_), .Y(new_n21206_));
  OAI21X1  g21014(.A0(new_n21199_), .A1(new_n21197_), .B0(\asqrt[47] ), .Y(new_n21207_));
  NAND2X1  g21015(.A(new_n21207_), .B(new_n1834_), .Y(new_n21208_));
  OAI21X1  g21016(.A0(new_n21208_), .A1(new_n21201_), .B0(new_n21206_), .Y(new_n21209_));
  AOI21X1  g21017(.A0(new_n21209_), .A1(new_n21191_), .B0(new_n1632_), .Y(new_n21210_));
  AOI21X1  g21018(.A0(new_n20524_), .A1(new_n20523_), .B0(new_n20485_), .Y(new_n21211_));
  AND2X1   g21019(.A(new_n21211_), .B(new_n20469_), .Y(new_n21212_));
  AOI22X1  g21020(.A0(new_n20524_), .A1(new_n20523_), .B0(new_n20496_), .B1(\asqrt[48] ), .Y(new_n21213_));
  AOI21X1  g21021(.A0(new_n21213_), .A1(\asqrt[7] ), .B0(new_n20484_), .Y(new_n21214_));
  AOI21X1  g21022(.A0(new_n21212_), .A1(\asqrt[7] ), .B0(new_n21214_), .Y(new_n21215_));
  OAI21X1  g21023(.A0(new_n21200_), .A1(new_n21187_), .B0(new_n21207_), .Y(new_n21216_));
  AOI21X1  g21024(.A0(new_n21216_), .A1(\asqrt[48] ), .B0(\asqrt[49] ), .Y(new_n21217_));
  AOI21X1  g21025(.A0(new_n21217_), .A1(new_n21209_), .B0(new_n21215_), .Y(new_n21218_));
  OAI21X1  g21026(.A0(new_n21218_), .A1(new_n21210_), .B0(\asqrt[50] ), .Y(new_n21219_));
  AND2X1   g21027(.A(new_n20497_), .B(new_n20488_), .Y(new_n21220_));
  NOR3X1   g21028(.A(new_n21220_), .B(new_n20494_), .C(new_n20489_), .Y(new_n21221_));
  NOR3X1   g21029(.A(new_n20676_), .B(new_n21220_), .C(new_n20489_), .Y(new_n21222_));
  NOR2X1   g21030(.A(new_n21222_), .B(new_n20495_), .Y(new_n21223_));
  AOI21X1  g21031(.A0(new_n21221_), .A1(\asqrt[7] ), .B0(new_n21223_), .Y(new_n21224_));
  NOR3X1   g21032(.A(new_n21218_), .B(new_n21210_), .C(\asqrt[50] ), .Y(new_n21225_));
  OAI21X1  g21033(.A0(new_n21225_), .A1(new_n21224_), .B0(new_n21219_), .Y(new_n21226_));
  AND2X1   g21034(.A(new_n21226_), .B(\asqrt[51] ), .Y(new_n21227_));
  OR2X1    g21035(.A(new_n21225_), .B(new_n21224_), .Y(new_n21228_));
  OR4X1    g21036(.A(new_n20676_), .B(new_n20504_), .C(new_n20530_), .D(new_n20529_), .Y(new_n21229_));
  OR2X1    g21037(.A(new_n20504_), .B(new_n20529_), .Y(new_n21230_));
  OAI21X1  g21038(.A0(new_n21230_), .A1(new_n20676_), .B0(new_n20530_), .Y(new_n21231_));
  AND2X1   g21039(.A(new_n21231_), .B(new_n21229_), .Y(new_n21232_));
  AND2X1   g21040(.A(new_n21219_), .B(new_n1277_), .Y(new_n21233_));
  AOI21X1  g21041(.A0(new_n21233_), .A1(new_n21228_), .B0(new_n21232_), .Y(new_n21234_));
  OAI21X1  g21042(.A0(new_n21234_), .A1(new_n21227_), .B0(\asqrt[52] ), .Y(new_n21235_));
  AND2X1   g21043(.A(new_n20513_), .B(new_n20507_), .Y(new_n21236_));
  NOR3X1   g21044(.A(new_n21236_), .B(new_n20546_), .C(new_n20506_), .Y(new_n21237_));
  NOR3X1   g21045(.A(new_n20676_), .B(new_n21236_), .C(new_n20506_), .Y(new_n21238_));
  NOR2X1   g21046(.A(new_n21238_), .B(new_n20512_), .Y(new_n21239_));
  AOI21X1  g21047(.A0(new_n21237_), .A1(\asqrt[7] ), .B0(new_n21239_), .Y(new_n21240_));
  INVX1    g21048(.A(new_n21240_), .Y(new_n21241_));
  AND2X1   g21049(.A(new_n21216_), .B(\asqrt[48] ), .Y(new_n21242_));
  OR2X1    g21050(.A(new_n21200_), .B(new_n21187_), .Y(new_n21243_));
  AND2X1   g21051(.A(new_n21207_), .B(new_n1834_), .Y(new_n21244_));
  AOI21X1  g21052(.A0(new_n21244_), .A1(new_n21243_), .B0(new_n21205_), .Y(new_n21245_));
  OAI21X1  g21053(.A0(new_n21245_), .A1(new_n21242_), .B0(\asqrt[49] ), .Y(new_n21246_));
  INVX1    g21054(.A(new_n21215_), .Y(new_n21247_));
  OAI21X1  g21055(.A0(new_n21190_), .A1(new_n1834_), .B0(new_n1632_), .Y(new_n21248_));
  OAI21X1  g21056(.A0(new_n21248_), .A1(new_n21245_), .B0(new_n21247_), .Y(new_n21249_));
  AOI21X1  g21057(.A0(new_n21249_), .A1(new_n21246_), .B0(new_n1469_), .Y(new_n21250_));
  INVX1    g21058(.A(new_n21224_), .Y(new_n21251_));
  NAND3X1  g21059(.A(new_n21249_), .B(new_n21246_), .C(new_n1469_), .Y(new_n21252_));
  AOI21X1  g21060(.A0(new_n21252_), .A1(new_n21251_), .B0(new_n21250_), .Y(new_n21253_));
  OAI21X1  g21061(.A0(new_n21253_), .A1(new_n1277_), .B0(new_n1111_), .Y(new_n21254_));
  OAI21X1  g21062(.A0(new_n21254_), .A1(new_n21234_), .B0(new_n21241_), .Y(new_n21255_));
  AOI21X1  g21063(.A0(new_n21255_), .A1(new_n21235_), .B0(new_n968_), .Y(new_n21256_));
  AND2X1   g21064(.A(new_n20550_), .B(new_n20548_), .Y(new_n21257_));
  NOR3X1   g21065(.A(new_n21257_), .B(new_n20521_), .C(new_n20549_), .Y(new_n21258_));
  NOR3X1   g21066(.A(new_n20676_), .B(new_n21257_), .C(new_n20549_), .Y(new_n21259_));
  NOR2X1   g21067(.A(new_n21259_), .B(new_n20520_), .Y(new_n21260_));
  AOI21X1  g21068(.A0(new_n21258_), .A1(\asqrt[7] ), .B0(new_n21260_), .Y(new_n21261_));
  INVX1    g21069(.A(new_n21261_), .Y(new_n21262_));
  NAND3X1  g21070(.A(new_n21255_), .B(new_n21235_), .C(new_n968_), .Y(new_n21263_));
  AOI21X1  g21071(.A0(new_n21263_), .A1(new_n21262_), .B0(new_n21256_), .Y(new_n21264_));
  OR2X1    g21072(.A(new_n21264_), .B(new_n902_), .Y(new_n21265_));
  OR2X1    g21073(.A(new_n21253_), .B(new_n1277_), .Y(new_n21266_));
  NOR2X1   g21074(.A(new_n21225_), .B(new_n21224_), .Y(new_n21267_));
  INVX1    g21075(.A(new_n21232_), .Y(new_n21268_));
  NAND2X1  g21076(.A(new_n21219_), .B(new_n1277_), .Y(new_n21269_));
  OAI21X1  g21077(.A0(new_n21269_), .A1(new_n21267_), .B0(new_n21268_), .Y(new_n21270_));
  AOI21X1  g21078(.A0(new_n21270_), .A1(new_n21266_), .B0(new_n1111_), .Y(new_n21271_));
  AOI21X1  g21079(.A0(new_n21226_), .A1(\asqrt[51] ), .B0(\asqrt[52] ), .Y(new_n21272_));
  AOI21X1  g21080(.A0(new_n21272_), .A1(new_n21270_), .B0(new_n21240_), .Y(new_n21273_));
  NOR3X1   g21081(.A(new_n21273_), .B(new_n21271_), .C(\asqrt[53] ), .Y(new_n21274_));
  NOR2X1   g21082(.A(new_n21274_), .B(new_n21261_), .Y(new_n21275_));
  OR4X1    g21083(.A(new_n20676_), .B(new_n20552_), .C(new_n20540_), .D(new_n20535_), .Y(new_n21276_));
  OR2X1    g21084(.A(new_n20552_), .B(new_n20535_), .Y(new_n21277_));
  OAI21X1  g21085(.A0(new_n21277_), .A1(new_n20676_), .B0(new_n20540_), .Y(new_n21278_));
  AND2X1   g21086(.A(new_n21278_), .B(new_n21276_), .Y(new_n21279_));
  INVX1    g21087(.A(new_n21279_), .Y(new_n21280_));
  OAI21X1  g21088(.A0(new_n21273_), .A1(new_n21271_), .B0(\asqrt[53] ), .Y(new_n21281_));
  NAND2X1  g21089(.A(new_n21281_), .B(new_n902_), .Y(new_n21282_));
  OAI21X1  g21090(.A0(new_n21282_), .A1(new_n21275_), .B0(new_n21280_), .Y(new_n21283_));
  AOI21X1  g21091(.A0(new_n21283_), .A1(new_n21265_), .B0(new_n697_), .Y(new_n21284_));
  AOI21X1  g21092(.A0(new_n20597_), .A1(new_n20596_), .B0(new_n20559_), .Y(new_n21285_));
  AND2X1   g21093(.A(new_n21285_), .B(new_n20543_), .Y(new_n21286_));
  AOI22X1  g21094(.A0(new_n20597_), .A1(new_n20596_), .B0(new_n20569_), .B1(\asqrt[54] ), .Y(new_n21287_));
  AOI21X1  g21095(.A0(new_n21287_), .A1(\asqrt[7] ), .B0(new_n20558_), .Y(new_n21288_));
  AOI21X1  g21096(.A0(new_n21286_), .A1(\asqrt[7] ), .B0(new_n21288_), .Y(new_n21289_));
  OAI21X1  g21097(.A0(new_n21274_), .A1(new_n21261_), .B0(new_n21281_), .Y(new_n21290_));
  AOI21X1  g21098(.A0(new_n21290_), .A1(\asqrt[54] ), .B0(\asqrt[55] ), .Y(new_n21291_));
  AOI21X1  g21099(.A0(new_n21291_), .A1(new_n21283_), .B0(new_n21289_), .Y(new_n21292_));
  OAI21X1  g21100(.A0(new_n21292_), .A1(new_n21284_), .B0(\asqrt[56] ), .Y(new_n21293_));
  AND2X1   g21101(.A(new_n20570_), .B(new_n20562_), .Y(new_n21294_));
  NOR3X1   g21102(.A(new_n21294_), .B(new_n20600_), .C(new_n20563_), .Y(new_n21295_));
  NOR3X1   g21103(.A(new_n20676_), .B(new_n21294_), .C(new_n20563_), .Y(new_n21296_));
  NOR2X1   g21104(.A(new_n21296_), .B(new_n20568_), .Y(new_n21297_));
  AOI21X1  g21105(.A0(new_n21295_), .A1(\asqrt[7] ), .B0(new_n21297_), .Y(new_n21298_));
  NOR3X1   g21106(.A(new_n21292_), .B(new_n21284_), .C(\asqrt[56] ), .Y(new_n21299_));
  OAI21X1  g21107(.A0(new_n21299_), .A1(new_n21298_), .B0(new_n21293_), .Y(new_n21300_));
  AND2X1   g21108(.A(new_n21300_), .B(\asqrt[57] ), .Y(new_n21301_));
  OR2X1    g21109(.A(new_n21299_), .B(new_n21298_), .Y(new_n21302_));
  OR4X1    g21110(.A(new_n20676_), .B(new_n20577_), .C(new_n20604_), .D(new_n20603_), .Y(new_n21303_));
  OR2X1    g21111(.A(new_n20577_), .B(new_n20603_), .Y(new_n21304_));
  OAI21X1  g21112(.A0(new_n21304_), .A1(new_n20676_), .B0(new_n20604_), .Y(new_n21305_));
  AND2X1   g21113(.A(new_n21305_), .B(new_n21303_), .Y(new_n21306_));
  AND2X1   g21114(.A(new_n21293_), .B(new_n481_), .Y(new_n21307_));
  AOI21X1  g21115(.A0(new_n21307_), .A1(new_n21302_), .B0(new_n21306_), .Y(new_n21308_));
  OAI21X1  g21116(.A0(new_n21308_), .A1(new_n21301_), .B0(\asqrt[58] ), .Y(new_n21309_));
  AND2X1   g21117(.A(new_n21290_), .B(\asqrt[54] ), .Y(new_n21310_));
  OR2X1    g21118(.A(new_n21274_), .B(new_n21261_), .Y(new_n21311_));
  AND2X1   g21119(.A(new_n21281_), .B(new_n902_), .Y(new_n21312_));
  AOI21X1  g21120(.A0(new_n21312_), .A1(new_n21311_), .B0(new_n21279_), .Y(new_n21313_));
  OAI21X1  g21121(.A0(new_n21313_), .A1(new_n21310_), .B0(\asqrt[55] ), .Y(new_n21314_));
  INVX1    g21122(.A(new_n21289_), .Y(new_n21315_));
  OAI21X1  g21123(.A0(new_n21264_), .A1(new_n902_), .B0(new_n697_), .Y(new_n21316_));
  OAI21X1  g21124(.A0(new_n21316_), .A1(new_n21313_), .B0(new_n21315_), .Y(new_n21317_));
  AOI21X1  g21125(.A0(new_n21317_), .A1(new_n21314_), .B0(new_n582_), .Y(new_n21318_));
  INVX1    g21126(.A(new_n21298_), .Y(new_n21319_));
  NAND3X1  g21127(.A(new_n21317_), .B(new_n21314_), .C(new_n582_), .Y(new_n21320_));
  AOI21X1  g21128(.A0(new_n21320_), .A1(new_n21319_), .B0(new_n21318_), .Y(new_n21321_));
  OAI21X1  g21129(.A0(new_n21321_), .A1(new_n481_), .B0(new_n399_), .Y(new_n21322_));
  AND2X1   g21130(.A(new_n20581_), .B(new_n20580_), .Y(new_n21323_));
  NOR3X1   g21131(.A(new_n20620_), .B(new_n21323_), .C(new_n20579_), .Y(new_n21324_));
  NOR3X1   g21132(.A(new_n20676_), .B(new_n21323_), .C(new_n20579_), .Y(new_n21325_));
  NOR2X1   g21133(.A(new_n21325_), .B(new_n20586_), .Y(new_n21326_));
  AOI21X1  g21134(.A0(new_n21324_), .A1(\asqrt[7] ), .B0(new_n21326_), .Y(new_n21327_));
  INVX1    g21135(.A(new_n21327_), .Y(new_n21328_));
  OAI21X1  g21136(.A0(new_n21322_), .A1(new_n21308_), .B0(new_n21328_), .Y(new_n21329_));
  AOI21X1  g21137(.A0(new_n21329_), .A1(new_n21309_), .B0(new_n328_), .Y(new_n21330_));
  AND2X1   g21138(.A(new_n20623_), .B(new_n20621_), .Y(new_n21331_));
  NOR3X1   g21139(.A(new_n21331_), .B(new_n20594_), .C(new_n20622_), .Y(new_n21332_));
  NOR3X1   g21140(.A(new_n20676_), .B(new_n21331_), .C(new_n20622_), .Y(new_n21333_));
  NOR2X1   g21141(.A(new_n21333_), .B(new_n20593_), .Y(new_n21334_));
  AOI21X1  g21142(.A0(new_n21332_), .A1(\asqrt[7] ), .B0(new_n21334_), .Y(new_n21335_));
  INVX1    g21143(.A(new_n21335_), .Y(new_n21336_));
  NAND3X1  g21144(.A(new_n21329_), .B(new_n21309_), .C(new_n328_), .Y(new_n21337_));
  AOI21X1  g21145(.A0(new_n21337_), .A1(new_n21336_), .B0(new_n21330_), .Y(new_n21338_));
  OR2X1    g21146(.A(new_n21338_), .B(new_n292_), .Y(new_n21339_));
  OR2X1    g21147(.A(new_n21321_), .B(new_n481_), .Y(new_n21340_));
  NOR2X1   g21148(.A(new_n21299_), .B(new_n21298_), .Y(new_n21341_));
  INVX1    g21149(.A(new_n21306_), .Y(new_n21342_));
  NAND2X1  g21150(.A(new_n21293_), .B(new_n481_), .Y(new_n21343_));
  OAI21X1  g21151(.A0(new_n21343_), .A1(new_n21341_), .B0(new_n21342_), .Y(new_n21344_));
  AOI21X1  g21152(.A0(new_n21344_), .A1(new_n21340_), .B0(new_n399_), .Y(new_n21345_));
  AOI21X1  g21153(.A0(new_n21300_), .A1(\asqrt[57] ), .B0(\asqrt[58] ), .Y(new_n21346_));
  AOI21X1  g21154(.A0(new_n21346_), .A1(new_n21344_), .B0(new_n21327_), .Y(new_n21347_));
  NOR3X1   g21155(.A(new_n21347_), .B(new_n21345_), .C(\asqrt[59] ), .Y(new_n21348_));
  NOR2X1   g21156(.A(new_n21348_), .B(new_n21335_), .Y(new_n21349_));
  OR4X1    g21157(.A(new_n20676_), .B(new_n20625_), .C(new_n20612_), .D(new_n20609_), .Y(new_n21350_));
  OR2X1    g21158(.A(new_n20625_), .B(new_n20609_), .Y(new_n21351_));
  OAI21X1  g21159(.A0(new_n21351_), .A1(new_n20676_), .B0(new_n20612_), .Y(new_n21352_));
  AND2X1   g21160(.A(new_n21352_), .B(new_n21350_), .Y(new_n21353_));
  INVX1    g21161(.A(new_n21353_), .Y(new_n21354_));
  OAI21X1  g21162(.A0(new_n21347_), .A1(new_n21345_), .B0(\asqrt[59] ), .Y(new_n21355_));
  NAND2X1  g21163(.A(new_n21355_), .B(new_n292_), .Y(new_n21356_));
  OAI21X1  g21164(.A0(new_n21356_), .A1(new_n21349_), .B0(new_n21354_), .Y(new_n21357_));
  AOI21X1  g21165(.A0(new_n21357_), .A1(new_n21339_), .B0(new_n217_), .Y(new_n21358_));
  AOI21X1  g21166(.A0(new_n20685_), .A1(new_n20684_), .B0(new_n20632_), .Y(new_n21359_));
  AND2X1   g21167(.A(new_n21359_), .B(new_n20615_), .Y(new_n21360_));
  AOI22X1  g21168(.A0(new_n20685_), .A1(new_n20684_), .B0(new_n20642_), .B1(\asqrt[60] ), .Y(new_n21361_));
  AOI21X1  g21169(.A0(new_n21361_), .A1(\asqrt[7] ), .B0(new_n20631_), .Y(new_n21362_));
  AOI21X1  g21170(.A0(new_n21360_), .A1(\asqrt[7] ), .B0(new_n21362_), .Y(new_n21363_));
  OAI21X1  g21171(.A0(new_n21348_), .A1(new_n21335_), .B0(new_n21355_), .Y(new_n21364_));
  AOI21X1  g21172(.A0(new_n21364_), .A1(\asqrt[60] ), .B0(\asqrt[61] ), .Y(new_n21365_));
  AOI21X1  g21173(.A0(new_n21365_), .A1(new_n21357_), .B0(new_n21363_), .Y(new_n21366_));
  OAI21X1  g21174(.A0(new_n21366_), .A1(new_n21358_), .B0(\asqrt[62] ), .Y(new_n21367_));
  AND2X1   g21175(.A(new_n20643_), .B(new_n20635_), .Y(new_n21368_));
  NOR3X1   g21176(.A(new_n21368_), .B(new_n20688_), .C(new_n20636_), .Y(new_n21369_));
  NOR3X1   g21177(.A(new_n20676_), .B(new_n21368_), .C(new_n20636_), .Y(new_n21370_));
  NOR2X1   g21178(.A(new_n21370_), .B(new_n20641_), .Y(new_n21371_));
  AOI21X1  g21179(.A0(new_n21369_), .A1(\asqrt[7] ), .B0(new_n21371_), .Y(new_n21372_));
  NOR3X1   g21180(.A(new_n21366_), .B(new_n21358_), .C(\asqrt[62] ), .Y(new_n21373_));
  OAI21X1  g21181(.A0(new_n21373_), .A1(new_n21372_), .B0(new_n21367_), .Y(new_n21374_));
  NAND4X1  g21182(.A(\asqrt[7] ), .B(new_n20693_), .C(new_n20649_), .D(new_n20645_), .Y(new_n21375_));
  NAND2X1  g21183(.A(new_n20693_), .B(new_n20645_), .Y(new_n21376_));
  OAI21X1  g21184(.A0(new_n21376_), .A1(new_n20676_), .B0(new_n20692_), .Y(new_n21377_));
  AND2X1   g21185(.A(new_n21377_), .B(new_n21375_), .Y(new_n21378_));
  INVX1    g21186(.A(new_n21378_), .Y(new_n21379_));
  AND2X1   g21187(.A(new_n20657_), .B(new_n20651_), .Y(new_n21380_));
  AOI21X1  g21188(.A0(new_n21380_), .A1(\asqrt[7] ), .B0(new_n20717_), .Y(new_n21381_));
  AND2X1   g21189(.A(new_n21381_), .B(new_n21379_), .Y(new_n21382_));
  AOI21X1  g21190(.A0(new_n21382_), .A1(new_n21374_), .B0(\asqrt[63] ), .Y(new_n21383_));
  NOR2X1   g21191(.A(new_n21373_), .B(new_n21372_), .Y(new_n21384_));
  NAND2X1  g21192(.A(new_n21378_), .B(new_n21367_), .Y(new_n21385_));
  AOI21X1  g21193(.A0(\asqrt[7] ), .A1(new_n20657_), .B0(new_n20651_), .Y(new_n21386_));
  NOR3X1   g21194(.A(new_n21386_), .B(new_n21380_), .C(new_n193_), .Y(new_n21387_));
  NOR4X1   g21195(.A(new_n20673_), .B(new_n20718_), .C(new_n20655_), .D(new_n20653_), .Y(new_n21388_));
  OAI21X1  g21196(.A0(new_n20664_), .A1(new_n20663_), .B0(new_n21388_), .Y(new_n21389_));
  NOR2X1   g21197(.A(new_n21389_), .B(new_n20662_), .Y(new_n21390_));
  NOR2X1   g21198(.A(new_n21390_), .B(new_n21387_), .Y(new_n21391_));
  OAI21X1  g21199(.A0(new_n21385_), .A1(new_n21384_), .B0(new_n21391_), .Y(new_n21392_));
  NOR2X1   g21200(.A(new_n21392_), .B(new_n21383_), .Y(new_n21393_));
  INVX1    g21201(.A(\a[12] ), .Y(new_n21394_));
  AND2X1   g21202(.A(new_n21364_), .B(\asqrt[60] ), .Y(new_n21395_));
  OR2X1    g21203(.A(new_n21348_), .B(new_n21335_), .Y(new_n21396_));
  AND2X1   g21204(.A(new_n21355_), .B(new_n292_), .Y(new_n21397_));
  AOI21X1  g21205(.A0(new_n21397_), .A1(new_n21396_), .B0(new_n21353_), .Y(new_n21398_));
  OAI21X1  g21206(.A0(new_n21398_), .A1(new_n21395_), .B0(\asqrt[61] ), .Y(new_n21399_));
  INVX1    g21207(.A(new_n21363_), .Y(new_n21400_));
  OAI21X1  g21208(.A0(new_n21338_), .A1(new_n292_), .B0(new_n217_), .Y(new_n21401_));
  OAI21X1  g21209(.A0(new_n21401_), .A1(new_n21398_), .B0(new_n21400_), .Y(new_n21402_));
  AOI21X1  g21210(.A0(new_n21402_), .A1(new_n21399_), .B0(new_n199_), .Y(new_n21403_));
  INVX1    g21211(.A(new_n21372_), .Y(new_n21404_));
  NAND3X1  g21212(.A(new_n21402_), .B(new_n21399_), .C(new_n199_), .Y(new_n21405_));
  AOI21X1  g21213(.A0(new_n21405_), .A1(new_n21404_), .B0(new_n21403_), .Y(new_n21406_));
  INVX1    g21214(.A(new_n21382_), .Y(new_n21407_));
  OAI21X1  g21215(.A0(new_n21407_), .A1(new_n21406_), .B0(new_n193_), .Y(new_n21408_));
  OR2X1    g21216(.A(new_n21373_), .B(new_n21372_), .Y(new_n21409_));
  AND2X1   g21217(.A(new_n21378_), .B(new_n21367_), .Y(new_n21410_));
  INVX1    g21218(.A(new_n21391_), .Y(new_n21411_));
  AOI21X1  g21219(.A0(new_n21410_), .A1(new_n21409_), .B0(new_n21411_), .Y(new_n21412_));
  AOI21X1  g21220(.A0(new_n21412_), .A1(new_n21408_), .B0(new_n21394_), .Y(new_n21413_));
  NOR3X1   g21221(.A(\a[12] ), .B(\a[11] ), .C(\a[10] ), .Y(new_n21414_));
  OAI21X1  g21222(.A0(new_n21414_), .A1(new_n21413_), .B0(\asqrt[7] ), .Y(new_n21415_));
  OAI21X1  g21223(.A0(new_n21392_), .A1(new_n21383_), .B0(\a[12] ), .Y(new_n21416_));
  INVX1    g21224(.A(new_n21414_), .Y(new_n21417_));
  OAI21X1  g21225(.A0(new_n20672_), .A1(new_n20668_), .B0(new_n21417_), .Y(new_n21418_));
  NOR4X1   g21226(.A(new_n21418_), .B(new_n20718_), .C(new_n20717_), .D(new_n20662_), .Y(new_n21419_));
  AND2X1   g21227(.A(new_n21419_), .B(new_n21416_), .Y(new_n21420_));
  INVX1    g21228(.A(\a[13] ), .Y(new_n21421_));
  AOI21X1  g21229(.A0(new_n21412_), .A1(new_n21408_), .B0(\a[12] ), .Y(new_n21422_));
  OAI21X1  g21230(.A0(new_n21392_), .A1(new_n21383_), .B0(new_n20680_), .Y(new_n21423_));
  OAI21X1  g21231(.A0(new_n21422_), .A1(new_n21421_), .B0(new_n21423_), .Y(new_n21424_));
  OAI21X1  g21232(.A0(new_n21424_), .A1(new_n21420_), .B0(new_n21415_), .Y(new_n21425_));
  AND2X1   g21233(.A(new_n21425_), .B(\asqrt[8] ), .Y(new_n21426_));
  NAND2X1  g21234(.A(new_n21419_), .B(new_n21416_), .Y(new_n21427_));
  OAI21X1  g21235(.A0(new_n21392_), .A1(new_n21383_), .B0(new_n21394_), .Y(new_n21428_));
  INVX1    g21236(.A(new_n20680_), .Y(new_n21429_));
  AOI21X1  g21237(.A0(new_n21412_), .A1(new_n21408_), .B0(new_n21429_), .Y(new_n21430_));
  AOI21X1  g21238(.A0(new_n21428_), .A1(\a[13] ), .B0(new_n21430_), .Y(new_n21431_));
  NAND2X1  g21239(.A(new_n21431_), .B(new_n21427_), .Y(new_n21432_));
  AND2X1   g21240(.A(new_n21415_), .B(new_n19976_), .Y(new_n21433_));
  NOR3X1   g21241(.A(new_n21390_), .B(new_n21387_), .C(new_n20676_), .Y(new_n21434_));
  OAI21X1  g21242(.A0(new_n21385_), .A1(new_n21384_), .B0(new_n21434_), .Y(new_n21435_));
  OR2X1    g21243(.A(new_n21435_), .B(new_n21383_), .Y(new_n21436_));
  AOI21X1  g21244(.A0(new_n21436_), .A1(new_n21423_), .B0(new_n20679_), .Y(new_n21437_));
  OAI21X1  g21245(.A0(new_n21435_), .A1(new_n21383_), .B0(new_n20679_), .Y(new_n21438_));
  NOR2X1   g21246(.A(new_n21438_), .B(new_n21430_), .Y(new_n21439_));
  NOR2X1   g21247(.A(new_n21439_), .B(new_n21437_), .Y(new_n21440_));
  AOI21X1  g21248(.A0(new_n21433_), .A1(new_n21432_), .B0(new_n21440_), .Y(new_n21441_));
  OAI21X1  g21249(.A0(new_n21441_), .A1(new_n21426_), .B0(\asqrt[9] ), .Y(new_n21442_));
  NOR3X1   g21250(.A(new_n20713_), .B(new_n20703_), .C(new_n20715_), .Y(new_n21443_));
  OAI21X1  g21251(.A0(new_n21392_), .A1(new_n21383_), .B0(new_n21443_), .Y(new_n21444_));
  NOR2X1   g21252(.A(new_n20703_), .B(new_n20715_), .Y(new_n21445_));
  OAI21X1  g21253(.A0(new_n21392_), .A1(new_n21383_), .B0(new_n21445_), .Y(new_n21446_));
  NAND2X1  g21254(.A(new_n21446_), .B(new_n20713_), .Y(new_n21447_));
  NAND2X1  g21255(.A(new_n21447_), .B(new_n21444_), .Y(new_n21448_));
  AOI21X1  g21256(.A0(new_n21417_), .A1(new_n21416_), .B0(new_n20676_), .Y(new_n21449_));
  AOI21X1  g21257(.A0(new_n21431_), .A1(new_n21427_), .B0(new_n21449_), .Y(new_n21450_));
  OAI21X1  g21258(.A0(new_n21450_), .A1(new_n19976_), .B0(new_n19273_), .Y(new_n21451_));
  OAI21X1  g21259(.A0(new_n21451_), .A1(new_n21441_), .B0(new_n21448_), .Y(new_n21452_));
  AOI21X1  g21260(.A0(new_n21452_), .A1(new_n21442_), .B0(new_n18591_), .Y(new_n21453_));
  AOI21X1  g21261(.A0(new_n20716_), .A1(new_n20714_), .B0(new_n20752_), .Y(new_n21454_));
  AND2X1   g21262(.A(new_n21454_), .B(new_n20749_), .Y(new_n21455_));
  OAI21X1  g21263(.A0(new_n21392_), .A1(new_n21383_), .B0(new_n21455_), .Y(new_n21456_));
  AOI22X1  g21264(.A0(new_n20716_), .A1(new_n20714_), .B0(new_n20708_), .B1(\asqrt[9] ), .Y(new_n21457_));
  OAI21X1  g21265(.A0(new_n21392_), .A1(new_n21383_), .B0(new_n21457_), .Y(new_n21458_));
  NAND2X1  g21266(.A(new_n21458_), .B(new_n20752_), .Y(new_n21459_));
  AND2X1   g21267(.A(new_n21459_), .B(new_n21456_), .Y(new_n21460_));
  INVX1    g21268(.A(new_n21460_), .Y(new_n21461_));
  NAND3X1  g21269(.A(new_n21452_), .B(new_n21442_), .C(new_n18591_), .Y(new_n21462_));
  AOI21X1  g21270(.A0(new_n21462_), .A1(new_n21461_), .B0(new_n21453_), .Y(new_n21463_));
  OR2X1    g21271(.A(new_n21463_), .B(new_n17927_), .Y(new_n21464_));
  OR2X1    g21272(.A(new_n21450_), .B(new_n19976_), .Y(new_n21465_));
  AND2X1   g21273(.A(new_n21431_), .B(new_n21427_), .Y(new_n21466_));
  OR2X1    g21274(.A(new_n21449_), .B(\asqrt[8] ), .Y(new_n21467_));
  OR2X1    g21275(.A(new_n21439_), .B(new_n21437_), .Y(new_n21468_));
  OAI21X1  g21276(.A0(new_n21467_), .A1(new_n21466_), .B0(new_n21468_), .Y(new_n21469_));
  AOI21X1  g21277(.A0(new_n21469_), .A1(new_n21465_), .B0(new_n19273_), .Y(new_n21470_));
  AND2X1   g21278(.A(new_n21447_), .B(new_n21444_), .Y(new_n21471_));
  AOI21X1  g21279(.A0(new_n21425_), .A1(\asqrt[8] ), .B0(\asqrt[9] ), .Y(new_n21472_));
  AOI21X1  g21280(.A0(new_n21472_), .A1(new_n21469_), .B0(new_n21471_), .Y(new_n21473_));
  NOR3X1   g21281(.A(new_n21473_), .B(new_n21470_), .C(\asqrt[10] ), .Y(new_n21474_));
  NOR2X1   g21282(.A(new_n21474_), .B(new_n21460_), .Y(new_n21475_));
  INVX1    g21283(.A(new_n21393_), .Y(\asqrt[6] ));
  AND2X1   g21284(.A(new_n20755_), .B(new_n20753_), .Y(new_n21477_));
  NOR3X1   g21285(.A(new_n21477_), .B(new_n20733_), .C(new_n20754_), .Y(new_n21478_));
  NOR2X1   g21286(.A(new_n21477_), .B(new_n20754_), .Y(new_n21479_));
  OAI21X1  g21287(.A0(new_n21392_), .A1(new_n21383_), .B0(new_n21479_), .Y(new_n21480_));
  AOI22X1  g21288(.A0(new_n21480_), .A1(new_n20733_), .B0(new_n21478_), .B1(\asqrt[6] ), .Y(new_n21481_));
  INVX1    g21289(.A(new_n21481_), .Y(new_n21482_));
  OAI21X1  g21290(.A0(new_n21473_), .A1(new_n21470_), .B0(\asqrt[10] ), .Y(new_n21483_));
  NAND2X1  g21291(.A(new_n21483_), .B(new_n17927_), .Y(new_n21484_));
  OAI21X1  g21292(.A0(new_n21484_), .A1(new_n21475_), .B0(new_n21482_), .Y(new_n21485_));
  AOI21X1  g21293(.A0(new_n21485_), .A1(new_n21464_), .B0(new_n17262_), .Y(new_n21486_));
  NAND4X1  g21294(.A(\asqrt[6] ), .B(new_n20746_), .C(new_n20744_), .D(new_n20771_), .Y(new_n21487_));
  NOR3X1   g21295(.A(new_n21393_), .B(new_n20757_), .C(new_n20737_), .Y(new_n21488_));
  OAI21X1  g21296(.A0(new_n21488_), .A1(new_n20744_), .B0(new_n21487_), .Y(new_n21489_));
  INVX1    g21297(.A(new_n21489_), .Y(new_n21490_));
  OAI21X1  g21298(.A0(new_n21474_), .A1(new_n21460_), .B0(new_n21483_), .Y(new_n21491_));
  AOI21X1  g21299(.A0(new_n21491_), .A1(\asqrt[11] ), .B0(\asqrt[12] ), .Y(new_n21492_));
  AOI21X1  g21300(.A0(new_n21492_), .A1(new_n21485_), .B0(new_n21490_), .Y(new_n21493_));
  OAI21X1  g21301(.A0(new_n21493_), .A1(new_n21486_), .B0(\asqrt[13] ), .Y(new_n21494_));
  AND2X1   g21302(.A(new_n20800_), .B(new_n20799_), .Y(new_n21495_));
  NOR3X1   g21303(.A(new_n21495_), .B(new_n20762_), .C(new_n20798_), .Y(new_n21496_));
  NOR3X1   g21304(.A(new_n21393_), .B(new_n21495_), .C(new_n20798_), .Y(new_n21497_));
  NOR2X1   g21305(.A(new_n21497_), .B(new_n20761_), .Y(new_n21498_));
  AOI21X1  g21306(.A0(new_n21496_), .A1(\asqrt[6] ), .B0(new_n21498_), .Y(new_n21499_));
  NOR3X1   g21307(.A(new_n21493_), .B(new_n21486_), .C(\asqrt[13] ), .Y(new_n21500_));
  OAI21X1  g21308(.A0(new_n21500_), .A1(new_n21499_), .B0(new_n21494_), .Y(new_n21501_));
  AND2X1   g21309(.A(new_n21501_), .B(\asqrt[14] ), .Y(new_n21502_));
  INVX1    g21310(.A(new_n21499_), .Y(new_n21503_));
  AND2X1   g21311(.A(new_n21491_), .B(\asqrt[11] ), .Y(new_n21504_));
  OR2X1    g21312(.A(new_n21474_), .B(new_n21460_), .Y(new_n21505_));
  AND2X1   g21313(.A(new_n21483_), .B(new_n17927_), .Y(new_n21506_));
  AOI21X1  g21314(.A0(new_n21506_), .A1(new_n21505_), .B0(new_n21481_), .Y(new_n21507_));
  OAI21X1  g21315(.A0(new_n21507_), .A1(new_n21504_), .B0(\asqrt[12] ), .Y(new_n21508_));
  OAI21X1  g21316(.A0(new_n21463_), .A1(new_n17927_), .B0(new_n17262_), .Y(new_n21509_));
  OAI21X1  g21317(.A0(new_n21509_), .A1(new_n21507_), .B0(new_n21489_), .Y(new_n21510_));
  NAND3X1  g21318(.A(new_n21510_), .B(new_n21508_), .C(new_n16617_), .Y(new_n21511_));
  NAND2X1  g21319(.A(new_n21511_), .B(new_n21503_), .Y(new_n21512_));
  AND2X1   g21320(.A(new_n20773_), .B(new_n20764_), .Y(new_n21513_));
  NOR3X1   g21321(.A(new_n21513_), .B(new_n20803_), .C(new_n20765_), .Y(new_n21514_));
  NOR3X1   g21322(.A(new_n21393_), .B(new_n21513_), .C(new_n20765_), .Y(new_n21515_));
  NOR2X1   g21323(.A(new_n21515_), .B(new_n20770_), .Y(new_n21516_));
  AOI21X1  g21324(.A0(new_n21514_), .A1(\asqrt[6] ), .B0(new_n21516_), .Y(new_n21517_));
  AND2X1   g21325(.A(new_n21494_), .B(new_n15990_), .Y(new_n21518_));
  AOI21X1  g21326(.A0(new_n21518_), .A1(new_n21512_), .B0(new_n21517_), .Y(new_n21519_));
  OAI21X1  g21327(.A0(new_n21519_), .A1(new_n21502_), .B0(\asqrt[15] ), .Y(new_n21520_));
  OR4X1    g21328(.A(new_n21393_), .B(new_n20781_), .C(new_n20807_), .D(new_n20806_), .Y(new_n21521_));
  OR2X1    g21329(.A(new_n20781_), .B(new_n20806_), .Y(new_n21522_));
  OAI21X1  g21330(.A0(new_n21522_), .A1(new_n21393_), .B0(new_n20807_), .Y(new_n21523_));
  AND2X1   g21331(.A(new_n21523_), .B(new_n21521_), .Y(new_n21524_));
  INVX1    g21332(.A(new_n21524_), .Y(new_n21525_));
  AOI21X1  g21333(.A0(new_n21510_), .A1(new_n21508_), .B0(new_n16617_), .Y(new_n21526_));
  AOI21X1  g21334(.A0(new_n21511_), .A1(new_n21503_), .B0(new_n21526_), .Y(new_n21527_));
  OAI21X1  g21335(.A0(new_n21527_), .A1(new_n15990_), .B0(new_n15362_), .Y(new_n21528_));
  OAI21X1  g21336(.A0(new_n21528_), .A1(new_n21519_), .B0(new_n21525_), .Y(new_n21529_));
  AOI21X1  g21337(.A0(new_n21529_), .A1(new_n21520_), .B0(new_n14754_), .Y(new_n21530_));
  OAI21X1  g21338(.A0(new_n20825_), .A1(new_n20823_), .B0(new_n20788_), .Y(new_n21531_));
  NOR2X1   g21339(.A(new_n21531_), .B(new_n20783_), .Y(new_n21532_));
  AOI22X1  g21340(.A0(new_n20789_), .A1(new_n20784_), .B0(new_n20782_), .B1(\asqrt[15] ), .Y(new_n21533_));
  AOI21X1  g21341(.A0(new_n21533_), .A1(\asqrt[6] ), .B0(new_n20788_), .Y(new_n21534_));
  AOI21X1  g21342(.A0(new_n21532_), .A1(\asqrt[6] ), .B0(new_n21534_), .Y(new_n21535_));
  INVX1    g21343(.A(new_n21535_), .Y(new_n21536_));
  NAND3X1  g21344(.A(new_n21529_), .B(new_n21520_), .C(new_n14754_), .Y(new_n21537_));
  AOI21X1  g21345(.A0(new_n21537_), .A1(new_n21536_), .B0(new_n21530_), .Y(new_n21538_));
  OR2X1    g21346(.A(new_n21538_), .B(new_n14165_), .Y(new_n21539_));
  AND2X1   g21347(.A(new_n21537_), .B(new_n21536_), .Y(new_n21540_));
  AND2X1   g21348(.A(new_n20828_), .B(new_n20826_), .Y(new_n21541_));
  NOR3X1   g21349(.A(new_n21541_), .B(new_n20797_), .C(new_n20827_), .Y(new_n21542_));
  NOR3X1   g21350(.A(new_n21393_), .B(new_n21541_), .C(new_n20827_), .Y(new_n21543_));
  NOR2X1   g21351(.A(new_n21543_), .B(new_n20796_), .Y(new_n21544_));
  AOI21X1  g21352(.A0(new_n21542_), .A1(\asqrt[6] ), .B0(new_n21544_), .Y(new_n21545_));
  INVX1    g21353(.A(new_n21545_), .Y(new_n21546_));
  OR2X1    g21354(.A(new_n21527_), .B(new_n15990_), .Y(new_n21547_));
  AND2X1   g21355(.A(new_n21511_), .B(new_n21503_), .Y(new_n21548_));
  INVX1    g21356(.A(new_n21517_), .Y(new_n21549_));
  NAND2X1  g21357(.A(new_n21494_), .B(new_n15990_), .Y(new_n21550_));
  OAI21X1  g21358(.A0(new_n21550_), .A1(new_n21548_), .B0(new_n21549_), .Y(new_n21551_));
  AOI21X1  g21359(.A0(new_n21551_), .A1(new_n21547_), .B0(new_n15362_), .Y(new_n21552_));
  AOI21X1  g21360(.A0(new_n21501_), .A1(\asqrt[14] ), .B0(\asqrt[15] ), .Y(new_n21553_));
  AOI21X1  g21361(.A0(new_n21553_), .A1(new_n21551_), .B0(new_n21524_), .Y(new_n21554_));
  OAI21X1  g21362(.A0(new_n21554_), .A1(new_n21552_), .B0(\asqrt[16] ), .Y(new_n21555_));
  NAND2X1  g21363(.A(new_n21555_), .B(new_n14165_), .Y(new_n21556_));
  OAI21X1  g21364(.A0(new_n21556_), .A1(new_n21540_), .B0(new_n21546_), .Y(new_n21557_));
  AOI21X1  g21365(.A0(new_n21557_), .A1(new_n21539_), .B0(new_n13571_), .Y(new_n21558_));
  OR4X1    g21366(.A(new_n21393_), .B(new_n20830_), .C(new_n20818_), .D(new_n20812_), .Y(new_n21559_));
  OR2X1    g21367(.A(new_n20830_), .B(new_n20812_), .Y(new_n21560_));
  OAI21X1  g21368(.A0(new_n21560_), .A1(new_n21393_), .B0(new_n20818_), .Y(new_n21561_));
  AND2X1   g21369(.A(new_n21561_), .B(new_n21559_), .Y(new_n21562_));
  NOR3X1   g21370(.A(new_n21554_), .B(new_n21552_), .C(\asqrt[16] ), .Y(new_n21563_));
  OAI21X1  g21371(.A0(new_n21563_), .A1(new_n21535_), .B0(new_n21555_), .Y(new_n21564_));
  AOI21X1  g21372(.A0(new_n21564_), .A1(\asqrt[17] ), .B0(\asqrt[18] ), .Y(new_n21565_));
  AOI21X1  g21373(.A0(new_n21565_), .A1(new_n21557_), .B0(new_n21562_), .Y(new_n21566_));
  OAI21X1  g21374(.A0(new_n21566_), .A1(new_n21558_), .B0(\asqrt[19] ), .Y(new_n21567_));
  AND2X1   g21375(.A(new_n20861_), .B(new_n20860_), .Y(new_n21568_));
  NOR3X1   g21376(.A(new_n21568_), .B(new_n20836_), .C(new_n20859_), .Y(new_n21569_));
  NOR3X1   g21377(.A(new_n21393_), .B(new_n21568_), .C(new_n20859_), .Y(new_n21570_));
  NOR2X1   g21378(.A(new_n21570_), .B(new_n20835_), .Y(new_n21571_));
  AOI21X1  g21379(.A0(new_n21569_), .A1(\asqrt[6] ), .B0(new_n21571_), .Y(new_n21572_));
  NOR3X1   g21380(.A(new_n21566_), .B(new_n21558_), .C(\asqrt[19] ), .Y(new_n21573_));
  OAI21X1  g21381(.A0(new_n21573_), .A1(new_n21572_), .B0(new_n21567_), .Y(new_n21574_));
  AND2X1   g21382(.A(new_n21574_), .B(\asqrt[20] ), .Y(new_n21575_));
  INVX1    g21383(.A(new_n21572_), .Y(new_n21576_));
  AND2X1   g21384(.A(new_n21564_), .B(\asqrt[17] ), .Y(new_n21577_));
  NAND2X1  g21385(.A(new_n21537_), .B(new_n21536_), .Y(new_n21578_));
  AND2X1   g21386(.A(new_n21555_), .B(new_n14165_), .Y(new_n21579_));
  AOI21X1  g21387(.A0(new_n21579_), .A1(new_n21578_), .B0(new_n21545_), .Y(new_n21580_));
  OAI21X1  g21388(.A0(new_n21580_), .A1(new_n21577_), .B0(\asqrt[18] ), .Y(new_n21581_));
  INVX1    g21389(.A(new_n21562_), .Y(new_n21582_));
  OAI21X1  g21390(.A0(new_n21538_), .A1(new_n14165_), .B0(new_n13571_), .Y(new_n21583_));
  OAI21X1  g21391(.A0(new_n21583_), .A1(new_n21580_), .B0(new_n21582_), .Y(new_n21584_));
  NAND3X1  g21392(.A(new_n21584_), .B(new_n21581_), .C(new_n13000_), .Y(new_n21585_));
  NAND2X1  g21393(.A(new_n21585_), .B(new_n21576_), .Y(new_n21586_));
  AND2X1   g21394(.A(new_n20847_), .B(new_n20839_), .Y(new_n21587_));
  NOR3X1   g21395(.A(new_n21587_), .B(new_n20864_), .C(new_n20840_), .Y(new_n21588_));
  NOR3X1   g21396(.A(new_n21393_), .B(new_n21587_), .C(new_n20840_), .Y(new_n21589_));
  NOR2X1   g21397(.A(new_n21589_), .B(new_n20845_), .Y(new_n21590_));
  AOI21X1  g21398(.A0(new_n21588_), .A1(\asqrt[6] ), .B0(new_n21590_), .Y(new_n21591_));
  AND2X1   g21399(.A(new_n21567_), .B(new_n12447_), .Y(new_n21592_));
  AOI21X1  g21400(.A0(new_n21592_), .A1(new_n21586_), .B0(new_n21591_), .Y(new_n21593_));
  OAI21X1  g21401(.A0(new_n21593_), .A1(new_n21575_), .B0(\asqrt[21] ), .Y(new_n21594_));
  NAND4X1  g21402(.A(\asqrt[6] ), .B(new_n20867_), .C(new_n20854_), .D(new_n20849_), .Y(new_n21595_));
  NAND2X1  g21403(.A(new_n20867_), .B(new_n20849_), .Y(new_n21596_));
  OAI21X1  g21404(.A0(new_n21596_), .A1(new_n21393_), .B0(new_n20858_), .Y(new_n21597_));
  AND2X1   g21405(.A(new_n21597_), .B(new_n21595_), .Y(new_n21598_));
  INVX1    g21406(.A(new_n21598_), .Y(new_n21599_));
  AOI21X1  g21407(.A0(new_n21584_), .A1(new_n21581_), .B0(new_n13000_), .Y(new_n21600_));
  AOI21X1  g21408(.A0(new_n21585_), .A1(new_n21576_), .B0(new_n21600_), .Y(new_n21601_));
  OAI21X1  g21409(.A0(new_n21601_), .A1(new_n12447_), .B0(new_n11896_), .Y(new_n21602_));
  OAI21X1  g21410(.A0(new_n21602_), .A1(new_n21593_), .B0(new_n21599_), .Y(new_n21603_));
  AOI21X1  g21411(.A0(new_n21603_), .A1(new_n21594_), .B0(new_n11362_), .Y(new_n21604_));
  AOI21X1  g21412(.A0(new_n20874_), .A1(new_n20868_), .B0(new_n20912_), .Y(new_n21605_));
  AND2X1   g21413(.A(new_n21605_), .B(new_n20910_), .Y(new_n21606_));
  AOI22X1  g21414(.A0(new_n20874_), .A1(new_n20868_), .B0(new_n20856_), .B1(\asqrt[21] ), .Y(new_n21607_));
  AOI21X1  g21415(.A0(new_n21607_), .A1(\asqrt[6] ), .B0(new_n20872_), .Y(new_n21608_));
  AOI21X1  g21416(.A0(new_n21606_), .A1(\asqrt[6] ), .B0(new_n21608_), .Y(new_n21609_));
  INVX1    g21417(.A(new_n21609_), .Y(new_n21610_));
  NAND3X1  g21418(.A(new_n21603_), .B(new_n21594_), .C(new_n11362_), .Y(new_n21611_));
  AOI21X1  g21419(.A0(new_n21611_), .A1(new_n21610_), .B0(new_n21604_), .Y(new_n21612_));
  OR2X1    g21420(.A(new_n21612_), .B(new_n10849_), .Y(new_n21613_));
  AND2X1   g21421(.A(new_n21611_), .B(new_n21610_), .Y(new_n21614_));
  AND2X1   g21422(.A(new_n20916_), .B(new_n20914_), .Y(new_n21615_));
  NOR3X1   g21423(.A(new_n21615_), .B(new_n20882_), .C(new_n20915_), .Y(new_n21616_));
  NOR3X1   g21424(.A(new_n21393_), .B(new_n21615_), .C(new_n20915_), .Y(new_n21617_));
  NOR2X1   g21425(.A(new_n21617_), .B(new_n20881_), .Y(new_n21618_));
  AOI21X1  g21426(.A0(new_n21616_), .A1(\asqrt[6] ), .B0(new_n21618_), .Y(new_n21619_));
  INVX1    g21427(.A(new_n21619_), .Y(new_n21620_));
  OR2X1    g21428(.A(new_n21601_), .B(new_n12447_), .Y(new_n21621_));
  AND2X1   g21429(.A(new_n21585_), .B(new_n21576_), .Y(new_n21622_));
  INVX1    g21430(.A(new_n21591_), .Y(new_n21623_));
  NAND2X1  g21431(.A(new_n21567_), .B(new_n12447_), .Y(new_n21624_));
  OAI21X1  g21432(.A0(new_n21624_), .A1(new_n21622_), .B0(new_n21623_), .Y(new_n21625_));
  AOI21X1  g21433(.A0(new_n21625_), .A1(new_n21621_), .B0(new_n11896_), .Y(new_n21626_));
  AOI21X1  g21434(.A0(new_n21574_), .A1(\asqrt[20] ), .B0(\asqrt[21] ), .Y(new_n21627_));
  AOI21X1  g21435(.A0(new_n21627_), .A1(new_n21625_), .B0(new_n21598_), .Y(new_n21628_));
  OAI21X1  g21436(.A0(new_n21628_), .A1(new_n21626_), .B0(\asqrt[22] ), .Y(new_n21629_));
  NAND2X1  g21437(.A(new_n21629_), .B(new_n10849_), .Y(new_n21630_));
  OAI21X1  g21438(.A0(new_n21630_), .A1(new_n21614_), .B0(new_n21620_), .Y(new_n21631_));
  AOI21X1  g21439(.A0(new_n21631_), .A1(new_n21613_), .B0(new_n10332_), .Y(new_n21632_));
  NAND4X1  g21440(.A(\asqrt[6] ), .B(new_n20893_), .C(new_n20891_), .D(new_n20918_), .Y(new_n21633_));
  NAND2X1  g21441(.A(new_n20893_), .B(new_n20918_), .Y(new_n21634_));
  OAI21X1  g21442(.A0(new_n21634_), .A1(new_n21393_), .B0(new_n20892_), .Y(new_n21635_));
  AND2X1   g21443(.A(new_n21635_), .B(new_n21633_), .Y(new_n21636_));
  NOR3X1   g21444(.A(new_n21628_), .B(new_n21626_), .C(\asqrt[22] ), .Y(new_n21637_));
  OAI21X1  g21445(.A0(new_n21637_), .A1(new_n21609_), .B0(new_n21629_), .Y(new_n21638_));
  AOI21X1  g21446(.A0(new_n21638_), .A1(\asqrt[23] ), .B0(\asqrt[24] ), .Y(new_n21639_));
  AOI21X1  g21447(.A0(new_n21639_), .A1(new_n21631_), .B0(new_n21636_), .Y(new_n21640_));
  OAI21X1  g21448(.A0(new_n21640_), .A1(new_n21632_), .B0(\asqrt[25] ), .Y(new_n21641_));
  AND2X1   g21449(.A(new_n20948_), .B(new_n20947_), .Y(new_n21642_));
  NOR3X1   g21450(.A(new_n21642_), .B(new_n20901_), .C(new_n20946_), .Y(new_n21643_));
  NOR3X1   g21451(.A(new_n21393_), .B(new_n21642_), .C(new_n20946_), .Y(new_n21644_));
  NOR2X1   g21452(.A(new_n21644_), .B(new_n20900_), .Y(new_n21645_));
  AOI21X1  g21453(.A0(new_n21643_), .A1(\asqrt[6] ), .B0(new_n21645_), .Y(new_n21646_));
  NOR3X1   g21454(.A(new_n21640_), .B(new_n21632_), .C(\asqrt[25] ), .Y(new_n21647_));
  OAI21X1  g21455(.A0(new_n21647_), .A1(new_n21646_), .B0(new_n21641_), .Y(new_n21648_));
  AND2X1   g21456(.A(new_n21648_), .B(\asqrt[26] ), .Y(new_n21649_));
  INVX1    g21457(.A(new_n21646_), .Y(new_n21650_));
  AND2X1   g21458(.A(new_n21638_), .B(\asqrt[23] ), .Y(new_n21651_));
  NAND2X1  g21459(.A(new_n21611_), .B(new_n21610_), .Y(new_n21652_));
  AND2X1   g21460(.A(new_n21629_), .B(new_n10849_), .Y(new_n21653_));
  AOI21X1  g21461(.A0(new_n21653_), .A1(new_n21652_), .B0(new_n21619_), .Y(new_n21654_));
  OAI21X1  g21462(.A0(new_n21654_), .A1(new_n21651_), .B0(\asqrt[24] ), .Y(new_n21655_));
  INVX1    g21463(.A(new_n21636_), .Y(new_n21656_));
  OAI21X1  g21464(.A0(new_n21612_), .A1(new_n10849_), .B0(new_n10332_), .Y(new_n21657_));
  OAI21X1  g21465(.A0(new_n21657_), .A1(new_n21654_), .B0(new_n21656_), .Y(new_n21658_));
  NAND3X1  g21466(.A(new_n21658_), .B(new_n21655_), .C(new_n9833_), .Y(new_n21659_));
  NAND2X1  g21467(.A(new_n21659_), .B(new_n21650_), .Y(new_n21660_));
  AND2X1   g21468(.A(new_n20921_), .B(new_n20903_), .Y(new_n21661_));
  NOR3X1   g21469(.A(new_n21661_), .B(new_n20951_), .C(new_n20904_), .Y(new_n21662_));
  NOR3X1   g21470(.A(new_n21393_), .B(new_n21661_), .C(new_n20904_), .Y(new_n21663_));
  NOR2X1   g21471(.A(new_n21663_), .B(new_n20909_), .Y(new_n21664_));
  AOI21X1  g21472(.A0(new_n21662_), .A1(\asqrt[6] ), .B0(new_n21664_), .Y(new_n21665_));
  AND2X1   g21473(.A(new_n21641_), .B(new_n9353_), .Y(new_n21666_));
  AOI21X1  g21474(.A0(new_n21666_), .A1(new_n21660_), .B0(new_n21665_), .Y(new_n21667_));
  OAI21X1  g21475(.A0(new_n21667_), .A1(new_n21649_), .B0(\asqrt[27] ), .Y(new_n21668_));
  NAND4X1  g21476(.A(\asqrt[6] ), .B(new_n20956_), .C(new_n20928_), .D(new_n20923_), .Y(new_n21669_));
  OR2X1    g21477(.A(new_n20929_), .B(new_n20954_), .Y(new_n21670_));
  OAI21X1  g21478(.A0(new_n21670_), .A1(new_n21393_), .B0(new_n20955_), .Y(new_n21671_));
  AND2X1   g21479(.A(new_n21671_), .B(new_n21669_), .Y(new_n21672_));
  INVX1    g21480(.A(new_n21672_), .Y(new_n21673_));
  AOI21X1  g21481(.A0(new_n21658_), .A1(new_n21655_), .B0(new_n9833_), .Y(new_n21674_));
  AOI21X1  g21482(.A0(new_n21659_), .A1(new_n21650_), .B0(new_n21674_), .Y(new_n21675_));
  OAI21X1  g21483(.A0(new_n21675_), .A1(new_n9353_), .B0(new_n8874_), .Y(new_n21676_));
  OAI21X1  g21484(.A0(new_n21676_), .A1(new_n21667_), .B0(new_n21673_), .Y(new_n21677_));
  AOI21X1  g21485(.A0(new_n21677_), .A1(new_n21668_), .B0(new_n8412_), .Y(new_n21678_));
  AOI21X1  g21486(.A0(new_n20937_), .A1(new_n20932_), .B0(new_n20972_), .Y(new_n21679_));
  AND2X1   g21487(.A(new_n21679_), .B(new_n20970_), .Y(new_n21680_));
  AOI22X1  g21488(.A0(new_n20937_), .A1(new_n20932_), .B0(new_n20930_), .B1(\asqrt[27] ), .Y(new_n21681_));
  AOI21X1  g21489(.A0(new_n21681_), .A1(\asqrt[6] ), .B0(new_n20936_), .Y(new_n21682_));
  AOI21X1  g21490(.A0(new_n21680_), .A1(\asqrt[6] ), .B0(new_n21682_), .Y(new_n21683_));
  INVX1    g21491(.A(new_n21683_), .Y(new_n21684_));
  NAND3X1  g21492(.A(new_n21677_), .B(new_n21668_), .C(new_n8412_), .Y(new_n21685_));
  AOI21X1  g21493(.A0(new_n21685_), .A1(new_n21684_), .B0(new_n21678_), .Y(new_n21686_));
  OR2X1    g21494(.A(new_n21686_), .B(new_n7970_), .Y(new_n21687_));
  AND2X1   g21495(.A(new_n21685_), .B(new_n21684_), .Y(new_n21688_));
  AND2X1   g21496(.A(new_n20976_), .B(new_n20974_), .Y(new_n21689_));
  NOR3X1   g21497(.A(new_n21689_), .B(new_n20945_), .C(new_n20975_), .Y(new_n21690_));
  NOR3X1   g21498(.A(new_n21393_), .B(new_n21689_), .C(new_n20975_), .Y(new_n21691_));
  NOR2X1   g21499(.A(new_n21691_), .B(new_n20944_), .Y(new_n21692_));
  AOI21X1  g21500(.A0(new_n21690_), .A1(\asqrt[6] ), .B0(new_n21692_), .Y(new_n21693_));
  INVX1    g21501(.A(new_n21693_), .Y(new_n21694_));
  OR2X1    g21502(.A(new_n21675_), .B(new_n9353_), .Y(new_n21695_));
  AND2X1   g21503(.A(new_n21659_), .B(new_n21650_), .Y(new_n21696_));
  INVX1    g21504(.A(new_n21665_), .Y(new_n21697_));
  NAND2X1  g21505(.A(new_n21641_), .B(new_n9353_), .Y(new_n21698_));
  OAI21X1  g21506(.A0(new_n21698_), .A1(new_n21696_), .B0(new_n21697_), .Y(new_n21699_));
  AOI21X1  g21507(.A0(new_n21699_), .A1(new_n21695_), .B0(new_n8874_), .Y(new_n21700_));
  AOI21X1  g21508(.A0(new_n21648_), .A1(\asqrt[26] ), .B0(\asqrt[27] ), .Y(new_n21701_));
  AOI21X1  g21509(.A0(new_n21701_), .A1(new_n21699_), .B0(new_n21672_), .Y(new_n21702_));
  OAI21X1  g21510(.A0(new_n21702_), .A1(new_n21700_), .B0(\asqrt[28] ), .Y(new_n21703_));
  NAND2X1  g21511(.A(new_n21703_), .B(new_n7970_), .Y(new_n21704_));
  OAI21X1  g21512(.A0(new_n21704_), .A1(new_n21688_), .B0(new_n21694_), .Y(new_n21705_));
  AOI21X1  g21513(.A0(new_n21705_), .A1(new_n21687_), .B0(new_n7527_), .Y(new_n21706_));
  OR4X1    g21514(.A(new_n21393_), .B(new_n20978_), .C(new_n20966_), .D(new_n20960_), .Y(new_n21707_));
  OR2X1    g21515(.A(new_n20978_), .B(new_n20960_), .Y(new_n21708_));
  OAI21X1  g21516(.A0(new_n21708_), .A1(new_n21393_), .B0(new_n20966_), .Y(new_n21709_));
  AND2X1   g21517(.A(new_n21709_), .B(new_n21707_), .Y(new_n21710_));
  NOR3X1   g21518(.A(new_n21702_), .B(new_n21700_), .C(\asqrt[28] ), .Y(new_n21711_));
  OAI21X1  g21519(.A0(new_n21711_), .A1(new_n21683_), .B0(new_n21703_), .Y(new_n21712_));
  AOI21X1  g21520(.A0(new_n21712_), .A1(\asqrt[29] ), .B0(\asqrt[30] ), .Y(new_n21713_));
  AOI21X1  g21521(.A0(new_n21713_), .A1(new_n21705_), .B0(new_n21710_), .Y(new_n21714_));
  OAI21X1  g21522(.A0(new_n21714_), .A1(new_n21706_), .B0(\asqrt[31] ), .Y(new_n21715_));
  AND2X1   g21523(.A(new_n21022_), .B(new_n21021_), .Y(new_n21716_));
  NOR3X1   g21524(.A(new_n21716_), .B(new_n20984_), .C(new_n21020_), .Y(new_n21717_));
  NOR3X1   g21525(.A(new_n21393_), .B(new_n21716_), .C(new_n21020_), .Y(new_n21718_));
  NOR2X1   g21526(.A(new_n21718_), .B(new_n20983_), .Y(new_n21719_));
  AOI21X1  g21527(.A0(new_n21717_), .A1(\asqrt[6] ), .B0(new_n21719_), .Y(new_n21720_));
  NOR3X1   g21528(.A(new_n21714_), .B(new_n21706_), .C(\asqrt[31] ), .Y(new_n21721_));
  OAI21X1  g21529(.A0(new_n21721_), .A1(new_n21720_), .B0(new_n21715_), .Y(new_n21722_));
  AND2X1   g21530(.A(new_n21722_), .B(\asqrt[32] ), .Y(new_n21723_));
  OR2X1    g21531(.A(new_n21721_), .B(new_n21720_), .Y(new_n21724_));
  AND2X1   g21532(.A(new_n20995_), .B(new_n20987_), .Y(new_n21725_));
  NOR3X1   g21533(.A(new_n21725_), .B(new_n21025_), .C(new_n20988_), .Y(new_n21726_));
  NOR3X1   g21534(.A(new_n21393_), .B(new_n21725_), .C(new_n20988_), .Y(new_n21727_));
  NOR2X1   g21535(.A(new_n21727_), .B(new_n20993_), .Y(new_n21728_));
  AOI21X1  g21536(.A0(new_n21726_), .A1(\asqrt[6] ), .B0(new_n21728_), .Y(new_n21729_));
  AND2X1   g21537(.A(new_n21715_), .B(new_n6699_), .Y(new_n21730_));
  AOI21X1  g21538(.A0(new_n21730_), .A1(new_n21724_), .B0(new_n21729_), .Y(new_n21731_));
  OAI21X1  g21539(.A0(new_n21731_), .A1(new_n21723_), .B0(\asqrt[33] ), .Y(new_n21732_));
  OR4X1    g21540(.A(new_n21393_), .B(new_n21003_), .C(new_n21029_), .D(new_n21028_), .Y(new_n21733_));
  OR2X1    g21541(.A(new_n21003_), .B(new_n21028_), .Y(new_n21734_));
  OAI21X1  g21542(.A0(new_n21734_), .A1(new_n21393_), .B0(new_n21029_), .Y(new_n21735_));
  AND2X1   g21543(.A(new_n21735_), .B(new_n21733_), .Y(new_n21736_));
  INVX1    g21544(.A(new_n21736_), .Y(new_n21737_));
  AND2X1   g21545(.A(new_n21712_), .B(\asqrt[29] ), .Y(new_n21738_));
  NAND2X1  g21546(.A(new_n21685_), .B(new_n21684_), .Y(new_n21739_));
  AND2X1   g21547(.A(new_n21703_), .B(new_n7970_), .Y(new_n21740_));
  AOI21X1  g21548(.A0(new_n21740_), .A1(new_n21739_), .B0(new_n21693_), .Y(new_n21741_));
  OAI21X1  g21549(.A0(new_n21741_), .A1(new_n21738_), .B0(\asqrt[30] ), .Y(new_n21742_));
  INVX1    g21550(.A(new_n21710_), .Y(new_n21743_));
  OAI21X1  g21551(.A0(new_n21686_), .A1(new_n7970_), .B0(new_n7527_), .Y(new_n21744_));
  OAI21X1  g21552(.A0(new_n21744_), .A1(new_n21741_), .B0(new_n21743_), .Y(new_n21745_));
  AOI21X1  g21553(.A0(new_n21745_), .A1(new_n21742_), .B0(new_n7103_), .Y(new_n21746_));
  INVX1    g21554(.A(new_n21720_), .Y(new_n21747_));
  NAND3X1  g21555(.A(new_n21745_), .B(new_n21742_), .C(new_n7103_), .Y(new_n21748_));
  AOI21X1  g21556(.A0(new_n21748_), .A1(new_n21747_), .B0(new_n21746_), .Y(new_n21749_));
  OAI21X1  g21557(.A0(new_n21749_), .A1(new_n6699_), .B0(new_n6294_), .Y(new_n21750_));
  OAI21X1  g21558(.A0(new_n21750_), .A1(new_n21731_), .B0(new_n21737_), .Y(new_n21751_));
  AOI21X1  g21559(.A0(new_n21751_), .A1(new_n21732_), .B0(new_n5941_), .Y(new_n21752_));
  AOI21X1  g21560(.A0(new_n21011_), .A1(new_n21006_), .B0(new_n21046_), .Y(new_n21753_));
  AND2X1   g21561(.A(new_n21753_), .B(new_n21044_), .Y(new_n21754_));
  AOI22X1  g21562(.A0(new_n21011_), .A1(new_n21006_), .B0(new_n21004_), .B1(\asqrt[33] ), .Y(new_n21755_));
  AOI21X1  g21563(.A0(new_n21755_), .A1(\asqrt[6] ), .B0(new_n21010_), .Y(new_n21756_));
  AOI21X1  g21564(.A0(new_n21754_), .A1(\asqrt[6] ), .B0(new_n21756_), .Y(new_n21757_));
  INVX1    g21565(.A(new_n21757_), .Y(new_n21758_));
  NAND3X1  g21566(.A(new_n21751_), .B(new_n21732_), .C(new_n5941_), .Y(new_n21759_));
  AOI21X1  g21567(.A0(new_n21759_), .A1(new_n21758_), .B0(new_n21752_), .Y(new_n21760_));
  OR2X1    g21568(.A(new_n21760_), .B(new_n5541_), .Y(new_n21761_));
  OR2X1    g21569(.A(new_n21749_), .B(new_n6699_), .Y(new_n21762_));
  NOR2X1   g21570(.A(new_n21721_), .B(new_n21720_), .Y(new_n21763_));
  INVX1    g21571(.A(new_n21729_), .Y(new_n21764_));
  NAND2X1  g21572(.A(new_n21715_), .B(new_n6699_), .Y(new_n21765_));
  OAI21X1  g21573(.A0(new_n21765_), .A1(new_n21763_), .B0(new_n21764_), .Y(new_n21766_));
  AOI21X1  g21574(.A0(new_n21766_), .A1(new_n21762_), .B0(new_n6294_), .Y(new_n21767_));
  AOI21X1  g21575(.A0(new_n21722_), .A1(\asqrt[32] ), .B0(\asqrt[33] ), .Y(new_n21768_));
  AOI21X1  g21576(.A0(new_n21768_), .A1(new_n21766_), .B0(new_n21736_), .Y(new_n21769_));
  NOR3X1   g21577(.A(new_n21769_), .B(new_n21767_), .C(\asqrt[34] ), .Y(new_n21770_));
  NOR2X1   g21578(.A(new_n21770_), .B(new_n21757_), .Y(new_n21771_));
  AND2X1   g21579(.A(new_n21050_), .B(new_n21048_), .Y(new_n21772_));
  NOR3X1   g21580(.A(new_n21772_), .B(new_n21019_), .C(new_n21049_), .Y(new_n21773_));
  NOR3X1   g21581(.A(new_n21393_), .B(new_n21772_), .C(new_n21049_), .Y(new_n21774_));
  NOR2X1   g21582(.A(new_n21774_), .B(new_n21018_), .Y(new_n21775_));
  AOI21X1  g21583(.A0(new_n21773_), .A1(\asqrt[6] ), .B0(new_n21775_), .Y(new_n21776_));
  INVX1    g21584(.A(new_n21776_), .Y(new_n21777_));
  OAI21X1  g21585(.A0(new_n21769_), .A1(new_n21767_), .B0(\asqrt[34] ), .Y(new_n21778_));
  NAND2X1  g21586(.A(new_n21778_), .B(new_n5541_), .Y(new_n21779_));
  OAI21X1  g21587(.A0(new_n21779_), .A1(new_n21771_), .B0(new_n21777_), .Y(new_n21780_));
  AOI21X1  g21588(.A0(new_n21780_), .A1(new_n21761_), .B0(new_n5176_), .Y(new_n21781_));
  OR4X1    g21589(.A(new_n21393_), .B(new_n21052_), .C(new_n21040_), .D(new_n21034_), .Y(new_n21782_));
  OR2X1    g21590(.A(new_n21052_), .B(new_n21034_), .Y(new_n21783_));
  OAI21X1  g21591(.A0(new_n21783_), .A1(new_n21393_), .B0(new_n21040_), .Y(new_n21784_));
  AND2X1   g21592(.A(new_n21784_), .B(new_n21782_), .Y(new_n21785_));
  OAI21X1  g21593(.A0(new_n21770_), .A1(new_n21757_), .B0(new_n21778_), .Y(new_n21786_));
  AOI21X1  g21594(.A0(new_n21786_), .A1(\asqrt[35] ), .B0(\asqrt[36] ), .Y(new_n21787_));
  AOI21X1  g21595(.A0(new_n21787_), .A1(new_n21780_), .B0(new_n21785_), .Y(new_n21788_));
  OAI21X1  g21596(.A0(new_n21788_), .A1(new_n21781_), .B0(\asqrt[37] ), .Y(new_n21789_));
  AND2X1   g21597(.A(new_n21096_), .B(new_n21095_), .Y(new_n21790_));
  NOR3X1   g21598(.A(new_n21790_), .B(new_n21058_), .C(new_n21094_), .Y(new_n21791_));
  NOR3X1   g21599(.A(new_n21393_), .B(new_n21790_), .C(new_n21094_), .Y(new_n21792_));
  NOR2X1   g21600(.A(new_n21792_), .B(new_n21057_), .Y(new_n21793_));
  AOI21X1  g21601(.A0(new_n21791_), .A1(\asqrt[6] ), .B0(new_n21793_), .Y(new_n21794_));
  NOR3X1   g21602(.A(new_n21788_), .B(new_n21781_), .C(\asqrt[37] ), .Y(new_n21795_));
  OAI21X1  g21603(.A0(new_n21795_), .A1(new_n21794_), .B0(new_n21789_), .Y(new_n21796_));
  AND2X1   g21604(.A(new_n21796_), .B(\asqrt[38] ), .Y(new_n21797_));
  OR2X1    g21605(.A(new_n21795_), .B(new_n21794_), .Y(new_n21798_));
  AND2X1   g21606(.A(new_n21069_), .B(new_n21061_), .Y(new_n21799_));
  NOR3X1   g21607(.A(new_n21799_), .B(new_n21099_), .C(new_n21062_), .Y(new_n21800_));
  NOR3X1   g21608(.A(new_n21393_), .B(new_n21799_), .C(new_n21062_), .Y(new_n21801_));
  NOR2X1   g21609(.A(new_n21801_), .B(new_n21067_), .Y(new_n21802_));
  AOI21X1  g21610(.A0(new_n21800_), .A1(\asqrt[6] ), .B0(new_n21802_), .Y(new_n21803_));
  AND2X1   g21611(.A(new_n21789_), .B(new_n4493_), .Y(new_n21804_));
  AOI21X1  g21612(.A0(new_n21804_), .A1(new_n21798_), .B0(new_n21803_), .Y(new_n21805_));
  OAI21X1  g21613(.A0(new_n21805_), .A1(new_n21797_), .B0(\asqrt[39] ), .Y(new_n21806_));
  OR4X1    g21614(.A(new_n21393_), .B(new_n21077_), .C(new_n21103_), .D(new_n21102_), .Y(new_n21807_));
  OR2X1    g21615(.A(new_n21077_), .B(new_n21102_), .Y(new_n21808_));
  OAI21X1  g21616(.A0(new_n21808_), .A1(new_n21393_), .B0(new_n21103_), .Y(new_n21809_));
  AND2X1   g21617(.A(new_n21809_), .B(new_n21807_), .Y(new_n21810_));
  INVX1    g21618(.A(new_n21810_), .Y(new_n21811_));
  AND2X1   g21619(.A(new_n21786_), .B(\asqrt[35] ), .Y(new_n21812_));
  OR2X1    g21620(.A(new_n21770_), .B(new_n21757_), .Y(new_n21813_));
  AND2X1   g21621(.A(new_n21778_), .B(new_n5541_), .Y(new_n21814_));
  AOI21X1  g21622(.A0(new_n21814_), .A1(new_n21813_), .B0(new_n21776_), .Y(new_n21815_));
  OAI21X1  g21623(.A0(new_n21815_), .A1(new_n21812_), .B0(\asqrt[36] ), .Y(new_n21816_));
  INVX1    g21624(.A(new_n21785_), .Y(new_n21817_));
  OAI21X1  g21625(.A0(new_n21760_), .A1(new_n5541_), .B0(new_n5176_), .Y(new_n21818_));
  OAI21X1  g21626(.A0(new_n21818_), .A1(new_n21815_), .B0(new_n21817_), .Y(new_n21819_));
  AOI21X1  g21627(.A0(new_n21819_), .A1(new_n21816_), .B0(new_n4826_), .Y(new_n21820_));
  INVX1    g21628(.A(new_n21794_), .Y(new_n21821_));
  NAND3X1  g21629(.A(new_n21819_), .B(new_n21816_), .C(new_n4826_), .Y(new_n21822_));
  AOI21X1  g21630(.A0(new_n21822_), .A1(new_n21821_), .B0(new_n21820_), .Y(new_n21823_));
  OAI21X1  g21631(.A0(new_n21823_), .A1(new_n4493_), .B0(new_n4165_), .Y(new_n21824_));
  OAI21X1  g21632(.A0(new_n21824_), .A1(new_n21805_), .B0(new_n21811_), .Y(new_n21825_));
  AOI21X1  g21633(.A0(new_n21825_), .A1(new_n21806_), .B0(new_n3863_), .Y(new_n21826_));
  AOI21X1  g21634(.A0(new_n21085_), .A1(new_n21080_), .B0(new_n21120_), .Y(new_n21827_));
  AND2X1   g21635(.A(new_n21827_), .B(new_n21118_), .Y(new_n21828_));
  AOI22X1  g21636(.A0(new_n21085_), .A1(new_n21080_), .B0(new_n21078_), .B1(\asqrt[39] ), .Y(new_n21829_));
  AOI21X1  g21637(.A0(new_n21829_), .A1(\asqrt[6] ), .B0(new_n21084_), .Y(new_n21830_));
  AOI21X1  g21638(.A0(new_n21828_), .A1(\asqrt[6] ), .B0(new_n21830_), .Y(new_n21831_));
  INVX1    g21639(.A(new_n21831_), .Y(new_n21832_));
  NAND3X1  g21640(.A(new_n21825_), .B(new_n21806_), .C(new_n3863_), .Y(new_n21833_));
  AOI21X1  g21641(.A0(new_n21833_), .A1(new_n21832_), .B0(new_n21826_), .Y(new_n21834_));
  OR2X1    g21642(.A(new_n21834_), .B(new_n3564_), .Y(new_n21835_));
  OR2X1    g21643(.A(new_n21823_), .B(new_n4493_), .Y(new_n21836_));
  NOR2X1   g21644(.A(new_n21795_), .B(new_n21794_), .Y(new_n21837_));
  INVX1    g21645(.A(new_n21803_), .Y(new_n21838_));
  NAND2X1  g21646(.A(new_n21789_), .B(new_n4493_), .Y(new_n21839_));
  OAI21X1  g21647(.A0(new_n21839_), .A1(new_n21837_), .B0(new_n21838_), .Y(new_n21840_));
  AOI21X1  g21648(.A0(new_n21840_), .A1(new_n21836_), .B0(new_n4165_), .Y(new_n21841_));
  AOI21X1  g21649(.A0(new_n21796_), .A1(\asqrt[38] ), .B0(\asqrt[39] ), .Y(new_n21842_));
  AOI21X1  g21650(.A0(new_n21842_), .A1(new_n21840_), .B0(new_n21810_), .Y(new_n21843_));
  NOR3X1   g21651(.A(new_n21843_), .B(new_n21841_), .C(\asqrt[40] ), .Y(new_n21844_));
  NOR2X1   g21652(.A(new_n21844_), .B(new_n21831_), .Y(new_n21845_));
  AND2X1   g21653(.A(new_n21124_), .B(new_n21122_), .Y(new_n21846_));
  NOR3X1   g21654(.A(new_n21846_), .B(new_n21093_), .C(new_n21123_), .Y(new_n21847_));
  NOR3X1   g21655(.A(new_n21393_), .B(new_n21846_), .C(new_n21123_), .Y(new_n21848_));
  NOR2X1   g21656(.A(new_n21848_), .B(new_n21092_), .Y(new_n21849_));
  AOI21X1  g21657(.A0(new_n21847_), .A1(\asqrt[6] ), .B0(new_n21849_), .Y(new_n21850_));
  INVX1    g21658(.A(new_n21850_), .Y(new_n21851_));
  OAI21X1  g21659(.A0(new_n21843_), .A1(new_n21841_), .B0(\asqrt[40] ), .Y(new_n21852_));
  NAND2X1  g21660(.A(new_n21852_), .B(new_n3564_), .Y(new_n21853_));
  OAI21X1  g21661(.A0(new_n21853_), .A1(new_n21845_), .B0(new_n21851_), .Y(new_n21854_));
  AOI21X1  g21662(.A0(new_n21854_), .A1(new_n21835_), .B0(new_n3276_), .Y(new_n21855_));
  OR4X1    g21663(.A(new_n21393_), .B(new_n21126_), .C(new_n21114_), .D(new_n21108_), .Y(new_n21856_));
  OR2X1    g21664(.A(new_n21126_), .B(new_n21108_), .Y(new_n21857_));
  OAI21X1  g21665(.A0(new_n21857_), .A1(new_n21393_), .B0(new_n21114_), .Y(new_n21858_));
  AND2X1   g21666(.A(new_n21858_), .B(new_n21856_), .Y(new_n21859_));
  OAI21X1  g21667(.A0(new_n21844_), .A1(new_n21831_), .B0(new_n21852_), .Y(new_n21860_));
  AOI21X1  g21668(.A0(new_n21860_), .A1(\asqrt[41] ), .B0(\asqrt[42] ), .Y(new_n21861_));
  AOI21X1  g21669(.A0(new_n21861_), .A1(new_n21854_), .B0(new_n21859_), .Y(new_n21862_));
  OAI21X1  g21670(.A0(new_n21862_), .A1(new_n21855_), .B0(\asqrt[43] ), .Y(new_n21863_));
  AND2X1   g21671(.A(new_n21170_), .B(new_n21169_), .Y(new_n21864_));
  NOR3X1   g21672(.A(new_n21864_), .B(new_n21132_), .C(new_n21168_), .Y(new_n21865_));
  NOR3X1   g21673(.A(new_n21393_), .B(new_n21864_), .C(new_n21168_), .Y(new_n21866_));
  NOR2X1   g21674(.A(new_n21866_), .B(new_n21131_), .Y(new_n21867_));
  AOI21X1  g21675(.A0(new_n21865_), .A1(\asqrt[6] ), .B0(new_n21867_), .Y(new_n21868_));
  NOR3X1   g21676(.A(new_n21862_), .B(new_n21855_), .C(\asqrt[43] ), .Y(new_n21869_));
  OAI21X1  g21677(.A0(new_n21869_), .A1(new_n21868_), .B0(new_n21863_), .Y(new_n21870_));
  AND2X1   g21678(.A(new_n21870_), .B(\asqrt[44] ), .Y(new_n21871_));
  OR2X1    g21679(.A(new_n21869_), .B(new_n21868_), .Y(new_n21872_));
  AND2X1   g21680(.A(new_n21143_), .B(new_n21135_), .Y(new_n21873_));
  NOR3X1   g21681(.A(new_n21873_), .B(new_n21173_), .C(new_n21136_), .Y(new_n21874_));
  NOR3X1   g21682(.A(new_n21393_), .B(new_n21873_), .C(new_n21136_), .Y(new_n21875_));
  NOR2X1   g21683(.A(new_n21875_), .B(new_n21141_), .Y(new_n21876_));
  AOI21X1  g21684(.A0(new_n21874_), .A1(\asqrt[6] ), .B0(new_n21876_), .Y(new_n21877_));
  AND2X1   g21685(.A(new_n21863_), .B(new_n2769_), .Y(new_n21878_));
  AOI21X1  g21686(.A0(new_n21878_), .A1(new_n21872_), .B0(new_n21877_), .Y(new_n21879_));
  OAI21X1  g21687(.A0(new_n21879_), .A1(new_n21871_), .B0(\asqrt[45] ), .Y(new_n21880_));
  OR4X1    g21688(.A(new_n21393_), .B(new_n21151_), .C(new_n21177_), .D(new_n21176_), .Y(new_n21881_));
  OR2X1    g21689(.A(new_n21151_), .B(new_n21176_), .Y(new_n21882_));
  OAI21X1  g21690(.A0(new_n21882_), .A1(new_n21393_), .B0(new_n21177_), .Y(new_n21883_));
  AND2X1   g21691(.A(new_n21883_), .B(new_n21881_), .Y(new_n21884_));
  INVX1    g21692(.A(new_n21884_), .Y(new_n21885_));
  AND2X1   g21693(.A(new_n21860_), .B(\asqrt[41] ), .Y(new_n21886_));
  OR2X1    g21694(.A(new_n21844_), .B(new_n21831_), .Y(new_n21887_));
  AND2X1   g21695(.A(new_n21852_), .B(new_n3564_), .Y(new_n21888_));
  AOI21X1  g21696(.A0(new_n21888_), .A1(new_n21887_), .B0(new_n21850_), .Y(new_n21889_));
  OAI21X1  g21697(.A0(new_n21889_), .A1(new_n21886_), .B0(\asqrt[42] ), .Y(new_n21890_));
  INVX1    g21698(.A(new_n21859_), .Y(new_n21891_));
  OAI21X1  g21699(.A0(new_n21834_), .A1(new_n3564_), .B0(new_n3276_), .Y(new_n21892_));
  OAI21X1  g21700(.A0(new_n21892_), .A1(new_n21889_), .B0(new_n21891_), .Y(new_n21893_));
  AOI21X1  g21701(.A0(new_n21893_), .A1(new_n21890_), .B0(new_n3008_), .Y(new_n21894_));
  INVX1    g21702(.A(new_n21868_), .Y(new_n21895_));
  NAND3X1  g21703(.A(new_n21893_), .B(new_n21890_), .C(new_n3008_), .Y(new_n21896_));
  AOI21X1  g21704(.A0(new_n21896_), .A1(new_n21895_), .B0(new_n21894_), .Y(new_n21897_));
  OAI21X1  g21705(.A0(new_n21897_), .A1(new_n2769_), .B0(new_n2570_), .Y(new_n21898_));
  OAI21X1  g21706(.A0(new_n21898_), .A1(new_n21879_), .B0(new_n21885_), .Y(new_n21899_));
  AOI21X1  g21707(.A0(new_n21899_), .A1(new_n21880_), .B0(new_n2263_), .Y(new_n21900_));
  AOI21X1  g21708(.A0(new_n21159_), .A1(new_n21154_), .B0(new_n21194_), .Y(new_n21901_));
  AND2X1   g21709(.A(new_n21901_), .B(new_n21192_), .Y(new_n21902_));
  AOI22X1  g21710(.A0(new_n21159_), .A1(new_n21154_), .B0(new_n21152_), .B1(\asqrt[45] ), .Y(new_n21903_));
  AOI21X1  g21711(.A0(new_n21903_), .A1(\asqrt[6] ), .B0(new_n21158_), .Y(new_n21904_));
  AOI21X1  g21712(.A0(new_n21902_), .A1(\asqrt[6] ), .B0(new_n21904_), .Y(new_n21905_));
  INVX1    g21713(.A(new_n21905_), .Y(new_n21906_));
  NAND3X1  g21714(.A(new_n21899_), .B(new_n21880_), .C(new_n2263_), .Y(new_n21907_));
  AOI21X1  g21715(.A0(new_n21907_), .A1(new_n21906_), .B0(new_n21900_), .Y(new_n21908_));
  OR2X1    g21716(.A(new_n21908_), .B(new_n2040_), .Y(new_n21909_));
  OR2X1    g21717(.A(new_n21897_), .B(new_n2769_), .Y(new_n21910_));
  NOR2X1   g21718(.A(new_n21869_), .B(new_n21868_), .Y(new_n21911_));
  INVX1    g21719(.A(new_n21877_), .Y(new_n21912_));
  NAND2X1  g21720(.A(new_n21863_), .B(new_n2769_), .Y(new_n21913_));
  OAI21X1  g21721(.A0(new_n21913_), .A1(new_n21911_), .B0(new_n21912_), .Y(new_n21914_));
  AOI21X1  g21722(.A0(new_n21914_), .A1(new_n21910_), .B0(new_n2570_), .Y(new_n21915_));
  AOI21X1  g21723(.A0(new_n21870_), .A1(\asqrt[44] ), .B0(\asqrt[45] ), .Y(new_n21916_));
  AOI21X1  g21724(.A0(new_n21916_), .A1(new_n21914_), .B0(new_n21884_), .Y(new_n21917_));
  NOR3X1   g21725(.A(new_n21917_), .B(new_n21915_), .C(\asqrt[46] ), .Y(new_n21918_));
  NOR2X1   g21726(.A(new_n21918_), .B(new_n21905_), .Y(new_n21919_));
  AND2X1   g21727(.A(new_n21198_), .B(new_n21196_), .Y(new_n21920_));
  NOR3X1   g21728(.A(new_n21920_), .B(new_n21167_), .C(new_n21197_), .Y(new_n21921_));
  NOR3X1   g21729(.A(new_n21393_), .B(new_n21920_), .C(new_n21197_), .Y(new_n21922_));
  NOR2X1   g21730(.A(new_n21922_), .B(new_n21166_), .Y(new_n21923_));
  AOI21X1  g21731(.A0(new_n21921_), .A1(\asqrt[6] ), .B0(new_n21923_), .Y(new_n21924_));
  INVX1    g21732(.A(new_n21924_), .Y(new_n21925_));
  OAI21X1  g21733(.A0(new_n21917_), .A1(new_n21915_), .B0(\asqrt[46] ), .Y(new_n21926_));
  NAND2X1  g21734(.A(new_n21926_), .B(new_n2040_), .Y(new_n21927_));
  OAI21X1  g21735(.A0(new_n21927_), .A1(new_n21919_), .B0(new_n21925_), .Y(new_n21928_));
  AOI21X1  g21736(.A0(new_n21928_), .A1(new_n21909_), .B0(new_n1834_), .Y(new_n21929_));
  OR4X1    g21737(.A(new_n21393_), .B(new_n21200_), .C(new_n21188_), .D(new_n21182_), .Y(new_n21930_));
  OR2X1    g21738(.A(new_n21200_), .B(new_n21182_), .Y(new_n21931_));
  OAI21X1  g21739(.A0(new_n21931_), .A1(new_n21393_), .B0(new_n21188_), .Y(new_n21932_));
  AND2X1   g21740(.A(new_n21932_), .B(new_n21930_), .Y(new_n21933_));
  OAI21X1  g21741(.A0(new_n21918_), .A1(new_n21905_), .B0(new_n21926_), .Y(new_n21934_));
  AOI21X1  g21742(.A0(new_n21934_), .A1(\asqrt[47] ), .B0(\asqrt[48] ), .Y(new_n21935_));
  AOI21X1  g21743(.A0(new_n21935_), .A1(new_n21928_), .B0(new_n21933_), .Y(new_n21936_));
  OAI21X1  g21744(.A0(new_n21936_), .A1(new_n21929_), .B0(\asqrt[49] ), .Y(new_n21937_));
  AND2X1   g21745(.A(new_n21244_), .B(new_n21243_), .Y(new_n21938_));
  NOR3X1   g21746(.A(new_n21938_), .B(new_n21206_), .C(new_n21242_), .Y(new_n21939_));
  NOR3X1   g21747(.A(new_n21393_), .B(new_n21938_), .C(new_n21242_), .Y(new_n21940_));
  NOR2X1   g21748(.A(new_n21940_), .B(new_n21205_), .Y(new_n21941_));
  AOI21X1  g21749(.A0(new_n21939_), .A1(\asqrt[6] ), .B0(new_n21941_), .Y(new_n21942_));
  NOR3X1   g21750(.A(new_n21936_), .B(new_n21929_), .C(\asqrt[49] ), .Y(new_n21943_));
  OAI21X1  g21751(.A0(new_n21943_), .A1(new_n21942_), .B0(new_n21937_), .Y(new_n21944_));
  AND2X1   g21752(.A(new_n21944_), .B(\asqrt[50] ), .Y(new_n21945_));
  OR2X1    g21753(.A(new_n21943_), .B(new_n21942_), .Y(new_n21946_));
  AND2X1   g21754(.A(new_n21217_), .B(new_n21209_), .Y(new_n21947_));
  NOR3X1   g21755(.A(new_n21947_), .B(new_n21247_), .C(new_n21210_), .Y(new_n21948_));
  NOR3X1   g21756(.A(new_n21393_), .B(new_n21947_), .C(new_n21210_), .Y(new_n21949_));
  NOR2X1   g21757(.A(new_n21949_), .B(new_n21215_), .Y(new_n21950_));
  AOI21X1  g21758(.A0(new_n21948_), .A1(\asqrt[6] ), .B0(new_n21950_), .Y(new_n21951_));
  AND2X1   g21759(.A(new_n21937_), .B(new_n1469_), .Y(new_n21952_));
  AOI21X1  g21760(.A0(new_n21952_), .A1(new_n21946_), .B0(new_n21951_), .Y(new_n21953_));
  OAI21X1  g21761(.A0(new_n21953_), .A1(new_n21945_), .B0(\asqrt[51] ), .Y(new_n21954_));
  OR4X1    g21762(.A(new_n21393_), .B(new_n21225_), .C(new_n21251_), .D(new_n21250_), .Y(new_n21955_));
  OR2X1    g21763(.A(new_n21225_), .B(new_n21250_), .Y(new_n21956_));
  OAI21X1  g21764(.A0(new_n21956_), .A1(new_n21393_), .B0(new_n21251_), .Y(new_n21957_));
  AND2X1   g21765(.A(new_n21957_), .B(new_n21955_), .Y(new_n21958_));
  INVX1    g21766(.A(new_n21958_), .Y(new_n21959_));
  AND2X1   g21767(.A(new_n21934_), .B(\asqrt[47] ), .Y(new_n21960_));
  OR2X1    g21768(.A(new_n21918_), .B(new_n21905_), .Y(new_n21961_));
  AND2X1   g21769(.A(new_n21926_), .B(new_n2040_), .Y(new_n21962_));
  AOI21X1  g21770(.A0(new_n21962_), .A1(new_n21961_), .B0(new_n21924_), .Y(new_n21963_));
  OAI21X1  g21771(.A0(new_n21963_), .A1(new_n21960_), .B0(\asqrt[48] ), .Y(new_n21964_));
  INVX1    g21772(.A(new_n21933_), .Y(new_n21965_));
  OAI21X1  g21773(.A0(new_n21908_), .A1(new_n2040_), .B0(new_n1834_), .Y(new_n21966_));
  OAI21X1  g21774(.A0(new_n21966_), .A1(new_n21963_), .B0(new_n21965_), .Y(new_n21967_));
  AOI21X1  g21775(.A0(new_n21967_), .A1(new_n21964_), .B0(new_n1632_), .Y(new_n21968_));
  INVX1    g21776(.A(new_n21942_), .Y(new_n21969_));
  NAND3X1  g21777(.A(new_n21967_), .B(new_n21964_), .C(new_n1632_), .Y(new_n21970_));
  AOI21X1  g21778(.A0(new_n21970_), .A1(new_n21969_), .B0(new_n21968_), .Y(new_n21971_));
  OAI21X1  g21779(.A0(new_n21971_), .A1(new_n1469_), .B0(new_n1277_), .Y(new_n21972_));
  OAI21X1  g21780(.A0(new_n21972_), .A1(new_n21953_), .B0(new_n21959_), .Y(new_n21973_));
  AOI21X1  g21781(.A0(new_n21973_), .A1(new_n21954_), .B0(new_n1111_), .Y(new_n21974_));
  AOI21X1  g21782(.A0(new_n21233_), .A1(new_n21228_), .B0(new_n21268_), .Y(new_n21975_));
  AND2X1   g21783(.A(new_n21975_), .B(new_n21266_), .Y(new_n21976_));
  AOI22X1  g21784(.A0(new_n21233_), .A1(new_n21228_), .B0(new_n21226_), .B1(\asqrt[51] ), .Y(new_n21977_));
  AOI21X1  g21785(.A0(new_n21977_), .A1(\asqrt[6] ), .B0(new_n21232_), .Y(new_n21978_));
  AOI21X1  g21786(.A0(new_n21976_), .A1(\asqrt[6] ), .B0(new_n21978_), .Y(new_n21979_));
  INVX1    g21787(.A(new_n21979_), .Y(new_n21980_));
  NAND3X1  g21788(.A(new_n21973_), .B(new_n21954_), .C(new_n1111_), .Y(new_n21981_));
  AOI21X1  g21789(.A0(new_n21981_), .A1(new_n21980_), .B0(new_n21974_), .Y(new_n21982_));
  OR2X1    g21790(.A(new_n21982_), .B(new_n968_), .Y(new_n21983_));
  OR2X1    g21791(.A(new_n21971_), .B(new_n1469_), .Y(new_n21984_));
  NOR2X1   g21792(.A(new_n21943_), .B(new_n21942_), .Y(new_n21985_));
  INVX1    g21793(.A(new_n21951_), .Y(new_n21986_));
  NAND2X1  g21794(.A(new_n21937_), .B(new_n1469_), .Y(new_n21987_));
  OAI21X1  g21795(.A0(new_n21987_), .A1(new_n21985_), .B0(new_n21986_), .Y(new_n21988_));
  AOI21X1  g21796(.A0(new_n21988_), .A1(new_n21984_), .B0(new_n1277_), .Y(new_n21989_));
  AOI21X1  g21797(.A0(new_n21944_), .A1(\asqrt[50] ), .B0(\asqrt[51] ), .Y(new_n21990_));
  AOI21X1  g21798(.A0(new_n21990_), .A1(new_n21988_), .B0(new_n21958_), .Y(new_n21991_));
  NOR3X1   g21799(.A(new_n21991_), .B(new_n21989_), .C(\asqrt[52] ), .Y(new_n21992_));
  NOR2X1   g21800(.A(new_n21992_), .B(new_n21979_), .Y(new_n21993_));
  AND2X1   g21801(.A(new_n21272_), .B(new_n21270_), .Y(new_n21994_));
  NOR3X1   g21802(.A(new_n21994_), .B(new_n21241_), .C(new_n21271_), .Y(new_n21995_));
  NOR3X1   g21803(.A(new_n21393_), .B(new_n21994_), .C(new_n21271_), .Y(new_n21996_));
  NOR2X1   g21804(.A(new_n21996_), .B(new_n21240_), .Y(new_n21997_));
  AOI21X1  g21805(.A0(new_n21995_), .A1(\asqrt[6] ), .B0(new_n21997_), .Y(new_n21998_));
  INVX1    g21806(.A(new_n21998_), .Y(new_n21999_));
  OAI21X1  g21807(.A0(new_n21991_), .A1(new_n21989_), .B0(\asqrt[52] ), .Y(new_n22000_));
  NAND2X1  g21808(.A(new_n22000_), .B(new_n968_), .Y(new_n22001_));
  OAI21X1  g21809(.A0(new_n22001_), .A1(new_n21993_), .B0(new_n21999_), .Y(new_n22002_));
  AOI21X1  g21810(.A0(new_n22002_), .A1(new_n21983_), .B0(new_n902_), .Y(new_n22003_));
  OR4X1    g21811(.A(new_n21393_), .B(new_n21274_), .C(new_n21262_), .D(new_n21256_), .Y(new_n22004_));
  OR2X1    g21812(.A(new_n21274_), .B(new_n21256_), .Y(new_n22005_));
  OAI21X1  g21813(.A0(new_n22005_), .A1(new_n21393_), .B0(new_n21262_), .Y(new_n22006_));
  AND2X1   g21814(.A(new_n22006_), .B(new_n22004_), .Y(new_n22007_));
  OAI21X1  g21815(.A0(new_n21992_), .A1(new_n21979_), .B0(new_n22000_), .Y(new_n22008_));
  AOI21X1  g21816(.A0(new_n22008_), .A1(\asqrt[53] ), .B0(\asqrt[54] ), .Y(new_n22009_));
  AOI21X1  g21817(.A0(new_n22009_), .A1(new_n22002_), .B0(new_n22007_), .Y(new_n22010_));
  OAI21X1  g21818(.A0(new_n22010_), .A1(new_n22003_), .B0(\asqrt[55] ), .Y(new_n22011_));
  AND2X1   g21819(.A(new_n21312_), .B(new_n21311_), .Y(new_n22012_));
  NOR3X1   g21820(.A(new_n22012_), .B(new_n21280_), .C(new_n21310_), .Y(new_n22013_));
  NOR3X1   g21821(.A(new_n21393_), .B(new_n22012_), .C(new_n21310_), .Y(new_n22014_));
  NOR2X1   g21822(.A(new_n22014_), .B(new_n21279_), .Y(new_n22015_));
  AOI21X1  g21823(.A0(new_n22013_), .A1(\asqrt[6] ), .B0(new_n22015_), .Y(new_n22016_));
  NOR3X1   g21824(.A(new_n22010_), .B(new_n22003_), .C(\asqrt[55] ), .Y(new_n22017_));
  OAI21X1  g21825(.A0(new_n22017_), .A1(new_n22016_), .B0(new_n22011_), .Y(new_n22018_));
  AND2X1   g21826(.A(new_n22018_), .B(\asqrt[56] ), .Y(new_n22019_));
  OR2X1    g21827(.A(new_n22017_), .B(new_n22016_), .Y(new_n22020_));
  AND2X1   g21828(.A(new_n21291_), .B(new_n21283_), .Y(new_n22021_));
  NOR3X1   g21829(.A(new_n22021_), .B(new_n21315_), .C(new_n21284_), .Y(new_n22022_));
  NOR3X1   g21830(.A(new_n21393_), .B(new_n22021_), .C(new_n21284_), .Y(new_n22023_));
  NOR2X1   g21831(.A(new_n22023_), .B(new_n21289_), .Y(new_n22024_));
  AOI21X1  g21832(.A0(new_n22022_), .A1(\asqrt[6] ), .B0(new_n22024_), .Y(new_n22025_));
  AND2X1   g21833(.A(new_n22011_), .B(new_n582_), .Y(new_n22026_));
  AOI21X1  g21834(.A0(new_n22026_), .A1(new_n22020_), .B0(new_n22025_), .Y(new_n22027_));
  OAI21X1  g21835(.A0(new_n22027_), .A1(new_n22019_), .B0(\asqrt[57] ), .Y(new_n22028_));
  OR4X1    g21836(.A(new_n21393_), .B(new_n21299_), .C(new_n21319_), .D(new_n21318_), .Y(new_n22029_));
  OR2X1    g21837(.A(new_n21299_), .B(new_n21318_), .Y(new_n22030_));
  OAI21X1  g21838(.A0(new_n22030_), .A1(new_n21393_), .B0(new_n21319_), .Y(new_n22031_));
  AND2X1   g21839(.A(new_n22031_), .B(new_n22029_), .Y(new_n22032_));
  INVX1    g21840(.A(new_n22032_), .Y(new_n22033_));
  AND2X1   g21841(.A(new_n22008_), .B(\asqrt[53] ), .Y(new_n22034_));
  OR2X1    g21842(.A(new_n21992_), .B(new_n21979_), .Y(new_n22035_));
  AND2X1   g21843(.A(new_n22000_), .B(new_n968_), .Y(new_n22036_));
  AOI21X1  g21844(.A0(new_n22036_), .A1(new_n22035_), .B0(new_n21998_), .Y(new_n22037_));
  OAI21X1  g21845(.A0(new_n22037_), .A1(new_n22034_), .B0(\asqrt[54] ), .Y(new_n22038_));
  INVX1    g21846(.A(new_n22007_), .Y(new_n22039_));
  OAI21X1  g21847(.A0(new_n21982_), .A1(new_n968_), .B0(new_n902_), .Y(new_n22040_));
  OAI21X1  g21848(.A0(new_n22040_), .A1(new_n22037_), .B0(new_n22039_), .Y(new_n22041_));
  AOI21X1  g21849(.A0(new_n22041_), .A1(new_n22038_), .B0(new_n697_), .Y(new_n22042_));
  INVX1    g21850(.A(new_n22016_), .Y(new_n22043_));
  NAND3X1  g21851(.A(new_n22041_), .B(new_n22038_), .C(new_n697_), .Y(new_n22044_));
  AOI21X1  g21852(.A0(new_n22044_), .A1(new_n22043_), .B0(new_n22042_), .Y(new_n22045_));
  OAI21X1  g21853(.A0(new_n22045_), .A1(new_n582_), .B0(new_n481_), .Y(new_n22046_));
  OAI21X1  g21854(.A0(new_n22046_), .A1(new_n22027_), .B0(new_n22033_), .Y(new_n22047_));
  AOI21X1  g21855(.A0(new_n22047_), .A1(new_n22028_), .B0(new_n399_), .Y(new_n22048_));
  AOI21X1  g21856(.A0(new_n21307_), .A1(new_n21302_), .B0(new_n21342_), .Y(new_n22049_));
  AND2X1   g21857(.A(new_n22049_), .B(new_n21340_), .Y(new_n22050_));
  AOI22X1  g21858(.A0(new_n21307_), .A1(new_n21302_), .B0(new_n21300_), .B1(\asqrt[57] ), .Y(new_n22051_));
  AOI21X1  g21859(.A0(new_n22051_), .A1(\asqrt[6] ), .B0(new_n21306_), .Y(new_n22052_));
  AOI21X1  g21860(.A0(new_n22050_), .A1(\asqrt[6] ), .B0(new_n22052_), .Y(new_n22053_));
  INVX1    g21861(.A(new_n22053_), .Y(new_n22054_));
  NAND3X1  g21862(.A(new_n22047_), .B(new_n22028_), .C(new_n399_), .Y(new_n22055_));
  AOI21X1  g21863(.A0(new_n22055_), .A1(new_n22054_), .B0(new_n22048_), .Y(new_n22056_));
  OR2X1    g21864(.A(new_n22056_), .B(new_n328_), .Y(new_n22057_));
  OR2X1    g21865(.A(new_n22045_), .B(new_n582_), .Y(new_n22058_));
  NOR2X1   g21866(.A(new_n22017_), .B(new_n22016_), .Y(new_n22059_));
  INVX1    g21867(.A(new_n22025_), .Y(new_n22060_));
  NAND2X1  g21868(.A(new_n22011_), .B(new_n582_), .Y(new_n22061_));
  OAI21X1  g21869(.A0(new_n22061_), .A1(new_n22059_), .B0(new_n22060_), .Y(new_n22062_));
  AOI21X1  g21870(.A0(new_n22062_), .A1(new_n22058_), .B0(new_n481_), .Y(new_n22063_));
  AOI21X1  g21871(.A0(new_n22018_), .A1(\asqrt[56] ), .B0(\asqrt[57] ), .Y(new_n22064_));
  AOI21X1  g21872(.A0(new_n22064_), .A1(new_n22062_), .B0(new_n22032_), .Y(new_n22065_));
  NOR3X1   g21873(.A(new_n22065_), .B(new_n22063_), .C(\asqrt[58] ), .Y(new_n22066_));
  NOR2X1   g21874(.A(new_n22066_), .B(new_n22053_), .Y(new_n22067_));
  OAI21X1  g21875(.A0(new_n22065_), .A1(new_n22063_), .B0(\asqrt[58] ), .Y(new_n22068_));
  NAND2X1  g21876(.A(new_n22068_), .B(new_n328_), .Y(new_n22069_));
  AND2X1   g21877(.A(new_n21346_), .B(new_n21344_), .Y(new_n22070_));
  NOR3X1   g21878(.A(new_n21328_), .B(new_n22070_), .C(new_n21345_), .Y(new_n22071_));
  NOR3X1   g21879(.A(new_n21393_), .B(new_n22070_), .C(new_n21345_), .Y(new_n22072_));
  NOR2X1   g21880(.A(new_n22072_), .B(new_n21327_), .Y(new_n22073_));
  AOI21X1  g21881(.A0(new_n22071_), .A1(\asqrt[6] ), .B0(new_n22073_), .Y(new_n22074_));
  INVX1    g21882(.A(new_n22074_), .Y(new_n22075_));
  OAI21X1  g21883(.A0(new_n22069_), .A1(new_n22067_), .B0(new_n22075_), .Y(new_n22076_));
  AOI21X1  g21884(.A0(new_n22076_), .A1(new_n22057_), .B0(new_n292_), .Y(new_n22077_));
  OR4X1    g21885(.A(new_n21393_), .B(new_n21348_), .C(new_n21336_), .D(new_n21330_), .Y(new_n22078_));
  OR2X1    g21886(.A(new_n21348_), .B(new_n21330_), .Y(new_n22079_));
  OAI21X1  g21887(.A0(new_n22079_), .A1(new_n21393_), .B0(new_n21336_), .Y(new_n22080_));
  AND2X1   g21888(.A(new_n22080_), .B(new_n22078_), .Y(new_n22081_));
  OAI21X1  g21889(.A0(new_n22066_), .A1(new_n22053_), .B0(new_n22068_), .Y(new_n22082_));
  AOI21X1  g21890(.A0(new_n22082_), .A1(\asqrt[59] ), .B0(\asqrt[60] ), .Y(new_n22083_));
  AOI21X1  g21891(.A0(new_n22083_), .A1(new_n22076_), .B0(new_n22081_), .Y(new_n22084_));
  OAI21X1  g21892(.A0(new_n22084_), .A1(new_n22077_), .B0(\asqrt[61] ), .Y(new_n22085_));
  AND2X1   g21893(.A(new_n21397_), .B(new_n21396_), .Y(new_n22086_));
  NOR3X1   g21894(.A(new_n22086_), .B(new_n21354_), .C(new_n21395_), .Y(new_n22087_));
  NOR3X1   g21895(.A(new_n21393_), .B(new_n22086_), .C(new_n21395_), .Y(new_n22088_));
  NOR2X1   g21896(.A(new_n22088_), .B(new_n21353_), .Y(new_n22089_));
  AOI21X1  g21897(.A0(new_n22087_), .A1(\asqrt[6] ), .B0(new_n22089_), .Y(new_n22090_));
  NOR3X1   g21898(.A(new_n22084_), .B(new_n22077_), .C(\asqrt[61] ), .Y(new_n22091_));
  OAI21X1  g21899(.A0(new_n22091_), .A1(new_n22090_), .B0(new_n22085_), .Y(new_n22092_));
  AND2X1   g21900(.A(new_n22092_), .B(\asqrt[62] ), .Y(new_n22093_));
  OR2X1    g21901(.A(new_n22091_), .B(new_n22090_), .Y(new_n22094_));
  AND2X1   g21902(.A(new_n21365_), .B(new_n21357_), .Y(new_n22095_));
  NOR3X1   g21903(.A(new_n22095_), .B(new_n21400_), .C(new_n21358_), .Y(new_n22096_));
  NOR3X1   g21904(.A(new_n21393_), .B(new_n22095_), .C(new_n21358_), .Y(new_n22097_));
  NOR2X1   g21905(.A(new_n22097_), .B(new_n21363_), .Y(new_n22098_));
  AOI21X1  g21906(.A0(new_n22096_), .A1(\asqrt[6] ), .B0(new_n22098_), .Y(new_n22099_));
  AND2X1   g21907(.A(new_n22085_), .B(new_n199_), .Y(new_n22100_));
  AOI21X1  g21908(.A0(new_n22100_), .A1(new_n22094_), .B0(new_n22099_), .Y(new_n22101_));
  NOR3X1   g21909(.A(new_n21373_), .B(new_n21404_), .C(new_n21403_), .Y(new_n22102_));
  NOR3X1   g21910(.A(new_n21393_), .B(new_n21373_), .C(new_n21403_), .Y(new_n22103_));
  NOR2X1   g21911(.A(new_n22103_), .B(new_n21372_), .Y(new_n22104_));
  AOI21X1  g21912(.A0(new_n22102_), .A1(\asqrt[6] ), .B0(new_n22104_), .Y(new_n22105_));
  INVX1    g21913(.A(new_n22105_), .Y(new_n22106_));
  NOR3X1   g21914(.A(new_n21393_), .B(new_n21378_), .C(new_n21406_), .Y(new_n22107_));
  AOI21X1  g21915(.A0(new_n21410_), .A1(new_n21409_), .B0(new_n22107_), .Y(new_n22108_));
  AND2X1   g21916(.A(new_n22108_), .B(new_n22106_), .Y(new_n22109_));
  OAI21X1  g21917(.A0(new_n22101_), .A1(new_n22093_), .B0(new_n22109_), .Y(new_n22110_));
  AND2X1   g21918(.A(new_n22082_), .B(\asqrt[59] ), .Y(new_n22111_));
  OR2X1    g21919(.A(new_n22066_), .B(new_n22053_), .Y(new_n22112_));
  AND2X1   g21920(.A(new_n22068_), .B(new_n328_), .Y(new_n22113_));
  AOI21X1  g21921(.A0(new_n22113_), .A1(new_n22112_), .B0(new_n22074_), .Y(new_n22114_));
  OAI21X1  g21922(.A0(new_n22114_), .A1(new_n22111_), .B0(\asqrt[60] ), .Y(new_n22115_));
  INVX1    g21923(.A(new_n22081_), .Y(new_n22116_));
  OAI21X1  g21924(.A0(new_n22056_), .A1(new_n328_), .B0(new_n292_), .Y(new_n22117_));
  OAI21X1  g21925(.A0(new_n22117_), .A1(new_n22114_), .B0(new_n22116_), .Y(new_n22118_));
  AOI21X1  g21926(.A0(new_n22118_), .A1(new_n22115_), .B0(new_n217_), .Y(new_n22119_));
  INVX1    g21927(.A(new_n22090_), .Y(new_n22120_));
  NAND3X1  g21928(.A(new_n22118_), .B(new_n22115_), .C(new_n217_), .Y(new_n22121_));
  AOI21X1  g21929(.A0(new_n22121_), .A1(new_n22120_), .B0(new_n22119_), .Y(new_n22122_));
  OAI21X1  g21930(.A0(new_n22122_), .A1(new_n199_), .B0(new_n22105_), .Y(new_n22123_));
  AOI21X1  g21931(.A0(new_n21412_), .A1(new_n21408_), .B0(new_n21378_), .Y(new_n22124_));
  AOI21X1  g21932(.A0(new_n21379_), .A1(new_n21374_), .B0(new_n193_), .Y(new_n22125_));
  OAI21X1  g21933(.A0(new_n22124_), .A1(new_n21374_), .B0(new_n22125_), .Y(new_n22126_));
  OAI21X1  g21934(.A0(new_n22123_), .A1(new_n22101_), .B0(new_n22126_), .Y(new_n22127_));
  AOI21X1  g21935(.A0(new_n22110_), .A1(new_n193_), .B0(new_n22127_), .Y(new_n22128_));
  OR2X1    g21936(.A(new_n22122_), .B(new_n199_), .Y(new_n22129_));
  NOR2X1   g21937(.A(new_n22091_), .B(new_n22090_), .Y(new_n22130_));
  INVX1    g21938(.A(new_n22099_), .Y(new_n22131_));
  NAND2X1  g21939(.A(new_n22085_), .B(new_n199_), .Y(new_n22132_));
  OAI21X1  g21940(.A0(new_n22132_), .A1(new_n22130_), .B0(new_n22131_), .Y(new_n22133_));
  INVX1    g21941(.A(new_n22109_), .Y(new_n22134_));
  AOI21X1  g21942(.A0(new_n22133_), .A1(new_n22129_), .B0(new_n22134_), .Y(new_n22135_));
  AOI21X1  g21943(.A0(new_n22092_), .A1(\asqrt[62] ), .B0(new_n22106_), .Y(new_n22136_));
  INVX1    g21944(.A(new_n22126_), .Y(new_n22137_));
  AOI21X1  g21945(.A0(new_n22136_), .A1(new_n22133_), .B0(new_n22137_), .Y(new_n22138_));
  OAI21X1  g21946(.A0(new_n22135_), .A1(\asqrt[63] ), .B0(new_n22138_), .Y(\asqrt[5] ));
  NOR2X1   g21947(.A(\a[9] ), .B(\a[8] ), .Y(new_n22140_));
  MX2X1    g21948(.A(new_n22140_), .B(\asqrt[5] ), .S0(\a[10] ), .Y(new_n22141_));
  AND2X1   g21949(.A(new_n22141_), .B(\asqrt[6] ), .Y(new_n22142_));
  OR2X1    g21950(.A(new_n21385_), .B(new_n21384_), .Y(new_n22143_));
  INVX1    g21951(.A(new_n22140_), .Y(new_n22144_));
  OAI22X1  g21952(.A0(new_n22144_), .A1(\a[10] ), .B0(new_n21389_), .B1(new_n20662_), .Y(new_n22145_));
  NOR2X1   g21953(.A(new_n22145_), .B(new_n21387_), .Y(new_n22146_));
  NAND3X1  g21954(.A(new_n22146_), .B(new_n22143_), .C(new_n21408_), .Y(new_n22147_));
  AOI21X1  g21955(.A0(\asqrt[5] ), .A1(\a[10] ), .B0(new_n22147_), .Y(new_n22148_));
  INVX1    g21956(.A(\a[10] ), .Y(new_n22149_));
  INVX1    g21957(.A(\a[11] ), .Y(new_n22150_));
  AOI21X1  g21958(.A0(\asqrt[5] ), .A1(new_n22149_), .B0(new_n22150_), .Y(new_n22151_));
  NOR2X1   g21959(.A(\a[11] ), .B(\a[10] ), .Y(new_n22152_));
  AND2X1   g21960(.A(\asqrt[5] ), .B(new_n22152_), .Y(new_n22153_));
  NOR3X1   g21961(.A(new_n22153_), .B(new_n22151_), .C(new_n22148_), .Y(new_n22154_));
  OAI21X1  g21962(.A0(new_n22154_), .A1(new_n22142_), .B0(\asqrt[7] ), .Y(new_n22155_));
  MX2X1    g21963(.A(new_n22144_), .B(new_n22128_), .S0(\a[10] ), .Y(new_n22156_));
  OAI21X1  g21964(.A0(new_n22156_), .A1(new_n21393_), .B0(new_n20676_), .Y(new_n22157_));
  AND2X1   g21965(.A(new_n22126_), .B(\asqrt[6] ), .Y(new_n22158_));
  OAI21X1  g21966(.A0(new_n22123_), .A1(new_n22101_), .B0(new_n22158_), .Y(new_n22159_));
  AOI21X1  g21967(.A0(new_n22110_), .A1(new_n193_), .B0(new_n22159_), .Y(new_n22160_));
  AOI21X1  g21968(.A0(\asqrt[5] ), .A1(new_n22152_), .B0(new_n22160_), .Y(new_n22161_));
  OR2X1    g21969(.A(new_n22160_), .B(\a[12] ), .Y(new_n22162_));
  OAI22X1  g21970(.A0(new_n22162_), .A1(new_n22153_), .B0(new_n22161_), .B1(new_n21394_), .Y(new_n22163_));
  OAI21X1  g21971(.A0(new_n22157_), .A1(new_n22154_), .B0(new_n22163_), .Y(new_n22164_));
  AOI21X1  g21972(.A0(new_n22164_), .A1(new_n22155_), .B0(new_n19976_), .Y(new_n22165_));
  AND2X1   g21973(.A(new_n21427_), .B(new_n21415_), .Y(new_n22166_));
  NAND3X1  g21974(.A(new_n22166_), .B(\asqrt[5] ), .C(new_n21424_), .Y(new_n22167_));
  INVX1    g21975(.A(new_n22166_), .Y(new_n22168_));
  OAI21X1  g21976(.A0(new_n22168_), .A1(new_n22128_), .B0(new_n21431_), .Y(new_n22169_));
  AND2X1   g21977(.A(new_n22169_), .B(new_n22167_), .Y(new_n22170_));
  INVX1    g21978(.A(new_n22170_), .Y(new_n22171_));
  NAND3X1  g21979(.A(new_n22164_), .B(new_n22155_), .C(new_n19976_), .Y(new_n22172_));
  AOI21X1  g21980(.A0(new_n22172_), .A1(new_n22171_), .B0(new_n22165_), .Y(new_n22173_));
  OR2X1    g21981(.A(new_n22173_), .B(new_n19273_), .Y(new_n22174_));
  AND2X1   g21982(.A(new_n22172_), .B(new_n22171_), .Y(new_n22175_));
  AOI21X1  g21983(.A0(new_n21433_), .A1(new_n21432_), .B0(new_n21468_), .Y(new_n22176_));
  NAND3X1  g21984(.A(new_n22176_), .B(\asqrt[5] ), .C(new_n21465_), .Y(new_n22177_));
  OAI22X1  g21985(.A0(new_n21467_), .A1(new_n21466_), .B0(new_n21450_), .B1(new_n19976_), .Y(new_n22178_));
  OAI21X1  g21986(.A0(new_n22178_), .A1(new_n22128_), .B0(new_n21468_), .Y(new_n22179_));
  AND2X1   g21987(.A(new_n22179_), .B(new_n22177_), .Y(new_n22180_));
  INVX1    g21988(.A(new_n22180_), .Y(new_n22181_));
  OR2X1    g21989(.A(new_n22165_), .B(\asqrt[9] ), .Y(new_n22182_));
  OAI21X1  g21990(.A0(new_n22182_), .A1(new_n22175_), .B0(new_n22181_), .Y(new_n22183_));
  AOI21X1  g21991(.A0(new_n22183_), .A1(new_n22174_), .B0(new_n18591_), .Y(new_n22184_));
  OR2X1    g21992(.A(new_n21451_), .B(new_n21441_), .Y(new_n22185_));
  NAND4X1  g21993(.A(\asqrt[5] ), .B(new_n22185_), .C(new_n21471_), .D(new_n21442_), .Y(new_n22186_));
  NAND2X1  g21994(.A(new_n22185_), .B(new_n21442_), .Y(new_n22187_));
  OAI21X1  g21995(.A0(new_n22187_), .A1(new_n22128_), .B0(new_n21448_), .Y(new_n22188_));
  AND2X1   g21996(.A(new_n22188_), .B(new_n22186_), .Y(new_n22189_));
  OR2X1    g21997(.A(new_n22156_), .B(new_n21393_), .Y(new_n22190_));
  INVX1    g21998(.A(new_n22147_), .Y(new_n22191_));
  OAI21X1  g21999(.A0(new_n22128_), .A1(new_n22149_), .B0(new_n22191_), .Y(new_n22192_));
  OAI21X1  g22000(.A0(new_n22128_), .A1(\a[10] ), .B0(\a[11] ), .Y(new_n22193_));
  INVX1    g22001(.A(new_n22152_), .Y(new_n22194_));
  OR2X1    g22002(.A(new_n22128_), .B(new_n22194_), .Y(new_n22195_));
  NAND3X1  g22003(.A(new_n22195_), .B(new_n22193_), .C(new_n22192_), .Y(new_n22196_));
  AOI21X1  g22004(.A0(new_n22196_), .A1(new_n22190_), .B0(new_n20676_), .Y(new_n22197_));
  AOI21X1  g22005(.A0(new_n22141_), .A1(\asqrt[6] ), .B0(\asqrt[7] ), .Y(new_n22198_));
  AND2X1   g22006(.A(new_n22110_), .B(new_n193_), .Y(new_n22199_));
  OAI22X1  g22007(.A0(new_n22159_), .A1(new_n22199_), .B0(new_n22128_), .B1(new_n22194_), .Y(new_n22200_));
  NOR2X1   g22008(.A(new_n22160_), .B(\a[12] ), .Y(new_n22201_));
  AOI22X1  g22009(.A0(new_n22201_), .A1(new_n22195_), .B0(new_n22200_), .B1(\a[12] ), .Y(new_n22202_));
  AOI21X1  g22010(.A0(new_n22198_), .A1(new_n22196_), .B0(new_n22202_), .Y(new_n22203_));
  OAI21X1  g22011(.A0(new_n22203_), .A1(new_n22197_), .B0(\asqrt[8] ), .Y(new_n22204_));
  NOR3X1   g22012(.A(new_n22203_), .B(new_n22197_), .C(\asqrt[8] ), .Y(new_n22205_));
  OAI21X1  g22013(.A0(new_n22205_), .A1(new_n22170_), .B0(new_n22204_), .Y(new_n22206_));
  AOI21X1  g22014(.A0(new_n22206_), .A1(\asqrt[9] ), .B0(\asqrt[10] ), .Y(new_n22207_));
  AOI21X1  g22015(.A0(new_n22207_), .A1(new_n22183_), .B0(new_n22189_), .Y(new_n22208_));
  OAI21X1  g22016(.A0(new_n22208_), .A1(new_n22184_), .B0(\asqrt[11] ), .Y(new_n22209_));
  OR4X1    g22017(.A(new_n22128_), .B(new_n21474_), .C(new_n21461_), .D(new_n21453_), .Y(new_n22210_));
  NAND2X1  g22018(.A(new_n21462_), .B(new_n21483_), .Y(new_n22211_));
  OAI21X1  g22019(.A0(new_n22211_), .A1(new_n22128_), .B0(new_n21461_), .Y(new_n22212_));
  AND2X1   g22020(.A(new_n22212_), .B(new_n22210_), .Y(new_n22213_));
  NOR3X1   g22021(.A(new_n22208_), .B(new_n22184_), .C(\asqrt[11] ), .Y(new_n22214_));
  OAI21X1  g22022(.A0(new_n22214_), .A1(new_n22213_), .B0(new_n22209_), .Y(new_n22215_));
  AND2X1   g22023(.A(new_n22215_), .B(\asqrt[12] ), .Y(new_n22216_));
  INVX1    g22024(.A(new_n22213_), .Y(new_n22217_));
  AND2X1   g22025(.A(new_n22206_), .B(\asqrt[9] ), .Y(new_n22218_));
  NAND2X1  g22026(.A(new_n22172_), .B(new_n22171_), .Y(new_n22219_));
  NOR2X1   g22027(.A(new_n22165_), .B(\asqrt[9] ), .Y(new_n22220_));
  AOI21X1  g22028(.A0(new_n22220_), .A1(new_n22219_), .B0(new_n22180_), .Y(new_n22221_));
  OAI21X1  g22029(.A0(new_n22221_), .A1(new_n22218_), .B0(\asqrt[10] ), .Y(new_n22222_));
  INVX1    g22030(.A(new_n22189_), .Y(new_n22223_));
  OAI21X1  g22031(.A0(new_n22173_), .A1(new_n19273_), .B0(new_n18591_), .Y(new_n22224_));
  OAI21X1  g22032(.A0(new_n22224_), .A1(new_n22221_), .B0(new_n22223_), .Y(new_n22225_));
  NAND3X1  g22033(.A(new_n22225_), .B(new_n22222_), .C(new_n17927_), .Y(new_n22226_));
  NAND2X1  g22034(.A(new_n22226_), .B(new_n22217_), .Y(new_n22227_));
  AND2X1   g22035(.A(new_n21506_), .B(new_n21505_), .Y(new_n22228_));
  NOR4X1   g22036(.A(new_n22128_), .B(new_n22228_), .C(new_n21482_), .D(new_n21504_), .Y(new_n22229_));
  AOI22X1  g22037(.A0(new_n21506_), .A1(new_n21505_), .B0(new_n21491_), .B1(\asqrt[11] ), .Y(new_n22230_));
  AOI21X1  g22038(.A0(new_n22230_), .A1(\asqrt[5] ), .B0(new_n21481_), .Y(new_n22231_));
  NOR2X1   g22039(.A(new_n22231_), .B(new_n22229_), .Y(new_n22232_));
  AOI21X1  g22040(.A0(new_n22225_), .A1(new_n22222_), .B0(new_n17927_), .Y(new_n22233_));
  NOR2X1   g22041(.A(new_n22233_), .B(\asqrt[12] ), .Y(new_n22234_));
  AOI21X1  g22042(.A0(new_n22234_), .A1(new_n22227_), .B0(new_n22232_), .Y(new_n22235_));
  OAI21X1  g22043(.A0(new_n22235_), .A1(new_n22216_), .B0(\asqrt[13] ), .Y(new_n22236_));
  AND2X1   g22044(.A(new_n21492_), .B(new_n21485_), .Y(new_n22237_));
  OR4X1    g22045(.A(new_n22128_), .B(new_n22237_), .C(new_n21489_), .D(new_n21486_), .Y(new_n22238_));
  OR2X1    g22046(.A(new_n22237_), .B(new_n21486_), .Y(new_n22239_));
  OAI21X1  g22047(.A0(new_n22239_), .A1(new_n22128_), .B0(new_n21489_), .Y(new_n22240_));
  AND2X1   g22048(.A(new_n22240_), .B(new_n22238_), .Y(new_n22241_));
  INVX1    g22049(.A(new_n22241_), .Y(new_n22242_));
  AOI21X1  g22050(.A0(new_n22226_), .A1(new_n22217_), .B0(new_n22233_), .Y(new_n22243_));
  OAI21X1  g22051(.A0(new_n22243_), .A1(new_n17262_), .B0(new_n16617_), .Y(new_n22244_));
  OAI21X1  g22052(.A0(new_n22244_), .A1(new_n22235_), .B0(new_n22242_), .Y(new_n22245_));
  AOI21X1  g22053(.A0(new_n22245_), .A1(new_n22236_), .B0(new_n15990_), .Y(new_n22246_));
  OR4X1    g22054(.A(new_n22128_), .B(new_n21500_), .C(new_n21503_), .D(new_n21526_), .Y(new_n22247_));
  NAND2X1  g22055(.A(new_n21511_), .B(new_n21494_), .Y(new_n22248_));
  OAI21X1  g22056(.A0(new_n22248_), .A1(new_n22128_), .B0(new_n21503_), .Y(new_n22249_));
  AND2X1   g22057(.A(new_n22249_), .B(new_n22247_), .Y(new_n22250_));
  INVX1    g22058(.A(new_n22250_), .Y(new_n22251_));
  NAND3X1  g22059(.A(new_n22245_), .B(new_n22236_), .C(new_n15990_), .Y(new_n22252_));
  AOI21X1  g22060(.A0(new_n22252_), .A1(new_n22251_), .B0(new_n22246_), .Y(new_n22253_));
  OR2X1    g22061(.A(new_n22253_), .B(new_n15362_), .Y(new_n22254_));
  AND2X1   g22062(.A(new_n22252_), .B(new_n22251_), .Y(new_n22255_));
  OAI21X1  g22063(.A0(new_n21550_), .A1(new_n21548_), .B0(new_n21517_), .Y(new_n22256_));
  NOR3X1   g22064(.A(new_n22256_), .B(new_n22128_), .C(new_n21502_), .Y(new_n22257_));
  AOI22X1  g22065(.A0(new_n21518_), .A1(new_n21512_), .B0(new_n21501_), .B1(\asqrt[14] ), .Y(new_n22258_));
  AOI21X1  g22066(.A0(new_n22258_), .A1(\asqrt[5] ), .B0(new_n21517_), .Y(new_n22259_));
  NOR2X1   g22067(.A(new_n22259_), .B(new_n22257_), .Y(new_n22260_));
  INVX1    g22068(.A(new_n22260_), .Y(new_n22261_));
  OR2X1    g22069(.A(new_n22246_), .B(\asqrt[15] ), .Y(new_n22262_));
  OAI21X1  g22070(.A0(new_n22262_), .A1(new_n22255_), .B0(new_n22261_), .Y(new_n22263_));
  AOI21X1  g22071(.A0(new_n22263_), .A1(new_n22254_), .B0(new_n14754_), .Y(new_n22264_));
  AND2X1   g22072(.A(new_n21553_), .B(new_n21551_), .Y(new_n22265_));
  OR4X1    g22073(.A(new_n22128_), .B(new_n22265_), .C(new_n21525_), .D(new_n21552_), .Y(new_n22266_));
  OR2X1    g22074(.A(new_n22265_), .B(new_n21552_), .Y(new_n22267_));
  OAI21X1  g22075(.A0(new_n22267_), .A1(new_n22128_), .B0(new_n21525_), .Y(new_n22268_));
  AND2X1   g22076(.A(new_n22268_), .B(new_n22266_), .Y(new_n22269_));
  OR2X1    g22077(.A(new_n22243_), .B(new_n17262_), .Y(new_n22270_));
  AND2X1   g22078(.A(new_n22226_), .B(new_n22217_), .Y(new_n22271_));
  INVX1    g22079(.A(new_n22232_), .Y(new_n22272_));
  OR2X1    g22080(.A(new_n22233_), .B(\asqrt[12] ), .Y(new_n22273_));
  OAI21X1  g22081(.A0(new_n22273_), .A1(new_n22271_), .B0(new_n22272_), .Y(new_n22274_));
  AOI21X1  g22082(.A0(new_n22274_), .A1(new_n22270_), .B0(new_n16617_), .Y(new_n22275_));
  AOI21X1  g22083(.A0(new_n22215_), .A1(\asqrt[12] ), .B0(\asqrt[13] ), .Y(new_n22276_));
  AOI21X1  g22084(.A0(new_n22276_), .A1(new_n22274_), .B0(new_n22241_), .Y(new_n22277_));
  OAI21X1  g22085(.A0(new_n22277_), .A1(new_n22275_), .B0(\asqrt[14] ), .Y(new_n22278_));
  NOR3X1   g22086(.A(new_n22277_), .B(new_n22275_), .C(\asqrt[14] ), .Y(new_n22279_));
  OAI21X1  g22087(.A0(new_n22279_), .A1(new_n22250_), .B0(new_n22278_), .Y(new_n22280_));
  AOI21X1  g22088(.A0(new_n22280_), .A1(\asqrt[15] ), .B0(\asqrt[16] ), .Y(new_n22281_));
  AOI21X1  g22089(.A0(new_n22281_), .A1(new_n22263_), .B0(new_n22269_), .Y(new_n22282_));
  OAI21X1  g22090(.A0(new_n22282_), .A1(new_n22264_), .B0(\asqrt[17] ), .Y(new_n22283_));
  OR4X1    g22091(.A(new_n22128_), .B(new_n21563_), .C(new_n21536_), .D(new_n21530_), .Y(new_n22284_));
  NAND2X1  g22092(.A(new_n21537_), .B(new_n21555_), .Y(new_n22285_));
  OAI21X1  g22093(.A0(new_n22285_), .A1(new_n22128_), .B0(new_n21536_), .Y(new_n22286_));
  AND2X1   g22094(.A(new_n22286_), .B(new_n22284_), .Y(new_n22287_));
  NOR3X1   g22095(.A(new_n22282_), .B(new_n22264_), .C(\asqrt[17] ), .Y(new_n22288_));
  OAI21X1  g22096(.A0(new_n22288_), .A1(new_n22287_), .B0(new_n22283_), .Y(new_n22289_));
  AND2X1   g22097(.A(new_n22289_), .B(\asqrt[18] ), .Y(new_n22290_));
  INVX1    g22098(.A(new_n22287_), .Y(new_n22291_));
  AND2X1   g22099(.A(new_n22280_), .B(\asqrt[15] ), .Y(new_n22292_));
  NAND2X1  g22100(.A(new_n22252_), .B(new_n22251_), .Y(new_n22293_));
  NOR2X1   g22101(.A(new_n22246_), .B(\asqrt[15] ), .Y(new_n22294_));
  AOI21X1  g22102(.A0(new_n22294_), .A1(new_n22293_), .B0(new_n22260_), .Y(new_n22295_));
  OAI21X1  g22103(.A0(new_n22295_), .A1(new_n22292_), .B0(\asqrt[16] ), .Y(new_n22296_));
  INVX1    g22104(.A(new_n22269_), .Y(new_n22297_));
  OAI21X1  g22105(.A0(new_n22253_), .A1(new_n15362_), .B0(new_n14754_), .Y(new_n22298_));
  OAI21X1  g22106(.A0(new_n22298_), .A1(new_n22295_), .B0(new_n22297_), .Y(new_n22299_));
  NAND3X1  g22107(.A(new_n22299_), .B(new_n22296_), .C(new_n14165_), .Y(new_n22300_));
  NAND2X1  g22108(.A(new_n22300_), .B(new_n22291_), .Y(new_n22301_));
  AND2X1   g22109(.A(new_n21579_), .B(new_n21578_), .Y(new_n22302_));
  NOR4X1   g22110(.A(new_n22128_), .B(new_n22302_), .C(new_n21546_), .D(new_n21577_), .Y(new_n22303_));
  AOI22X1  g22111(.A0(new_n21579_), .A1(new_n21578_), .B0(new_n21564_), .B1(\asqrt[17] ), .Y(new_n22304_));
  AOI21X1  g22112(.A0(new_n22304_), .A1(\asqrt[5] ), .B0(new_n21545_), .Y(new_n22305_));
  NOR2X1   g22113(.A(new_n22305_), .B(new_n22303_), .Y(new_n22306_));
  AOI21X1  g22114(.A0(new_n22299_), .A1(new_n22296_), .B0(new_n14165_), .Y(new_n22307_));
  NOR2X1   g22115(.A(new_n22307_), .B(\asqrt[18] ), .Y(new_n22308_));
  AOI21X1  g22116(.A0(new_n22308_), .A1(new_n22301_), .B0(new_n22306_), .Y(new_n22309_));
  OAI21X1  g22117(.A0(new_n22309_), .A1(new_n22290_), .B0(\asqrt[19] ), .Y(new_n22310_));
  AND2X1   g22118(.A(new_n21565_), .B(new_n21557_), .Y(new_n22311_));
  OR4X1    g22119(.A(new_n22128_), .B(new_n22311_), .C(new_n21582_), .D(new_n21558_), .Y(new_n22312_));
  OR2X1    g22120(.A(new_n22311_), .B(new_n21558_), .Y(new_n22313_));
  OAI21X1  g22121(.A0(new_n22313_), .A1(new_n22128_), .B0(new_n21582_), .Y(new_n22314_));
  AND2X1   g22122(.A(new_n22314_), .B(new_n22312_), .Y(new_n22315_));
  INVX1    g22123(.A(new_n22315_), .Y(new_n22316_));
  AOI21X1  g22124(.A0(new_n22300_), .A1(new_n22291_), .B0(new_n22307_), .Y(new_n22317_));
  OAI21X1  g22125(.A0(new_n22317_), .A1(new_n13571_), .B0(new_n13000_), .Y(new_n22318_));
  OAI21X1  g22126(.A0(new_n22318_), .A1(new_n22309_), .B0(new_n22316_), .Y(new_n22319_));
  AOI21X1  g22127(.A0(new_n22319_), .A1(new_n22310_), .B0(new_n12447_), .Y(new_n22320_));
  OR4X1    g22128(.A(new_n22128_), .B(new_n21573_), .C(new_n21576_), .D(new_n21600_), .Y(new_n22321_));
  NAND2X1  g22129(.A(new_n21585_), .B(new_n21567_), .Y(new_n22322_));
  OAI21X1  g22130(.A0(new_n22322_), .A1(new_n22128_), .B0(new_n21576_), .Y(new_n22323_));
  AND2X1   g22131(.A(new_n22323_), .B(new_n22321_), .Y(new_n22324_));
  INVX1    g22132(.A(new_n22324_), .Y(new_n22325_));
  NAND3X1  g22133(.A(new_n22319_), .B(new_n22310_), .C(new_n12447_), .Y(new_n22326_));
  AOI21X1  g22134(.A0(new_n22326_), .A1(new_n22325_), .B0(new_n22320_), .Y(new_n22327_));
  OR2X1    g22135(.A(new_n22327_), .B(new_n11896_), .Y(new_n22328_));
  AND2X1   g22136(.A(new_n22326_), .B(new_n22325_), .Y(new_n22329_));
  OAI21X1  g22137(.A0(new_n21624_), .A1(new_n21622_), .B0(new_n21591_), .Y(new_n22330_));
  NOR3X1   g22138(.A(new_n22330_), .B(new_n22128_), .C(new_n21575_), .Y(new_n22331_));
  AOI22X1  g22139(.A0(new_n21592_), .A1(new_n21586_), .B0(new_n21574_), .B1(\asqrt[20] ), .Y(new_n22332_));
  AOI21X1  g22140(.A0(new_n22332_), .A1(\asqrt[5] ), .B0(new_n21591_), .Y(new_n22333_));
  NOR2X1   g22141(.A(new_n22333_), .B(new_n22331_), .Y(new_n22334_));
  INVX1    g22142(.A(new_n22334_), .Y(new_n22335_));
  OR2X1    g22143(.A(new_n22320_), .B(\asqrt[21] ), .Y(new_n22336_));
  OAI21X1  g22144(.A0(new_n22336_), .A1(new_n22329_), .B0(new_n22335_), .Y(new_n22337_));
  AOI21X1  g22145(.A0(new_n22337_), .A1(new_n22328_), .B0(new_n11362_), .Y(new_n22338_));
  AND2X1   g22146(.A(new_n21627_), .B(new_n21625_), .Y(new_n22339_));
  OR4X1    g22147(.A(new_n22128_), .B(new_n22339_), .C(new_n21599_), .D(new_n21626_), .Y(new_n22340_));
  OR2X1    g22148(.A(new_n22339_), .B(new_n21626_), .Y(new_n22341_));
  OAI21X1  g22149(.A0(new_n22341_), .A1(new_n22128_), .B0(new_n21599_), .Y(new_n22342_));
  AND2X1   g22150(.A(new_n22342_), .B(new_n22340_), .Y(new_n22343_));
  OR2X1    g22151(.A(new_n22317_), .B(new_n13571_), .Y(new_n22344_));
  AND2X1   g22152(.A(new_n22300_), .B(new_n22291_), .Y(new_n22345_));
  INVX1    g22153(.A(new_n22306_), .Y(new_n22346_));
  OR2X1    g22154(.A(new_n22307_), .B(\asqrt[18] ), .Y(new_n22347_));
  OAI21X1  g22155(.A0(new_n22347_), .A1(new_n22345_), .B0(new_n22346_), .Y(new_n22348_));
  AOI21X1  g22156(.A0(new_n22348_), .A1(new_n22344_), .B0(new_n13000_), .Y(new_n22349_));
  AOI21X1  g22157(.A0(new_n22289_), .A1(\asqrt[18] ), .B0(\asqrt[19] ), .Y(new_n22350_));
  AOI21X1  g22158(.A0(new_n22350_), .A1(new_n22348_), .B0(new_n22315_), .Y(new_n22351_));
  OAI21X1  g22159(.A0(new_n22351_), .A1(new_n22349_), .B0(\asqrt[20] ), .Y(new_n22352_));
  NOR3X1   g22160(.A(new_n22351_), .B(new_n22349_), .C(\asqrt[20] ), .Y(new_n22353_));
  OAI21X1  g22161(.A0(new_n22353_), .A1(new_n22324_), .B0(new_n22352_), .Y(new_n22354_));
  AOI21X1  g22162(.A0(new_n22354_), .A1(\asqrt[21] ), .B0(\asqrt[22] ), .Y(new_n22355_));
  AOI21X1  g22163(.A0(new_n22355_), .A1(new_n22337_), .B0(new_n22343_), .Y(new_n22356_));
  OAI21X1  g22164(.A0(new_n22356_), .A1(new_n22338_), .B0(\asqrt[23] ), .Y(new_n22357_));
  OR4X1    g22165(.A(new_n22128_), .B(new_n21637_), .C(new_n21610_), .D(new_n21604_), .Y(new_n22358_));
  NAND2X1  g22166(.A(new_n21611_), .B(new_n21629_), .Y(new_n22359_));
  OAI21X1  g22167(.A0(new_n22359_), .A1(new_n22128_), .B0(new_n21610_), .Y(new_n22360_));
  AND2X1   g22168(.A(new_n22360_), .B(new_n22358_), .Y(new_n22361_));
  NOR3X1   g22169(.A(new_n22356_), .B(new_n22338_), .C(\asqrt[23] ), .Y(new_n22362_));
  OAI21X1  g22170(.A0(new_n22362_), .A1(new_n22361_), .B0(new_n22357_), .Y(new_n22363_));
  AND2X1   g22171(.A(new_n22363_), .B(\asqrt[24] ), .Y(new_n22364_));
  INVX1    g22172(.A(new_n22361_), .Y(new_n22365_));
  AND2X1   g22173(.A(new_n22354_), .B(\asqrt[21] ), .Y(new_n22366_));
  NAND2X1  g22174(.A(new_n22326_), .B(new_n22325_), .Y(new_n22367_));
  NOR2X1   g22175(.A(new_n22320_), .B(\asqrt[21] ), .Y(new_n22368_));
  AOI21X1  g22176(.A0(new_n22368_), .A1(new_n22367_), .B0(new_n22334_), .Y(new_n22369_));
  OAI21X1  g22177(.A0(new_n22369_), .A1(new_n22366_), .B0(\asqrt[22] ), .Y(new_n22370_));
  INVX1    g22178(.A(new_n22343_), .Y(new_n22371_));
  OAI21X1  g22179(.A0(new_n22327_), .A1(new_n11896_), .B0(new_n11362_), .Y(new_n22372_));
  OAI21X1  g22180(.A0(new_n22372_), .A1(new_n22369_), .B0(new_n22371_), .Y(new_n22373_));
  NAND3X1  g22181(.A(new_n22373_), .B(new_n22370_), .C(new_n10849_), .Y(new_n22374_));
  NAND2X1  g22182(.A(new_n22374_), .B(new_n22365_), .Y(new_n22375_));
  AND2X1   g22183(.A(new_n21653_), .B(new_n21652_), .Y(new_n22376_));
  NOR4X1   g22184(.A(new_n22128_), .B(new_n22376_), .C(new_n21620_), .D(new_n21651_), .Y(new_n22377_));
  AOI22X1  g22185(.A0(new_n21653_), .A1(new_n21652_), .B0(new_n21638_), .B1(\asqrt[23] ), .Y(new_n22378_));
  AOI21X1  g22186(.A0(new_n22378_), .A1(\asqrt[5] ), .B0(new_n21619_), .Y(new_n22379_));
  NOR2X1   g22187(.A(new_n22379_), .B(new_n22377_), .Y(new_n22380_));
  AOI21X1  g22188(.A0(new_n22373_), .A1(new_n22370_), .B0(new_n10849_), .Y(new_n22381_));
  NOR2X1   g22189(.A(new_n22381_), .B(\asqrt[24] ), .Y(new_n22382_));
  AOI21X1  g22190(.A0(new_n22382_), .A1(new_n22375_), .B0(new_n22380_), .Y(new_n22383_));
  OAI21X1  g22191(.A0(new_n22383_), .A1(new_n22364_), .B0(\asqrt[25] ), .Y(new_n22384_));
  AND2X1   g22192(.A(new_n21639_), .B(new_n21631_), .Y(new_n22385_));
  OR4X1    g22193(.A(new_n22128_), .B(new_n22385_), .C(new_n21656_), .D(new_n21632_), .Y(new_n22386_));
  OR2X1    g22194(.A(new_n22385_), .B(new_n21632_), .Y(new_n22387_));
  OAI21X1  g22195(.A0(new_n22387_), .A1(new_n22128_), .B0(new_n21656_), .Y(new_n22388_));
  AND2X1   g22196(.A(new_n22388_), .B(new_n22386_), .Y(new_n22389_));
  INVX1    g22197(.A(new_n22389_), .Y(new_n22390_));
  AOI21X1  g22198(.A0(new_n22374_), .A1(new_n22365_), .B0(new_n22381_), .Y(new_n22391_));
  OAI21X1  g22199(.A0(new_n22391_), .A1(new_n10332_), .B0(new_n9833_), .Y(new_n22392_));
  OAI21X1  g22200(.A0(new_n22392_), .A1(new_n22383_), .B0(new_n22390_), .Y(new_n22393_));
  AOI21X1  g22201(.A0(new_n22393_), .A1(new_n22384_), .B0(new_n9353_), .Y(new_n22394_));
  NAND3X1  g22202(.A(new_n21659_), .B(new_n21646_), .C(new_n21641_), .Y(new_n22395_));
  NOR3X1   g22203(.A(new_n22128_), .B(new_n21647_), .C(new_n21674_), .Y(new_n22396_));
  OAI22X1  g22204(.A0(new_n22396_), .A1(new_n21646_), .B0(new_n22395_), .B1(new_n22128_), .Y(new_n22397_));
  NAND3X1  g22205(.A(new_n22393_), .B(new_n22384_), .C(new_n9353_), .Y(new_n22398_));
  AOI21X1  g22206(.A0(new_n22398_), .A1(new_n22397_), .B0(new_n22394_), .Y(new_n22399_));
  OR2X1    g22207(.A(new_n22399_), .B(new_n8874_), .Y(new_n22400_));
  AND2X1   g22208(.A(new_n22398_), .B(new_n22397_), .Y(new_n22401_));
  OAI21X1  g22209(.A0(new_n21698_), .A1(new_n21696_), .B0(new_n21665_), .Y(new_n22402_));
  NOR3X1   g22210(.A(new_n22402_), .B(new_n22128_), .C(new_n21649_), .Y(new_n22403_));
  AOI22X1  g22211(.A0(new_n21666_), .A1(new_n21660_), .B0(new_n21648_), .B1(\asqrt[26] ), .Y(new_n22404_));
  AOI21X1  g22212(.A0(new_n22404_), .A1(\asqrt[5] ), .B0(new_n21665_), .Y(new_n22405_));
  NOR2X1   g22213(.A(new_n22405_), .B(new_n22403_), .Y(new_n22406_));
  INVX1    g22214(.A(new_n22406_), .Y(new_n22407_));
  OR2X1    g22215(.A(new_n22394_), .B(\asqrt[27] ), .Y(new_n22408_));
  OAI21X1  g22216(.A0(new_n22408_), .A1(new_n22401_), .B0(new_n22407_), .Y(new_n22409_));
  AOI21X1  g22217(.A0(new_n22409_), .A1(new_n22400_), .B0(new_n8412_), .Y(new_n22410_));
  AND2X1   g22218(.A(new_n21701_), .B(new_n21699_), .Y(new_n22411_));
  OR4X1    g22219(.A(new_n22128_), .B(new_n22411_), .C(new_n21673_), .D(new_n21700_), .Y(new_n22412_));
  OR2X1    g22220(.A(new_n22411_), .B(new_n21700_), .Y(new_n22413_));
  OAI21X1  g22221(.A0(new_n22413_), .A1(new_n22128_), .B0(new_n21673_), .Y(new_n22414_));
  AND2X1   g22222(.A(new_n22414_), .B(new_n22412_), .Y(new_n22415_));
  OR2X1    g22223(.A(new_n22391_), .B(new_n10332_), .Y(new_n22416_));
  AND2X1   g22224(.A(new_n22374_), .B(new_n22365_), .Y(new_n22417_));
  INVX1    g22225(.A(new_n22380_), .Y(new_n22418_));
  OR2X1    g22226(.A(new_n22381_), .B(\asqrt[24] ), .Y(new_n22419_));
  OAI21X1  g22227(.A0(new_n22419_), .A1(new_n22417_), .B0(new_n22418_), .Y(new_n22420_));
  AOI21X1  g22228(.A0(new_n22420_), .A1(new_n22416_), .B0(new_n9833_), .Y(new_n22421_));
  AOI21X1  g22229(.A0(new_n22363_), .A1(\asqrt[24] ), .B0(\asqrt[25] ), .Y(new_n22422_));
  AOI21X1  g22230(.A0(new_n22422_), .A1(new_n22420_), .B0(new_n22389_), .Y(new_n22423_));
  OAI21X1  g22231(.A0(new_n22423_), .A1(new_n22421_), .B0(\asqrt[26] ), .Y(new_n22424_));
  INVX1    g22232(.A(new_n22397_), .Y(new_n22425_));
  NOR3X1   g22233(.A(new_n22423_), .B(new_n22421_), .C(\asqrt[26] ), .Y(new_n22426_));
  OAI21X1  g22234(.A0(new_n22426_), .A1(new_n22425_), .B0(new_n22424_), .Y(new_n22427_));
  AOI21X1  g22235(.A0(new_n22427_), .A1(\asqrt[27] ), .B0(\asqrt[28] ), .Y(new_n22428_));
  AOI21X1  g22236(.A0(new_n22428_), .A1(new_n22409_), .B0(new_n22415_), .Y(new_n22429_));
  OAI21X1  g22237(.A0(new_n22429_), .A1(new_n22410_), .B0(\asqrt[29] ), .Y(new_n22430_));
  OR4X1    g22238(.A(new_n22128_), .B(new_n21711_), .C(new_n21684_), .D(new_n21678_), .Y(new_n22431_));
  NAND2X1  g22239(.A(new_n21685_), .B(new_n21703_), .Y(new_n22432_));
  OAI21X1  g22240(.A0(new_n22432_), .A1(new_n22128_), .B0(new_n21684_), .Y(new_n22433_));
  AND2X1   g22241(.A(new_n22433_), .B(new_n22431_), .Y(new_n22434_));
  NOR3X1   g22242(.A(new_n22429_), .B(new_n22410_), .C(\asqrt[29] ), .Y(new_n22435_));
  OAI21X1  g22243(.A0(new_n22435_), .A1(new_n22434_), .B0(new_n22430_), .Y(new_n22436_));
  AND2X1   g22244(.A(new_n22436_), .B(\asqrt[30] ), .Y(new_n22437_));
  INVX1    g22245(.A(new_n22434_), .Y(new_n22438_));
  AND2X1   g22246(.A(new_n22427_), .B(\asqrt[27] ), .Y(new_n22439_));
  NAND2X1  g22247(.A(new_n22398_), .B(new_n22397_), .Y(new_n22440_));
  NOR2X1   g22248(.A(new_n22394_), .B(\asqrt[27] ), .Y(new_n22441_));
  AOI21X1  g22249(.A0(new_n22441_), .A1(new_n22440_), .B0(new_n22406_), .Y(new_n22442_));
  OAI21X1  g22250(.A0(new_n22442_), .A1(new_n22439_), .B0(\asqrt[28] ), .Y(new_n22443_));
  INVX1    g22251(.A(new_n22415_), .Y(new_n22444_));
  OAI21X1  g22252(.A0(new_n22399_), .A1(new_n8874_), .B0(new_n8412_), .Y(new_n22445_));
  OAI21X1  g22253(.A0(new_n22445_), .A1(new_n22442_), .B0(new_n22444_), .Y(new_n22446_));
  NAND3X1  g22254(.A(new_n22446_), .B(new_n22443_), .C(new_n7970_), .Y(new_n22447_));
  NAND2X1  g22255(.A(new_n22447_), .B(new_n22438_), .Y(new_n22448_));
  AND2X1   g22256(.A(new_n21740_), .B(new_n21739_), .Y(new_n22449_));
  NOR4X1   g22257(.A(new_n22128_), .B(new_n22449_), .C(new_n21694_), .D(new_n21738_), .Y(new_n22450_));
  AOI22X1  g22258(.A0(new_n21740_), .A1(new_n21739_), .B0(new_n21712_), .B1(\asqrt[29] ), .Y(new_n22451_));
  AOI21X1  g22259(.A0(new_n22451_), .A1(\asqrt[5] ), .B0(new_n21693_), .Y(new_n22452_));
  NOR2X1   g22260(.A(new_n22452_), .B(new_n22450_), .Y(new_n22453_));
  AOI21X1  g22261(.A0(new_n22446_), .A1(new_n22443_), .B0(new_n7970_), .Y(new_n22454_));
  NOR2X1   g22262(.A(new_n22454_), .B(\asqrt[30] ), .Y(new_n22455_));
  AOI21X1  g22263(.A0(new_n22455_), .A1(new_n22448_), .B0(new_n22453_), .Y(new_n22456_));
  OAI21X1  g22264(.A0(new_n22456_), .A1(new_n22437_), .B0(\asqrt[31] ), .Y(new_n22457_));
  AND2X1   g22265(.A(new_n21713_), .B(new_n21705_), .Y(new_n22458_));
  OR4X1    g22266(.A(new_n22128_), .B(new_n22458_), .C(new_n21743_), .D(new_n21706_), .Y(new_n22459_));
  OR2X1    g22267(.A(new_n22458_), .B(new_n21706_), .Y(new_n22460_));
  OAI21X1  g22268(.A0(new_n22460_), .A1(new_n22128_), .B0(new_n21743_), .Y(new_n22461_));
  AND2X1   g22269(.A(new_n22461_), .B(new_n22459_), .Y(new_n22462_));
  INVX1    g22270(.A(new_n22462_), .Y(new_n22463_));
  AOI21X1  g22271(.A0(new_n22447_), .A1(new_n22438_), .B0(new_n22454_), .Y(new_n22464_));
  OAI21X1  g22272(.A0(new_n22464_), .A1(new_n7527_), .B0(new_n7103_), .Y(new_n22465_));
  OAI21X1  g22273(.A0(new_n22465_), .A1(new_n22456_), .B0(new_n22463_), .Y(new_n22466_));
  AOI21X1  g22274(.A0(new_n22466_), .A1(new_n22457_), .B0(new_n6699_), .Y(new_n22467_));
  OR4X1    g22275(.A(new_n22128_), .B(new_n21721_), .C(new_n21747_), .D(new_n21746_), .Y(new_n22468_));
  OR2X1    g22276(.A(new_n21721_), .B(new_n21746_), .Y(new_n22469_));
  OAI21X1  g22277(.A0(new_n22469_), .A1(new_n22128_), .B0(new_n21747_), .Y(new_n22470_));
  AND2X1   g22278(.A(new_n22470_), .B(new_n22468_), .Y(new_n22471_));
  INVX1    g22279(.A(new_n22471_), .Y(new_n22472_));
  NAND3X1  g22280(.A(new_n22466_), .B(new_n22457_), .C(new_n6699_), .Y(new_n22473_));
  AOI21X1  g22281(.A0(new_n22473_), .A1(new_n22472_), .B0(new_n22467_), .Y(new_n22474_));
  OR2X1    g22282(.A(new_n22474_), .B(new_n6294_), .Y(new_n22475_));
  AND2X1   g22283(.A(new_n22473_), .B(new_n22472_), .Y(new_n22476_));
  OAI21X1  g22284(.A0(new_n21765_), .A1(new_n21763_), .B0(new_n21729_), .Y(new_n22477_));
  NOR3X1   g22285(.A(new_n22477_), .B(new_n22128_), .C(new_n21723_), .Y(new_n22478_));
  AOI22X1  g22286(.A0(new_n21730_), .A1(new_n21724_), .B0(new_n21722_), .B1(\asqrt[32] ), .Y(new_n22479_));
  AOI21X1  g22287(.A0(new_n22479_), .A1(\asqrt[5] ), .B0(new_n21729_), .Y(new_n22480_));
  NOR2X1   g22288(.A(new_n22480_), .B(new_n22478_), .Y(new_n22481_));
  INVX1    g22289(.A(new_n22481_), .Y(new_n22482_));
  OR2X1    g22290(.A(new_n22467_), .B(\asqrt[33] ), .Y(new_n22483_));
  OAI21X1  g22291(.A0(new_n22483_), .A1(new_n22476_), .B0(new_n22482_), .Y(new_n22484_));
  AOI21X1  g22292(.A0(new_n22484_), .A1(new_n22475_), .B0(new_n5941_), .Y(new_n22485_));
  AND2X1   g22293(.A(new_n21768_), .B(new_n21766_), .Y(new_n22486_));
  OR4X1    g22294(.A(new_n22128_), .B(new_n22486_), .C(new_n21737_), .D(new_n21767_), .Y(new_n22487_));
  OR2X1    g22295(.A(new_n22486_), .B(new_n21767_), .Y(new_n22488_));
  OAI21X1  g22296(.A0(new_n22488_), .A1(new_n22128_), .B0(new_n21737_), .Y(new_n22489_));
  AND2X1   g22297(.A(new_n22489_), .B(new_n22487_), .Y(new_n22490_));
  OR2X1    g22298(.A(new_n22464_), .B(new_n7527_), .Y(new_n22491_));
  AND2X1   g22299(.A(new_n22447_), .B(new_n22438_), .Y(new_n22492_));
  INVX1    g22300(.A(new_n22453_), .Y(new_n22493_));
  OR2X1    g22301(.A(new_n22454_), .B(\asqrt[30] ), .Y(new_n22494_));
  OAI21X1  g22302(.A0(new_n22494_), .A1(new_n22492_), .B0(new_n22493_), .Y(new_n22495_));
  AOI21X1  g22303(.A0(new_n22495_), .A1(new_n22491_), .B0(new_n7103_), .Y(new_n22496_));
  AOI21X1  g22304(.A0(new_n22436_), .A1(\asqrt[30] ), .B0(\asqrt[31] ), .Y(new_n22497_));
  AOI21X1  g22305(.A0(new_n22497_), .A1(new_n22495_), .B0(new_n22462_), .Y(new_n22498_));
  OAI21X1  g22306(.A0(new_n22498_), .A1(new_n22496_), .B0(\asqrt[32] ), .Y(new_n22499_));
  NOR3X1   g22307(.A(new_n22498_), .B(new_n22496_), .C(\asqrt[32] ), .Y(new_n22500_));
  OAI21X1  g22308(.A0(new_n22500_), .A1(new_n22471_), .B0(new_n22499_), .Y(new_n22501_));
  AOI21X1  g22309(.A0(new_n22501_), .A1(\asqrt[33] ), .B0(\asqrt[34] ), .Y(new_n22502_));
  AOI21X1  g22310(.A0(new_n22502_), .A1(new_n22484_), .B0(new_n22490_), .Y(new_n22503_));
  OAI21X1  g22311(.A0(new_n22503_), .A1(new_n22485_), .B0(\asqrt[35] ), .Y(new_n22504_));
  OR4X1    g22312(.A(new_n22128_), .B(new_n21770_), .C(new_n21758_), .D(new_n21752_), .Y(new_n22505_));
  OR2X1    g22313(.A(new_n21770_), .B(new_n21752_), .Y(new_n22506_));
  OAI21X1  g22314(.A0(new_n22506_), .A1(new_n22128_), .B0(new_n21758_), .Y(new_n22507_));
  AND2X1   g22315(.A(new_n22507_), .B(new_n22505_), .Y(new_n22508_));
  NOR3X1   g22316(.A(new_n22503_), .B(new_n22485_), .C(\asqrt[35] ), .Y(new_n22509_));
  OAI21X1  g22317(.A0(new_n22509_), .A1(new_n22508_), .B0(new_n22504_), .Y(new_n22510_));
  AND2X1   g22318(.A(new_n22510_), .B(\asqrt[36] ), .Y(new_n22511_));
  OR2X1    g22319(.A(new_n22509_), .B(new_n22508_), .Y(new_n22512_));
  AND2X1   g22320(.A(new_n21814_), .B(new_n21813_), .Y(new_n22513_));
  NOR4X1   g22321(.A(new_n22128_), .B(new_n22513_), .C(new_n21777_), .D(new_n21812_), .Y(new_n22514_));
  AOI22X1  g22322(.A0(new_n21814_), .A1(new_n21813_), .B0(new_n21786_), .B1(\asqrt[35] ), .Y(new_n22515_));
  AOI21X1  g22323(.A0(new_n22515_), .A1(\asqrt[5] ), .B0(new_n21776_), .Y(new_n22516_));
  NOR2X1   g22324(.A(new_n22516_), .B(new_n22514_), .Y(new_n22517_));
  AND2X1   g22325(.A(new_n22504_), .B(new_n5176_), .Y(new_n22518_));
  AOI21X1  g22326(.A0(new_n22518_), .A1(new_n22512_), .B0(new_n22517_), .Y(new_n22519_));
  OAI21X1  g22327(.A0(new_n22519_), .A1(new_n22511_), .B0(\asqrt[37] ), .Y(new_n22520_));
  AND2X1   g22328(.A(new_n21787_), .B(new_n21780_), .Y(new_n22521_));
  OR4X1    g22329(.A(new_n22128_), .B(new_n22521_), .C(new_n21817_), .D(new_n21781_), .Y(new_n22522_));
  OR2X1    g22330(.A(new_n22521_), .B(new_n21781_), .Y(new_n22523_));
  OAI21X1  g22331(.A0(new_n22523_), .A1(new_n22128_), .B0(new_n21817_), .Y(new_n22524_));
  AND2X1   g22332(.A(new_n22524_), .B(new_n22522_), .Y(new_n22525_));
  INVX1    g22333(.A(new_n22525_), .Y(new_n22526_));
  AND2X1   g22334(.A(new_n22501_), .B(\asqrt[33] ), .Y(new_n22527_));
  NAND2X1  g22335(.A(new_n22473_), .B(new_n22472_), .Y(new_n22528_));
  NOR2X1   g22336(.A(new_n22467_), .B(\asqrt[33] ), .Y(new_n22529_));
  AOI21X1  g22337(.A0(new_n22529_), .A1(new_n22528_), .B0(new_n22481_), .Y(new_n22530_));
  OAI21X1  g22338(.A0(new_n22530_), .A1(new_n22527_), .B0(\asqrt[34] ), .Y(new_n22531_));
  INVX1    g22339(.A(new_n22490_), .Y(new_n22532_));
  OAI21X1  g22340(.A0(new_n22474_), .A1(new_n6294_), .B0(new_n5941_), .Y(new_n22533_));
  OAI21X1  g22341(.A0(new_n22533_), .A1(new_n22530_), .B0(new_n22532_), .Y(new_n22534_));
  AOI21X1  g22342(.A0(new_n22534_), .A1(new_n22531_), .B0(new_n5541_), .Y(new_n22535_));
  INVX1    g22343(.A(new_n22508_), .Y(new_n22536_));
  NAND3X1  g22344(.A(new_n22534_), .B(new_n22531_), .C(new_n5541_), .Y(new_n22537_));
  AOI21X1  g22345(.A0(new_n22537_), .A1(new_n22536_), .B0(new_n22535_), .Y(new_n22538_));
  OAI21X1  g22346(.A0(new_n22538_), .A1(new_n5176_), .B0(new_n4826_), .Y(new_n22539_));
  OAI21X1  g22347(.A0(new_n22539_), .A1(new_n22519_), .B0(new_n22526_), .Y(new_n22540_));
  AOI21X1  g22348(.A0(new_n22540_), .A1(new_n22520_), .B0(new_n4493_), .Y(new_n22541_));
  OR4X1    g22349(.A(new_n22128_), .B(new_n21795_), .C(new_n21821_), .D(new_n21820_), .Y(new_n22542_));
  OR2X1    g22350(.A(new_n21795_), .B(new_n21820_), .Y(new_n22543_));
  OAI21X1  g22351(.A0(new_n22543_), .A1(new_n22128_), .B0(new_n21821_), .Y(new_n22544_));
  AND2X1   g22352(.A(new_n22544_), .B(new_n22542_), .Y(new_n22545_));
  INVX1    g22353(.A(new_n22545_), .Y(new_n22546_));
  NAND3X1  g22354(.A(new_n22540_), .B(new_n22520_), .C(new_n4493_), .Y(new_n22547_));
  AOI21X1  g22355(.A0(new_n22547_), .A1(new_n22546_), .B0(new_n22541_), .Y(new_n22548_));
  OR2X1    g22356(.A(new_n22548_), .B(new_n4165_), .Y(new_n22549_));
  OR2X1    g22357(.A(new_n22538_), .B(new_n5176_), .Y(new_n22550_));
  NOR2X1   g22358(.A(new_n22509_), .B(new_n22508_), .Y(new_n22551_));
  INVX1    g22359(.A(new_n22517_), .Y(new_n22552_));
  NAND2X1  g22360(.A(new_n22504_), .B(new_n5176_), .Y(new_n22553_));
  OAI21X1  g22361(.A0(new_n22553_), .A1(new_n22551_), .B0(new_n22552_), .Y(new_n22554_));
  AOI21X1  g22362(.A0(new_n22554_), .A1(new_n22550_), .B0(new_n4826_), .Y(new_n22555_));
  AOI21X1  g22363(.A0(new_n22510_), .A1(\asqrt[36] ), .B0(\asqrt[37] ), .Y(new_n22556_));
  AOI21X1  g22364(.A0(new_n22556_), .A1(new_n22554_), .B0(new_n22525_), .Y(new_n22557_));
  NOR3X1   g22365(.A(new_n22557_), .B(new_n22555_), .C(\asqrt[38] ), .Y(new_n22558_));
  NOR2X1   g22366(.A(new_n22558_), .B(new_n22545_), .Y(new_n22559_));
  OAI21X1  g22367(.A0(new_n21839_), .A1(new_n21837_), .B0(new_n21803_), .Y(new_n22560_));
  NOR3X1   g22368(.A(new_n22560_), .B(new_n22128_), .C(new_n21797_), .Y(new_n22561_));
  AOI22X1  g22369(.A0(new_n21804_), .A1(new_n21798_), .B0(new_n21796_), .B1(\asqrt[38] ), .Y(new_n22562_));
  AOI21X1  g22370(.A0(new_n22562_), .A1(\asqrt[5] ), .B0(new_n21803_), .Y(new_n22563_));
  NOR2X1   g22371(.A(new_n22563_), .B(new_n22561_), .Y(new_n22564_));
  INVX1    g22372(.A(new_n22564_), .Y(new_n22565_));
  OAI21X1  g22373(.A0(new_n22557_), .A1(new_n22555_), .B0(\asqrt[38] ), .Y(new_n22566_));
  NAND2X1  g22374(.A(new_n22566_), .B(new_n4165_), .Y(new_n22567_));
  OAI21X1  g22375(.A0(new_n22567_), .A1(new_n22559_), .B0(new_n22565_), .Y(new_n22568_));
  AOI21X1  g22376(.A0(new_n22568_), .A1(new_n22549_), .B0(new_n3863_), .Y(new_n22569_));
  AND2X1   g22377(.A(new_n21842_), .B(new_n21840_), .Y(new_n22570_));
  OR4X1    g22378(.A(new_n22128_), .B(new_n22570_), .C(new_n21811_), .D(new_n21841_), .Y(new_n22571_));
  OR2X1    g22379(.A(new_n22570_), .B(new_n21841_), .Y(new_n22572_));
  OAI21X1  g22380(.A0(new_n22572_), .A1(new_n22128_), .B0(new_n21811_), .Y(new_n22573_));
  AND2X1   g22381(.A(new_n22573_), .B(new_n22571_), .Y(new_n22574_));
  OAI21X1  g22382(.A0(new_n22558_), .A1(new_n22545_), .B0(new_n22566_), .Y(new_n22575_));
  AOI21X1  g22383(.A0(new_n22575_), .A1(\asqrt[39] ), .B0(\asqrt[40] ), .Y(new_n22576_));
  AOI21X1  g22384(.A0(new_n22576_), .A1(new_n22568_), .B0(new_n22574_), .Y(new_n22577_));
  OAI21X1  g22385(.A0(new_n22577_), .A1(new_n22569_), .B0(\asqrt[41] ), .Y(new_n22578_));
  OR4X1    g22386(.A(new_n22128_), .B(new_n21844_), .C(new_n21832_), .D(new_n21826_), .Y(new_n22579_));
  OR2X1    g22387(.A(new_n21844_), .B(new_n21826_), .Y(new_n22580_));
  OAI21X1  g22388(.A0(new_n22580_), .A1(new_n22128_), .B0(new_n21832_), .Y(new_n22581_));
  AND2X1   g22389(.A(new_n22581_), .B(new_n22579_), .Y(new_n22582_));
  NOR3X1   g22390(.A(new_n22577_), .B(new_n22569_), .C(\asqrt[41] ), .Y(new_n22583_));
  OAI21X1  g22391(.A0(new_n22583_), .A1(new_n22582_), .B0(new_n22578_), .Y(new_n22584_));
  AND2X1   g22392(.A(new_n22584_), .B(\asqrt[42] ), .Y(new_n22585_));
  OR2X1    g22393(.A(new_n22583_), .B(new_n22582_), .Y(new_n22586_));
  AND2X1   g22394(.A(new_n21888_), .B(new_n21887_), .Y(new_n22587_));
  NOR4X1   g22395(.A(new_n22128_), .B(new_n22587_), .C(new_n21851_), .D(new_n21886_), .Y(new_n22588_));
  AOI22X1  g22396(.A0(new_n21888_), .A1(new_n21887_), .B0(new_n21860_), .B1(\asqrt[41] ), .Y(new_n22589_));
  AOI21X1  g22397(.A0(new_n22589_), .A1(\asqrt[5] ), .B0(new_n21850_), .Y(new_n22590_));
  NOR2X1   g22398(.A(new_n22590_), .B(new_n22588_), .Y(new_n22591_));
  AND2X1   g22399(.A(new_n22578_), .B(new_n3276_), .Y(new_n22592_));
  AOI21X1  g22400(.A0(new_n22592_), .A1(new_n22586_), .B0(new_n22591_), .Y(new_n22593_));
  OAI21X1  g22401(.A0(new_n22593_), .A1(new_n22585_), .B0(\asqrt[43] ), .Y(new_n22594_));
  AND2X1   g22402(.A(new_n21861_), .B(new_n21854_), .Y(new_n22595_));
  OR4X1    g22403(.A(new_n22128_), .B(new_n22595_), .C(new_n21891_), .D(new_n21855_), .Y(new_n22596_));
  OR2X1    g22404(.A(new_n22595_), .B(new_n21855_), .Y(new_n22597_));
  OAI21X1  g22405(.A0(new_n22597_), .A1(new_n22128_), .B0(new_n21891_), .Y(new_n22598_));
  AND2X1   g22406(.A(new_n22598_), .B(new_n22596_), .Y(new_n22599_));
  INVX1    g22407(.A(new_n22599_), .Y(new_n22600_));
  AND2X1   g22408(.A(new_n22575_), .B(\asqrt[39] ), .Y(new_n22601_));
  OR2X1    g22409(.A(new_n22558_), .B(new_n22545_), .Y(new_n22602_));
  AND2X1   g22410(.A(new_n22566_), .B(new_n4165_), .Y(new_n22603_));
  AOI21X1  g22411(.A0(new_n22603_), .A1(new_n22602_), .B0(new_n22564_), .Y(new_n22604_));
  OAI21X1  g22412(.A0(new_n22604_), .A1(new_n22601_), .B0(\asqrt[40] ), .Y(new_n22605_));
  INVX1    g22413(.A(new_n22574_), .Y(new_n22606_));
  OAI21X1  g22414(.A0(new_n22548_), .A1(new_n4165_), .B0(new_n3863_), .Y(new_n22607_));
  OAI21X1  g22415(.A0(new_n22607_), .A1(new_n22604_), .B0(new_n22606_), .Y(new_n22608_));
  AOI21X1  g22416(.A0(new_n22608_), .A1(new_n22605_), .B0(new_n3564_), .Y(new_n22609_));
  INVX1    g22417(.A(new_n22582_), .Y(new_n22610_));
  NAND3X1  g22418(.A(new_n22608_), .B(new_n22605_), .C(new_n3564_), .Y(new_n22611_));
  AOI21X1  g22419(.A0(new_n22611_), .A1(new_n22610_), .B0(new_n22609_), .Y(new_n22612_));
  OAI21X1  g22420(.A0(new_n22612_), .A1(new_n3276_), .B0(new_n3008_), .Y(new_n22613_));
  OAI21X1  g22421(.A0(new_n22613_), .A1(new_n22593_), .B0(new_n22600_), .Y(new_n22614_));
  AOI21X1  g22422(.A0(new_n22614_), .A1(new_n22594_), .B0(new_n2769_), .Y(new_n22615_));
  OR4X1    g22423(.A(new_n22128_), .B(new_n21869_), .C(new_n21895_), .D(new_n21894_), .Y(new_n22616_));
  OR2X1    g22424(.A(new_n21869_), .B(new_n21894_), .Y(new_n22617_));
  OAI21X1  g22425(.A0(new_n22617_), .A1(new_n22128_), .B0(new_n21895_), .Y(new_n22618_));
  AND2X1   g22426(.A(new_n22618_), .B(new_n22616_), .Y(new_n22619_));
  INVX1    g22427(.A(new_n22619_), .Y(new_n22620_));
  NAND3X1  g22428(.A(new_n22614_), .B(new_n22594_), .C(new_n2769_), .Y(new_n22621_));
  AOI21X1  g22429(.A0(new_n22621_), .A1(new_n22620_), .B0(new_n22615_), .Y(new_n22622_));
  OR2X1    g22430(.A(new_n22622_), .B(new_n2570_), .Y(new_n22623_));
  OR2X1    g22431(.A(new_n22612_), .B(new_n3276_), .Y(new_n22624_));
  NOR2X1   g22432(.A(new_n22583_), .B(new_n22582_), .Y(new_n22625_));
  INVX1    g22433(.A(new_n22591_), .Y(new_n22626_));
  NAND2X1  g22434(.A(new_n22578_), .B(new_n3276_), .Y(new_n22627_));
  OAI21X1  g22435(.A0(new_n22627_), .A1(new_n22625_), .B0(new_n22626_), .Y(new_n22628_));
  AOI21X1  g22436(.A0(new_n22628_), .A1(new_n22624_), .B0(new_n3008_), .Y(new_n22629_));
  AOI21X1  g22437(.A0(new_n22584_), .A1(\asqrt[42] ), .B0(\asqrt[43] ), .Y(new_n22630_));
  AOI21X1  g22438(.A0(new_n22630_), .A1(new_n22628_), .B0(new_n22599_), .Y(new_n22631_));
  NOR3X1   g22439(.A(new_n22631_), .B(new_n22629_), .C(\asqrt[44] ), .Y(new_n22632_));
  NOR2X1   g22440(.A(new_n22632_), .B(new_n22619_), .Y(new_n22633_));
  OAI21X1  g22441(.A0(new_n21913_), .A1(new_n21911_), .B0(new_n21877_), .Y(new_n22634_));
  NOR3X1   g22442(.A(new_n22634_), .B(new_n22128_), .C(new_n21871_), .Y(new_n22635_));
  AOI22X1  g22443(.A0(new_n21878_), .A1(new_n21872_), .B0(new_n21870_), .B1(\asqrt[44] ), .Y(new_n22636_));
  AOI21X1  g22444(.A0(new_n22636_), .A1(\asqrt[5] ), .B0(new_n21877_), .Y(new_n22637_));
  NOR2X1   g22445(.A(new_n22637_), .B(new_n22635_), .Y(new_n22638_));
  INVX1    g22446(.A(new_n22638_), .Y(new_n22639_));
  OAI21X1  g22447(.A0(new_n22631_), .A1(new_n22629_), .B0(\asqrt[44] ), .Y(new_n22640_));
  NAND2X1  g22448(.A(new_n22640_), .B(new_n2570_), .Y(new_n22641_));
  OAI21X1  g22449(.A0(new_n22641_), .A1(new_n22633_), .B0(new_n22639_), .Y(new_n22642_));
  AOI21X1  g22450(.A0(new_n22642_), .A1(new_n22623_), .B0(new_n2263_), .Y(new_n22643_));
  AND2X1   g22451(.A(new_n21916_), .B(new_n21914_), .Y(new_n22644_));
  OR4X1    g22452(.A(new_n22128_), .B(new_n22644_), .C(new_n21885_), .D(new_n21915_), .Y(new_n22645_));
  OR2X1    g22453(.A(new_n22644_), .B(new_n21915_), .Y(new_n22646_));
  OAI21X1  g22454(.A0(new_n22646_), .A1(new_n22128_), .B0(new_n21885_), .Y(new_n22647_));
  AND2X1   g22455(.A(new_n22647_), .B(new_n22645_), .Y(new_n22648_));
  OAI21X1  g22456(.A0(new_n22632_), .A1(new_n22619_), .B0(new_n22640_), .Y(new_n22649_));
  AOI21X1  g22457(.A0(new_n22649_), .A1(\asqrt[45] ), .B0(\asqrt[46] ), .Y(new_n22650_));
  AOI21X1  g22458(.A0(new_n22650_), .A1(new_n22642_), .B0(new_n22648_), .Y(new_n22651_));
  OAI21X1  g22459(.A0(new_n22651_), .A1(new_n22643_), .B0(\asqrt[47] ), .Y(new_n22652_));
  OR4X1    g22460(.A(new_n22128_), .B(new_n21918_), .C(new_n21906_), .D(new_n21900_), .Y(new_n22653_));
  OR2X1    g22461(.A(new_n21918_), .B(new_n21900_), .Y(new_n22654_));
  OAI21X1  g22462(.A0(new_n22654_), .A1(new_n22128_), .B0(new_n21906_), .Y(new_n22655_));
  AND2X1   g22463(.A(new_n22655_), .B(new_n22653_), .Y(new_n22656_));
  NOR3X1   g22464(.A(new_n22651_), .B(new_n22643_), .C(\asqrt[47] ), .Y(new_n22657_));
  OAI21X1  g22465(.A0(new_n22657_), .A1(new_n22656_), .B0(new_n22652_), .Y(new_n22658_));
  AND2X1   g22466(.A(new_n22658_), .B(\asqrt[48] ), .Y(new_n22659_));
  OR2X1    g22467(.A(new_n22657_), .B(new_n22656_), .Y(new_n22660_));
  AND2X1   g22468(.A(new_n21962_), .B(new_n21961_), .Y(new_n22661_));
  NOR4X1   g22469(.A(new_n22128_), .B(new_n22661_), .C(new_n21925_), .D(new_n21960_), .Y(new_n22662_));
  AOI22X1  g22470(.A0(new_n21962_), .A1(new_n21961_), .B0(new_n21934_), .B1(\asqrt[47] ), .Y(new_n22663_));
  AOI21X1  g22471(.A0(new_n22663_), .A1(\asqrt[5] ), .B0(new_n21924_), .Y(new_n22664_));
  NOR2X1   g22472(.A(new_n22664_), .B(new_n22662_), .Y(new_n22665_));
  AND2X1   g22473(.A(new_n22652_), .B(new_n1834_), .Y(new_n22666_));
  AOI21X1  g22474(.A0(new_n22666_), .A1(new_n22660_), .B0(new_n22665_), .Y(new_n22667_));
  OAI21X1  g22475(.A0(new_n22667_), .A1(new_n22659_), .B0(\asqrt[49] ), .Y(new_n22668_));
  AND2X1   g22476(.A(new_n21935_), .B(new_n21928_), .Y(new_n22669_));
  OR4X1    g22477(.A(new_n22128_), .B(new_n22669_), .C(new_n21965_), .D(new_n21929_), .Y(new_n22670_));
  OR2X1    g22478(.A(new_n22669_), .B(new_n21929_), .Y(new_n22671_));
  OAI21X1  g22479(.A0(new_n22671_), .A1(new_n22128_), .B0(new_n21965_), .Y(new_n22672_));
  AND2X1   g22480(.A(new_n22672_), .B(new_n22670_), .Y(new_n22673_));
  INVX1    g22481(.A(new_n22673_), .Y(new_n22674_));
  AND2X1   g22482(.A(new_n22649_), .B(\asqrt[45] ), .Y(new_n22675_));
  OR2X1    g22483(.A(new_n22632_), .B(new_n22619_), .Y(new_n22676_));
  AND2X1   g22484(.A(new_n22640_), .B(new_n2570_), .Y(new_n22677_));
  AOI21X1  g22485(.A0(new_n22677_), .A1(new_n22676_), .B0(new_n22638_), .Y(new_n22678_));
  OAI21X1  g22486(.A0(new_n22678_), .A1(new_n22675_), .B0(\asqrt[46] ), .Y(new_n22679_));
  INVX1    g22487(.A(new_n22648_), .Y(new_n22680_));
  OAI21X1  g22488(.A0(new_n22622_), .A1(new_n2570_), .B0(new_n2263_), .Y(new_n22681_));
  OAI21X1  g22489(.A0(new_n22681_), .A1(new_n22678_), .B0(new_n22680_), .Y(new_n22682_));
  AOI21X1  g22490(.A0(new_n22682_), .A1(new_n22679_), .B0(new_n2040_), .Y(new_n22683_));
  INVX1    g22491(.A(new_n22656_), .Y(new_n22684_));
  NAND3X1  g22492(.A(new_n22682_), .B(new_n22679_), .C(new_n2040_), .Y(new_n22685_));
  AOI21X1  g22493(.A0(new_n22685_), .A1(new_n22684_), .B0(new_n22683_), .Y(new_n22686_));
  OAI21X1  g22494(.A0(new_n22686_), .A1(new_n1834_), .B0(new_n1632_), .Y(new_n22687_));
  OAI21X1  g22495(.A0(new_n22687_), .A1(new_n22667_), .B0(new_n22674_), .Y(new_n22688_));
  AOI21X1  g22496(.A0(new_n22688_), .A1(new_n22668_), .B0(new_n1469_), .Y(new_n22689_));
  OR4X1    g22497(.A(new_n22128_), .B(new_n21943_), .C(new_n21969_), .D(new_n21968_), .Y(new_n22690_));
  OR2X1    g22498(.A(new_n21943_), .B(new_n21968_), .Y(new_n22691_));
  OAI21X1  g22499(.A0(new_n22691_), .A1(new_n22128_), .B0(new_n21969_), .Y(new_n22692_));
  AND2X1   g22500(.A(new_n22692_), .B(new_n22690_), .Y(new_n22693_));
  INVX1    g22501(.A(new_n22693_), .Y(new_n22694_));
  NAND3X1  g22502(.A(new_n22688_), .B(new_n22668_), .C(new_n1469_), .Y(new_n22695_));
  AOI21X1  g22503(.A0(new_n22695_), .A1(new_n22694_), .B0(new_n22689_), .Y(new_n22696_));
  OR2X1    g22504(.A(new_n22696_), .B(new_n1277_), .Y(new_n22697_));
  OR2X1    g22505(.A(new_n22686_), .B(new_n1834_), .Y(new_n22698_));
  NOR2X1   g22506(.A(new_n22657_), .B(new_n22656_), .Y(new_n22699_));
  INVX1    g22507(.A(new_n22665_), .Y(new_n22700_));
  NAND2X1  g22508(.A(new_n22652_), .B(new_n1834_), .Y(new_n22701_));
  OAI21X1  g22509(.A0(new_n22701_), .A1(new_n22699_), .B0(new_n22700_), .Y(new_n22702_));
  AOI21X1  g22510(.A0(new_n22702_), .A1(new_n22698_), .B0(new_n1632_), .Y(new_n22703_));
  AOI21X1  g22511(.A0(new_n22658_), .A1(\asqrt[48] ), .B0(\asqrt[49] ), .Y(new_n22704_));
  AOI21X1  g22512(.A0(new_n22704_), .A1(new_n22702_), .B0(new_n22673_), .Y(new_n22705_));
  NOR3X1   g22513(.A(new_n22705_), .B(new_n22703_), .C(\asqrt[50] ), .Y(new_n22706_));
  NOR2X1   g22514(.A(new_n22706_), .B(new_n22693_), .Y(new_n22707_));
  OAI21X1  g22515(.A0(new_n21987_), .A1(new_n21985_), .B0(new_n21951_), .Y(new_n22708_));
  NOR3X1   g22516(.A(new_n22708_), .B(new_n22128_), .C(new_n21945_), .Y(new_n22709_));
  AOI22X1  g22517(.A0(new_n21952_), .A1(new_n21946_), .B0(new_n21944_), .B1(\asqrt[50] ), .Y(new_n22710_));
  AOI21X1  g22518(.A0(new_n22710_), .A1(\asqrt[5] ), .B0(new_n21951_), .Y(new_n22711_));
  NOR2X1   g22519(.A(new_n22711_), .B(new_n22709_), .Y(new_n22712_));
  INVX1    g22520(.A(new_n22712_), .Y(new_n22713_));
  OAI21X1  g22521(.A0(new_n22705_), .A1(new_n22703_), .B0(\asqrt[50] ), .Y(new_n22714_));
  NAND2X1  g22522(.A(new_n22714_), .B(new_n1277_), .Y(new_n22715_));
  OAI21X1  g22523(.A0(new_n22715_), .A1(new_n22707_), .B0(new_n22713_), .Y(new_n22716_));
  AOI21X1  g22524(.A0(new_n22716_), .A1(new_n22697_), .B0(new_n1111_), .Y(new_n22717_));
  AND2X1   g22525(.A(new_n21990_), .B(new_n21988_), .Y(new_n22718_));
  OR4X1    g22526(.A(new_n22128_), .B(new_n22718_), .C(new_n21959_), .D(new_n21989_), .Y(new_n22719_));
  OR2X1    g22527(.A(new_n22718_), .B(new_n21989_), .Y(new_n22720_));
  OAI21X1  g22528(.A0(new_n22720_), .A1(new_n22128_), .B0(new_n21959_), .Y(new_n22721_));
  AND2X1   g22529(.A(new_n22721_), .B(new_n22719_), .Y(new_n22722_));
  OAI21X1  g22530(.A0(new_n22706_), .A1(new_n22693_), .B0(new_n22714_), .Y(new_n22723_));
  AOI21X1  g22531(.A0(new_n22723_), .A1(\asqrt[51] ), .B0(\asqrt[52] ), .Y(new_n22724_));
  AOI21X1  g22532(.A0(new_n22724_), .A1(new_n22716_), .B0(new_n22722_), .Y(new_n22725_));
  OAI21X1  g22533(.A0(new_n22725_), .A1(new_n22717_), .B0(\asqrt[53] ), .Y(new_n22726_));
  OR4X1    g22534(.A(new_n22128_), .B(new_n21992_), .C(new_n21980_), .D(new_n21974_), .Y(new_n22727_));
  OR2X1    g22535(.A(new_n21992_), .B(new_n21974_), .Y(new_n22728_));
  OAI21X1  g22536(.A0(new_n22728_), .A1(new_n22128_), .B0(new_n21980_), .Y(new_n22729_));
  AND2X1   g22537(.A(new_n22729_), .B(new_n22727_), .Y(new_n22730_));
  NOR3X1   g22538(.A(new_n22725_), .B(new_n22717_), .C(\asqrt[53] ), .Y(new_n22731_));
  OAI21X1  g22539(.A0(new_n22731_), .A1(new_n22730_), .B0(new_n22726_), .Y(new_n22732_));
  AND2X1   g22540(.A(new_n22732_), .B(\asqrt[54] ), .Y(new_n22733_));
  OR2X1    g22541(.A(new_n22731_), .B(new_n22730_), .Y(new_n22734_));
  AND2X1   g22542(.A(new_n22036_), .B(new_n22035_), .Y(new_n22735_));
  NOR4X1   g22543(.A(new_n22128_), .B(new_n22735_), .C(new_n21999_), .D(new_n22034_), .Y(new_n22736_));
  AOI22X1  g22544(.A0(new_n22036_), .A1(new_n22035_), .B0(new_n22008_), .B1(\asqrt[53] ), .Y(new_n22737_));
  AOI21X1  g22545(.A0(new_n22737_), .A1(\asqrt[5] ), .B0(new_n21998_), .Y(new_n22738_));
  NOR2X1   g22546(.A(new_n22738_), .B(new_n22736_), .Y(new_n22739_));
  AND2X1   g22547(.A(new_n22726_), .B(new_n902_), .Y(new_n22740_));
  AOI21X1  g22548(.A0(new_n22740_), .A1(new_n22734_), .B0(new_n22739_), .Y(new_n22741_));
  OAI21X1  g22549(.A0(new_n22741_), .A1(new_n22733_), .B0(\asqrt[55] ), .Y(new_n22742_));
  AND2X1   g22550(.A(new_n22009_), .B(new_n22002_), .Y(new_n22743_));
  OR4X1    g22551(.A(new_n22128_), .B(new_n22743_), .C(new_n22039_), .D(new_n22003_), .Y(new_n22744_));
  OR2X1    g22552(.A(new_n22743_), .B(new_n22003_), .Y(new_n22745_));
  OAI21X1  g22553(.A0(new_n22745_), .A1(new_n22128_), .B0(new_n22039_), .Y(new_n22746_));
  AND2X1   g22554(.A(new_n22746_), .B(new_n22744_), .Y(new_n22747_));
  INVX1    g22555(.A(new_n22747_), .Y(new_n22748_));
  AND2X1   g22556(.A(new_n22723_), .B(\asqrt[51] ), .Y(new_n22749_));
  OR2X1    g22557(.A(new_n22706_), .B(new_n22693_), .Y(new_n22750_));
  AND2X1   g22558(.A(new_n22714_), .B(new_n1277_), .Y(new_n22751_));
  AOI21X1  g22559(.A0(new_n22751_), .A1(new_n22750_), .B0(new_n22712_), .Y(new_n22752_));
  OAI21X1  g22560(.A0(new_n22752_), .A1(new_n22749_), .B0(\asqrt[52] ), .Y(new_n22753_));
  INVX1    g22561(.A(new_n22722_), .Y(new_n22754_));
  OAI21X1  g22562(.A0(new_n22696_), .A1(new_n1277_), .B0(new_n1111_), .Y(new_n22755_));
  OAI21X1  g22563(.A0(new_n22755_), .A1(new_n22752_), .B0(new_n22754_), .Y(new_n22756_));
  AOI21X1  g22564(.A0(new_n22756_), .A1(new_n22753_), .B0(new_n968_), .Y(new_n22757_));
  INVX1    g22565(.A(new_n22730_), .Y(new_n22758_));
  NAND3X1  g22566(.A(new_n22756_), .B(new_n22753_), .C(new_n968_), .Y(new_n22759_));
  AOI21X1  g22567(.A0(new_n22759_), .A1(new_n22758_), .B0(new_n22757_), .Y(new_n22760_));
  OAI21X1  g22568(.A0(new_n22760_), .A1(new_n902_), .B0(new_n697_), .Y(new_n22761_));
  OAI21X1  g22569(.A0(new_n22761_), .A1(new_n22741_), .B0(new_n22748_), .Y(new_n22762_));
  AOI21X1  g22570(.A0(new_n22762_), .A1(new_n22742_), .B0(new_n582_), .Y(new_n22763_));
  OR4X1    g22571(.A(new_n22128_), .B(new_n22017_), .C(new_n22043_), .D(new_n22042_), .Y(new_n22764_));
  OR2X1    g22572(.A(new_n22017_), .B(new_n22042_), .Y(new_n22765_));
  OAI21X1  g22573(.A0(new_n22765_), .A1(new_n22128_), .B0(new_n22043_), .Y(new_n22766_));
  AND2X1   g22574(.A(new_n22766_), .B(new_n22764_), .Y(new_n22767_));
  INVX1    g22575(.A(new_n22767_), .Y(new_n22768_));
  NAND3X1  g22576(.A(new_n22762_), .B(new_n22742_), .C(new_n582_), .Y(new_n22769_));
  AOI21X1  g22577(.A0(new_n22769_), .A1(new_n22768_), .B0(new_n22763_), .Y(new_n22770_));
  OR2X1    g22578(.A(new_n22770_), .B(new_n481_), .Y(new_n22771_));
  OR2X1    g22579(.A(new_n22760_), .B(new_n902_), .Y(new_n22772_));
  NOR2X1   g22580(.A(new_n22731_), .B(new_n22730_), .Y(new_n22773_));
  INVX1    g22581(.A(new_n22739_), .Y(new_n22774_));
  NAND2X1  g22582(.A(new_n22726_), .B(new_n902_), .Y(new_n22775_));
  OAI21X1  g22583(.A0(new_n22775_), .A1(new_n22773_), .B0(new_n22774_), .Y(new_n22776_));
  AOI21X1  g22584(.A0(new_n22776_), .A1(new_n22772_), .B0(new_n697_), .Y(new_n22777_));
  AOI21X1  g22585(.A0(new_n22732_), .A1(\asqrt[54] ), .B0(\asqrt[55] ), .Y(new_n22778_));
  AOI21X1  g22586(.A0(new_n22778_), .A1(new_n22776_), .B0(new_n22747_), .Y(new_n22779_));
  NOR3X1   g22587(.A(new_n22779_), .B(new_n22777_), .C(\asqrt[56] ), .Y(new_n22780_));
  NOR2X1   g22588(.A(new_n22780_), .B(new_n22767_), .Y(new_n22781_));
  OAI21X1  g22589(.A0(new_n22061_), .A1(new_n22059_), .B0(new_n22025_), .Y(new_n22782_));
  NOR3X1   g22590(.A(new_n22782_), .B(new_n22128_), .C(new_n22019_), .Y(new_n22783_));
  AOI22X1  g22591(.A0(new_n22026_), .A1(new_n22020_), .B0(new_n22018_), .B1(\asqrt[56] ), .Y(new_n22784_));
  AOI21X1  g22592(.A0(new_n22784_), .A1(\asqrt[5] ), .B0(new_n22025_), .Y(new_n22785_));
  NOR2X1   g22593(.A(new_n22785_), .B(new_n22783_), .Y(new_n22786_));
  INVX1    g22594(.A(new_n22786_), .Y(new_n22787_));
  OAI21X1  g22595(.A0(new_n22779_), .A1(new_n22777_), .B0(\asqrt[56] ), .Y(new_n22788_));
  NAND2X1  g22596(.A(new_n22788_), .B(new_n481_), .Y(new_n22789_));
  OAI21X1  g22597(.A0(new_n22789_), .A1(new_n22781_), .B0(new_n22787_), .Y(new_n22790_));
  AOI21X1  g22598(.A0(new_n22790_), .A1(new_n22771_), .B0(new_n399_), .Y(new_n22791_));
  AND2X1   g22599(.A(new_n22064_), .B(new_n22062_), .Y(new_n22792_));
  OR4X1    g22600(.A(new_n22128_), .B(new_n22792_), .C(new_n22033_), .D(new_n22063_), .Y(new_n22793_));
  OR2X1    g22601(.A(new_n22792_), .B(new_n22063_), .Y(new_n22794_));
  OAI21X1  g22602(.A0(new_n22794_), .A1(new_n22128_), .B0(new_n22033_), .Y(new_n22795_));
  AND2X1   g22603(.A(new_n22795_), .B(new_n22793_), .Y(new_n22796_));
  OAI21X1  g22604(.A0(new_n22780_), .A1(new_n22767_), .B0(new_n22788_), .Y(new_n22797_));
  AOI21X1  g22605(.A0(new_n22797_), .A1(\asqrt[57] ), .B0(\asqrt[58] ), .Y(new_n22798_));
  AOI21X1  g22606(.A0(new_n22798_), .A1(new_n22790_), .B0(new_n22796_), .Y(new_n22799_));
  OAI21X1  g22607(.A0(new_n22799_), .A1(new_n22791_), .B0(\asqrt[59] ), .Y(new_n22800_));
  OR4X1    g22608(.A(new_n22128_), .B(new_n22066_), .C(new_n22054_), .D(new_n22048_), .Y(new_n22801_));
  OR2X1    g22609(.A(new_n22066_), .B(new_n22048_), .Y(new_n22802_));
  OAI21X1  g22610(.A0(new_n22802_), .A1(new_n22128_), .B0(new_n22054_), .Y(new_n22803_));
  AND2X1   g22611(.A(new_n22803_), .B(new_n22801_), .Y(new_n22804_));
  NOR3X1   g22612(.A(new_n22799_), .B(new_n22791_), .C(\asqrt[59] ), .Y(new_n22805_));
  OAI21X1  g22613(.A0(new_n22805_), .A1(new_n22804_), .B0(new_n22800_), .Y(new_n22806_));
  AND2X1   g22614(.A(new_n22806_), .B(\asqrt[60] ), .Y(new_n22807_));
  OR2X1    g22615(.A(new_n22805_), .B(new_n22804_), .Y(new_n22808_));
  AND2X1   g22616(.A(new_n22800_), .B(new_n292_), .Y(new_n22809_));
  AND2X1   g22617(.A(new_n22113_), .B(new_n22112_), .Y(new_n22810_));
  NOR4X1   g22618(.A(new_n22128_), .B(new_n22075_), .C(new_n22810_), .D(new_n22111_), .Y(new_n22811_));
  AOI22X1  g22619(.A0(new_n22113_), .A1(new_n22112_), .B0(new_n22082_), .B1(\asqrt[59] ), .Y(new_n22812_));
  AOI21X1  g22620(.A0(new_n22812_), .A1(\asqrt[5] ), .B0(new_n22074_), .Y(new_n22813_));
  NOR2X1   g22621(.A(new_n22813_), .B(new_n22811_), .Y(new_n22814_));
  AOI21X1  g22622(.A0(new_n22809_), .A1(new_n22808_), .B0(new_n22814_), .Y(new_n22815_));
  OAI21X1  g22623(.A0(new_n22815_), .A1(new_n22807_), .B0(\asqrt[61] ), .Y(new_n22816_));
  AND2X1   g22624(.A(new_n22083_), .B(new_n22076_), .Y(new_n22817_));
  OR4X1    g22625(.A(new_n22128_), .B(new_n22817_), .C(new_n22116_), .D(new_n22077_), .Y(new_n22818_));
  OR2X1    g22626(.A(new_n22817_), .B(new_n22077_), .Y(new_n22819_));
  OAI21X1  g22627(.A0(new_n22819_), .A1(new_n22128_), .B0(new_n22116_), .Y(new_n22820_));
  AND2X1   g22628(.A(new_n22820_), .B(new_n22818_), .Y(new_n22821_));
  INVX1    g22629(.A(new_n22821_), .Y(new_n22822_));
  AND2X1   g22630(.A(new_n22797_), .B(\asqrt[57] ), .Y(new_n22823_));
  OR2X1    g22631(.A(new_n22780_), .B(new_n22767_), .Y(new_n22824_));
  AND2X1   g22632(.A(new_n22788_), .B(new_n481_), .Y(new_n22825_));
  AOI21X1  g22633(.A0(new_n22825_), .A1(new_n22824_), .B0(new_n22786_), .Y(new_n22826_));
  OAI21X1  g22634(.A0(new_n22826_), .A1(new_n22823_), .B0(\asqrt[58] ), .Y(new_n22827_));
  INVX1    g22635(.A(new_n22796_), .Y(new_n22828_));
  OAI21X1  g22636(.A0(new_n22770_), .A1(new_n481_), .B0(new_n399_), .Y(new_n22829_));
  OAI21X1  g22637(.A0(new_n22829_), .A1(new_n22826_), .B0(new_n22828_), .Y(new_n22830_));
  AOI21X1  g22638(.A0(new_n22830_), .A1(new_n22827_), .B0(new_n328_), .Y(new_n22831_));
  INVX1    g22639(.A(new_n22804_), .Y(new_n22832_));
  NAND3X1  g22640(.A(new_n22830_), .B(new_n22827_), .C(new_n328_), .Y(new_n22833_));
  AOI21X1  g22641(.A0(new_n22833_), .A1(new_n22832_), .B0(new_n22831_), .Y(new_n22834_));
  OAI21X1  g22642(.A0(new_n22834_), .A1(new_n292_), .B0(new_n217_), .Y(new_n22835_));
  OAI21X1  g22643(.A0(new_n22835_), .A1(new_n22815_), .B0(new_n22822_), .Y(new_n22836_));
  AOI21X1  g22644(.A0(new_n22836_), .A1(new_n22816_), .B0(new_n199_), .Y(new_n22837_));
  OR4X1    g22645(.A(new_n22128_), .B(new_n22091_), .C(new_n22120_), .D(new_n22119_), .Y(new_n22838_));
  NAND2X1  g22646(.A(new_n22121_), .B(new_n22085_), .Y(new_n22839_));
  OAI21X1  g22647(.A0(new_n22839_), .A1(new_n22128_), .B0(new_n22120_), .Y(new_n22840_));
  AND2X1   g22648(.A(new_n22840_), .B(new_n22838_), .Y(new_n22841_));
  INVX1    g22649(.A(new_n22841_), .Y(new_n22842_));
  NAND3X1  g22650(.A(new_n22836_), .B(new_n22816_), .C(new_n199_), .Y(new_n22843_));
  AOI21X1  g22651(.A0(new_n22843_), .A1(new_n22842_), .B0(new_n22837_), .Y(new_n22844_));
  AOI21X1  g22652(.A0(new_n22100_), .A1(new_n22094_), .B0(new_n22131_), .Y(new_n22845_));
  NAND3X1  g22653(.A(new_n22845_), .B(\asqrt[5] ), .C(new_n22129_), .Y(new_n22846_));
  OAI22X1  g22654(.A0(new_n22132_), .A1(new_n22130_), .B0(new_n22122_), .B1(new_n199_), .Y(new_n22847_));
  OAI21X1  g22655(.A0(new_n22847_), .A1(new_n22128_), .B0(new_n22131_), .Y(new_n22848_));
  AND2X1   g22656(.A(new_n22848_), .B(new_n22846_), .Y(new_n22849_));
  INVX1    g22657(.A(new_n22849_), .Y(new_n22850_));
  AND2X1   g22658(.A(new_n22136_), .B(new_n22133_), .Y(new_n22851_));
  AOI21X1  g22659(.A0(new_n22133_), .A1(new_n22129_), .B0(new_n22105_), .Y(new_n22852_));
  AOI21X1  g22660(.A0(new_n22852_), .A1(\asqrt[5] ), .B0(new_n22851_), .Y(new_n22853_));
  AND2X1   g22661(.A(new_n22853_), .B(new_n22850_), .Y(new_n22854_));
  INVX1    g22662(.A(new_n22854_), .Y(new_n22855_));
  OAI21X1  g22663(.A0(new_n22855_), .A1(new_n22844_), .B0(new_n193_), .Y(new_n22856_));
  OR2X1    g22664(.A(new_n22834_), .B(new_n292_), .Y(new_n22857_));
  NOR2X1   g22665(.A(new_n22805_), .B(new_n22804_), .Y(new_n22858_));
  NAND2X1  g22666(.A(new_n22800_), .B(new_n292_), .Y(new_n22859_));
  INVX1    g22667(.A(new_n22814_), .Y(new_n22860_));
  OAI21X1  g22668(.A0(new_n22859_), .A1(new_n22858_), .B0(new_n22860_), .Y(new_n22861_));
  AOI21X1  g22669(.A0(new_n22861_), .A1(new_n22857_), .B0(new_n217_), .Y(new_n22862_));
  AOI21X1  g22670(.A0(new_n22806_), .A1(\asqrt[60] ), .B0(\asqrt[61] ), .Y(new_n22863_));
  AOI21X1  g22671(.A0(new_n22863_), .A1(new_n22861_), .B0(new_n22821_), .Y(new_n22864_));
  NOR3X1   g22672(.A(new_n22864_), .B(new_n22862_), .C(\asqrt[62] ), .Y(new_n22865_));
  OR2X1    g22673(.A(new_n22865_), .B(new_n22841_), .Y(new_n22866_));
  OAI21X1  g22674(.A0(new_n22864_), .A1(new_n22862_), .B0(\asqrt[62] ), .Y(new_n22867_));
  AND2X1   g22675(.A(new_n22849_), .B(new_n22867_), .Y(new_n22868_));
  NAND2X1  g22676(.A(new_n22133_), .B(new_n22129_), .Y(new_n22869_));
  AOI21X1  g22677(.A0(\asqrt[5] ), .A1(new_n22106_), .B0(new_n22869_), .Y(new_n22870_));
  OR2X1    g22678(.A(new_n22852_), .B(new_n193_), .Y(new_n22871_));
  NOR2X1   g22679(.A(new_n22871_), .B(new_n22870_), .Y(new_n22872_));
  AOI21X1  g22680(.A0(new_n22868_), .A1(new_n22866_), .B0(new_n22872_), .Y(new_n22873_));
  AND2X1   g22681(.A(new_n22873_), .B(new_n22856_), .Y(new_n22874_));
  INVX1    g22682(.A(new_n22874_), .Y(\asqrt[4] ));
  INVX1    g22683(.A(\a[8] ), .Y(new_n22876_));
  AOI21X1  g22684(.A0(new_n22873_), .A1(new_n22856_), .B0(new_n22876_), .Y(new_n22877_));
  NOR3X1   g22685(.A(\a[8] ), .B(\a[7] ), .C(\a[6] ), .Y(new_n22878_));
  OAI21X1  g22686(.A0(new_n22878_), .A1(new_n22877_), .B0(\asqrt[5] ), .Y(new_n22879_));
  INVX1    g22687(.A(new_n22878_), .Y(new_n22880_));
  NAND2X1  g22688(.A(new_n22880_), .B(new_n22126_), .Y(new_n22881_));
  NOR4X1   g22689(.A(new_n22881_), .B(new_n22877_), .C(new_n22851_), .D(new_n22199_), .Y(new_n22882_));
  INVX1    g22690(.A(\a[9] ), .Y(new_n22883_));
  AOI21X1  g22691(.A0(new_n22873_), .A1(new_n22856_), .B0(\a[8] ), .Y(new_n22884_));
  OAI21X1  g22692(.A0(new_n22865_), .A1(new_n22841_), .B0(new_n22867_), .Y(new_n22885_));
  AOI21X1  g22693(.A0(new_n22854_), .A1(new_n22885_), .B0(\asqrt[63] ), .Y(new_n22886_));
  NOR2X1   g22694(.A(new_n22865_), .B(new_n22841_), .Y(new_n22887_));
  NAND2X1  g22695(.A(new_n22849_), .B(new_n22867_), .Y(new_n22888_));
  OAI22X1  g22696(.A0(new_n22871_), .A1(new_n22870_), .B0(new_n22888_), .B1(new_n22887_), .Y(new_n22889_));
  OAI21X1  g22697(.A0(new_n22889_), .A1(new_n22886_), .B0(new_n22140_), .Y(new_n22890_));
  OAI21X1  g22698(.A0(new_n22884_), .A1(new_n22883_), .B0(new_n22890_), .Y(new_n22891_));
  OAI21X1  g22699(.A0(new_n22891_), .A1(new_n22882_), .B0(new_n22879_), .Y(new_n22892_));
  AND2X1   g22700(.A(new_n22892_), .B(\asqrt[6] ), .Y(new_n22893_));
  OR2X1    g22701(.A(new_n22891_), .B(new_n22882_), .Y(new_n22894_));
  AND2X1   g22702(.A(new_n22879_), .B(new_n21393_), .Y(new_n22895_));
  AND2X1   g22703(.A(new_n22868_), .B(new_n22866_), .Y(new_n22896_));
  OR4X1    g22704(.A(new_n22872_), .B(new_n22896_), .C(new_n22886_), .D(new_n22128_), .Y(new_n22897_));
  AOI21X1  g22705(.A0(new_n22897_), .A1(new_n22890_), .B0(new_n22149_), .Y(new_n22898_));
  AOI21X1  g22706(.A0(new_n22873_), .A1(new_n22856_), .B0(new_n22144_), .Y(new_n22899_));
  NOR4X1   g22707(.A(new_n22872_), .B(new_n22896_), .C(new_n22886_), .D(new_n22128_), .Y(new_n22900_));
  NOR3X1   g22708(.A(new_n22900_), .B(new_n22899_), .C(\a[10] ), .Y(new_n22901_));
  NOR2X1   g22709(.A(new_n22901_), .B(new_n22898_), .Y(new_n22902_));
  AOI21X1  g22710(.A0(new_n22895_), .A1(new_n22894_), .B0(new_n22902_), .Y(new_n22903_));
  OAI21X1  g22711(.A0(new_n22903_), .A1(new_n22893_), .B0(\asqrt[7] ), .Y(new_n22904_));
  AND2X1   g22712(.A(new_n22195_), .B(new_n22193_), .Y(new_n22905_));
  NOR3X1   g22713(.A(new_n22905_), .B(new_n22148_), .C(new_n22142_), .Y(new_n22906_));
  OAI21X1  g22714(.A0(new_n22889_), .A1(new_n22886_), .B0(new_n22906_), .Y(new_n22907_));
  AOI21X1  g22715(.A0(new_n22141_), .A1(\asqrt[6] ), .B0(new_n22148_), .Y(new_n22908_));
  OAI21X1  g22716(.A0(new_n22889_), .A1(new_n22886_), .B0(new_n22908_), .Y(new_n22909_));
  NAND2X1  g22717(.A(new_n22909_), .B(new_n22905_), .Y(new_n22910_));
  NAND2X1  g22718(.A(new_n22910_), .B(new_n22907_), .Y(new_n22911_));
  OAI21X1  g22719(.A0(new_n22889_), .A1(new_n22886_), .B0(\a[8] ), .Y(new_n22912_));
  AOI21X1  g22720(.A0(new_n22880_), .A1(new_n22912_), .B0(new_n22128_), .Y(new_n22913_));
  OR4X1    g22721(.A(new_n22881_), .B(new_n22877_), .C(new_n22851_), .D(new_n22199_), .Y(new_n22914_));
  OAI21X1  g22722(.A0(new_n22889_), .A1(new_n22886_), .B0(new_n22876_), .Y(new_n22915_));
  AOI21X1  g22723(.A0(new_n22915_), .A1(\a[9] ), .B0(new_n22899_), .Y(new_n22916_));
  AOI21X1  g22724(.A0(new_n22916_), .A1(new_n22914_), .B0(new_n22913_), .Y(new_n22917_));
  OAI21X1  g22725(.A0(new_n22917_), .A1(new_n21393_), .B0(new_n20676_), .Y(new_n22918_));
  OAI21X1  g22726(.A0(new_n22918_), .A1(new_n22903_), .B0(new_n22911_), .Y(new_n22919_));
  AOI21X1  g22727(.A0(new_n22919_), .A1(new_n22904_), .B0(new_n19976_), .Y(new_n22920_));
  AND2X1   g22728(.A(new_n22198_), .B(new_n22196_), .Y(new_n22921_));
  NOR3X1   g22729(.A(new_n22163_), .B(new_n22921_), .C(new_n22197_), .Y(new_n22922_));
  OAI21X1  g22730(.A0(new_n22889_), .A1(new_n22886_), .B0(new_n22922_), .Y(new_n22923_));
  NOR2X1   g22731(.A(new_n22921_), .B(new_n22197_), .Y(new_n22924_));
  OAI21X1  g22732(.A0(new_n22889_), .A1(new_n22886_), .B0(new_n22924_), .Y(new_n22925_));
  NAND2X1  g22733(.A(new_n22925_), .B(new_n22163_), .Y(new_n22926_));
  AND2X1   g22734(.A(new_n22926_), .B(new_n22923_), .Y(new_n22927_));
  INVX1    g22735(.A(new_n22927_), .Y(new_n22928_));
  NAND3X1  g22736(.A(new_n22919_), .B(new_n22904_), .C(new_n19976_), .Y(new_n22929_));
  AOI21X1  g22737(.A0(new_n22929_), .A1(new_n22928_), .B0(new_n22920_), .Y(new_n22930_));
  OR2X1    g22738(.A(new_n22930_), .B(new_n19273_), .Y(new_n22931_));
  OR2X1    g22739(.A(new_n22917_), .B(new_n21393_), .Y(new_n22932_));
  NOR2X1   g22740(.A(new_n22891_), .B(new_n22882_), .Y(new_n22933_));
  OR2X1    g22741(.A(new_n22913_), .B(\asqrt[6] ), .Y(new_n22934_));
  OR2X1    g22742(.A(new_n22901_), .B(new_n22898_), .Y(new_n22935_));
  OAI21X1  g22743(.A0(new_n22934_), .A1(new_n22933_), .B0(new_n22935_), .Y(new_n22936_));
  AOI21X1  g22744(.A0(new_n22936_), .A1(new_n22932_), .B0(new_n20676_), .Y(new_n22937_));
  AOI21X1  g22745(.A0(new_n22892_), .A1(\asqrt[6] ), .B0(\asqrt[7] ), .Y(new_n22938_));
  AOI22X1  g22746(.A0(new_n22938_), .A1(new_n22936_), .B0(new_n22910_), .B1(new_n22907_), .Y(new_n22939_));
  NOR3X1   g22747(.A(new_n22939_), .B(new_n22937_), .C(\asqrt[8] ), .Y(new_n22940_));
  NOR2X1   g22748(.A(new_n22940_), .B(new_n22927_), .Y(new_n22941_));
  NAND4X1  g22749(.A(\asqrt[4] ), .B(new_n22172_), .C(new_n22170_), .D(new_n22204_), .Y(new_n22942_));
  NOR3X1   g22750(.A(new_n22874_), .B(new_n22205_), .C(new_n22165_), .Y(new_n22943_));
  OAI21X1  g22751(.A0(new_n22943_), .A1(new_n22170_), .B0(new_n22942_), .Y(new_n22944_));
  OR2X1    g22752(.A(new_n22920_), .B(\asqrt[9] ), .Y(new_n22945_));
  OAI21X1  g22753(.A0(new_n22945_), .A1(new_n22941_), .B0(new_n22944_), .Y(new_n22946_));
  AOI21X1  g22754(.A0(new_n22946_), .A1(new_n22931_), .B0(new_n18591_), .Y(new_n22947_));
  AOI21X1  g22755(.A0(new_n22220_), .A1(new_n22219_), .B0(new_n22181_), .Y(new_n22948_));
  NAND3X1  g22756(.A(new_n22948_), .B(\asqrt[4] ), .C(new_n22174_), .Y(new_n22949_));
  OAI22X1  g22757(.A0(new_n22182_), .A1(new_n22175_), .B0(new_n22173_), .B1(new_n19273_), .Y(new_n22950_));
  OAI21X1  g22758(.A0(new_n22950_), .A1(new_n22874_), .B0(new_n22181_), .Y(new_n22951_));
  AND2X1   g22759(.A(new_n22951_), .B(new_n22949_), .Y(new_n22952_));
  OAI21X1  g22760(.A0(new_n22939_), .A1(new_n22937_), .B0(\asqrt[8] ), .Y(new_n22953_));
  OAI21X1  g22761(.A0(new_n22940_), .A1(new_n22927_), .B0(new_n22953_), .Y(new_n22954_));
  AOI21X1  g22762(.A0(new_n22954_), .A1(\asqrt[9] ), .B0(\asqrt[10] ), .Y(new_n22955_));
  AOI21X1  g22763(.A0(new_n22955_), .A1(new_n22946_), .B0(new_n22952_), .Y(new_n22956_));
  OAI21X1  g22764(.A0(new_n22956_), .A1(new_n22947_), .B0(\asqrt[11] ), .Y(new_n22957_));
  AND2X1   g22765(.A(new_n22207_), .B(new_n22183_), .Y(new_n22958_));
  NOR3X1   g22766(.A(new_n22958_), .B(new_n22223_), .C(new_n22184_), .Y(new_n22959_));
  OAI21X1  g22767(.A0(new_n22889_), .A1(new_n22886_), .B0(new_n22959_), .Y(new_n22960_));
  OR2X1    g22768(.A(new_n22958_), .B(new_n22184_), .Y(new_n22961_));
  OAI21X1  g22769(.A0(new_n22961_), .A1(new_n22874_), .B0(new_n22223_), .Y(new_n22962_));
  AND2X1   g22770(.A(new_n22962_), .B(new_n22960_), .Y(new_n22963_));
  NOR3X1   g22771(.A(new_n22956_), .B(new_n22947_), .C(\asqrt[11] ), .Y(new_n22964_));
  OAI21X1  g22772(.A0(new_n22964_), .A1(new_n22963_), .B0(new_n22957_), .Y(new_n22965_));
  AND2X1   g22773(.A(new_n22965_), .B(\asqrt[12] ), .Y(new_n22966_));
  OR2X1    g22774(.A(new_n22964_), .B(new_n22963_), .Y(new_n22967_));
  NAND4X1  g22775(.A(\asqrt[4] ), .B(new_n22226_), .C(new_n22213_), .D(new_n22209_), .Y(new_n22968_));
  NAND2X1  g22776(.A(new_n22226_), .B(new_n22209_), .Y(new_n22969_));
  OAI21X1  g22777(.A0(new_n22969_), .A1(new_n22874_), .B0(new_n22217_), .Y(new_n22970_));
  AND2X1   g22778(.A(new_n22970_), .B(new_n22968_), .Y(new_n22971_));
  AND2X1   g22779(.A(new_n22957_), .B(new_n17262_), .Y(new_n22972_));
  AOI21X1  g22780(.A0(new_n22972_), .A1(new_n22967_), .B0(new_n22971_), .Y(new_n22973_));
  OAI21X1  g22781(.A0(new_n22973_), .A1(new_n22966_), .B0(\asqrt[13] ), .Y(new_n22974_));
  AND2X1   g22782(.A(new_n22234_), .B(new_n22227_), .Y(new_n22975_));
  OR4X1    g22783(.A(new_n22874_), .B(new_n22975_), .C(new_n22272_), .D(new_n22216_), .Y(new_n22976_));
  OAI22X1  g22784(.A0(new_n22273_), .A1(new_n22271_), .B0(new_n22243_), .B1(new_n17262_), .Y(new_n22977_));
  OAI21X1  g22785(.A0(new_n22977_), .A1(new_n22874_), .B0(new_n22272_), .Y(new_n22978_));
  AND2X1   g22786(.A(new_n22978_), .B(new_n22976_), .Y(new_n22979_));
  INVX1    g22787(.A(new_n22979_), .Y(new_n22980_));
  AND2X1   g22788(.A(new_n22954_), .B(\asqrt[9] ), .Y(new_n22981_));
  OR2X1    g22789(.A(new_n22940_), .B(new_n22927_), .Y(new_n22982_));
  INVX1    g22790(.A(new_n22944_), .Y(new_n22983_));
  NOR2X1   g22791(.A(new_n22920_), .B(\asqrt[9] ), .Y(new_n22984_));
  AOI21X1  g22792(.A0(new_n22984_), .A1(new_n22982_), .B0(new_n22983_), .Y(new_n22985_));
  OAI21X1  g22793(.A0(new_n22985_), .A1(new_n22981_), .B0(\asqrt[10] ), .Y(new_n22986_));
  INVX1    g22794(.A(new_n22952_), .Y(new_n22987_));
  OAI21X1  g22795(.A0(new_n22930_), .A1(new_n19273_), .B0(new_n18591_), .Y(new_n22988_));
  OAI21X1  g22796(.A0(new_n22988_), .A1(new_n22985_), .B0(new_n22987_), .Y(new_n22989_));
  AOI21X1  g22797(.A0(new_n22989_), .A1(new_n22986_), .B0(new_n17927_), .Y(new_n22990_));
  INVX1    g22798(.A(new_n22963_), .Y(new_n22991_));
  NAND3X1  g22799(.A(new_n22989_), .B(new_n22986_), .C(new_n17927_), .Y(new_n22992_));
  AOI21X1  g22800(.A0(new_n22992_), .A1(new_n22991_), .B0(new_n22990_), .Y(new_n22993_));
  OAI21X1  g22801(.A0(new_n22993_), .A1(new_n17262_), .B0(new_n16617_), .Y(new_n22994_));
  OAI21X1  g22802(.A0(new_n22994_), .A1(new_n22973_), .B0(new_n22980_), .Y(new_n22995_));
  AOI21X1  g22803(.A0(new_n22995_), .A1(new_n22974_), .B0(new_n15990_), .Y(new_n22996_));
  AND2X1   g22804(.A(new_n22276_), .B(new_n22274_), .Y(new_n22997_));
  NOR3X1   g22805(.A(new_n22997_), .B(new_n22242_), .C(new_n22275_), .Y(new_n22998_));
  NOR3X1   g22806(.A(new_n22874_), .B(new_n22997_), .C(new_n22275_), .Y(new_n22999_));
  NOR2X1   g22807(.A(new_n22999_), .B(new_n22241_), .Y(new_n23000_));
  AOI21X1  g22808(.A0(new_n22998_), .A1(\asqrt[4] ), .B0(new_n23000_), .Y(new_n23001_));
  INVX1    g22809(.A(new_n23001_), .Y(new_n23002_));
  NAND3X1  g22810(.A(new_n22995_), .B(new_n22974_), .C(new_n15990_), .Y(new_n23003_));
  AOI21X1  g22811(.A0(new_n23003_), .A1(new_n23002_), .B0(new_n22996_), .Y(new_n23004_));
  OR2X1    g22812(.A(new_n23004_), .B(new_n15362_), .Y(new_n23005_));
  OR2X1    g22813(.A(new_n22993_), .B(new_n17262_), .Y(new_n23006_));
  NOR2X1   g22814(.A(new_n22964_), .B(new_n22963_), .Y(new_n23007_));
  INVX1    g22815(.A(new_n22971_), .Y(new_n23008_));
  NAND2X1  g22816(.A(new_n22957_), .B(new_n17262_), .Y(new_n23009_));
  OAI21X1  g22817(.A0(new_n23009_), .A1(new_n23007_), .B0(new_n23008_), .Y(new_n23010_));
  AOI21X1  g22818(.A0(new_n23010_), .A1(new_n23006_), .B0(new_n16617_), .Y(new_n23011_));
  AOI21X1  g22819(.A0(new_n22965_), .A1(\asqrt[12] ), .B0(\asqrt[13] ), .Y(new_n23012_));
  AOI21X1  g22820(.A0(new_n23012_), .A1(new_n23010_), .B0(new_n22979_), .Y(new_n23013_));
  NOR3X1   g22821(.A(new_n23013_), .B(new_n23011_), .C(\asqrt[14] ), .Y(new_n23014_));
  NOR2X1   g22822(.A(new_n23014_), .B(new_n23001_), .Y(new_n23015_));
  NAND4X1  g22823(.A(\asqrt[4] ), .B(new_n22252_), .C(new_n22250_), .D(new_n22278_), .Y(new_n23016_));
  NAND2X1  g22824(.A(new_n22252_), .B(new_n22278_), .Y(new_n23017_));
  OAI21X1  g22825(.A0(new_n23017_), .A1(new_n22874_), .B0(new_n22251_), .Y(new_n23018_));
  AND2X1   g22826(.A(new_n23018_), .B(new_n23016_), .Y(new_n23019_));
  INVX1    g22827(.A(new_n23019_), .Y(new_n23020_));
  OAI21X1  g22828(.A0(new_n23013_), .A1(new_n23011_), .B0(\asqrt[14] ), .Y(new_n23021_));
  NAND2X1  g22829(.A(new_n23021_), .B(new_n15362_), .Y(new_n23022_));
  OAI21X1  g22830(.A0(new_n23022_), .A1(new_n23015_), .B0(new_n23020_), .Y(new_n23023_));
  AOI21X1  g22831(.A0(new_n23023_), .A1(new_n23005_), .B0(new_n14754_), .Y(new_n23024_));
  AND2X1   g22832(.A(new_n22294_), .B(new_n22293_), .Y(new_n23025_));
  OR4X1    g22833(.A(new_n22874_), .B(new_n23025_), .C(new_n22261_), .D(new_n22292_), .Y(new_n23026_));
  OAI22X1  g22834(.A0(new_n22262_), .A1(new_n22255_), .B0(new_n22253_), .B1(new_n15362_), .Y(new_n23027_));
  OAI21X1  g22835(.A0(new_n23027_), .A1(new_n22874_), .B0(new_n22261_), .Y(new_n23028_));
  AND2X1   g22836(.A(new_n23028_), .B(new_n23026_), .Y(new_n23029_));
  OAI21X1  g22837(.A0(new_n23014_), .A1(new_n23001_), .B0(new_n23021_), .Y(new_n23030_));
  AOI21X1  g22838(.A0(new_n23030_), .A1(\asqrt[15] ), .B0(\asqrt[16] ), .Y(new_n23031_));
  AOI21X1  g22839(.A0(new_n23031_), .A1(new_n23023_), .B0(new_n23029_), .Y(new_n23032_));
  OAI21X1  g22840(.A0(new_n23032_), .A1(new_n23024_), .B0(\asqrt[17] ), .Y(new_n23033_));
  AND2X1   g22841(.A(new_n22281_), .B(new_n22263_), .Y(new_n23034_));
  NOR3X1   g22842(.A(new_n23034_), .B(new_n22297_), .C(new_n22264_), .Y(new_n23035_));
  NOR3X1   g22843(.A(new_n22874_), .B(new_n23034_), .C(new_n22264_), .Y(new_n23036_));
  NOR2X1   g22844(.A(new_n23036_), .B(new_n22269_), .Y(new_n23037_));
  AOI21X1  g22845(.A0(new_n23035_), .A1(\asqrt[4] ), .B0(new_n23037_), .Y(new_n23038_));
  NOR3X1   g22846(.A(new_n23032_), .B(new_n23024_), .C(\asqrt[17] ), .Y(new_n23039_));
  OAI21X1  g22847(.A0(new_n23039_), .A1(new_n23038_), .B0(new_n23033_), .Y(new_n23040_));
  AND2X1   g22848(.A(new_n23040_), .B(\asqrt[18] ), .Y(new_n23041_));
  INVX1    g22849(.A(new_n23038_), .Y(new_n23042_));
  AND2X1   g22850(.A(new_n23030_), .B(\asqrt[15] ), .Y(new_n23043_));
  OR2X1    g22851(.A(new_n23014_), .B(new_n23001_), .Y(new_n23044_));
  AND2X1   g22852(.A(new_n23021_), .B(new_n15362_), .Y(new_n23045_));
  AOI21X1  g22853(.A0(new_n23045_), .A1(new_n23044_), .B0(new_n23019_), .Y(new_n23046_));
  OAI21X1  g22854(.A0(new_n23046_), .A1(new_n23043_), .B0(\asqrt[16] ), .Y(new_n23047_));
  INVX1    g22855(.A(new_n23029_), .Y(new_n23048_));
  OAI21X1  g22856(.A0(new_n23004_), .A1(new_n15362_), .B0(new_n14754_), .Y(new_n23049_));
  OAI21X1  g22857(.A0(new_n23049_), .A1(new_n23046_), .B0(new_n23048_), .Y(new_n23050_));
  NAND3X1  g22858(.A(new_n23050_), .B(new_n23047_), .C(new_n14165_), .Y(new_n23051_));
  NAND2X1  g22859(.A(new_n23051_), .B(new_n23042_), .Y(new_n23052_));
  NAND4X1  g22860(.A(\asqrt[4] ), .B(new_n22300_), .C(new_n22287_), .D(new_n22283_), .Y(new_n23053_));
  NAND2X1  g22861(.A(new_n22300_), .B(new_n22283_), .Y(new_n23054_));
  OAI21X1  g22862(.A0(new_n23054_), .A1(new_n22874_), .B0(new_n22291_), .Y(new_n23055_));
  AND2X1   g22863(.A(new_n23055_), .B(new_n23053_), .Y(new_n23056_));
  AOI21X1  g22864(.A0(new_n23050_), .A1(new_n23047_), .B0(new_n14165_), .Y(new_n23057_));
  NOR2X1   g22865(.A(new_n23057_), .B(\asqrt[18] ), .Y(new_n23058_));
  AOI21X1  g22866(.A0(new_n23058_), .A1(new_n23052_), .B0(new_n23056_), .Y(new_n23059_));
  OAI21X1  g22867(.A0(new_n23059_), .A1(new_n23041_), .B0(\asqrt[19] ), .Y(new_n23060_));
  AND2X1   g22868(.A(new_n22308_), .B(new_n22301_), .Y(new_n23061_));
  NOR3X1   g22869(.A(new_n23061_), .B(new_n22346_), .C(new_n22290_), .Y(new_n23062_));
  NOR3X1   g22870(.A(new_n22874_), .B(new_n23061_), .C(new_n22290_), .Y(new_n23063_));
  NOR2X1   g22871(.A(new_n23063_), .B(new_n22306_), .Y(new_n23064_));
  AOI21X1  g22872(.A0(new_n23062_), .A1(\asqrt[4] ), .B0(new_n23064_), .Y(new_n23065_));
  INVX1    g22873(.A(new_n23065_), .Y(new_n23066_));
  AOI21X1  g22874(.A0(new_n23051_), .A1(new_n23042_), .B0(new_n23057_), .Y(new_n23067_));
  OAI21X1  g22875(.A0(new_n23067_), .A1(new_n13571_), .B0(new_n13000_), .Y(new_n23068_));
  OAI21X1  g22876(.A0(new_n23068_), .A1(new_n23059_), .B0(new_n23066_), .Y(new_n23069_));
  AOI21X1  g22877(.A0(new_n23069_), .A1(new_n23060_), .B0(new_n12447_), .Y(new_n23070_));
  AND2X1   g22878(.A(new_n22350_), .B(new_n22348_), .Y(new_n23071_));
  NOR3X1   g22879(.A(new_n23071_), .B(new_n22316_), .C(new_n22349_), .Y(new_n23072_));
  NOR3X1   g22880(.A(new_n22874_), .B(new_n23071_), .C(new_n22349_), .Y(new_n23073_));
  NOR2X1   g22881(.A(new_n23073_), .B(new_n22315_), .Y(new_n23074_));
  AOI21X1  g22882(.A0(new_n23072_), .A1(\asqrt[4] ), .B0(new_n23074_), .Y(new_n23075_));
  INVX1    g22883(.A(new_n23075_), .Y(new_n23076_));
  NAND3X1  g22884(.A(new_n23069_), .B(new_n23060_), .C(new_n12447_), .Y(new_n23077_));
  AOI21X1  g22885(.A0(new_n23077_), .A1(new_n23076_), .B0(new_n23070_), .Y(new_n23078_));
  OR2X1    g22886(.A(new_n23078_), .B(new_n11896_), .Y(new_n23079_));
  AND2X1   g22887(.A(new_n23077_), .B(new_n23076_), .Y(new_n23080_));
  NAND4X1  g22888(.A(\asqrt[4] ), .B(new_n22326_), .C(new_n22324_), .D(new_n22352_), .Y(new_n23081_));
  NAND2X1  g22889(.A(new_n22326_), .B(new_n22352_), .Y(new_n23082_));
  OAI21X1  g22890(.A0(new_n23082_), .A1(new_n22874_), .B0(new_n22325_), .Y(new_n23083_));
  AND2X1   g22891(.A(new_n23083_), .B(new_n23081_), .Y(new_n23084_));
  INVX1    g22892(.A(new_n23084_), .Y(new_n23085_));
  OR2X1    g22893(.A(new_n23070_), .B(\asqrt[21] ), .Y(new_n23086_));
  OAI21X1  g22894(.A0(new_n23086_), .A1(new_n23080_), .B0(new_n23085_), .Y(new_n23087_));
  AOI21X1  g22895(.A0(new_n23087_), .A1(new_n23079_), .B0(new_n11362_), .Y(new_n23088_));
  AOI21X1  g22896(.A0(new_n22368_), .A1(new_n22367_), .B0(new_n22335_), .Y(new_n23089_));
  AND2X1   g22897(.A(new_n23089_), .B(new_n22328_), .Y(new_n23090_));
  AOI22X1  g22898(.A0(new_n22368_), .A1(new_n22367_), .B0(new_n22354_), .B1(\asqrt[21] ), .Y(new_n23091_));
  AOI21X1  g22899(.A0(new_n23091_), .A1(\asqrt[4] ), .B0(new_n22334_), .Y(new_n23092_));
  AOI21X1  g22900(.A0(new_n23090_), .A1(\asqrt[4] ), .B0(new_n23092_), .Y(new_n23093_));
  OR2X1    g22901(.A(new_n23067_), .B(new_n13571_), .Y(new_n23094_));
  AND2X1   g22902(.A(new_n23051_), .B(new_n23042_), .Y(new_n23095_));
  INVX1    g22903(.A(new_n23056_), .Y(new_n23096_));
  OR2X1    g22904(.A(new_n23057_), .B(\asqrt[18] ), .Y(new_n23097_));
  OAI21X1  g22905(.A0(new_n23097_), .A1(new_n23095_), .B0(new_n23096_), .Y(new_n23098_));
  AOI21X1  g22906(.A0(new_n23098_), .A1(new_n23094_), .B0(new_n13000_), .Y(new_n23099_));
  AOI21X1  g22907(.A0(new_n23040_), .A1(\asqrt[18] ), .B0(\asqrt[19] ), .Y(new_n23100_));
  AOI21X1  g22908(.A0(new_n23100_), .A1(new_n23098_), .B0(new_n23065_), .Y(new_n23101_));
  OAI21X1  g22909(.A0(new_n23101_), .A1(new_n23099_), .B0(\asqrt[20] ), .Y(new_n23102_));
  NOR3X1   g22910(.A(new_n23101_), .B(new_n23099_), .C(\asqrt[20] ), .Y(new_n23103_));
  OAI21X1  g22911(.A0(new_n23103_), .A1(new_n23075_), .B0(new_n23102_), .Y(new_n23104_));
  AOI21X1  g22912(.A0(new_n23104_), .A1(\asqrt[21] ), .B0(\asqrt[22] ), .Y(new_n23105_));
  AOI21X1  g22913(.A0(new_n23105_), .A1(new_n23087_), .B0(new_n23093_), .Y(new_n23106_));
  OAI21X1  g22914(.A0(new_n23106_), .A1(new_n23088_), .B0(\asqrt[23] ), .Y(new_n23107_));
  AND2X1   g22915(.A(new_n22355_), .B(new_n22337_), .Y(new_n23108_));
  NOR3X1   g22916(.A(new_n23108_), .B(new_n22371_), .C(new_n22338_), .Y(new_n23109_));
  NOR3X1   g22917(.A(new_n22874_), .B(new_n23108_), .C(new_n22338_), .Y(new_n23110_));
  NOR2X1   g22918(.A(new_n23110_), .B(new_n22343_), .Y(new_n23111_));
  AOI21X1  g22919(.A0(new_n23109_), .A1(\asqrt[4] ), .B0(new_n23111_), .Y(new_n23112_));
  NOR3X1   g22920(.A(new_n23106_), .B(new_n23088_), .C(\asqrt[23] ), .Y(new_n23113_));
  OAI21X1  g22921(.A0(new_n23113_), .A1(new_n23112_), .B0(new_n23107_), .Y(new_n23114_));
  AND2X1   g22922(.A(new_n23114_), .B(\asqrt[24] ), .Y(new_n23115_));
  INVX1    g22923(.A(new_n23112_), .Y(new_n23116_));
  AND2X1   g22924(.A(new_n23104_), .B(\asqrt[21] ), .Y(new_n23117_));
  NAND2X1  g22925(.A(new_n23077_), .B(new_n23076_), .Y(new_n23118_));
  NOR2X1   g22926(.A(new_n23070_), .B(\asqrt[21] ), .Y(new_n23119_));
  AOI21X1  g22927(.A0(new_n23119_), .A1(new_n23118_), .B0(new_n23084_), .Y(new_n23120_));
  OAI21X1  g22928(.A0(new_n23120_), .A1(new_n23117_), .B0(\asqrt[22] ), .Y(new_n23121_));
  INVX1    g22929(.A(new_n23093_), .Y(new_n23122_));
  OAI21X1  g22930(.A0(new_n23078_), .A1(new_n11896_), .B0(new_n11362_), .Y(new_n23123_));
  OAI21X1  g22931(.A0(new_n23123_), .A1(new_n23120_), .B0(new_n23122_), .Y(new_n23124_));
  NAND3X1  g22932(.A(new_n23124_), .B(new_n23121_), .C(new_n10849_), .Y(new_n23125_));
  NAND2X1  g22933(.A(new_n23125_), .B(new_n23116_), .Y(new_n23126_));
  NAND4X1  g22934(.A(\asqrt[4] ), .B(new_n22374_), .C(new_n22361_), .D(new_n22357_), .Y(new_n23127_));
  NAND2X1  g22935(.A(new_n22374_), .B(new_n22357_), .Y(new_n23128_));
  OAI21X1  g22936(.A0(new_n23128_), .A1(new_n22874_), .B0(new_n22365_), .Y(new_n23129_));
  AND2X1   g22937(.A(new_n23129_), .B(new_n23127_), .Y(new_n23130_));
  AOI21X1  g22938(.A0(new_n23124_), .A1(new_n23121_), .B0(new_n10849_), .Y(new_n23131_));
  NOR2X1   g22939(.A(new_n23131_), .B(\asqrt[24] ), .Y(new_n23132_));
  AOI21X1  g22940(.A0(new_n23132_), .A1(new_n23126_), .B0(new_n23130_), .Y(new_n23133_));
  OAI21X1  g22941(.A0(new_n23133_), .A1(new_n23115_), .B0(\asqrt[25] ), .Y(new_n23134_));
  AND2X1   g22942(.A(new_n22382_), .B(new_n22375_), .Y(new_n23135_));
  NOR3X1   g22943(.A(new_n23135_), .B(new_n22418_), .C(new_n22364_), .Y(new_n23136_));
  NOR3X1   g22944(.A(new_n22874_), .B(new_n23135_), .C(new_n22364_), .Y(new_n23137_));
  NOR2X1   g22945(.A(new_n23137_), .B(new_n22380_), .Y(new_n23138_));
  AOI21X1  g22946(.A0(new_n23136_), .A1(\asqrt[4] ), .B0(new_n23138_), .Y(new_n23139_));
  INVX1    g22947(.A(new_n23139_), .Y(new_n23140_));
  AOI21X1  g22948(.A0(new_n23125_), .A1(new_n23116_), .B0(new_n23131_), .Y(new_n23141_));
  OAI21X1  g22949(.A0(new_n23141_), .A1(new_n10332_), .B0(new_n9833_), .Y(new_n23142_));
  OAI21X1  g22950(.A0(new_n23142_), .A1(new_n23133_), .B0(new_n23140_), .Y(new_n23143_));
  AOI21X1  g22951(.A0(new_n23143_), .A1(new_n23134_), .B0(new_n9353_), .Y(new_n23144_));
  AND2X1   g22952(.A(new_n22422_), .B(new_n22420_), .Y(new_n23145_));
  NOR3X1   g22953(.A(new_n23145_), .B(new_n22390_), .C(new_n22421_), .Y(new_n23146_));
  NOR3X1   g22954(.A(new_n22874_), .B(new_n23145_), .C(new_n22421_), .Y(new_n23147_));
  NOR2X1   g22955(.A(new_n23147_), .B(new_n22389_), .Y(new_n23148_));
  AOI21X1  g22956(.A0(new_n23146_), .A1(\asqrt[4] ), .B0(new_n23148_), .Y(new_n23149_));
  INVX1    g22957(.A(new_n23149_), .Y(new_n23150_));
  NAND3X1  g22958(.A(new_n23143_), .B(new_n23134_), .C(new_n9353_), .Y(new_n23151_));
  AOI21X1  g22959(.A0(new_n23151_), .A1(new_n23150_), .B0(new_n23144_), .Y(new_n23152_));
  OR2X1    g22960(.A(new_n23152_), .B(new_n8874_), .Y(new_n23153_));
  AND2X1   g22961(.A(new_n23151_), .B(new_n23150_), .Y(new_n23154_));
  OR4X1    g22962(.A(new_n22874_), .B(new_n22426_), .C(new_n22397_), .D(new_n22394_), .Y(new_n23155_));
  NAND2X1  g22963(.A(new_n22398_), .B(new_n22424_), .Y(new_n23156_));
  OAI21X1  g22964(.A0(new_n23156_), .A1(new_n22874_), .B0(new_n22397_), .Y(new_n23157_));
  AND2X1   g22965(.A(new_n23157_), .B(new_n23155_), .Y(new_n23158_));
  INVX1    g22966(.A(new_n23158_), .Y(new_n23159_));
  OR2X1    g22967(.A(new_n23144_), .B(\asqrt[27] ), .Y(new_n23160_));
  OAI21X1  g22968(.A0(new_n23160_), .A1(new_n23154_), .B0(new_n23159_), .Y(new_n23161_));
  AOI21X1  g22969(.A0(new_n23161_), .A1(new_n23153_), .B0(new_n8412_), .Y(new_n23162_));
  AOI21X1  g22970(.A0(new_n22441_), .A1(new_n22440_), .B0(new_n22407_), .Y(new_n23163_));
  AND2X1   g22971(.A(new_n23163_), .B(new_n22400_), .Y(new_n23164_));
  AOI22X1  g22972(.A0(new_n22441_), .A1(new_n22440_), .B0(new_n22427_), .B1(\asqrt[27] ), .Y(new_n23165_));
  AOI21X1  g22973(.A0(new_n23165_), .A1(\asqrt[4] ), .B0(new_n22406_), .Y(new_n23166_));
  AOI21X1  g22974(.A0(new_n23164_), .A1(\asqrt[4] ), .B0(new_n23166_), .Y(new_n23167_));
  OR2X1    g22975(.A(new_n23141_), .B(new_n10332_), .Y(new_n23168_));
  AND2X1   g22976(.A(new_n23125_), .B(new_n23116_), .Y(new_n23169_));
  INVX1    g22977(.A(new_n23130_), .Y(new_n23170_));
  OR2X1    g22978(.A(new_n23131_), .B(\asqrt[24] ), .Y(new_n23171_));
  OAI21X1  g22979(.A0(new_n23171_), .A1(new_n23169_), .B0(new_n23170_), .Y(new_n23172_));
  AOI21X1  g22980(.A0(new_n23172_), .A1(new_n23168_), .B0(new_n9833_), .Y(new_n23173_));
  AOI21X1  g22981(.A0(new_n23114_), .A1(\asqrt[24] ), .B0(\asqrt[25] ), .Y(new_n23174_));
  AOI21X1  g22982(.A0(new_n23174_), .A1(new_n23172_), .B0(new_n23139_), .Y(new_n23175_));
  OAI21X1  g22983(.A0(new_n23175_), .A1(new_n23173_), .B0(\asqrt[26] ), .Y(new_n23176_));
  NOR3X1   g22984(.A(new_n23175_), .B(new_n23173_), .C(\asqrt[26] ), .Y(new_n23177_));
  OAI21X1  g22985(.A0(new_n23177_), .A1(new_n23149_), .B0(new_n23176_), .Y(new_n23178_));
  AOI21X1  g22986(.A0(new_n23178_), .A1(\asqrt[27] ), .B0(\asqrt[28] ), .Y(new_n23179_));
  AOI21X1  g22987(.A0(new_n23179_), .A1(new_n23161_), .B0(new_n23167_), .Y(new_n23180_));
  OAI21X1  g22988(.A0(new_n23180_), .A1(new_n23162_), .B0(\asqrt[29] ), .Y(new_n23181_));
  AND2X1   g22989(.A(new_n22428_), .B(new_n22409_), .Y(new_n23182_));
  NOR3X1   g22990(.A(new_n23182_), .B(new_n22444_), .C(new_n22410_), .Y(new_n23183_));
  NOR3X1   g22991(.A(new_n22874_), .B(new_n23182_), .C(new_n22410_), .Y(new_n23184_));
  NOR2X1   g22992(.A(new_n23184_), .B(new_n22415_), .Y(new_n23185_));
  AOI21X1  g22993(.A0(new_n23183_), .A1(\asqrt[4] ), .B0(new_n23185_), .Y(new_n23186_));
  NOR3X1   g22994(.A(new_n23180_), .B(new_n23162_), .C(\asqrt[29] ), .Y(new_n23187_));
  OAI21X1  g22995(.A0(new_n23187_), .A1(new_n23186_), .B0(new_n23181_), .Y(new_n23188_));
  AND2X1   g22996(.A(new_n23188_), .B(\asqrt[30] ), .Y(new_n23189_));
  INVX1    g22997(.A(new_n23186_), .Y(new_n23190_));
  AND2X1   g22998(.A(new_n23178_), .B(\asqrt[27] ), .Y(new_n23191_));
  NAND2X1  g22999(.A(new_n23151_), .B(new_n23150_), .Y(new_n23192_));
  NOR2X1   g23000(.A(new_n23144_), .B(\asqrt[27] ), .Y(new_n23193_));
  AOI21X1  g23001(.A0(new_n23193_), .A1(new_n23192_), .B0(new_n23158_), .Y(new_n23194_));
  OAI21X1  g23002(.A0(new_n23194_), .A1(new_n23191_), .B0(\asqrt[28] ), .Y(new_n23195_));
  INVX1    g23003(.A(new_n23167_), .Y(new_n23196_));
  OAI21X1  g23004(.A0(new_n23152_), .A1(new_n8874_), .B0(new_n8412_), .Y(new_n23197_));
  OAI21X1  g23005(.A0(new_n23197_), .A1(new_n23194_), .B0(new_n23196_), .Y(new_n23198_));
  NAND3X1  g23006(.A(new_n23198_), .B(new_n23195_), .C(new_n7970_), .Y(new_n23199_));
  NAND2X1  g23007(.A(new_n23199_), .B(new_n23190_), .Y(new_n23200_));
  NAND4X1  g23008(.A(\asqrt[4] ), .B(new_n22447_), .C(new_n22434_), .D(new_n22430_), .Y(new_n23201_));
  NAND2X1  g23009(.A(new_n22447_), .B(new_n22430_), .Y(new_n23202_));
  OAI21X1  g23010(.A0(new_n23202_), .A1(new_n22874_), .B0(new_n22438_), .Y(new_n23203_));
  AND2X1   g23011(.A(new_n23203_), .B(new_n23201_), .Y(new_n23204_));
  AOI21X1  g23012(.A0(new_n23198_), .A1(new_n23195_), .B0(new_n7970_), .Y(new_n23205_));
  NOR2X1   g23013(.A(new_n23205_), .B(\asqrt[30] ), .Y(new_n23206_));
  AOI21X1  g23014(.A0(new_n23206_), .A1(new_n23200_), .B0(new_n23204_), .Y(new_n23207_));
  OAI21X1  g23015(.A0(new_n23207_), .A1(new_n23189_), .B0(\asqrt[31] ), .Y(new_n23208_));
  AND2X1   g23016(.A(new_n22455_), .B(new_n22448_), .Y(new_n23209_));
  NOR3X1   g23017(.A(new_n23209_), .B(new_n22493_), .C(new_n22437_), .Y(new_n23210_));
  NOR3X1   g23018(.A(new_n22874_), .B(new_n23209_), .C(new_n22437_), .Y(new_n23211_));
  NOR2X1   g23019(.A(new_n23211_), .B(new_n22453_), .Y(new_n23212_));
  AOI21X1  g23020(.A0(new_n23210_), .A1(\asqrt[4] ), .B0(new_n23212_), .Y(new_n23213_));
  INVX1    g23021(.A(new_n23213_), .Y(new_n23214_));
  AOI21X1  g23022(.A0(new_n23199_), .A1(new_n23190_), .B0(new_n23205_), .Y(new_n23215_));
  OAI21X1  g23023(.A0(new_n23215_), .A1(new_n7527_), .B0(new_n7103_), .Y(new_n23216_));
  OAI21X1  g23024(.A0(new_n23216_), .A1(new_n23207_), .B0(new_n23214_), .Y(new_n23217_));
  AOI21X1  g23025(.A0(new_n23217_), .A1(new_n23208_), .B0(new_n6699_), .Y(new_n23218_));
  AND2X1   g23026(.A(new_n22497_), .B(new_n22495_), .Y(new_n23219_));
  NOR3X1   g23027(.A(new_n23219_), .B(new_n22463_), .C(new_n22496_), .Y(new_n23220_));
  NOR3X1   g23028(.A(new_n22874_), .B(new_n23219_), .C(new_n22496_), .Y(new_n23221_));
  NOR2X1   g23029(.A(new_n23221_), .B(new_n22462_), .Y(new_n23222_));
  AOI21X1  g23030(.A0(new_n23220_), .A1(\asqrt[4] ), .B0(new_n23222_), .Y(new_n23223_));
  INVX1    g23031(.A(new_n23223_), .Y(new_n23224_));
  NAND3X1  g23032(.A(new_n23217_), .B(new_n23208_), .C(new_n6699_), .Y(new_n23225_));
  AOI21X1  g23033(.A0(new_n23225_), .A1(new_n23224_), .B0(new_n23218_), .Y(new_n23226_));
  OR2X1    g23034(.A(new_n23226_), .B(new_n6294_), .Y(new_n23227_));
  AND2X1   g23035(.A(new_n23225_), .B(new_n23224_), .Y(new_n23228_));
  OR4X1    g23036(.A(new_n22874_), .B(new_n22500_), .C(new_n22472_), .D(new_n22467_), .Y(new_n23229_));
  NAND2X1  g23037(.A(new_n22473_), .B(new_n22499_), .Y(new_n23230_));
  OAI21X1  g23038(.A0(new_n23230_), .A1(new_n22874_), .B0(new_n22472_), .Y(new_n23231_));
  AND2X1   g23039(.A(new_n23231_), .B(new_n23229_), .Y(new_n23232_));
  INVX1    g23040(.A(new_n23232_), .Y(new_n23233_));
  OR2X1    g23041(.A(new_n23218_), .B(\asqrt[33] ), .Y(new_n23234_));
  OAI21X1  g23042(.A0(new_n23234_), .A1(new_n23228_), .B0(new_n23233_), .Y(new_n23235_));
  AOI21X1  g23043(.A0(new_n23235_), .A1(new_n23227_), .B0(new_n5941_), .Y(new_n23236_));
  AOI21X1  g23044(.A0(new_n22529_), .A1(new_n22528_), .B0(new_n22482_), .Y(new_n23237_));
  AND2X1   g23045(.A(new_n23237_), .B(new_n22475_), .Y(new_n23238_));
  AOI22X1  g23046(.A0(new_n22529_), .A1(new_n22528_), .B0(new_n22501_), .B1(\asqrt[33] ), .Y(new_n23239_));
  AOI21X1  g23047(.A0(new_n23239_), .A1(\asqrt[4] ), .B0(new_n22481_), .Y(new_n23240_));
  AOI21X1  g23048(.A0(new_n23238_), .A1(\asqrt[4] ), .B0(new_n23240_), .Y(new_n23241_));
  OR2X1    g23049(.A(new_n23215_), .B(new_n7527_), .Y(new_n23242_));
  AND2X1   g23050(.A(new_n23199_), .B(new_n23190_), .Y(new_n23243_));
  INVX1    g23051(.A(new_n23204_), .Y(new_n23244_));
  OR2X1    g23052(.A(new_n23205_), .B(\asqrt[30] ), .Y(new_n23245_));
  OAI21X1  g23053(.A0(new_n23245_), .A1(new_n23243_), .B0(new_n23244_), .Y(new_n23246_));
  AOI21X1  g23054(.A0(new_n23246_), .A1(new_n23242_), .B0(new_n7103_), .Y(new_n23247_));
  AOI21X1  g23055(.A0(new_n23188_), .A1(\asqrt[30] ), .B0(\asqrt[31] ), .Y(new_n23248_));
  AOI21X1  g23056(.A0(new_n23248_), .A1(new_n23246_), .B0(new_n23213_), .Y(new_n23249_));
  OAI21X1  g23057(.A0(new_n23249_), .A1(new_n23247_), .B0(\asqrt[32] ), .Y(new_n23250_));
  NOR3X1   g23058(.A(new_n23249_), .B(new_n23247_), .C(\asqrt[32] ), .Y(new_n23251_));
  OAI21X1  g23059(.A0(new_n23251_), .A1(new_n23223_), .B0(new_n23250_), .Y(new_n23252_));
  AOI21X1  g23060(.A0(new_n23252_), .A1(\asqrt[33] ), .B0(\asqrt[34] ), .Y(new_n23253_));
  AOI21X1  g23061(.A0(new_n23253_), .A1(new_n23235_), .B0(new_n23241_), .Y(new_n23254_));
  OAI21X1  g23062(.A0(new_n23254_), .A1(new_n23236_), .B0(\asqrt[35] ), .Y(new_n23255_));
  AND2X1   g23063(.A(new_n22502_), .B(new_n22484_), .Y(new_n23256_));
  NOR3X1   g23064(.A(new_n23256_), .B(new_n22532_), .C(new_n22485_), .Y(new_n23257_));
  NOR3X1   g23065(.A(new_n22874_), .B(new_n23256_), .C(new_n22485_), .Y(new_n23258_));
  NOR2X1   g23066(.A(new_n23258_), .B(new_n22490_), .Y(new_n23259_));
  AOI21X1  g23067(.A0(new_n23257_), .A1(\asqrt[4] ), .B0(new_n23259_), .Y(new_n23260_));
  NOR3X1   g23068(.A(new_n23254_), .B(new_n23236_), .C(\asqrt[35] ), .Y(new_n23261_));
  OAI21X1  g23069(.A0(new_n23261_), .A1(new_n23260_), .B0(new_n23255_), .Y(new_n23262_));
  AND2X1   g23070(.A(new_n23262_), .B(\asqrt[36] ), .Y(new_n23263_));
  OR2X1    g23071(.A(new_n23261_), .B(new_n23260_), .Y(new_n23264_));
  OR4X1    g23072(.A(new_n22874_), .B(new_n22509_), .C(new_n22536_), .D(new_n22535_), .Y(new_n23265_));
  OR2X1    g23073(.A(new_n22509_), .B(new_n22535_), .Y(new_n23266_));
  OAI21X1  g23074(.A0(new_n23266_), .A1(new_n22874_), .B0(new_n22536_), .Y(new_n23267_));
  AND2X1   g23075(.A(new_n23267_), .B(new_n23265_), .Y(new_n23268_));
  AND2X1   g23076(.A(new_n23255_), .B(new_n5176_), .Y(new_n23269_));
  AOI21X1  g23077(.A0(new_n23269_), .A1(new_n23264_), .B0(new_n23268_), .Y(new_n23270_));
  OAI21X1  g23078(.A0(new_n23270_), .A1(new_n23263_), .B0(\asqrt[37] ), .Y(new_n23271_));
  AND2X1   g23079(.A(new_n22518_), .B(new_n22512_), .Y(new_n23272_));
  NOR3X1   g23080(.A(new_n23272_), .B(new_n22552_), .C(new_n22511_), .Y(new_n23273_));
  NOR3X1   g23081(.A(new_n22874_), .B(new_n23272_), .C(new_n22511_), .Y(new_n23274_));
  NOR2X1   g23082(.A(new_n23274_), .B(new_n22517_), .Y(new_n23275_));
  AOI21X1  g23083(.A0(new_n23273_), .A1(\asqrt[4] ), .B0(new_n23275_), .Y(new_n23276_));
  INVX1    g23084(.A(new_n23276_), .Y(new_n23277_));
  AND2X1   g23085(.A(new_n23252_), .B(\asqrt[33] ), .Y(new_n23278_));
  NAND2X1  g23086(.A(new_n23225_), .B(new_n23224_), .Y(new_n23279_));
  NOR2X1   g23087(.A(new_n23218_), .B(\asqrt[33] ), .Y(new_n23280_));
  AOI21X1  g23088(.A0(new_n23280_), .A1(new_n23279_), .B0(new_n23232_), .Y(new_n23281_));
  OAI21X1  g23089(.A0(new_n23281_), .A1(new_n23278_), .B0(\asqrt[34] ), .Y(new_n23282_));
  INVX1    g23090(.A(new_n23241_), .Y(new_n23283_));
  OAI21X1  g23091(.A0(new_n23226_), .A1(new_n6294_), .B0(new_n5941_), .Y(new_n23284_));
  OAI21X1  g23092(.A0(new_n23284_), .A1(new_n23281_), .B0(new_n23283_), .Y(new_n23285_));
  AOI21X1  g23093(.A0(new_n23285_), .A1(new_n23282_), .B0(new_n5541_), .Y(new_n23286_));
  INVX1    g23094(.A(new_n23260_), .Y(new_n23287_));
  NAND3X1  g23095(.A(new_n23285_), .B(new_n23282_), .C(new_n5541_), .Y(new_n23288_));
  AOI21X1  g23096(.A0(new_n23288_), .A1(new_n23287_), .B0(new_n23286_), .Y(new_n23289_));
  OAI21X1  g23097(.A0(new_n23289_), .A1(new_n5176_), .B0(new_n4826_), .Y(new_n23290_));
  OAI21X1  g23098(.A0(new_n23290_), .A1(new_n23270_), .B0(new_n23277_), .Y(new_n23291_));
  AOI21X1  g23099(.A0(new_n23291_), .A1(new_n23271_), .B0(new_n4493_), .Y(new_n23292_));
  AND2X1   g23100(.A(new_n22556_), .B(new_n22554_), .Y(new_n23293_));
  NOR3X1   g23101(.A(new_n23293_), .B(new_n22526_), .C(new_n22555_), .Y(new_n23294_));
  NOR3X1   g23102(.A(new_n22874_), .B(new_n23293_), .C(new_n22555_), .Y(new_n23295_));
  NOR2X1   g23103(.A(new_n23295_), .B(new_n22525_), .Y(new_n23296_));
  AOI21X1  g23104(.A0(new_n23294_), .A1(\asqrt[4] ), .B0(new_n23296_), .Y(new_n23297_));
  INVX1    g23105(.A(new_n23297_), .Y(new_n23298_));
  NAND3X1  g23106(.A(new_n23291_), .B(new_n23271_), .C(new_n4493_), .Y(new_n23299_));
  AOI21X1  g23107(.A0(new_n23299_), .A1(new_n23298_), .B0(new_n23292_), .Y(new_n23300_));
  OR2X1    g23108(.A(new_n23300_), .B(new_n4165_), .Y(new_n23301_));
  OR2X1    g23109(.A(new_n23289_), .B(new_n5176_), .Y(new_n23302_));
  NOR2X1   g23110(.A(new_n23261_), .B(new_n23260_), .Y(new_n23303_));
  INVX1    g23111(.A(new_n23268_), .Y(new_n23304_));
  NAND2X1  g23112(.A(new_n23255_), .B(new_n5176_), .Y(new_n23305_));
  OAI21X1  g23113(.A0(new_n23305_), .A1(new_n23303_), .B0(new_n23304_), .Y(new_n23306_));
  AOI21X1  g23114(.A0(new_n23306_), .A1(new_n23302_), .B0(new_n4826_), .Y(new_n23307_));
  AOI21X1  g23115(.A0(new_n23262_), .A1(\asqrt[36] ), .B0(\asqrt[37] ), .Y(new_n23308_));
  AOI21X1  g23116(.A0(new_n23308_), .A1(new_n23306_), .B0(new_n23276_), .Y(new_n23309_));
  NOR3X1   g23117(.A(new_n23309_), .B(new_n23307_), .C(\asqrt[38] ), .Y(new_n23310_));
  NOR2X1   g23118(.A(new_n23310_), .B(new_n23297_), .Y(new_n23311_));
  OR4X1    g23119(.A(new_n22874_), .B(new_n22558_), .C(new_n22546_), .D(new_n22541_), .Y(new_n23312_));
  OR2X1    g23120(.A(new_n22558_), .B(new_n22541_), .Y(new_n23313_));
  OAI21X1  g23121(.A0(new_n23313_), .A1(new_n22874_), .B0(new_n22546_), .Y(new_n23314_));
  AND2X1   g23122(.A(new_n23314_), .B(new_n23312_), .Y(new_n23315_));
  INVX1    g23123(.A(new_n23315_), .Y(new_n23316_));
  OAI21X1  g23124(.A0(new_n23309_), .A1(new_n23307_), .B0(\asqrt[38] ), .Y(new_n23317_));
  NAND2X1  g23125(.A(new_n23317_), .B(new_n4165_), .Y(new_n23318_));
  OAI21X1  g23126(.A0(new_n23318_), .A1(new_n23311_), .B0(new_n23316_), .Y(new_n23319_));
  AOI21X1  g23127(.A0(new_n23319_), .A1(new_n23301_), .B0(new_n3863_), .Y(new_n23320_));
  AOI21X1  g23128(.A0(new_n22603_), .A1(new_n22602_), .B0(new_n22565_), .Y(new_n23321_));
  AND2X1   g23129(.A(new_n23321_), .B(new_n22549_), .Y(new_n23322_));
  AOI22X1  g23130(.A0(new_n22603_), .A1(new_n22602_), .B0(new_n22575_), .B1(\asqrt[39] ), .Y(new_n23323_));
  AOI21X1  g23131(.A0(new_n23323_), .A1(\asqrt[4] ), .B0(new_n22564_), .Y(new_n23324_));
  AOI21X1  g23132(.A0(new_n23322_), .A1(\asqrt[4] ), .B0(new_n23324_), .Y(new_n23325_));
  OAI21X1  g23133(.A0(new_n23310_), .A1(new_n23297_), .B0(new_n23317_), .Y(new_n23326_));
  AOI21X1  g23134(.A0(new_n23326_), .A1(\asqrt[39] ), .B0(\asqrt[40] ), .Y(new_n23327_));
  AOI21X1  g23135(.A0(new_n23327_), .A1(new_n23319_), .B0(new_n23325_), .Y(new_n23328_));
  OAI21X1  g23136(.A0(new_n23328_), .A1(new_n23320_), .B0(\asqrt[41] ), .Y(new_n23329_));
  AND2X1   g23137(.A(new_n22576_), .B(new_n22568_), .Y(new_n23330_));
  NOR3X1   g23138(.A(new_n23330_), .B(new_n22606_), .C(new_n22569_), .Y(new_n23331_));
  NOR3X1   g23139(.A(new_n22874_), .B(new_n23330_), .C(new_n22569_), .Y(new_n23332_));
  NOR2X1   g23140(.A(new_n23332_), .B(new_n22574_), .Y(new_n23333_));
  AOI21X1  g23141(.A0(new_n23331_), .A1(\asqrt[4] ), .B0(new_n23333_), .Y(new_n23334_));
  NOR3X1   g23142(.A(new_n23328_), .B(new_n23320_), .C(\asqrt[41] ), .Y(new_n23335_));
  OAI21X1  g23143(.A0(new_n23335_), .A1(new_n23334_), .B0(new_n23329_), .Y(new_n23336_));
  AND2X1   g23144(.A(new_n23336_), .B(\asqrt[42] ), .Y(new_n23337_));
  OR2X1    g23145(.A(new_n23335_), .B(new_n23334_), .Y(new_n23338_));
  OR4X1    g23146(.A(new_n22874_), .B(new_n22583_), .C(new_n22610_), .D(new_n22609_), .Y(new_n23339_));
  OR2X1    g23147(.A(new_n22583_), .B(new_n22609_), .Y(new_n23340_));
  OAI21X1  g23148(.A0(new_n23340_), .A1(new_n22874_), .B0(new_n22610_), .Y(new_n23341_));
  AND2X1   g23149(.A(new_n23341_), .B(new_n23339_), .Y(new_n23342_));
  AND2X1   g23150(.A(new_n23329_), .B(new_n3276_), .Y(new_n23343_));
  AOI21X1  g23151(.A0(new_n23343_), .A1(new_n23338_), .B0(new_n23342_), .Y(new_n23344_));
  OAI21X1  g23152(.A0(new_n23344_), .A1(new_n23337_), .B0(\asqrt[43] ), .Y(new_n23345_));
  AND2X1   g23153(.A(new_n22592_), .B(new_n22586_), .Y(new_n23346_));
  NOR3X1   g23154(.A(new_n23346_), .B(new_n22626_), .C(new_n22585_), .Y(new_n23347_));
  NOR3X1   g23155(.A(new_n22874_), .B(new_n23346_), .C(new_n22585_), .Y(new_n23348_));
  NOR2X1   g23156(.A(new_n23348_), .B(new_n22591_), .Y(new_n23349_));
  AOI21X1  g23157(.A0(new_n23347_), .A1(\asqrt[4] ), .B0(new_n23349_), .Y(new_n23350_));
  INVX1    g23158(.A(new_n23350_), .Y(new_n23351_));
  AND2X1   g23159(.A(new_n23326_), .B(\asqrt[39] ), .Y(new_n23352_));
  OR2X1    g23160(.A(new_n23310_), .B(new_n23297_), .Y(new_n23353_));
  AND2X1   g23161(.A(new_n23317_), .B(new_n4165_), .Y(new_n23354_));
  AOI21X1  g23162(.A0(new_n23354_), .A1(new_n23353_), .B0(new_n23315_), .Y(new_n23355_));
  OAI21X1  g23163(.A0(new_n23355_), .A1(new_n23352_), .B0(\asqrt[40] ), .Y(new_n23356_));
  INVX1    g23164(.A(new_n23325_), .Y(new_n23357_));
  OAI21X1  g23165(.A0(new_n23300_), .A1(new_n4165_), .B0(new_n3863_), .Y(new_n23358_));
  OAI21X1  g23166(.A0(new_n23358_), .A1(new_n23355_), .B0(new_n23357_), .Y(new_n23359_));
  AOI21X1  g23167(.A0(new_n23359_), .A1(new_n23356_), .B0(new_n3564_), .Y(new_n23360_));
  INVX1    g23168(.A(new_n23334_), .Y(new_n23361_));
  NAND3X1  g23169(.A(new_n23359_), .B(new_n23356_), .C(new_n3564_), .Y(new_n23362_));
  AOI21X1  g23170(.A0(new_n23362_), .A1(new_n23361_), .B0(new_n23360_), .Y(new_n23363_));
  OAI21X1  g23171(.A0(new_n23363_), .A1(new_n3276_), .B0(new_n3008_), .Y(new_n23364_));
  OAI21X1  g23172(.A0(new_n23364_), .A1(new_n23344_), .B0(new_n23351_), .Y(new_n23365_));
  AOI21X1  g23173(.A0(new_n23365_), .A1(new_n23345_), .B0(new_n2769_), .Y(new_n23366_));
  AND2X1   g23174(.A(new_n22630_), .B(new_n22628_), .Y(new_n23367_));
  NOR3X1   g23175(.A(new_n23367_), .B(new_n22600_), .C(new_n22629_), .Y(new_n23368_));
  NOR3X1   g23176(.A(new_n22874_), .B(new_n23367_), .C(new_n22629_), .Y(new_n23369_));
  NOR2X1   g23177(.A(new_n23369_), .B(new_n22599_), .Y(new_n23370_));
  AOI21X1  g23178(.A0(new_n23368_), .A1(\asqrt[4] ), .B0(new_n23370_), .Y(new_n23371_));
  INVX1    g23179(.A(new_n23371_), .Y(new_n23372_));
  NAND3X1  g23180(.A(new_n23365_), .B(new_n23345_), .C(new_n2769_), .Y(new_n23373_));
  AOI21X1  g23181(.A0(new_n23373_), .A1(new_n23372_), .B0(new_n23366_), .Y(new_n23374_));
  OR2X1    g23182(.A(new_n23374_), .B(new_n2570_), .Y(new_n23375_));
  OR2X1    g23183(.A(new_n23363_), .B(new_n3276_), .Y(new_n23376_));
  NOR2X1   g23184(.A(new_n23335_), .B(new_n23334_), .Y(new_n23377_));
  INVX1    g23185(.A(new_n23342_), .Y(new_n23378_));
  NAND2X1  g23186(.A(new_n23329_), .B(new_n3276_), .Y(new_n23379_));
  OAI21X1  g23187(.A0(new_n23379_), .A1(new_n23377_), .B0(new_n23378_), .Y(new_n23380_));
  AOI21X1  g23188(.A0(new_n23380_), .A1(new_n23376_), .B0(new_n3008_), .Y(new_n23381_));
  AOI21X1  g23189(.A0(new_n23336_), .A1(\asqrt[42] ), .B0(\asqrt[43] ), .Y(new_n23382_));
  AOI21X1  g23190(.A0(new_n23382_), .A1(new_n23380_), .B0(new_n23350_), .Y(new_n23383_));
  NOR3X1   g23191(.A(new_n23383_), .B(new_n23381_), .C(\asqrt[44] ), .Y(new_n23384_));
  NOR2X1   g23192(.A(new_n23384_), .B(new_n23371_), .Y(new_n23385_));
  OR4X1    g23193(.A(new_n22874_), .B(new_n22632_), .C(new_n22620_), .D(new_n22615_), .Y(new_n23386_));
  OR2X1    g23194(.A(new_n22632_), .B(new_n22615_), .Y(new_n23387_));
  OAI21X1  g23195(.A0(new_n23387_), .A1(new_n22874_), .B0(new_n22620_), .Y(new_n23388_));
  AND2X1   g23196(.A(new_n23388_), .B(new_n23386_), .Y(new_n23389_));
  INVX1    g23197(.A(new_n23389_), .Y(new_n23390_));
  OAI21X1  g23198(.A0(new_n23383_), .A1(new_n23381_), .B0(\asqrt[44] ), .Y(new_n23391_));
  NAND2X1  g23199(.A(new_n23391_), .B(new_n2570_), .Y(new_n23392_));
  OAI21X1  g23200(.A0(new_n23392_), .A1(new_n23385_), .B0(new_n23390_), .Y(new_n23393_));
  AOI21X1  g23201(.A0(new_n23393_), .A1(new_n23375_), .B0(new_n2263_), .Y(new_n23394_));
  AOI21X1  g23202(.A0(new_n22677_), .A1(new_n22676_), .B0(new_n22639_), .Y(new_n23395_));
  AND2X1   g23203(.A(new_n23395_), .B(new_n22623_), .Y(new_n23396_));
  AOI22X1  g23204(.A0(new_n22677_), .A1(new_n22676_), .B0(new_n22649_), .B1(\asqrt[45] ), .Y(new_n23397_));
  AOI21X1  g23205(.A0(new_n23397_), .A1(\asqrt[4] ), .B0(new_n22638_), .Y(new_n23398_));
  AOI21X1  g23206(.A0(new_n23396_), .A1(\asqrt[4] ), .B0(new_n23398_), .Y(new_n23399_));
  OAI21X1  g23207(.A0(new_n23384_), .A1(new_n23371_), .B0(new_n23391_), .Y(new_n23400_));
  AOI21X1  g23208(.A0(new_n23400_), .A1(\asqrt[45] ), .B0(\asqrt[46] ), .Y(new_n23401_));
  AOI21X1  g23209(.A0(new_n23401_), .A1(new_n23393_), .B0(new_n23399_), .Y(new_n23402_));
  OAI21X1  g23210(.A0(new_n23402_), .A1(new_n23394_), .B0(\asqrt[47] ), .Y(new_n23403_));
  AND2X1   g23211(.A(new_n22650_), .B(new_n22642_), .Y(new_n23404_));
  NOR3X1   g23212(.A(new_n23404_), .B(new_n22680_), .C(new_n22643_), .Y(new_n23405_));
  NOR3X1   g23213(.A(new_n22874_), .B(new_n23404_), .C(new_n22643_), .Y(new_n23406_));
  NOR2X1   g23214(.A(new_n23406_), .B(new_n22648_), .Y(new_n23407_));
  AOI21X1  g23215(.A0(new_n23405_), .A1(\asqrt[4] ), .B0(new_n23407_), .Y(new_n23408_));
  NOR3X1   g23216(.A(new_n23402_), .B(new_n23394_), .C(\asqrt[47] ), .Y(new_n23409_));
  OAI21X1  g23217(.A0(new_n23409_), .A1(new_n23408_), .B0(new_n23403_), .Y(new_n23410_));
  AND2X1   g23218(.A(new_n23410_), .B(\asqrt[48] ), .Y(new_n23411_));
  OR2X1    g23219(.A(new_n23409_), .B(new_n23408_), .Y(new_n23412_));
  OR4X1    g23220(.A(new_n22874_), .B(new_n22657_), .C(new_n22684_), .D(new_n22683_), .Y(new_n23413_));
  OR2X1    g23221(.A(new_n22657_), .B(new_n22683_), .Y(new_n23414_));
  OAI21X1  g23222(.A0(new_n23414_), .A1(new_n22874_), .B0(new_n22684_), .Y(new_n23415_));
  AND2X1   g23223(.A(new_n23415_), .B(new_n23413_), .Y(new_n23416_));
  AND2X1   g23224(.A(new_n23403_), .B(new_n1834_), .Y(new_n23417_));
  AOI21X1  g23225(.A0(new_n23417_), .A1(new_n23412_), .B0(new_n23416_), .Y(new_n23418_));
  OAI21X1  g23226(.A0(new_n23418_), .A1(new_n23411_), .B0(\asqrt[49] ), .Y(new_n23419_));
  AND2X1   g23227(.A(new_n22666_), .B(new_n22660_), .Y(new_n23420_));
  NOR3X1   g23228(.A(new_n23420_), .B(new_n22700_), .C(new_n22659_), .Y(new_n23421_));
  NOR3X1   g23229(.A(new_n22874_), .B(new_n23420_), .C(new_n22659_), .Y(new_n23422_));
  NOR2X1   g23230(.A(new_n23422_), .B(new_n22665_), .Y(new_n23423_));
  AOI21X1  g23231(.A0(new_n23421_), .A1(\asqrt[4] ), .B0(new_n23423_), .Y(new_n23424_));
  INVX1    g23232(.A(new_n23424_), .Y(new_n23425_));
  AND2X1   g23233(.A(new_n23400_), .B(\asqrt[45] ), .Y(new_n23426_));
  OR2X1    g23234(.A(new_n23384_), .B(new_n23371_), .Y(new_n23427_));
  AND2X1   g23235(.A(new_n23391_), .B(new_n2570_), .Y(new_n23428_));
  AOI21X1  g23236(.A0(new_n23428_), .A1(new_n23427_), .B0(new_n23389_), .Y(new_n23429_));
  OAI21X1  g23237(.A0(new_n23429_), .A1(new_n23426_), .B0(\asqrt[46] ), .Y(new_n23430_));
  INVX1    g23238(.A(new_n23399_), .Y(new_n23431_));
  OAI21X1  g23239(.A0(new_n23374_), .A1(new_n2570_), .B0(new_n2263_), .Y(new_n23432_));
  OAI21X1  g23240(.A0(new_n23432_), .A1(new_n23429_), .B0(new_n23431_), .Y(new_n23433_));
  AOI21X1  g23241(.A0(new_n23433_), .A1(new_n23430_), .B0(new_n2040_), .Y(new_n23434_));
  INVX1    g23242(.A(new_n23408_), .Y(new_n23435_));
  NAND3X1  g23243(.A(new_n23433_), .B(new_n23430_), .C(new_n2040_), .Y(new_n23436_));
  AOI21X1  g23244(.A0(new_n23436_), .A1(new_n23435_), .B0(new_n23434_), .Y(new_n23437_));
  OAI21X1  g23245(.A0(new_n23437_), .A1(new_n1834_), .B0(new_n1632_), .Y(new_n23438_));
  OAI21X1  g23246(.A0(new_n23438_), .A1(new_n23418_), .B0(new_n23425_), .Y(new_n23439_));
  AOI21X1  g23247(.A0(new_n23439_), .A1(new_n23419_), .B0(new_n1469_), .Y(new_n23440_));
  AND2X1   g23248(.A(new_n22704_), .B(new_n22702_), .Y(new_n23441_));
  NOR3X1   g23249(.A(new_n23441_), .B(new_n22674_), .C(new_n22703_), .Y(new_n23442_));
  NOR3X1   g23250(.A(new_n22874_), .B(new_n23441_), .C(new_n22703_), .Y(new_n23443_));
  NOR2X1   g23251(.A(new_n23443_), .B(new_n22673_), .Y(new_n23444_));
  AOI21X1  g23252(.A0(new_n23442_), .A1(\asqrt[4] ), .B0(new_n23444_), .Y(new_n23445_));
  INVX1    g23253(.A(new_n23445_), .Y(new_n23446_));
  NAND3X1  g23254(.A(new_n23439_), .B(new_n23419_), .C(new_n1469_), .Y(new_n23447_));
  AOI21X1  g23255(.A0(new_n23447_), .A1(new_n23446_), .B0(new_n23440_), .Y(new_n23448_));
  OR2X1    g23256(.A(new_n23448_), .B(new_n1277_), .Y(new_n23449_));
  OR2X1    g23257(.A(new_n23437_), .B(new_n1834_), .Y(new_n23450_));
  NOR2X1   g23258(.A(new_n23409_), .B(new_n23408_), .Y(new_n23451_));
  INVX1    g23259(.A(new_n23416_), .Y(new_n23452_));
  NAND2X1  g23260(.A(new_n23403_), .B(new_n1834_), .Y(new_n23453_));
  OAI21X1  g23261(.A0(new_n23453_), .A1(new_n23451_), .B0(new_n23452_), .Y(new_n23454_));
  AOI21X1  g23262(.A0(new_n23454_), .A1(new_n23450_), .B0(new_n1632_), .Y(new_n23455_));
  AOI21X1  g23263(.A0(new_n23410_), .A1(\asqrt[48] ), .B0(\asqrt[49] ), .Y(new_n23456_));
  AOI21X1  g23264(.A0(new_n23456_), .A1(new_n23454_), .B0(new_n23424_), .Y(new_n23457_));
  NOR3X1   g23265(.A(new_n23457_), .B(new_n23455_), .C(\asqrt[50] ), .Y(new_n23458_));
  NOR2X1   g23266(.A(new_n23458_), .B(new_n23445_), .Y(new_n23459_));
  OR4X1    g23267(.A(new_n22874_), .B(new_n22706_), .C(new_n22694_), .D(new_n22689_), .Y(new_n23460_));
  OR2X1    g23268(.A(new_n22706_), .B(new_n22689_), .Y(new_n23461_));
  OAI21X1  g23269(.A0(new_n23461_), .A1(new_n22874_), .B0(new_n22694_), .Y(new_n23462_));
  AND2X1   g23270(.A(new_n23462_), .B(new_n23460_), .Y(new_n23463_));
  INVX1    g23271(.A(new_n23463_), .Y(new_n23464_));
  OAI21X1  g23272(.A0(new_n23457_), .A1(new_n23455_), .B0(\asqrt[50] ), .Y(new_n23465_));
  NAND2X1  g23273(.A(new_n23465_), .B(new_n1277_), .Y(new_n23466_));
  OAI21X1  g23274(.A0(new_n23466_), .A1(new_n23459_), .B0(new_n23464_), .Y(new_n23467_));
  AOI21X1  g23275(.A0(new_n23467_), .A1(new_n23449_), .B0(new_n1111_), .Y(new_n23468_));
  AOI21X1  g23276(.A0(new_n22751_), .A1(new_n22750_), .B0(new_n22713_), .Y(new_n23469_));
  AND2X1   g23277(.A(new_n23469_), .B(new_n22697_), .Y(new_n23470_));
  AOI22X1  g23278(.A0(new_n22751_), .A1(new_n22750_), .B0(new_n22723_), .B1(\asqrt[51] ), .Y(new_n23471_));
  AOI21X1  g23279(.A0(new_n23471_), .A1(\asqrt[4] ), .B0(new_n22712_), .Y(new_n23472_));
  AOI21X1  g23280(.A0(new_n23470_), .A1(\asqrt[4] ), .B0(new_n23472_), .Y(new_n23473_));
  OAI21X1  g23281(.A0(new_n23458_), .A1(new_n23445_), .B0(new_n23465_), .Y(new_n23474_));
  AOI21X1  g23282(.A0(new_n23474_), .A1(\asqrt[51] ), .B0(\asqrt[52] ), .Y(new_n23475_));
  AOI21X1  g23283(.A0(new_n23475_), .A1(new_n23467_), .B0(new_n23473_), .Y(new_n23476_));
  OAI21X1  g23284(.A0(new_n23476_), .A1(new_n23468_), .B0(\asqrt[53] ), .Y(new_n23477_));
  AND2X1   g23285(.A(new_n22724_), .B(new_n22716_), .Y(new_n23478_));
  NOR3X1   g23286(.A(new_n23478_), .B(new_n22754_), .C(new_n22717_), .Y(new_n23479_));
  NOR3X1   g23287(.A(new_n22874_), .B(new_n23478_), .C(new_n22717_), .Y(new_n23480_));
  NOR2X1   g23288(.A(new_n23480_), .B(new_n22722_), .Y(new_n23481_));
  AOI21X1  g23289(.A0(new_n23479_), .A1(\asqrt[4] ), .B0(new_n23481_), .Y(new_n23482_));
  NOR3X1   g23290(.A(new_n23476_), .B(new_n23468_), .C(\asqrt[53] ), .Y(new_n23483_));
  OAI21X1  g23291(.A0(new_n23483_), .A1(new_n23482_), .B0(new_n23477_), .Y(new_n23484_));
  AND2X1   g23292(.A(new_n23484_), .B(\asqrt[54] ), .Y(new_n23485_));
  OR2X1    g23293(.A(new_n23483_), .B(new_n23482_), .Y(new_n23486_));
  OR4X1    g23294(.A(new_n22874_), .B(new_n22731_), .C(new_n22758_), .D(new_n22757_), .Y(new_n23487_));
  OR2X1    g23295(.A(new_n22731_), .B(new_n22757_), .Y(new_n23488_));
  OAI21X1  g23296(.A0(new_n23488_), .A1(new_n22874_), .B0(new_n22758_), .Y(new_n23489_));
  AND2X1   g23297(.A(new_n23489_), .B(new_n23487_), .Y(new_n23490_));
  AND2X1   g23298(.A(new_n23477_), .B(new_n902_), .Y(new_n23491_));
  AOI21X1  g23299(.A0(new_n23491_), .A1(new_n23486_), .B0(new_n23490_), .Y(new_n23492_));
  OAI21X1  g23300(.A0(new_n23492_), .A1(new_n23485_), .B0(\asqrt[55] ), .Y(new_n23493_));
  AND2X1   g23301(.A(new_n22740_), .B(new_n22734_), .Y(new_n23494_));
  NOR3X1   g23302(.A(new_n23494_), .B(new_n22774_), .C(new_n22733_), .Y(new_n23495_));
  NOR3X1   g23303(.A(new_n22874_), .B(new_n23494_), .C(new_n22733_), .Y(new_n23496_));
  NOR2X1   g23304(.A(new_n23496_), .B(new_n22739_), .Y(new_n23497_));
  AOI21X1  g23305(.A0(new_n23495_), .A1(\asqrt[4] ), .B0(new_n23497_), .Y(new_n23498_));
  INVX1    g23306(.A(new_n23498_), .Y(new_n23499_));
  AND2X1   g23307(.A(new_n23474_), .B(\asqrt[51] ), .Y(new_n23500_));
  OR2X1    g23308(.A(new_n23458_), .B(new_n23445_), .Y(new_n23501_));
  AND2X1   g23309(.A(new_n23465_), .B(new_n1277_), .Y(new_n23502_));
  AOI21X1  g23310(.A0(new_n23502_), .A1(new_n23501_), .B0(new_n23463_), .Y(new_n23503_));
  OAI21X1  g23311(.A0(new_n23503_), .A1(new_n23500_), .B0(\asqrt[52] ), .Y(new_n23504_));
  INVX1    g23312(.A(new_n23473_), .Y(new_n23505_));
  OAI21X1  g23313(.A0(new_n23448_), .A1(new_n1277_), .B0(new_n1111_), .Y(new_n23506_));
  OAI21X1  g23314(.A0(new_n23506_), .A1(new_n23503_), .B0(new_n23505_), .Y(new_n23507_));
  AOI21X1  g23315(.A0(new_n23507_), .A1(new_n23504_), .B0(new_n968_), .Y(new_n23508_));
  INVX1    g23316(.A(new_n23482_), .Y(new_n23509_));
  NAND3X1  g23317(.A(new_n23507_), .B(new_n23504_), .C(new_n968_), .Y(new_n23510_));
  AOI21X1  g23318(.A0(new_n23510_), .A1(new_n23509_), .B0(new_n23508_), .Y(new_n23511_));
  OAI21X1  g23319(.A0(new_n23511_), .A1(new_n902_), .B0(new_n697_), .Y(new_n23512_));
  OAI21X1  g23320(.A0(new_n23512_), .A1(new_n23492_), .B0(new_n23499_), .Y(new_n23513_));
  AOI21X1  g23321(.A0(new_n23513_), .A1(new_n23493_), .B0(new_n582_), .Y(new_n23514_));
  AND2X1   g23322(.A(new_n22778_), .B(new_n22776_), .Y(new_n23515_));
  NOR3X1   g23323(.A(new_n23515_), .B(new_n22748_), .C(new_n22777_), .Y(new_n23516_));
  NOR3X1   g23324(.A(new_n22874_), .B(new_n23515_), .C(new_n22777_), .Y(new_n23517_));
  NOR2X1   g23325(.A(new_n23517_), .B(new_n22747_), .Y(new_n23518_));
  AOI21X1  g23326(.A0(new_n23516_), .A1(\asqrt[4] ), .B0(new_n23518_), .Y(new_n23519_));
  INVX1    g23327(.A(new_n23519_), .Y(new_n23520_));
  NAND3X1  g23328(.A(new_n23513_), .B(new_n23493_), .C(new_n582_), .Y(new_n23521_));
  AOI21X1  g23329(.A0(new_n23521_), .A1(new_n23520_), .B0(new_n23514_), .Y(new_n23522_));
  OR2X1    g23330(.A(new_n23522_), .B(new_n481_), .Y(new_n23523_));
  OR2X1    g23331(.A(new_n23511_), .B(new_n902_), .Y(new_n23524_));
  NOR2X1   g23332(.A(new_n23483_), .B(new_n23482_), .Y(new_n23525_));
  INVX1    g23333(.A(new_n23490_), .Y(new_n23526_));
  NAND2X1  g23334(.A(new_n23477_), .B(new_n902_), .Y(new_n23527_));
  OAI21X1  g23335(.A0(new_n23527_), .A1(new_n23525_), .B0(new_n23526_), .Y(new_n23528_));
  AOI21X1  g23336(.A0(new_n23528_), .A1(new_n23524_), .B0(new_n697_), .Y(new_n23529_));
  AOI21X1  g23337(.A0(new_n23484_), .A1(\asqrt[54] ), .B0(\asqrt[55] ), .Y(new_n23530_));
  AOI21X1  g23338(.A0(new_n23530_), .A1(new_n23528_), .B0(new_n23498_), .Y(new_n23531_));
  NOR3X1   g23339(.A(new_n23531_), .B(new_n23529_), .C(\asqrt[56] ), .Y(new_n23532_));
  NOR2X1   g23340(.A(new_n23532_), .B(new_n23519_), .Y(new_n23533_));
  OR4X1    g23341(.A(new_n22874_), .B(new_n22780_), .C(new_n22768_), .D(new_n22763_), .Y(new_n23534_));
  OR2X1    g23342(.A(new_n22780_), .B(new_n22763_), .Y(new_n23535_));
  OAI21X1  g23343(.A0(new_n23535_), .A1(new_n22874_), .B0(new_n22768_), .Y(new_n23536_));
  AND2X1   g23344(.A(new_n23536_), .B(new_n23534_), .Y(new_n23537_));
  INVX1    g23345(.A(new_n23537_), .Y(new_n23538_));
  OAI21X1  g23346(.A0(new_n23531_), .A1(new_n23529_), .B0(\asqrt[56] ), .Y(new_n23539_));
  NAND2X1  g23347(.A(new_n23539_), .B(new_n481_), .Y(new_n23540_));
  OAI21X1  g23348(.A0(new_n23540_), .A1(new_n23533_), .B0(new_n23538_), .Y(new_n23541_));
  AOI21X1  g23349(.A0(new_n23541_), .A1(new_n23523_), .B0(new_n399_), .Y(new_n23542_));
  AOI21X1  g23350(.A0(new_n22825_), .A1(new_n22824_), .B0(new_n22787_), .Y(new_n23543_));
  AND2X1   g23351(.A(new_n23543_), .B(new_n22771_), .Y(new_n23544_));
  AOI22X1  g23352(.A0(new_n22825_), .A1(new_n22824_), .B0(new_n22797_), .B1(\asqrt[57] ), .Y(new_n23545_));
  AOI21X1  g23353(.A0(new_n23545_), .A1(\asqrt[4] ), .B0(new_n22786_), .Y(new_n23546_));
  AOI21X1  g23354(.A0(new_n23544_), .A1(\asqrt[4] ), .B0(new_n23546_), .Y(new_n23547_));
  OAI21X1  g23355(.A0(new_n23532_), .A1(new_n23519_), .B0(new_n23539_), .Y(new_n23548_));
  AOI21X1  g23356(.A0(new_n23548_), .A1(\asqrt[57] ), .B0(\asqrt[58] ), .Y(new_n23549_));
  AOI21X1  g23357(.A0(new_n23549_), .A1(new_n23541_), .B0(new_n23547_), .Y(new_n23550_));
  OAI21X1  g23358(.A0(new_n23550_), .A1(new_n23542_), .B0(\asqrt[59] ), .Y(new_n23551_));
  AND2X1   g23359(.A(new_n22798_), .B(new_n22790_), .Y(new_n23552_));
  NOR3X1   g23360(.A(new_n23552_), .B(new_n22828_), .C(new_n22791_), .Y(new_n23553_));
  NOR3X1   g23361(.A(new_n22874_), .B(new_n23552_), .C(new_n22791_), .Y(new_n23554_));
  NOR2X1   g23362(.A(new_n23554_), .B(new_n22796_), .Y(new_n23555_));
  AOI21X1  g23363(.A0(new_n23553_), .A1(\asqrt[4] ), .B0(new_n23555_), .Y(new_n23556_));
  NOR3X1   g23364(.A(new_n23550_), .B(new_n23542_), .C(\asqrt[59] ), .Y(new_n23557_));
  OAI21X1  g23365(.A0(new_n23557_), .A1(new_n23556_), .B0(new_n23551_), .Y(new_n23558_));
  AND2X1   g23366(.A(new_n23558_), .B(\asqrt[60] ), .Y(new_n23559_));
  OR2X1    g23367(.A(new_n23557_), .B(new_n23556_), .Y(new_n23560_));
  OR4X1    g23368(.A(new_n22874_), .B(new_n22805_), .C(new_n22832_), .D(new_n22831_), .Y(new_n23561_));
  OR2X1    g23369(.A(new_n22805_), .B(new_n22831_), .Y(new_n23562_));
  OAI21X1  g23370(.A0(new_n23562_), .A1(new_n22874_), .B0(new_n22832_), .Y(new_n23563_));
  AND2X1   g23371(.A(new_n23563_), .B(new_n23561_), .Y(new_n23564_));
  AND2X1   g23372(.A(new_n23551_), .B(new_n292_), .Y(new_n23565_));
  AOI21X1  g23373(.A0(new_n23565_), .A1(new_n23560_), .B0(new_n23564_), .Y(new_n23566_));
  OAI21X1  g23374(.A0(new_n23566_), .A1(new_n23559_), .B0(\asqrt[61] ), .Y(new_n23567_));
  AND2X1   g23375(.A(new_n23548_), .B(\asqrt[57] ), .Y(new_n23568_));
  OR2X1    g23376(.A(new_n23532_), .B(new_n23519_), .Y(new_n23569_));
  AND2X1   g23377(.A(new_n23539_), .B(new_n481_), .Y(new_n23570_));
  AOI21X1  g23378(.A0(new_n23570_), .A1(new_n23569_), .B0(new_n23537_), .Y(new_n23571_));
  OAI21X1  g23379(.A0(new_n23571_), .A1(new_n23568_), .B0(\asqrt[58] ), .Y(new_n23572_));
  INVX1    g23380(.A(new_n23547_), .Y(new_n23573_));
  OAI21X1  g23381(.A0(new_n23522_), .A1(new_n481_), .B0(new_n399_), .Y(new_n23574_));
  OAI21X1  g23382(.A0(new_n23574_), .A1(new_n23571_), .B0(new_n23573_), .Y(new_n23575_));
  AOI21X1  g23383(.A0(new_n23575_), .A1(new_n23572_), .B0(new_n328_), .Y(new_n23576_));
  INVX1    g23384(.A(new_n23556_), .Y(new_n23577_));
  NAND3X1  g23385(.A(new_n23575_), .B(new_n23572_), .C(new_n328_), .Y(new_n23578_));
  AOI21X1  g23386(.A0(new_n23578_), .A1(new_n23577_), .B0(new_n23576_), .Y(new_n23579_));
  OAI21X1  g23387(.A0(new_n23579_), .A1(new_n292_), .B0(new_n217_), .Y(new_n23580_));
  AND2X1   g23388(.A(new_n22809_), .B(new_n22808_), .Y(new_n23581_));
  NOR3X1   g23389(.A(new_n22860_), .B(new_n23581_), .C(new_n22807_), .Y(new_n23582_));
  NOR3X1   g23390(.A(new_n22874_), .B(new_n23581_), .C(new_n22807_), .Y(new_n23583_));
  NOR2X1   g23391(.A(new_n23583_), .B(new_n22814_), .Y(new_n23584_));
  AOI21X1  g23392(.A0(new_n23582_), .A1(\asqrt[4] ), .B0(new_n23584_), .Y(new_n23585_));
  INVX1    g23393(.A(new_n23585_), .Y(new_n23586_));
  OAI21X1  g23394(.A0(new_n23580_), .A1(new_n23566_), .B0(new_n23586_), .Y(new_n23587_));
  AOI21X1  g23395(.A0(new_n23587_), .A1(new_n23567_), .B0(new_n199_), .Y(new_n23588_));
  AND2X1   g23396(.A(new_n22863_), .B(new_n22861_), .Y(new_n23589_));
  NOR3X1   g23397(.A(new_n23589_), .B(new_n22822_), .C(new_n22862_), .Y(new_n23590_));
  NOR3X1   g23398(.A(new_n22874_), .B(new_n23589_), .C(new_n22862_), .Y(new_n23591_));
  NOR2X1   g23399(.A(new_n23591_), .B(new_n22821_), .Y(new_n23592_));
  AOI21X1  g23400(.A0(new_n23590_), .A1(\asqrt[4] ), .B0(new_n23592_), .Y(new_n23593_));
  INVX1    g23401(.A(new_n23593_), .Y(new_n23594_));
  NAND3X1  g23402(.A(new_n23587_), .B(new_n23567_), .C(new_n199_), .Y(new_n23595_));
  AOI21X1  g23403(.A0(new_n23595_), .A1(new_n23594_), .B0(new_n23588_), .Y(new_n23596_));
  NAND4X1  g23404(.A(\asqrt[4] ), .B(new_n22843_), .C(new_n22841_), .D(new_n22867_), .Y(new_n23597_));
  NAND2X1  g23405(.A(new_n22843_), .B(new_n22867_), .Y(new_n23598_));
  OAI21X1  g23406(.A0(new_n23598_), .A1(new_n22874_), .B0(new_n22842_), .Y(new_n23599_));
  AND2X1   g23407(.A(new_n23599_), .B(new_n23597_), .Y(new_n23600_));
  NOR3X1   g23408(.A(new_n22874_), .B(new_n22849_), .C(new_n22844_), .Y(new_n23601_));
  NOR3X1   g23409(.A(new_n23601_), .B(new_n23600_), .C(new_n22896_), .Y(new_n23602_));
  INVX1    g23410(.A(new_n23602_), .Y(new_n23603_));
  OAI21X1  g23411(.A0(new_n23603_), .A1(new_n23596_), .B0(new_n193_), .Y(new_n23604_));
  OR2X1    g23412(.A(new_n23579_), .B(new_n292_), .Y(new_n23605_));
  NOR2X1   g23413(.A(new_n23557_), .B(new_n23556_), .Y(new_n23606_));
  INVX1    g23414(.A(new_n23564_), .Y(new_n23607_));
  NAND2X1  g23415(.A(new_n23551_), .B(new_n292_), .Y(new_n23608_));
  OAI21X1  g23416(.A0(new_n23608_), .A1(new_n23606_), .B0(new_n23607_), .Y(new_n23609_));
  AOI21X1  g23417(.A0(new_n23609_), .A1(new_n23605_), .B0(new_n217_), .Y(new_n23610_));
  AOI21X1  g23418(.A0(new_n23558_), .A1(\asqrt[60] ), .B0(\asqrt[61] ), .Y(new_n23611_));
  AOI21X1  g23419(.A0(new_n23611_), .A1(new_n23609_), .B0(new_n23585_), .Y(new_n23612_));
  NOR3X1   g23420(.A(new_n23612_), .B(new_n23610_), .C(\asqrt[62] ), .Y(new_n23613_));
  OR2X1    g23421(.A(new_n23613_), .B(new_n23593_), .Y(new_n23614_));
  OAI21X1  g23422(.A0(new_n23612_), .A1(new_n23610_), .B0(\asqrt[62] ), .Y(new_n23615_));
  AND2X1   g23423(.A(new_n23600_), .B(new_n23615_), .Y(new_n23616_));
  AOI21X1  g23424(.A0(new_n22873_), .A1(new_n22856_), .B0(new_n22849_), .Y(new_n23617_));
  AOI21X1  g23425(.A0(new_n22850_), .A1(new_n22885_), .B0(new_n193_), .Y(new_n23618_));
  OAI21X1  g23426(.A0(new_n23617_), .A1(new_n22885_), .B0(new_n23618_), .Y(new_n23619_));
  INVX1    g23427(.A(new_n23619_), .Y(new_n23620_));
  AOI21X1  g23428(.A0(new_n23616_), .A1(new_n23614_), .B0(new_n23620_), .Y(new_n23621_));
  AND2X1   g23429(.A(new_n23621_), .B(new_n23604_), .Y(new_n23622_));
  INVX1    g23430(.A(new_n23622_), .Y(\asqrt[3] ));
  INVX1    g23431(.A(\a[4] ), .Y(new_n23624_));
  NOR2X1   g23432(.A(\a[3] ), .B(\a[2] ), .Y(new_n23625_));
  INVX1    g23433(.A(\a[6] ), .Y(new_n23626_));
  AOI21X1  g23434(.A0(new_n23621_), .A1(new_n23604_), .B0(new_n23626_), .Y(new_n23627_));
  NOR3X1   g23435(.A(\a[6] ), .B(\a[5] ), .C(\a[4] ), .Y(new_n23628_));
  OAI21X1  g23436(.A0(new_n23628_), .A1(new_n23627_), .B0(\asqrt[4] ), .Y(new_n23629_));
  OAI21X1  g23437(.A0(new_n23613_), .A1(new_n23593_), .B0(new_n23615_), .Y(new_n23630_));
  AOI21X1  g23438(.A0(new_n23602_), .A1(new_n23630_), .B0(\asqrt[63] ), .Y(new_n23631_));
  NOR2X1   g23439(.A(new_n23613_), .B(new_n23593_), .Y(new_n23632_));
  NAND2X1  g23440(.A(new_n23600_), .B(new_n23615_), .Y(new_n23633_));
  OAI21X1  g23441(.A0(new_n23633_), .A1(new_n23632_), .B0(new_n23619_), .Y(new_n23634_));
  OAI21X1  g23442(.A0(new_n23634_), .A1(new_n23631_), .B0(\a[6] ), .Y(new_n23635_));
  NOR4X1   g23443(.A(new_n23628_), .B(new_n22872_), .C(new_n22896_), .D(new_n22886_), .Y(new_n23636_));
  AND2X1   g23444(.A(new_n23636_), .B(new_n23635_), .Y(new_n23637_));
  INVX1    g23445(.A(\a[7] ), .Y(new_n23638_));
  AOI21X1  g23446(.A0(new_n23621_), .A1(new_n23604_), .B0(\a[6] ), .Y(new_n23639_));
  NOR2X1   g23447(.A(\a[7] ), .B(\a[6] ), .Y(new_n23640_));
  OAI21X1  g23448(.A0(new_n23634_), .A1(new_n23631_), .B0(new_n23640_), .Y(new_n23641_));
  OAI21X1  g23449(.A0(new_n23639_), .A1(new_n23638_), .B0(new_n23641_), .Y(new_n23642_));
  OAI21X1  g23450(.A0(new_n23642_), .A1(new_n23637_), .B0(new_n23629_), .Y(new_n23643_));
  AND2X1   g23451(.A(new_n23643_), .B(\asqrt[5] ), .Y(new_n23644_));
  OR2X1    g23452(.A(new_n23642_), .B(new_n23637_), .Y(new_n23645_));
  AND2X1   g23453(.A(new_n23629_), .B(new_n22128_), .Y(new_n23646_));
  AND2X1   g23454(.A(new_n23616_), .B(new_n23614_), .Y(new_n23647_));
  OR4X1    g23455(.A(new_n23620_), .B(new_n23647_), .C(new_n23631_), .D(new_n22874_), .Y(new_n23648_));
  AOI21X1  g23456(.A0(new_n23648_), .A1(new_n23641_), .B0(new_n22876_), .Y(new_n23649_));
  INVX1    g23457(.A(new_n23640_), .Y(new_n23650_));
  AOI21X1  g23458(.A0(new_n23621_), .A1(new_n23604_), .B0(new_n23650_), .Y(new_n23651_));
  NOR4X1   g23459(.A(new_n23620_), .B(new_n23647_), .C(new_n23631_), .D(new_n22874_), .Y(new_n23652_));
  NOR3X1   g23460(.A(new_n23652_), .B(new_n23651_), .C(\a[8] ), .Y(new_n23653_));
  NOR2X1   g23461(.A(new_n23653_), .B(new_n23649_), .Y(new_n23654_));
  AOI21X1  g23462(.A0(new_n23646_), .A1(new_n23645_), .B0(new_n23654_), .Y(new_n23655_));
  OAI21X1  g23463(.A0(new_n23655_), .A1(new_n23644_), .B0(\asqrt[6] ), .Y(new_n23656_));
  OR4X1    g23464(.A(new_n23622_), .B(new_n22916_), .C(new_n22882_), .D(new_n22913_), .Y(new_n23657_));
  OR2X1    g23465(.A(new_n22882_), .B(new_n22913_), .Y(new_n23658_));
  OAI21X1  g23466(.A0(new_n23658_), .A1(new_n23622_), .B0(new_n22916_), .Y(new_n23659_));
  NAND2X1  g23467(.A(new_n23659_), .B(new_n23657_), .Y(new_n23660_));
  INVX1    g23468(.A(new_n23628_), .Y(new_n23661_));
  AOI21X1  g23469(.A0(new_n23661_), .A1(new_n23635_), .B0(new_n22874_), .Y(new_n23662_));
  NAND2X1  g23470(.A(new_n23636_), .B(new_n23635_), .Y(new_n23663_));
  OAI21X1  g23471(.A0(new_n23634_), .A1(new_n23631_), .B0(new_n23626_), .Y(new_n23664_));
  AOI21X1  g23472(.A0(new_n23664_), .A1(\a[7] ), .B0(new_n23651_), .Y(new_n23665_));
  AOI21X1  g23473(.A0(new_n23665_), .A1(new_n23663_), .B0(new_n23662_), .Y(new_n23666_));
  OAI21X1  g23474(.A0(new_n23666_), .A1(new_n22128_), .B0(new_n21393_), .Y(new_n23667_));
  OAI21X1  g23475(.A0(new_n23667_), .A1(new_n23655_), .B0(new_n23660_), .Y(new_n23668_));
  AOI21X1  g23476(.A0(new_n23668_), .A1(new_n23656_), .B0(new_n20676_), .Y(new_n23669_));
  AOI21X1  g23477(.A0(new_n22895_), .A1(new_n22894_), .B0(new_n22935_), .Y(new_n23670_));
  AND2X1   g23478(.A(new_n23670_), .B(new_n22932_), .Y(new_n23671_));
  OAI21X1  g23479(.A0(new_n23634_), .A1(new_n23631_), .B0(new_n23671_), .Y(new_n23672_));
  AOI22X1  g23480(.A0(new_n22895_), .A1(new_n22894_), .B0(new_n22892_), .B1(\asqrt[6] ), .Y(new_n23673_));
  OAI21X1  g23481(.A0(new_n23634_), .A1(new_n23631_), .B0(new_n23673_), .Y(new_n23674_));
  NAND2X1  g23482(.A(new_n23674_), .B(new_n22935_), .Y(new_n23675_));
  AND2X1   g23483(.A(new_n23675_), .B(new_n23672_), .Y(new_n23676_));
  INVX1    g23484(.A(new_n23676_), .Y(new_n23677_));
  NAND3X1  g23485(.A(new_n23668_), .B(new_n23656_), .C(new_n20676_), .Y(new_n23678_));
  AOI21X1  g23486(.A0(new_n23678_), .A1(new_n23677_), .B0(new_n23669_), .Y(new_n23679_));
  OR2X1    g23487(.A(new_n23679_), .B(new_n19976_), .Y(new_n23680_));
  AND2X1   g23488(.A(new_n23678_), .B(new_n23677_), .Y(new_n23681_));
  AND2X1   g23489(.A(new_n22938_), .B(new_n22936_), .Y(new_n23682_));
  NOR3X1   g23490(.A(new_n23682_), .B(new_n22911_), .C(new_n22937_), .Y(new_n23683_));
  NOR2X1   g23491(.A(new_n23682_), .B(new_n22937_), .Y(new_n23684_));
  OAI21X1  g23492(.A0(new_n23634_), .A1(new_n23631_), .B0(new_n23684_), .Y(new_n23685_));
  AOI22X1  g23493(.A0(new_n23685_), .A1(new_n22911_), .B0(new_n23683_), .B1(\asqrt[3] ), .Y(new_n23686_));
  INVX1    g23494(.A(new_n23686_), .Y(new_n23687_));
  OR2X1    g23495(.A(new_n23666_), .B(new_n22128_), .Y(new_n23688_));
  NOR2X1   g23496(.A(new_n23642_), .B(new_n23637_), .Y(new_n23689_));
  OR2X1    g23497(.A(new_n23662_), .B(\asqrt[5] ), .Y(new_n23690_));
  OR2X1    g23498(.A(new_n23653_), .B(new_n23649_), .Y(new_n23691_));
  OAI21X1  g23499(.A0(new_n23690_), .A1(new_n23689_), .B0(new_n23691_), .Y(new_n23692_));
  AOI21X1  g23500(.A0(new_n23692_), .A1(new_n23688_), .B0(new_n21393_), .Y(new_n23693_));
  AOI21X1  g23501(.A0(new_n23643_), .A1(\asqrt[5] ), .B0(\asqrt[6] ), .Y(new_n23694_));
  AOI22X1  g23502(.A0(new_n23694_), .A1(new_n23692_), .B0(new_n23659_), .B1(new_n23657_), .Y(new_n23695_));
  OAI21X1  g23503(.A0(new_n23695_), .A1(new_n23693_), .B0(\asqrt[7] ), .Y(new_n23696_));
  NAND2X1  g23504(.A(new_n23696_), .B(new_n19976_), .Y(new_n23697_));
  OAI21X1  g23505(.A0(new_n23697_), .A1(new_n23681_), .B0(new_n23687_), .Y(new_n23698_));
  AOI21X1  g23506(.A0(new_n23698_), .A1(new_n23680_), .B0(new_n19273_), .Y(new_n23699_));
  NOR3X1   g23507(.A(new_n22940_), .B(new_n22928_), .C(new_n22920_), .Y(new_n23700_));
  NOR3X1   g23508(.A(new_n23622_), .B(new_n22940_), .C(new_n22920_), .Y(new_n23701_));
  NOR2X1   g23509(.A(new_n23701_), .B(new_n22927_), .Y(new_n23702_));
  AOI21X1  g23510(.A0(new_n23700_), .A1(\asqrt[3] ), .B0(new_n23702_), .Y(new_n23703_));
  NOR3X1   g23511(.A(new_n23695_), .B(new_n23693_), .C(\asqrt[7] ), .Y(new_n23704_));
  OAI21X1  g23512(.A0(new_n23704_), .A1(new_n23676_), .B0(new_n23696_), .Y(new_n23705_));
  AOI21X1  g23513(.A0(new_n23705_), .A1(\asqrt[8] ), .B0(\asqrt[9] ), .Y(new_n23706_));
  AOI21X1  g23514(.A0(new_n23706_), .A1(new_n23698_), .B0(new_n23703_), .Y(new_n23707_));
  OAI21X1  g23515(.A0(new_n23707_), .A1(new_n23699_), .B0(\asqrt[10] ), .Y(new_n23708_));
  AND2X1   g23516(.A(new_n22984_), .B(new_n22982_), .Y(new_n23709_));
  NOR3X1   g23517(.A(new_n23709_), .B(new_n22944_), .C(new_n22981_), .Y(new_n23710_));
  NOR3X1   g23518(.A(new_n23622_), .B(new_n23709_), .C(new_n22981_), .Y(new_n23711_));
  NOR2X1   g23519(.A(new_n23711_), .B(new_n22983_), .Y(new_n23712_));
  AOI21X1  g23520(.A0(new_n23710_), .A1(\asqrt[3] ), .B0(new_n23712_), .Y(new_n23713_));
  NOR3X1   g23521(.A(new_n23707_), .B(new_n23699_), .C(\asqrt[10] ), .Y(new_n23714_));
  OAI21X1  g23522(.A0(new_n23714_), .A1(new_n23713_), .B0(new_n23708_), .Y(new_n23715_));
  AND2X1   g23523(.A(new_n23715_), .B(\asqrt[11] ), .Y(new_n23716_));
  INVX1    g23524(.A(new_n23713_), .Y(new_n23717_));
  AND2X1   g23525(.A(new_n23705_), .B(\asqrt[8] ), .Y(new_n23718_));
  NAND2X1  g23526(.A(new_n23678_), .B(new_n23677_), .Y(new_n23719_));
  AND2X1   g23527(.A(new_n23696_), .B(new_n19976_), .Y(new_n23720_));
  AOI21X1  g23528(.A0(new_n23720_), .A1(new_n23719_), .B0(new_n23686_), .Y(new_n23721_));
  OAI21X1  g23529(.A0(new_n23721_), .A1(new_n23718_), .B0(\asqrt[9] ), .Y(new_n23722_));
  INVX1    g23530(.A(new_n23703_), .Y(new_n23723_));
  OAI21X1  g23531(.A0(new_n23679_), .A1(new_n19976_), .B0(new_n19273_), .Y(new_n23724_));
  OAI21X1  g23532(.A0(new_n23724_), .A1(new_n23721_), .B0(new_n23723_), .Y(new_n23725_));
  NAND3X1  g23533(.A(new_n23725_), .B(new_n23722_), .C(new_n18591_), .Y(new_n23726_));
  NAND2X1  g23534(.A(new_n23726_), .B(new_n23717_), .Y(new_n23727_));
  AND2X1   g23535(.A(new_n22955_), .B(new_n22946_), .Y(new_n23728_));
  NOR3X1   g23536(.A(new_n23728_), .B(new_n22987_), .C(new_n22947_), .Y(new_n23729_));
  NOR3X1   g23537(.A(new_n23622_), .B(new_n23728_), .C(new_n22947_), .Y(new_n23730_));
  NOR2X1   g23538(.A(new_n23730_), .B(new_n22952_), .Y(new_n23731_));
  AOI21X1  g23539(.A0(new_n23729_), .A1(\asqrt[3] ), .B0(new_n23731_), .Y(new_n23732_));
  AOI21X1  g23540(.A0(new_n23725_), .A1(new_n23722_), .B0(new_n18591_), .Y(new_n23733_));
  NOR2X1   g23541(.A(new_n23733_), .B(\asqrt[11] ), .Y(new_n23734_));
  AOI21X1  g23542(.A0(new_n23734_), .A1(new_n23727_), .B0(new_n23732_), .Y(new_n23735_));
  OAI21X1  g23543(.A0(new_n23735_), .A1(new_n23716_), .B0(\asqrt[12] ), .Y(new_n23736_));
  OR4X1    g23544(.A(new_n23622_), .B(new_n22964_), .C(new_n22991_), .D(new_n22990_), .Y(new_n23737_));
  OR2X1    g23545(.A(new_n22964_), .B(new_n22990_), .Y(new_n23738_));
  OAI21X1  g23546(.A0(new_n23738_), .A1(new_n23622_), .B0(new_n22991_), .Y(new_n23739_));
  AND2X1   g23547(.A(new_n23739_), .B(new_n23737_), .Y(new_n23740_));
  INVX1    g23548(.A(new_n23740_), .Y(new_n23741_));
  AOI21X1  g23549(.A0(new_n23726_), .A1(new_n23717_), .B0(new_n23733_), .Y(new_n23742_));
  OAI21X1  g23550(.A0(new_n23742_), .A1(new_n17927_), .B0(new_n17262_), .Y(new_n23743_));
  OAI21X1  g23551(.A0(new_n23743_), .A1(new_n23735_), .B0(new_n23741_), .Y(new_n23744_));
  AOI21X1  g23552(.A0(new_n23744_), .A1(new_n23736_), .B0(new_n16617_), .Y(new_n23745_));
  OAI21X1  g23553(.A0(new_n23009_), .A1(new_n23007_), .B0(new_n22971_), .Y(new_n23746_));
  NOR2X1   g23554(.A(new_n23746_), .B(new_n22966_), .Y(new_n23747_));
  AOI22X1  g23555(.A0(new_n22972_), .A1(new_n22967_), .B0(new_n22965_), .B1(\asqrt[12] ), .Y(new_n23748_));
  AOI21X1  g23556(.A0(new_n23748_), .A1(\asqrt[3] ), .B0(new_n22971_), .Y(new_n23749_));
  AOI21X1  g23557(.A0(new_n23747_), .A1(\asqrt[3] ), .B0(new_n23749_), .Y(new_n23750_));
  INVX1    g23558(.A(new_n23750_), .Y(new_n23751_));
  NAND3X1  g23559(.A(new_n23744_), .B(new_n23736_), .C(new_n16617_), .Y(new_n23752_));
  AOI21X1  g23560(.A0(new_n23752_), .A1(new_n23751_), .B0(new_n23745_), .Y(new_n23753_));
  OR2X1    g23561(.A(new_n23753_), .B(new_n15990_), .Y(new_n23754_));
  AND2X1   g23562(.A(new_n23752_), .B(new_n23751_), .Y(new_n23755_));
  AND2X1   g23563(.A(new_n23012_), .B(new_n23010_), .Y(new_n23756_));
  NOR3X1   g23564(.A(new_n23756_), .B(new_n22980_), .C(new_n23011_), .Y(new_n23757_));
  NOR3X1   g23565(.A(new_n23622_), .B(new_n23756_), .C(new_n23011_), .Y(new_n23758_));
  NOR2X1   g23566(.A(new_n23758_), .B(new_n22979_), .Y(new_n23759_));
  AOI21X1  g23567(.A0(new_n23757_), .A1(\asqrt[3] ), .B0(new_n23759_), .Y(new_n23760_));
  INVX1    g23568(.A(new_n23760_), .Y(new_n23761_));
  OR2X1    g23569(.A(new_n23742_), .B(new_n17927_), .Y(new_n23762_));
  AND2X1   g23570(.A(new_n23726_), .B(new_n23717_), .Y(new_n23763_));
  INVX1    g23571(.A(new_n23732_), .Y(new_n23764_));
  OR2X1    g23572(.A(new_n23733_), .B(\asqrt[11] ), .Y(new_n23765_));
  OAI21X1  g23573(.A0(new_n23765_), .A1(new_n23763_), .B0(new_n23764_), .Y(new_n23766_));
  AOI21X1  g23574(.A0(new_n23766_), .A1(new_n23762_), .B0(new_n17262_), .Y(new_n23767_));
  AOI21X1  g23575(.A0(new_n23715_), .A1(\asqrt[11] ), .B0(\asqrt[12] ), .Y(new_n23768_));
  AOI21X1  g23576(.A0(new_n23768_), .A1(new_n23766_), .B0(new_n23740_), .Y(new_n23769_));
  OAI21X1  g23577(.A0(new_n23769_), .A1(new_n23767_), .B0(\asqrt[13] ), .Y(new_n23770_));
  NAND2X1  g23578(.A(new_n23770_), .B(new_n15990_), .Y(new_n23771_));
  OAI21X1  g23579(.A0(new_n23771_), .A1(new_n23755_), .B0(new_n23761_), .Y(new_n23772_));
  AOI21X1  g23580(.A0(new_n23772_), .A1(new_n23754_), .B0(new_n15362_), .Y(new_n23773_));
  OR4X1    g23581(.A(new_n23622_), .B(new_n23014_), .C(new_n23002_), .D(new_n22996_), .Y(new_n23774_));
  OR2X1    g23582(.A(new_n23014_), .B(new_n22996_), .Y(new_n23775_));
  OAI21X1  g23583(.A0(new_n23775_), .A1(new_n23622_), .B0(new_n23002_), .Y(new_n23776_));
  AND2X1   g23584(.A(new_n23776_), .B(new_n23774_), .Y(new_n23777_));
  NOR3X1   g23585(.A(new_n23769_), .B(new_n23767_), .C(\asqrt[13] ), .Y(new_n23778_));
  OAI21X1  g23586(.A0(new_n23778_), .A1(new_n23750_), .B0(new_n23770_), .Y(new_n23779_));
  AOI21X1  g23587(.A0(new_n23779_), .A1(\asqrt[14] ), .B0(\asqrt[15] ), .Y(new_n23780_));
  AOI21X1  g23588(.A0(new_n23780_), .A1(new_n23772_), .B0(new_n23777_), .Y(new_n23781_));
  OAI21X1  g23589(.A0(new_n23781_), .A1(new_n23773_), .B0(\asqrt[16] ), .Y(new_n23782_));
  AND2X1   g23590(.A(new_n23045_), .B(new_n23044_), .Y(new_n23783_));
  NOR3X1   g23591(.A(new_n23783_), .B(new_n23020_), .C(new_n23043_), .Y(new_n23784_));
  NOR3X1   g23592(.A(new_n23622_), .B(new_n23783_), .C(new_n23043_), .Y(new_n23785_));
  NOR2X1   g23593(.A(new_n23785_), .B(new_n23019_), .Y(new_n23786_));
  AOI21X1  g23594(.A0(new_n23784_), .A1(\asqrt[3] ), .B0(new_n23786_), .Y(new_n23787_));
  NOR3X1   g23595(.A(new_n23781_), .B(new_n23773_), .C(\asqrt[16] ), .Y(new_n23788_));
  OAI21X1  g23596(.A0(new_n23788_), .A1(new_n23787_), .B0(new_n23782_), .Y(new_n23789_));
  AND2X1   g23597(.A(new_n23789_), .B(\asqrt[17] ), .Y(new_n23790_));
  INVX1    g23598(.A(new_n23787_), .Y(new_n23791_));
  AND2X1   g23599(.A(new_n23779_), .B(\asqrt[14] ), .Y(new_n23792_));
  NAND2X1  g23600(.A(new_n23752_), .B(new_n23751_), .Y(new_n23793_));
  AND2X1   g23601(.A(new_n23770_), .B(new_n15990_), .Y(new_n23794_));
  AOI21X1  g23602(.A0(new_n23794_), .A1(new_n23793_), .B0(new_n23760_), .Y(new_n23795_));
  OAI21X1  g23603(.A0(new_n23795_), .A1(new_n23792_), .B0(\asqrt[15] ), .Y(new_n23796_));
  INVX1    g23604(.A(new_n23777_), .Y(new_n23797_));
  OAI21X1  g23605(.A0(new_n23753_), .A1(new_n15990_), .B0(new_n15362_), .Y(new_n23798_));
  OAI21X1  g23606(.A0(new_n23798_), .A1(new_n23795_), .B0(new_n23797_), .Y(new_n23799_));
  NAND3X1  g23607(.A(new_n23799_), .B(new_n23796_), .C(new_n14754_), .Y(new_n23800_));
  NAND2X1  g23608(.A(new_n23800_), .B(new_n23791_), .Y(new_n23801_));
  AND2X1   g23609(.A(new_n23031_), .B(new_n23023_), .Y(new_n23802_));
  NOR3X1   g23610(.A(new_n23802_), .B(new_n23048_), .C(new_n23024_), .Y(new_n23803_));
  NOR3X1   g23611(.A(new_n23622_), .B(new_n23802_), .C(new_n23024_), .Y(new_n23804_));
  NOR2X1   g23612(.A(new_n23804_), .B(new_n23029_), .Y(new_n23805_));
  AOI21X1  g23613(.A0(new_n23803_), .A1(\asqrt[3] ), .B0(new_n23805_), .Y(new_n23806_));
  AND2X1   g23614(.A(new_n23782_), .B(new_n14165_), .Y(new_n23807_));
  AOI21X1  g23615(.A0(new_n23807_), .A1(new_n23801_), .B0(new_n23806_), .Y(new_n23808_));
  OAI21X1  g23616(.A0(new_n23808_), .A1(new_n23790_), .B0(\asqrt[18] ), .Y(new_n23809_));
  NAND4X1  g23617(.A(\asqrt[3] ), .B(new_n23051_), .C(new_n23038_), .D(new_n23033_), .Y(new_n23810_));
  NAND2X1  g23618(.A(new_n23051_), .B(new_n23033_), .Y(new_n23811_));
  OAI21X1  g23619(.A0(new_n23811_), .A1(new_n23622_), .B0(new_n23042_), .Y(new_n23812_));
  AND2X1   g23620(.A(new_n23812_), .B(new_n23810_), .Y(new_n23813_));
  INVX1    g23621(.A(new_n23813_), .Y(new_n23814_));
  AOI21X1  g23622(.A0(new_n23799_), .A1(new_n23796_), .B0(new_n14754_), .Y(new_n23815_));
  AOI21X1  g23623(.A0(new_n23800_), .A1(new_n23791_), .B0(new_n23815_), .Y(new_n23816_));
  OAI21X1  g23624(.A0(new_n23816_), .A1(new_n14165_), .B0(new_n13571_), .Y(new_n23817_));
  OAI21X1  g23625(.A0(new_n23817_), .A1(new_n23808_), .B0(new_n23814_), .Y(new_n23818_));
  AOI21X1  g23626(.A0(new_n23818_), .A1(new_n23809_), .B0(new_n13000_), .Y(new_n23819_));
  AOI21X1  g23627(.A0(new_n23058_), .A1(new_n23052_), .B0(new_n23096_), .Y(new_n23820_));
  AND2X1   g23628(.A(new_n23820_), .B(new_n23094_), .Y(new_n23821_));
  AOI22X1  g23629(.A0(new_n23058_), .A1(new_n23052_), .B0(new_n23040_), .B1(\asqrt[18] ), .Y(new_n23822_));
  AOI21X1  g23630(.A0(new_n23822_), .A1(\asqrt[3] ), .B0(new_n23056_), .Y(new_n23823_));
  AOI21X1  g23631(.A0(new_n23821_), .A1(\asqrt[3] ), .B0(new_n23823_), .Y(new_n23824_));
  INVX1    g23632(.A(new_n23824_), .Y(new_n23825_));
  NAND3X1  g23633(.A(new_n23818_), .B(new_n23809_), .C(new_n13000_), .Y(new_n23826_));
  AOI21X1  g23634(.A0(new_n23826_), .A1(new_n23825_), .B0(new_n23819_), .Y(new_n23827_));
  OR2X1    g23635(.A(new_n23827_), .B(new_n12447_), .Y(new_n23828_));
  AND2X1   g23636(.A(new_n23826_), .B(new_n23825_), .Y(new_n23829_));
  AND2X1   g23637(.A(new_n23100_), .B(new_n23098_), .Y(new_n23830_));
  NOR3X1   g23638(.A(new_n23830_), .B(new_n23066_), .C(new_n23099_), .Y(new_n23831_));
  NOR3X1   g23639(.A(new_n23622_), .B(new_n23830_), .C(new_n23099_), .Y(new_n23832_));
  NOR2X1   g23640(.A(new_n23832_), .B(new_n23065_), .Y(new_n23833_));
  AOI21X1  g23641(.A0(new_n23831_), .A1(\asqrt[3] ), .B0(new_n23833_), .Y(new_n23834_));
  INVX1    g23642(.A(new_n23834_), .Y(new_n23835_));
  OR2X1    g23643(.A(new_n23816_), .B(new_n14165_), .Y(new_n23836_));
  AND2X1   g23644(.A(new_n23800_), .B(new_n23791_), .Y(new_n23837_));
  INVX1    g23645(.A(new_n23806_), .Y(new_n23838_));
  NAND2X1  g23646(.A(new_n23782_), .B(new_n14165_), .Y(new_n23839_));
  OAI21X1  g23647(.A0(new_n23839_), .A1(new_n23837_), .B0(new_n23838_), .Y(new_n23840_));
  AOI21X1  g23648(.A0(new_n23840_), .A1(new_n23836_), .B0(new_n13571_), .Y(new_n23841_));
  AOI21X1  g23649(.A0(new_n23789_), .A1(\asqrt[17] ), .B0(\asqrt[18] ), .Y(new_n23842_));
  AOI21X1  g23650(.A0(new_n23842_), .A1(new_n23840_), .B0(new_n23813_), .Y(new_n23843_));
  OAI21X1  g23651(.A0(new_n23843_), .A1(new_n23841_), .B0(\asqrt[19] ), .Y(new_n23844_));
  NAND2X1  g23652(.A(new_n23844_), .B(new_n12447_), .Y(new_n23845_));
  OAI21X1  g23653(.A0(new_n23845_), .A1(new_n23829_), .B0(new_n23835_), .Y(new_n23846_));
  AOI21X1  g23654(.A0(new_n23846_), .A1(new_n23828_), .B0(new_n11896_), .Y(new_n23847_));
  NAND4X1  g23655(.A(\asqrt[3] ), .B(new_n23077_), .C(new_n23075_), .D(new_n23102_), .Y(new_n23848_));
  NAND2X1  g23656(.A(new_n23077_), .B(new_n23102_), .Y(new_n23849_));
  OAI21X1  g23657(.A0(new_n23849_), .A1(new_n23622_), .B0(new_n23076_), .Y(new_n23850_));
  AND2X1   g23658(.A(new_n23850_), .B(new_n23848_), .Y(new_n23851_));
  NOR3X1   g23659(.A(new_n23843_), .B(new_n23841_), .C(\asqrt[19] ), .Y(new_n23852_));
  OAI21X1  g23660(.A0(new_n23852_), .A1(new_n23824_), .B0(new_n23844_), .Y(new_n23853_));
  AOI21X1  g23661(.A0(new_n23853_), .A1(\asqrt[20] ), .B0(\asqrt[21] ), .Y(new_n23854_));
  AOI21X1  g23662(.A0(new_n23854_), .A1(new_n23846_), .B0(new_n23851_), .Y(new_n23855_));
  OAI21X1  g23663(.A0(new_n23855_), .A1(new_n23847_), .B0(\asqrt[22] ), .Y(new_n23856_));
  AND2X1   g23664(.A(new_n23119_), .B(new_n23118_), .Y(new_n23857_));
  NOR3X1   g23665(.A(new_n23857_), .B(new_n23085_), .C(new_n23117_), .Y(new_n23858_));
  NOR3X1   g23666(.A(new_n23622_), .B(new_n23857_), .C(new_n23117_), .Y(new_n23859_));
  NOR2X1   g23667(.A(new_n23859_), .B(new_n23084_), .Y(new_n23860_));
  AOI21X1  g23668(.A0(new_n23858_), .A1(\asqrt[3] ), .B0(new_n23860_), .Y(new_n23861_));
  NOR3X1   g23669(.A(new_n23855_), .B(new_n23847_), .C(\asqrt[22] ), .Y(new_n23862_));
  OAI21X1  g23670(.A0(new_n23862_), .A1(new_n23861_), .B0(new_n23856_), .Y(new_n23863_));
  AND2X1   g23671(.A(new_n23863_), .B(\asqrt[23] ), .Y(new_n23864_));
  INVX1    g23672(.A(new_n23861_), .Y(new_n23865_));
  AND2X1   g23673(.A(new_n23853_), .B(\asqrt[20] ), .Y(new_n23866_));
  NAND2X1  g23674(.A(new_n23826_), .B(new_n23825_), .Y(new_n23867_));
  AND2X1   g23675(.A(new_n23844_), .B(new_n12447_), .Y(new_n23868_));
  AOI21X1  g23676(.A0(new_n23868_), .A1(new_n23867_), .B0(new_n23834_), .Y(new_n23869_));
  OAI21X1  g23677(.A0(new_n23869_), .A1(new_n23866_), .B0(\asqrt[21] ), .Y(new_n23870_));
  INVX1    g23678(.A(new_n23851_), .Y(new_n23871_));
  OAI21X1  g23679(.A0(new_n23827_), .A1(new_n12447_), .B0(new_n11896_), .Y(new_n23872_));
  OAI21X1  g23680(.A0(new_n23872_), .A1(new_n23869_), .B0(new_n23871_), .Y(new_n23873_));
  NAND3X1  g23681(.A(new_n23873_), .B(new_n23870_), .C(new_n11362_), .Y(new_n23874_));
  NAND2X1  g23682(.A(new_n23874_), .B(new_n23865_), .Y(new_n23875_));
  AND2X1   g23683(.A(new_n23105_), .B(new_n23087_), .Y(new_n23876_));
  NOR3X1   g23684(.A(new_n23876_), .B(new_n23122_), .C(new_n23088_), .Y(new_n23877_));
  NOR3X1   g23685(.A(new_n23622_), .B(new_n23876_), .C(new_n23088_), .Y(new_n23878_));
  NOR2X1   g23686(.A(new_n23878_), .B(new_n23093_), .Y(new_n23879_));
  AOI21X1  g23687(.A0(new_n23877_), .A1(\asqrt[3] ), .B0(new_n23879_), .Y(new_n23880_));
  AND2X1   g23688(.A(new_n23856_), .B(new_n10849_), .Y(new_n23881_));
  AOI21X1  g23689(.A0(new_n23881_), .A1(new_n23875_), .B0(new_n23880_), .Y(new_n23882_));
  OAI21X1  g23690(.A0(new_n23882_), .A1(new_n23864_), .B0(\asqrt[24] ), .Y(new_n23883_));
  NAND4X1  g23691(.A(\asqrt[3] ), .B(new_n23125_), .C(new_n23112_), .D(new_n23107_), .Y(new_n23884_));
  NAND2X1  g23692(.A(new_n23125_), .B(new_n23107_), .Y(new_n23885_));
  OAI21X1  g23693(.A0(new_n23885_), .A1(new_n23622_), .B0(new_n23116_), .Y(new_n23886_));
  AND2X1   g23694(.A(new_n23886_), .B(new_n23884_), .Y(new_n23887_));
  INVX1    g23695(.A(new_n23887_), .Y(new_n23888_));
  AOI21X1  g23696(.A0(new_n23873_), .A1(new_n23870_), .B0(new_n11362_), .Y(new_n23889_));
  AOI21X1  g23697(.A0(new_n23874_), .A1(new_n23865_), .B0(new_n23889_), .Y(new_n23890_));
  OAI21X1  g23698(.A0(new_n23890_), .A1(new_n10849_), .B0(new_n10332_), .Y(new_n23891_));
  OAI21X1  g23699(.A0(new_n23891_), .A1(new_n23882_), .B0(new_n23888_), .Y(new_n23892_));
  AOI21X1  g23700(.A0(new_n23892_), .A1(new_n23883_), .B0(new_n9833_), .Y(new_n23893_));
  AOI21X1  g23701(.A0(new_n23132_), .A1(new_n23126_), .B0(new_n23170_), .Y(new_n23894_));
  AND2X1   g23702(.A(new_n23894_), .B(new_n23168_), .Y(new_n23895_));
  AOI22X1  g23703(.A0(new_n23132_), .A1(new_n23126_), .B0(new_n23114_), .B1(\asqrt[24] ), .Y(new_n23896_));
  AOI21X1  g23704(.A0(new_n23896_), .A1(\asqrt[3] ), .B0(new_n23130_), .Y(new_n23897_));
  AOI21X1  g23705(.A0(new_n23895_), .A1(\asqrt[3] ), .B0(new_n23897_), .Y(new_n23898_));
  INVX1    g23706(.A(new_n23898_), .Y(new_n23899_));
  NAND3X1  g23707(.A(new_n23892_), .B(new_n23883_), .C(new_n9833_), .Y(new_n23900_));
  AOI21X1  g23708(.A0(new_n23900_), .A1(new_n23899_), .B0(new_n23893_), .Y(new_n23901_));
  OR2X1    g23709(.A(new_n23901_), .B(new_n9353_), .Y(new_n23902_));
  AND2X1   g23710(.A(new_n23900_), .B(new_n23899_), .Y(new_n23903_));
  AND2X1   g23711(.A(new_n23174_), .B(new_n23172_), .Y(new_n23904_));
  NOR3X1   g23712(.A(new_n23904_), .B(new_n23140_), .C(new_n23173_), .Y(new_n23905_));
  NOR3X1   g23713(.A(new_n23622_), .B(new_n23904_), .C(new_n23173_), .Y(new_n23906_));
  NOR2X1   g23714(.A(new_n23906_), .B(new_n23139_), .Y(new_n23907_));
  AOI21X1  g23715(.A0(new_n23905_), .A1(\asqrt[3] ), .B0(new_n23907_), .Y(new_n23908_));
  INVX1    g23716(.A(new_n23908_), .Y(new_n23909_));
  OR2X1    g23717(.A(new_n23890_), .B(new_n10849_), .Y(new_n23910_));
  AND2X1   g23718(.A(new_n23874_), .B(new_n23865_), .Y(new_n23911_));
  INVX1    g23719(.A(new_n23880_), .Y(new_n23912_));
  NAND2X1  g23720(.A(new_n23856_), .B(new_n10849_), .Y(new_n23913_));
  OAI21X1  g23721(.A0(new_n23913_), .A1(new_n23911_), .B0(new_n23912_), .Y(new_n23914_));
  AOI21X1  g23722(.A0(new_n23914_), .A1(new_n23910_), .B0(new_n10332_), .Y(new_n23915_));
  AOI21X1  g23723(.A0(new_n23863_), .A1(\asqrt[23] ), .B0(\asqrt[24] ), .Y(new_n23916_));
  AOI21X1  g23724(.A0(new_n23916_), .A1(new_n23914_), .B0(new_n23887_), .Y(new_n23917_));
  OAI21X1  g23725(.A0(new_n23917_), .A1(new_n23915_), .B0(\asqrt[25] ), .Y(new_n23918_));
  NAND2X1  g23726(.A(new_n23918_), .B(new_n9353_), .Y(new_n23919_));
  OAI21X1  g23727(.A0(new_n23919_), .A1(new_n23903_), .B0(new_n23909_), .Y(new_n23920_));
  AOI21X1  g23728(.A0(new_n23920_), .A1(new_n23902_), .B0(new_n8874_), .Y(new_n23921_));
  NAND4X1  g23729(.A(\asqrt[3] ), .B(new_n23151_), .C(new_n23149_), .D(new_n23176_), .Y(new_n23922_));
  NAND2X1  g23730(.A(new_n23151_), .B(new_n23176_), .Y(new_n23923_));
  OAI21X1  g23731(.A0(new_n23923_), .A1(new_n23622_), .B0(new_n23150_), .Y(new_n23924_));
  AND2X1   g23732(.A(new_n23924_), .B(new_n23922_), .Y(new_n23925_));
  NOR3X1   g23733(.A(new_n23917_), .B(new_n23915_), .C(\asqrt[25] ), .Y(new_n23926_));
  OAI21X1  g23734(.A0(new_n23926_), .A1(new_n23898_), .B0(new_n23918_), .Y(new_n23927_));
  AOI21X1  g23735(.A0(new_n23927_), .A1(\asqrt[26] ), .B0(\asqrt[27] ), .Y(new_n23928_));
  AOI21X1  g23736(.A0(new_n23928_), .A1(new_n23920_), .B0(new_n23925_), .Y(new_n23929_));
  OAI21X1  g23737(.A0(new_n23929_), .A1(new_n23921_), .B0(\asqrt[28] ), .Y(new_n23930_));
  AND2X1   g23738(.A(new_n23193_), .B(new_n23192_), .Y(new_n23931_));
  NOR3X1   g23739(.A(new_n23931_), .B(new_n23159_), .C(new_n23191_), .Y(new_n23932_));
  NOR3X1   g23740(.A(new_n23622_), .B(new_n23931_), .C(new_n23191_), .Y(new_n23933_));
  NOR2X1   g23741(.A(new_n23933_), .B(new_n23158_), .Y(new_n23934_));
  AOI21X1  g23742(.A0(new_n23932_), .A1(\asqrt[3] ), .B0(new_n23934_), .Y(new_n23935_));
  NOR3X1   g23743(.A(new_n23929_), .B(new_n23921_), .C(\asqrt[28] ), .Y(new_n23936_));
  OAI21X1  g23744(.A0(new_n23936_), .A1(new_n23935_), .B0(new_n23930_), .Y(new_n23937_));
  AND2X1   g23745(.A(new_n23937_), .B(\asqrt[29] ), .Y(new_n23938_));
  INVX1    g23746(.A(new_n23935_), .Y(new_n23939_));
  AND2X1   g23747(.A(new_n23927_), .B(\asqrt[26] ), .Y(new_n23940_));
  NAND2X1  g23748(.A(new_n23900_), .B(new_n23899_), .Y(new_n23941_));
  AND2X1   g23749(.A(new_n23918_), .B(new_n9353_), .Y(new_n23942_));
  AOI21X1  g23750(.A0(new_n23942_), .A1(new_n23941_), .B0(new_n23908_), .Y(new_n23943_));
  OAI21X1  g23751(.A0(new_n23943_), .A1(new_n23940_), .B0(\asqrt[27] ), .Y(new_n23944_));
  INVX1    g23752(.A(new_n23925_), .Y(new_n23945_));
  OAI21X1  g23753(.A0(new_n23901_), .A1(new_n9353_), .B0(new_n8874_), .Y(new_n23946_));
  OAI21X1  g23754(.A0(new_n23946_), .A1(new_n23943_), .B0(new_n23945_), .Y(new_n23947_));
  NAND3X1  g23755(.A(new_n23947_), .B(new_n23944_), .C(new_n8412_), .Y(new_n23948_));
  NAND2X1  g23756(.A(new_n23948_), .B(new_n23939_), .Y(new_n23949_));
  AND2X1   g23757(.A(new_n23179_), .B(new_n23161_), .Y(new_n23950_));
  NOR3X1   g23758(.A(new_n23950_), .B(new_n23196_), .C(new_n23162_), .Y(new_n23951_));
  NOR3X1   g23759(.A(new_n23622_), .B(new_n23950_), .C(new_n23162_), .Y(new_n23952_));
  NOR2X1   g23760(.A(new_n23952_), .B(new_n23167_), .Y(new_n23953_));
  AOI21X1  g23761(.A0(new_n23951_), .A1(\asqrt[3] ), .B0(new_n23953_), .Y(new_n23954_));
  AND2X1   g23762(.A(new_n23930_), .B(new_n7970_), .Y(new_n23955_));
  AOI21X1  g23763(.A0(new_n23955_), .A1(new_n23949_), .B0(new_n23954_), .Y(new_n23956_));
  OAI21X1  g23764(.A0(new_n23956_), .A1(new_n23938_), .B0(\asqrt[30] ), .Y(new_n23957_));
  NAND4X1  g23765(.A(\asqrt[3] ), .B(new_n23199_), .C(new_n23186_), .D(new_n23181_), .Y(new_n23958_));
  NAND2X1  g23766(.A(new_n23199_), .B(new_n23181_), .Y(new_n23959_));
  OAI21X1  g23767(.A0(new_n23959_), .A1(new_n23622_), .B0(new_n23190_), .Y(new_n23960_));
  AND2X1   g23768(.A(new_n23960_), .B(new_n23958_), .Y(new_n23961_));
  INVX1    g23769(.A(new_n23961_), .Y(new_n23962_));
  AOI21X1  g23770(.A0(new_n23947_), .A1(new_n23944_), .B0(new_n8412_), .Y(new_n23963_));
  AOI21X1  g23771(.A0(new_n23948_), .A1(new_n23939_), .B0(new_n23963_), .Y(new_n23964_));
  OAI21X1  g23772(.A0(new_n23964_), .A1(new_n7970_), .B0(new_n7527_), .Y(new_n23965_));
  OAI21X1  g23773(.A0(new_n23965_), .A1(new_n23956_), .B0(new_n23962_), .Y(new_n23966_));
  AOI21X1  g23774(.A0(new_n23966_), .A1(new_n23957_), .B0(new_n7103_), .Y(new_n23967_));
  AOI21X1  g23775(.A0(new_n23206_), .A1(new_n23200_), .B0(new_n23244_), .Y(new_n23968_));
  AND2X1   g23776(.A(new_n23968_), .B(new_n23242_), .Y(new_n23969_));
  AOI22X1  g23777(.A0(new_n23206_), .A1(new_n23200_), .B0(new_n23188_), .B1(\asqrt[30] ), .Y(new_n23970_));
  AOI21X1  g23778(.A0(new_n23970_), .A1(\asqrt[3] ), .B0(new_n23204_), .Y(new_n23971_));
  AOI21X1  g23779(.A0(new_n23969_), .A1(\asqrt[3] ), .B0(new_n23971_), .Y(new_n23972_));
  INVX1    g23780(.A(new_n23972_), .Y(new_n23973_));
  NAND3X1  g23781(.A(new_n23966_), .B(new_n23957_), .C(new_n7103_), .Y(new_n23974_));
  AOI21X1  g23782(.A0(new_n23974_), .A1(new_n23973_), .B0(new_n23967_), .Y(new_n23975_));
  OR2X1    g23783(.A(new_n23975_), .B(new_n6699_), .Y(new_n23976_));
  AND2X1   g23784(.A(new_n23974_), .B(new_n23973_), .Y(new_n23977_));
  AND2X1   g23785(.A(new_n23248_), .B(new_n23246_), .Y(new_n23978_));
  NOR3X1   g23786(.A(new_n23978_), .B(new_n23214_), .C(new_n23247_), .Y(new_n23979_));
  NOR3X1   g23787(.A(new_n23622_), .B(new_n23978_), .C(new_n23247_), .Y(new_n23980_));
  NOR2X1   g23788(.A(new_n23980_), .B(new_n23213_), .Y(new_n23981_));
  AOI21X1  g23789(.A0(new_n23979_), .A1(\asqrt[3] ), .B0(new_n23981_), .Y(new_n23982_));
  INVX1    g23790(.A(new_n23982_), .Y(new_n23983_));
  OR2X1    g23791(.A(new_n23964_), .B(new_n7970_), .Y(new_n23984_));
  AND2X1   g23792(.A(new_n23948_), .B(new_n23939_), .Y(new_n23985_));
  INVX1    g23793(.A(new_n23954_), .Y(new_n23986_));
  NAND2X1  g23794(.A(new_n23930_), .B(new_n7970_), .Y(new_n23987_));
  OAI21X1  g23795(.A0(new_n23987_), .A1(new_n23985_), .B0(new_n23986_), .Y(new_n23988_));
  AOI21X1  g23796(.A0(new_n23988_), .A1(new_n23984_), .B0(new_n7527_), .Y(new_n23989_));
  AOI21X1  g23797(.A0(new_n23937_), .A1(\asqrt[29] ), .B0(\asqrt[30] ), .Y(new_n23990_));
  AOI21X1  g23798(.A0(new_n23990_), .A1(new_n23988_), .B0(new_n23961_), .Y(new_n23991_));
  OAI21X1  g23799(.A0(new_n23991_), .A1(new_n23989_), .B0(\asqrt[31] ), .Y(new_n23992_));
  NAND2X1  g23800(.A(new_n23992_), .B(new_n6699_), .Y(new_n23993_));
  OAI21X1  g23801(.A0(new_n23993_), .A1(new_n23977_), .B0(new_n23983_), .Y(new_n23994_));
  AOI21X1  g23802(.A0(new_n23994_), .A1(new_n23976_), .B0(new_n6294_), .Y(new_n23995_));
  NAND4X1  g23803(.A(\asqrt[3] ), .B(new_n23225_), .C(new_n23223_), .D(new_n23250_), .Y(new_n23996_));
  NAND2X1  g23804(.A(new_n23225_), .B(new_n23250_), .Y(new_n23997_));
  OAI21X1  g23805(.A0(new_n23997_), .A1(new_n23622_), .B0(new_n23224_), .Y(new_n23998_));
  AND2X1   g23806(.A(new_n23998_), .B(new_n23996_), .Y(new_n23999_));
  NOR3X1   g23807(.A(new_n23991_), .B(new_n23989_), .C(\asqrt[31] ), .Y(new_n24000_));
  OAI21X1  g23808(.A0(new_n24000_), .A1(new_n23972_), .B0(new_n23992_), .Y(new_n24001_));
  AOI21X1  g23809(.A0(new_n24001_), .A1(\asqrt[32] ), .B0(\asqrt[33] ), .Y(new_n24002_));
  AOI21X1  g23810(.A0(new_n24002_), .A1(new_n23994_), .B0(new_n23999_), .Y(new_n24003_));
  OAI21X1  g23811(.A0(new_n24003_), .A1(new_n23995_), .B0(\asqrt[34] ), .Y(new_n24004_));
  AND2X1   g23812(.A(new_n23280_), .B(new_n23279_), .Y(new_n24005_));
  NOR3X1   g23813(.A(new_n24005_), .B(new_n23233_), .C(new_n23278_), .Y(new_n24006_));
  NOR3X1   g23814(.A(new_n23622_), .B(new_n24005_), .C(new_n23278_), .Y(new_n24007_));
  NOR2X1   g23815(.A(new_n24007_), .B(new_n23232_), .Y(new_n24008_));
  AOI21X1  g23816(.A0(new_n24006_), .A1(\asqrt[3] ), .B0(new_n24008_), .Y(new_n24009_));
  NOR3X1   g23817(.A(new_n24003_), .B(new_n23995_), .C(\asqrt[34] ), .Y(new_n24010_));
  OAI21X1  g23818(.A0(new_n24010_), .A1(new_n24009_), .B0(new_n24004_), .Y(new_n24011_));
  AND2X1   g23819(.A(new_n24011_), .B(\asqrt[35] ), .Y(new_n24012_));
  INVX1    g23820(.A(new_n24009_), .Y(new_n24013_));
  AND2X1   g23821(.A(new_n24001_), .B(\asqrt[32] ), .Y(new_n24014_));
  NAND2X1  g23822(.A(new_n23974_), .B(new_n23973_), .Y(new_n24015_));
  AND2X1   g23823(.A(new_n23992_), .B(new_n6699_), .Y(new_n24016_));
  AOI21X1  g23824(.A0(new_n24016_), .A1(new_n24015_), .B0(new_n23982_), .Y(new_n24017_));
  OAI21X1  g23825(.A0(new_n24017_), .A1(new_n24014_), .B0(\asqrt[33] ), .Y(new_n24018_));
  INVX1    g23826(.A(new_n23999_), .Y(new_n24019_));
  OAI21X1  g23827(.A0(new_n23975_), .A1(new_n6699_), .B0(new_n6294_), .Y(new_n24020_));
  OAI21X1  g23828(.A0(new_n24020_), .A1(new_n24017_), .B0(new_n24019_), .Y(new_n24021_));
  NAND3X1  g23829(.A(new_n24021_), .B(new_n24018_), .C(new_n5941_), .Y(new_n24022_));
  NAND2X1  g23830(.A(new_n24022_), .B(new_n24013_), .Y(new_n24023_));
  AND2X1   g23831(.A(new_n23253_), .B(new_n23235_), .Y(new_n24024_));
  NOR3X1   g23832(.A(new_n24024_), .B(new_n23283_), .C(new_n23236_), .Y(new_n24025_));
  NOR3X1   g23833(.A(new_n23622_), .B(new_n24024_), .C(new_n23236_), .Y(new_n24026_));
  NOR2X1   g23834(.A(new_n24026_), .B(new_n23241_), .Y(new_n24027_));
  AOI21X1  g23835(.A0(new_n24025_), .A1(\asqrt[3] ), .B0(new_n24027_), .Y(new_n24028_));
  AND2X1   g23836(.A(new_n24004_), .B(new_n5541_), .Y(new_n24029_));
  AOI21X1  g23837(.A0(new_n24029_), .A1(new_n24023_), .B0(new_n24028_), .Y(new_n24030_));
  OAI21X1  g23838(.A0(new_n24030_), .A1(new_n24012_), .B0(\asqrt[36] ), .Y(new_n24031_));
  NAND4X1  g23839(.A(\asqrt[3] ), .B(new_n23288_), .C(new_n23260_), .D(new_n23255_), .Y(new_n24032_));
  OR2X1    g23840(.A(new_n23261_), .B(new_n23286_), .Y(new_n24033_));
  OAI21X1  g23841(.A0(new_n24033_), .A1(new_n23622_), .B0(new_n23287_), .Y(new_n24034_));
  AND2X1   g23842(.A(new_n24034_), .B(new_n24032_), .Y(new_n24035_));
  INVX1    g23843(.A(new_n24035_), .Y(new_n24036_));
  AOI21X1  g23844(.A0(new_n24021_), .A1(new_n24018_), .B0(new_n5941_), .Y(new_n24037_));
  AOI21X1  g23845(.A0(new_n24022_), .A1(new_n24013_), .B0(new_n24037_), .Y(new_n24038_));
  OAI21X1  g23846(.A0(new_n24038_), .A1(new_n5541_), .B0(new_n5176_), .Y(new_n24039_));
  OAI21X1  g23847(.A0(new_n24039_), .A1(new_n24030_), .B0(new_n24036_), .Y(new_n24040_));
  AOI21X1  g23848(.A0(new_n24040_), .A1(new_n24031_), .B0(new_n4826_), .Y(new_n24041_));
  AOI21X1  g23849(.A0(new_n23269_), .A1(new_n23264_), .B0(new_n23304_), .Y(new_n24042_));
  AND2X1   g23850(.A(new_n24042_), .B(new_n23302_), .Y(new_n24043_));
  AOI22X1  g23851(.A0(new_n23269_), .A1(new_n23264_), .B0(new_n23262_), .B1(\asqrt[36] ), .Y(new_n24044_));
  AOI21X1  g23852(.A0(new_n24044_), .A1(\asqrt[3] ), .B0(new_n23268_), .Y(new_n24045_));
  AOI21X1  g23853(.A0(new_n24043_), .A1(\asqrt[3] ), .B0(new_n24045_), .Y(new_n24046_));
  INVX1    g23854(.A(new_n24046_), .Y(new_n24047_));
  NAND3X1  g23855(.A(new_n24040_), .B(new_n24031_), .C(new_n4826_), .Y(new_n24048_));
  AOI21X1  g23856(.A0(new_n24048_), .A1(new_n24047_), .B0(new_n24041_), .Y(new_n24049_));
  OR2X1    g23857(.A(new_n24049_), .B(new_n4493_), .Y(new_n24050_));
  OR2X1    g23858(.A(new_n24038_), .B(new_n5541_), .Y(new_n24051_));
  AND2X1   g23859(.A(new_n24022_), .B(new_n24013_), .Y(new_n24052_));
  INVX1    g23860(.A(new_n24028_), .Y(new_n24053_));
  NAND2X1  g23861(.A(new_n24004_), .B(new_n5541_), .Y(new_n24054_));
  OAI21X1  g23862(.A0(new_n24054_), .A1(new_n24052_), .B0(new_n24053_), .Y(new_n24055_));
  AOI21X1  g23863(.A0(new_n24055_), .A1(new_n24051_), .B0(new_n5176_), .Y(new_n24056_));
  AOI21X1  g23864(.A0(new_n24011_), .A1(\asqrt[35] ), .B0(\asqrt[36] ), .Y(new_n24057_));
  AOI21X1  g23865(.A0(new_n24057_), .A1(new_n24055_), .B0(new_n24035_), .Y(new_n24058_));
  NOR3X1   g23866(.A(new_n24058_), .B(new_n24056_), .C(\asqrt[37] ), .Y(new_n24059_));
  NOR2X1   g23867(.A(new_n24059_), .B(new_n24046_), .Y(new_n24060_));
  AND2X1   g23868(.A(new_n23308_), .B(new_n23306_), .Y(new_n24061_));
  NOR3X1   g23869(.A(new_n24061_), .B(new_n23277_), .C(new_n23307_), .Y(new_n24062_));
  NOR3X1   g23870(.A(new_n23622_), .B(new_n24061_), .C(new_n23307_), .Y(new_n24063_));
  NOR2X1   g23871(.A(new_n24063_), .B(new_n23276_), .Y(new_n24064_));
  AOI21X1  g23872(.A0(new_n24062_), .A1(\asqrt[3] ), .B0(new_n24064_), .Y(new_n24065_));
  INVX1    g23873(.A(new_n24065_), .Y(new_n24066_));
  OAI21X1  g23874(.A0(new_n24058_), .A1(new_n24056_), .B0(\asqrt[37] ), .Y(new_n24067_));
  NAND2X1  g23875(.A(new_n24067_), .B(new_n4493_), .Y(new_n24068_));
  OAI21X1  g23876(.A0(new_n24068_), .A1(new_n24060_), .B0(new_n24066_), .Y(new_n24069_));
  AOI21X1  g23877(.A0(new_n24069_), .A1(new_n24050_), .B0(new_n4165_), .Y(new_n24070_));
  NAND4X1  g23878(.A(\asqrt[3] ), .B(new_n23299_), .C(new_n23297_), .D(new_n23317_), .Y(new_n24071_));
  OR2X1    g23879(.A(new_n23310_), .B(new_n23292_), .Y(new_n24072_));
  OAI21X1  g23880(.A0(new_n24072_), .A1(new_n23622_), .B0(new_n23298_), .Y(new_n24073_));
  AND2X1   g23881(.A(new_n24073_), .B(new_n24071_), .Y(new_n24074_));
  OAI21X1  g23882(.A0(new_n24059_), .A1(new_n24046_), .B0(new_n24067_), .Y(new_n24075_));
  AOI21X1  g23883(.A0(new_n24075_), .A1(\asqrt[38] ), .B0(\asqrt[39] ), .Y(new_n24076_));
  AOI21X1  g23884(.A0(new_n24076_), .A1(new_n24069_), .B0(new_n24074_), .Y(new_n24077_));
  OAI21X1  g23885(.A0(new_n24077_), .A1(new_n24070_), .B0(\asqrt[40] ), .Y(new_n24078_));
  AND2X1   g23886(.A(new_n23354_), .B(new_n23353_), .Y(new_n24079_));
  NOR3X1   g23887(.A(new_n24079_), .B(new_n23316_), .C(new_n23352_), .Y(new_n24080_));
  NOR3X1   g23888(.A(new_n23622_), .B(new_n24079_), .C(new_n23352_), .Y(new_n24081_));
  NOR2X1   g23889(.A(new_n24081_), .B(new_n23315_), .Y(new_n24082_));
  AOI21X1  g23890(.A0(new_n24080_), .A1(\asqrt[3] ), .B0(new_n24082_), .Y(new_n24083_));
  NOR3X1   g23891(.A(new_n24077_), .B(new_n24070_), .C(\asqrt[40] ), .Y(new_n24084_));
  OAI21X1  g23892(.A0(new_n24084_), .A1(new_n24083_), .B0(new_n24078_), .Y(new_n24085_));
  AND2X1   g23893(.A(new_n24085_), .B(\asqrt[41] ), .Y(new_n24086_));
  OR2X1    g23894(.A(new_n24084_), .B(new_n24083_), .Y(new_n24087_));
  AND2X1   g23895(.A(new_n23327_), .B(new_n23319_), .Y(new_n24088_));
  NOR3X1   g23896(.A(new_n24088_), .B(new_n23357_), .C(new_n23320_), .Y(new_n24089_));
  NOR3X1   g23897(.A(new_n23622_), .B(new_n24088_), .C(new_n23320_), .Y(new_n24090_));
  NOR2X1   g23898(.A(new_n24090_), .B(new_n23325_), .Y(new_n24091_));
  AOI21X1  g23899(.A0(new_n24089_), .A1(\asqrt[3] ), .B0(new_n24091_), .Y(new_n24092_));
  AND2X1   g23900(.A(new_n24078_), .B(new_n3564_), .Y(new_n24093_));
  AOI21X1  g23901(.A0(new_n24093_), .A1(new_n24087_), .B0(new_n24092_), .Y(new_n24094_));
  OAI21X1  g23902(.A0(new_n24094_), .A1(new_n24086_), .B0(\asqrt[42] ), .Y(new_n24095_));
  NAND4X1  g23903(.A(\asqrt[3] ), .B(new_n23362_), .C(new_n23334_), .D(new_n23329_), .Y(new_n24096_));
  OR2X1    g23904(.A(new_n23335_), .B(new_n23360_), .Y(new_n24097_));
  OAI21X1  g23905(.A0(new_n24097_), .A1(new_n23622_), .B0(new_n23361_), .Y(new_n24098_));
  AND2X1   g23906(.A(new_n24098_), .B(new_n24096_), .Y(new_n24099_));
  INVX1    g23907(.A(new_n24099_), .Y(new_n24100_));
  AND2X1   g23908(.A(new_n24075_), .B(\asqrt[38] ), .Y(new_n24101_));
  OR2X1    g23909(.A(new_n24059_), .B(new_n24046_), .Y(new_n24102_));
  AND2X1   g23910(.A(new_n24067_), .B(new_n4493_), .Y(new_n24103_));
  AOI21X1  g23911(.A0(new_n24103_), .A1(new_n24102_), .B0(new_n24065_), .Y(new_n24104_));
  OAI21X1  g23912(.A0(new_n24104_), .A1(new_n24101_), .B0(\asqrt[39] ), .Y(new_n24105_));
  INVX1    g23913(.A(new_n24074_), .Y(new_n24106_));
  OAI21X1  g23914(.A0(new_n24049_), .A1(new_n4493_), .B0(new_n4165_), .Y(new_n24107_));
  OAI21X1  g23915(.A0(new_n24107_), .A1(new_n24104_), .B0(new_n24106_), .Y(new_n24108_));
  AOI21X1  g23916(.A0(new_n24108_), .A1(new_n24105_), .B0(new_n3863_), .Y(new_n24109_));
  INVX1    g23917(.A(new_n24083_), .Y(new_n24110_));
  NAND3X1  g23918(.A(new_n24108_), .B(new_n24105_), .C(new_n3863_), .Y(new_n24111_));
  AOI21X1  g23919(.A0(new_n24111_), .A1(new_n24110_), .B0(new_n24109_), .Y(new_n24112_));
  OAI21X1  g23920(.A0(new_n24112_), .A1(new_n3564_), .B0(new_n3276_), .Y(new_n24113_));
  OAI21X1  g23921(.A0(new_n24113_), .A1(new_n24094_), .B0(new_n24100_), .Y(new_n24114_));
  AOI21X1  g23922(.A0(new_n24114_), .A1(new_n24095_), .B0(new_n3008_), .Y(new_n24115_));
  AOI21X1  g23923(.A0(new_n23343_), .A1(new_n23338_), .B0(new_n23378_), .Y(new_n24116_));
  AND2X1   g23924(.A(new_n24116_), .B(new_n23376_), .Y(new_n24117_));
  AOI22X1  g23925(.A0(new_n23343_), .A1(new_n23338_), .B0(new_n23336_), .B1(\asqrt[42] ), .Y(new_n24118_));
  AOI21X1  g23926(.A0(new_n24118_), .A1(\asqrt[3] ), .B0(new_n23342_), .Y(new_n24119_));
  AOI21X1  g23927(.A0(new_n24117_), .A1(\asqrt[3] ), .B0(new_n24119_), .Y(new_n24120_));
  INVX1    g23928(.A(new_n24120_), .Y(new_n24121_));
  NAND3X1  g23929(.A(new_n24114_), .B(new_n24095_), .C(new_n3008_), .Y(new_n24122_));
  AOI21X1  g23930(.A0(new_n24122_), .A1(new_n24121_), .B0(new_n24115_), .Y(new_n24123_));
  OR2X1    g23931(.A(new_n24123_), .B(new_n2769_), .Y(new_n24124_));
  OR2X1    g23932(.A(new_n24112_), .B(new_n3564_), .Y(new_n24125_));
  NOR2X1   g23933(.A(new_n24084_), .B(new_n24083_), .Y(new_n24126_));
  INVX1    g23934(.A(new_n24092_), .Y(new_n24127_));
  NAND2X1  g23935(.A(new_n24078_), .B(new_n3564_), .Y(new_n24128_));
  OAI21X1  g23936(.A0(new_n24128_), .A1(new_n24126_), .B0(new_n24127_), .Y(new_n24129_));
  AOI21X1  g23937(.A0(new_n24129_), .A1(new_n24125_), .B0(new_n3276_), .Y(new_n24130_));
  AOI21X1  g23938(.A0(new_n24085_), .A1(\asqrt[41] ), .B0(\asqrt[42] ), .Y(new_n24131_));
  AOI21X1  g23939(.A0(new_n24131_), .A1(new_n24129_), .B0(new_n24099_), .Y(new_n24132_));
  NOR3X1   g23940(.A(new_n24132_), .B(new_n24130_), .C(\asqrt[43] ), .Y(new_n24133_));
  NOR2X1   g23941(.A(new_n24133_), .B(new_n24120_), .Y(new_n24134_));
  AND2X1   g23942(.A(new_n23382_), .B(new_n23380_), .Y(new_n24135_));
  NOR3X1   g23943(.A(new_n24135_), .B(new_n23351_), .C(new_n23381_), .Y(new_n24136_));
  NOR3X1   g23944(.A(new_n23622_), .B(new_n24135_), .C(new_n23381_), .Y(new_n24137_));
  NOR2X1   g23945(.A(new_n24137_), .B(new_n23350_), .Y(new_n24138_));
  AOI21X1  g23946(.A0(new_n24136_), .A1(\asqrt[3] ), .B0(new_n24138_), .Y(new_n24139_));
  INVX1    g23947(.A(new_n24139_), .Y(new_n24140_));
  OAI21X1  g23948(.A0(new_n24132_), .A1(new_n24130_), .B0(\asqrt[43] ), .Y(new_n24141_));
  NAND2X1  g23949(.A(new_n24141_), .B(new_n2769_), .Y(new_n24142_));
  OAI21X1  g23950(.A0(new_n24142_), .A1(new_n24134_), .B0(new_n24140_), .Y(new_n24143_));
  AOI21X1  g23951(.A0(new_n24143_), .A1(new_n24124_), .B0(new_n2570_), .Y(new_n24144_));
  NAND4X1  g23952(.A(\asqrt[3] ), .B(new_n23373_), .C(new_n23371_), .D(new_n23391_), .Y(new_n24145_));
  OR2X1    g23953(.A(new_n23384_), .B(new_n23366_), .Y(new_n24146_));
  OAI21X1  g23954(.A0(new_n24146_), .A1(new_n23622_), .B0(new_n23372_), .Y(new_n24147_));
  AND2X1   g23955(.A(new_n24147_), .B(new_n24145_), .Y(new_n24148_));
  OAI21X1  g23956(.A0(new_n24133_), .A1(new_n24120_), .B0(new_n24141_), .Y(new_n24149_));
  AOI21X1  g23957(.A0(new_n24149_), .A1(\asqrt[44] ), .B0(\asqrt[45] ), .Y(new_n24150_));
  AOI21X1  g23958(.A0(new_n24150_), .A1(new_n24143_), .B0(new_n24148_), .Y(new_n24151_));
  OAI21X1  g23959(.A0(new_n24151_), .A1(new_n24144_), .B0(\asqrt[46] ), .Y(new_n24152_));
  AND2X1   g23960(.A(new_n23428_), .B(new_n23427_), .Y(new_n24153_));
  NOR3X1   g23961(.A(new_n24153_), .B(new_n23390_), .C(new_n23426_), .Y(new_n24154_));
  NOR3X1   g23962(.A(new_n23622_), .B(new_n24153_), .C(new_n23426_), .Y(new_n24155_));
  NOR2X1   g23963(.A(new_n24155_), .B(new_n23389_), .Y(new_n24156_));
  AOI21X1  g23964(.A0(new_n24154_), .A1(\asqrt[3] ), .B0(new_n24156_), .Y(new_n24157_));
  NOR3X1   g23965(.A(new_n24151_), .B(new_n24144_), .C(\asqrt[46] ), .Y(new_n24158_));
  OAI21X1  g23966(.A0(new_n24158_), .A1(new_n24157_), .B0(new_n24152_), .Y(new_n24159_));
  AND2X1   g23967(.A(new_n24159_), .B(\asqrt[47] ), .Y(new_n24160_));
  OR2X1    g23968(.A(new_n24158_), .B(new_n24157_), .Y(new_n24161_));
  AND2X1   g23969(.A(new_n23401_), .B(new_n23393_), .Y(new_n24162_));
  NOR3X1   g23970(.A(new_n24162_), .B(new_n23431_), .C(new_n23394_), .Y(new_n24163_));
  NOR3X1   g23971(.A(new_n23622_), .B(new_n24162_), .C(new_n23394_), .Y(new_n24164_));
  NOR2X1   g23972(.A(new_n24164_), .B(new_n23399_), .Y(new_n24165_));
  AOI21X1  g23973(.A0(new_n24163_), .A1(\asqrt[3] ), .B0(new_n24165_), .Y(new_n24166_));
  AND2X1   g23974(.A(new_n24152_), .B(new_n2040_), .Y(new_n24167_));
  AOI21X1  g23975(.A0(new_n24167_), .A1(new_n24161_), .B0(new_n24166_), .Y(new_n24168_));
  OAI21X1  g23976(.A0(new_n24168_), .A1(new_n24160_), .B0(\asqrt[48] ), .Y(new_n24169_));
  OR4X1    g23977(.A(new_n23622_), .B(new_n23409_), .C(new_n23435_), .D(new_n23434_), .Y(new_n24170_));
  OR2X1    g23978(.A(new_n23409_), .B(new_n23434_), .Y(new_n24171_));
  OAI21X1  g23979(.A0(new_n24171_), .A1(new_n23622_), .B0(new_n23435_), .Y(new_n24172_));
  AND2X1   g23980(.A(new_n24172_), .B(new_n24170_), .Y(new_n24173_));
  INVX1    g23981(.A(new_n24173_), .Y(new_n24174_));
  AND2X1   g23982(.A(new_n24149_), .B(\asqrt[44] ), .Y(new_n24175_));
  OR2X1    g23983(.A(new_n24133_), .B(new_n24120_), .Y(new_n24176_));
  AND2X1   g23984(.A(new_n24141_), .B(new_n2769_), .Y(new_n24177_));
  AOI21X1  g23985(.A0(new_n24177_), .A1(new_n24176_), .B0(new_n24139_), .Y(new_n24178_));
  OAI21X1  g23986(.A0(new_n24178_), .A1(new_n24175_), .B0(\asqrt[45] ), .Y(new_n24179_));
  INVX1    g23987(.A(new_n24148_), .Y(new_n24180_));
  OAI21X1  g23988(.A0(new_n24123_), .A1(new_n2769_), .B0(new_n2570_), .Y(new_n24181_));
  OAI21X1  g23989(.A0(new_n24181_), .A1(new_n24178_), .B0(new_n24180_), .Y(new_n24182_));
  AOI21X1  g23990(.A0(new_n24182_), .A1(new_n24179_), .B0(new_n2263_), .Y(new_n24183_));
  INVX1    g23991(.A(new_n24157_), .Y(new_n24184_));
  NAND3X1  g23992(.A(new_n24182_), .B(new_n24179_), .C(new_n2263_), .Y(new_n24185_));
  AOI21X1  g23993(.A0(new_n24185_), .A1(new_n24184_), .B0(new_n24183_), .Y(new_n24186_));
  OAI21X1  g23994(.A0(new_n24186_), .A1(new_n2040_), .B0(new_n1834_), .Y(new_n24187_));
  OAI21X1  g23995(.A0(new_n24187_), .A1(new_n24168_), .B0(new_n24174_), .Y(new_n24188_));
  AOI21X1  g23996(.A0(new_n24188_), .A1(new_n24169_), .B0(new_n1632_), .Y(new_n24189_));
  AOI21X1  g23997(.A0(new_n23417_), .A1(new_n23412_), .B0(new_n23452_), .Y(new_n24190_));
  AND2X1   g23998(.A(new_n24190_), .B(new_n23450_), .Y(new_n24191_));
  AOI22X1  g23999(.A0(new_n23417_), .A1(new_n23412_), .B0(new_n23410_), .B1(\asqrt[48] ), .Y(new_n24192_));
  AOI21X1  g24000(.A0(new_n24192_), .A1(\asqrt[3] ), .B0(new_n23416_), .Y(new_n24193_));
  AOI21X1  g24001(.A0(new_n24191_), .A1(\asqrt[3] ), .B0(new_n24193_), .Y(new_n24194_));
  INVX1    g24002(.A(new_n24194_), .Y(new_n24195_));
  NAND3X1  g24003(.A(new_n24188_), .B(new_n24169_), .C(new_n1632_), .Y(new_n24196_));
  AOI21X1  g24004(.A0(new_n24196_), .A1(new_n24195_), .B0(new_n24189_), .Y(new_n24197_));
  OR2X1    g24005(.A(new_n24197_), .B(new_n1469_), .Y(new_n24198_));
  OR2X1    g24006(.A(new_n24186_), .B(new_n2040_), .Y(new_n24199_));
  NOR2X1   g24007(.A(new_n24158_), .B(new_n24157_), .Y(new_n24200_));
  INVX1    g24008(.A(new_n24166_), .Y(new_n24201_));
  NAND2X1  g24009(.A(new_n24152_), .B(new_n2040_), .Y(new_n24202_));
  OAI21X1  g24010(.A0(new_n24202_), .A1(new_n24200_), .B0(new_n24201_), .Y(new_n24203_));
  AOI21X1  g24011(.A0(new_n24203_), .A1(new_n24199_), .B0(new_n1834_), .Y(new_n24204_));
  AOI21X1  g24012(.A0(new_n24159_), .A1(\asqrt[47] ), .B0(\asqrt[48] ), .Y(new_n24205_));
  AOI21X1  g24013(.A0(new_n24205_), .A1(new_n24203_), .B0(new_n24173_), .Y(new_n24206_));
  NOR3X1   g24014(.A(new_n24206_), .B(new_n24204_), .C(\asqrt[49] ), .Y(new_n24207_));
  NOR2X1   g24015(.A(new_n24207_), .B(new_n24194_), .Y(new_n24208_));
  AND2X1   g24016(.A(new_n23456_), .B(new_n23454_), .Y(new_n24209_));
  NOR3X1   g24017(.A(new_n24209_), .B(new_n23425_), .C(new_n23455_), .Y(new_n24210_));
  NOR3X1   g24018(.A(new_n23622_), .B(new_n24209_), .C(new_n23455_), .Y(new_n24211_));
  NOR2X1   g24019(.A(new_n24211_), .B(new_n23424_), .Y(new_n24212_));
  AOI21X1  g24020(.A0(new_n24210_), .A1(\asqrt[3] ), .B0(new_n24212_), .Y(new_n24213_));
  INVX1    g24021(.A(new_n24213_), .Y(new_n24214_));
  OAI21X1  g24022(.A0(new_n24206_), .A1(new_n24204_), .B0(\asqrt[49] ), .Y(new_n24215_));
  NAND2X1  g24023(.A(new_n24215_), .B(new_n1469_), .Y(new_n24216_));
  OAI21X1  g24024(.A0(new_n24216_), .A1(new_n24208_), .B0(new_n24214_), .Y(new_n24217_));
  AOI21X1  g24025(.A0(new_n24217_), .A1(new_n24198_), .B0(new_n1277_), .Y(new_n24218_));
  OR4X1    g24026(.A(new_n23622_), .B(new_n23458_), .C(new_n23446_), .D(new_n23440_), .Y(new_n24219_));
  OR2X1    g24027(.A(new_n23458_), .B(new_n23440_), .Y(new_n24220_));
  OAI21X1  g24028(.A0(new_n24220_), .A1(new_n23622_), .B0(new_n23446_), .Y(new_n24221_));
  AND2X1   g24029(.A(new_n24221_), .B(new_n24219_), .Y(new_n24222_));
  OAI21X1  g24030(.A0(new_n24207_), .A1(new_n24194_), .B0(new_n24215_), .Y(new_n24223_));
  AOI21X1  g24031(.A0(new_n24223_), .A1(\asqrt[50] ), .B0(\asqrt[51] ), .Y(new_n24224_));
  AOI21X1  g24032(.A0(new_n24224_), .A1(new_n24217_), .B0(new_n24222_), .Y(new_n24225_));
  OAI21X1  g24033(.A0(new_n24225_), .A1(new_n24218_), .B0(\asqrt[52] ), .Y(new_n24226_));
  AND2X1   g24034(.A(new_n23502_), .B(new_n23501_), .Y(new_n24227_));
  NOR3X1   g24035(.A(new_n24227_), .B(new_n23464_), .C(new_n23500_), .Y(new_n24228_));
  NOR3X1   g24036(.A(new_n23622_), .B(new_n24227_), .C(new_n23500_), .Y(new_n24229_));
  NOR2X1   g24037(.A(new_n24229_), .B(new_n23463_), .Y(new_n24230_));
  AOI21X1  g24038(.A0(new_n24228_), .A1(\asqrt[3] ), .B0(new_n24230_), .Y(new_n24231_));
  NOR3X1   g24039(.A(new_n24225_), .B(new_n24218_), .C(\asqrt[52] ), .Y(new_n24232_));
  OAI21X1  g24040(.A0(new_n24232_), .A1(new_n24231_), .B0(new_n24226_), .Y(new_n24233_));
  AND2X1   g24041(.A(new_n24233_), .B(\asqrt[53] ), .Y(new_n24234_));
  OR2X1    g24042(.A(new_n24232_), .B(new_n24231_), .Y(new_n24235_));
  AND2X1   g24043(.A(new_n23475_), .B(new_n23467_), .Y(new_n24236_));
  NOR3X1   g24044(.A(new_n24236_), .B(new_n23505_), .C(new_n23468_), .Y(new_n24237_));
  NOR3X1   g24045(.A(new_n23622_), .B(new_n24236_), .C(new_n23468_), .Y(new_n24238_));
  NOR2X1   g24046(.A(new_n24238_), .B(new_n23473_), .Y(new_n24239_));
  AOI21X1  g24047(.A0(new_n24237_), .A1(\asqrt[3] ), .B0(new_n24239_), .Y(new_n24240_));
  AND2X1   g24048(.A(new_n24226_), .B(new_n968_), .Y(new_n24241_));
  AOI21X1  g24049(.A0(new_n24241_), .A1(new_n24235_), .B0(new_n24240_), .Y(new_n24242_));
  OAI21X1  g24050(.A0(new_n24242_), .A1(new_n24234_), .B0(\asqrt[54] ), .Y(new_n24243_));
  OR4X1    g24051(.A(new_n23622_), .B(new_n23483_), .C(new_n23509_), .D(new_n23508_), .Y(new_n24244_));
  OR2X1    g24052(.A(new_n23483_), .B(new_n23508_), .Y(new_n24245_));
  OAI21X1  g24053(.A0(new_n24245_), .A1(new_n23622_), .B0(new_n23509_), .Y(new_n24246_));
  AND2X1   g24054(.A(new_n24246_), .B(new_n24244_), .Y(new_n24247_));
  INVX1    g24055(.A(new_n24247_), .Y(new_n24248_));
  AND2X1   g24056(.A(new_n24223_), .B(\asqrt[50] ), .Y(new_n24249_));
  OR2X1    g24057(.A(new_n24207_), .B(new_n24194_), .Y(new_n24250_));
  AND2X1   g24058(.A(new_n24215_), .B(new_n1469_), .Y(new_n24251_));
  AOI21X1  g24059(.A0(new_n24251_), .A1(new_n24250_), .B0(new_n24213_), .Y(new_n24252_));
  OAI21X1  g24060(.A0(new_n24252_), .A1(new_n24249_), .B0(\asqrt[51] ), .Y(new_n24253_));
  INVX1    g24061(.A(new_n24222_), .Y(new_n24254_));
  OAI21X1  g24062(.A0(new_n24197_), .A1(new_n1469_), .B0(new_n1277_), .Y(new_n24255_));
  OAI21X1  g24063(.A0(new_n24255_), .A1(new_n24252_), .B0(new_n24254_), .Y(new_n24256_));
  AOI21X1  g24064(.A0(new_n24256_), .A1(new_n24253_), .B0(new_n1111_), .Y(new_n24257_));
  INVX1    g24065(.A(new_n24231_), .Y(new_n24258_));
  NAND3X1  g24066(.A(new_n24256_), .B(new_n24253_), .C(new_n1111_), .Y(new_n24259_));
  AOI21X1  g24067(.A0(new_n24259_), .A1(new_n24258_), .B0(new_n24257_), .Y(new_n24260_));
  OAI21X1  g24068(.A0(new_n24260_), .A1(new_n968_), .B0(new_n902_), .Y(new_n24261_));
  OAI21X1  g24069(.A0(new_n24261_), .A1(new_n24242_), .B0(new_n24248_), .Y(new_n24262_));
  AOI21X1  g24070(.A0(new_n24262_), .A1(new_n24243_), .B0(new_n697_), .Y(new_n24263_));
  AOI21X1  g24071(.A0(new_n23491_), .A1(new_n23486_), .B0(new_n23526_), .Y(new_n24264_));
  AND2X1   g24072(.A(new_n24264_), .B(new_n23524_), .Y(new_n24265_));
  AOI22X1  g24073(.A0(new_n23491_), .A1(new_n23486_), .B0(new_n23484_), .B1(\asqrt[54] ), .Y(new_n24266_));
  AOI21X1  g24074(.A0(new_n24266_), .A1(\asqrt[3] ), .B0(new_n23490_), .Y(new_n24267_));
  AOI21X1  g24075(.A0(new_n24265_), .A1(\asqrt[3] ), .B0(new_n24267_), .Y(new_n24268_));
  INVX1    g24076(.A(new_n24268_), .Y(new_n24269_));
  NAND3X1  g24077(.A(new_n24262_), .B(new_n24243_), .C(new_n697_), .Y(new_n24270_));
  AOI21X1  g24078(.A0(new_n24270_), .A1(new_n24269_), .B0(new_n24263_), .Y(new_n24271_));
  OR2X1    g24079(.A(new_n24271_), .B(new_n582_), .Y(new_n24272_));
  OR2X1    g24080(.A(new_n24260_), .B(new_n968_), .Y(new_n24273_));
  NOR2X1   g24081(.A(new_n24232_), .B(new_n24231_), .Y(new_n24274_));
  INVX1    g24082(.A(new_n24240_), .Y(new_n24275_));
  NAND2X1  g24083(.A(new_n24226_), .B(new_n968_), .Y(new_n24276_));
  OAI21X1  g24084(.A0(new_n24276_), .A1(new_n24274_), .B0(new_n24275_), .Y(new_n24277_));
  AOI21X1  g24085(.A0(new_n24277_), .A1(new_n24273_), .B0(new_n902_), .Y(new_n24278_));
  AOI21X1  g24086(.A0(new_n24233_), .A1(\asqrt[53] ), .B0(\asqrt[54] ), .Y(new_n24279_));
  AOI21X1  g24087(.A0(new_n24279_), .A1(new_n24277_), .B0(new_n24247_), .Y(new_n24280_));
  NOR3X1   g24088(.A(new_n24280_), .B(new_n24278_), .C(\asqrt[55] ), .Y(new_n24281_));
  NOR2X1   g24089(.A(new_n24281_), .B(new_n24268_), .Y(new_n24282_));
  AND2X1   g24090(.A(new_n23530_), .B(new_n23528_), .Y(new_n24283_));
  NOR3X1   g24091(.A(new_n24283_), .B(new_n23499_), .C(new_n23529_), .Y(new_n24284_));
  NOR3X1   g24092(.A(new_n23622_), .B(new_n24283_), .C(new_n23529_), .Y(new_n24285_));
  NOR2X1   g24093(.A(new_n24285_), .B(new_n23498_), .Y(new_n24286_));
  AOI21X1  g24094(.A0(new_n24284_), .A1(\asqrt[3] ), .B0(new_n24286_), .Y(new_n24287_));
  INVX1    g24095(.A(new_n24287_), .Y(new_n24288_));
  OAI21X1  g24096(.A0(new_n24280_), .A1(new_n24278_), .B0(\asqrt[55] ), .Y(new_n24289_));
  NAND2X1  g24097(.A(new_n24289_), .B(new_n582_), .Y(new_n24290_));
  OAI21X1  g24098(.A0(new_n24290_), .A1(new_n24282_), .B0(new_n24288_), .Y(new_n24291_));
  AOI21X1  g24099(.A0(new_n24291_), .A1(new_n24272_), .B0(new_n481_), .Y(new_n24292_));
  OR4X1    g24100(.A(new_n23622_), .B(new_n23532_), .C(new_n23520_), .D(new_n23514_), .Y(new_n24293_));
  OR2X1    g24101(.A(new_n23532_), .B(new_n23514_), .Y(new_n24294_));
  OAI21X1  g24102(.A0(new_n24294_), .A1(new_n23622_), .B0(new_n23520_), .Y(new_n24295_));
  AND2X1   g24103(.A(new_n24295_), .B(new_n24293_), .Y(new_n24296_));
  OAI21X1  g24104(.A0(new_n24281_), .A1(new_n24268_), .B0(new_n24289_), .Y(new_n24297_));
  AOI21X1  g24105(.A0(new_n24297_), .A1(\asqrt[56] ), .B0(\asqrt[57] ), .Y(new_n24298_));
  AOI21X1  g24106(.A0(new_n24298_), .A1(new_n24291_), .B0(new_n24296_), .Y(new_n24299_));
  OAI21X1  g24107(.A0(new_n24299_), .A1(new_n24292_), .B0(\asqrt[58] ), .Y(new_n24300_));
  AND2X1   g24108(.A(new_n23570_), .B(new_n23569_), .Y(new_n24301_));
  NOR3X1   g24109(.A(new_n24301_), .B(new_n23538_), .C(new_n23568_), .Y(new_n24302_));
  NOR3X1   g24110(.A(new_n23622_), .B(new_n24301_), .C(new_n23568_), .Y(new_n24303_));
  NOR2X1   g24111(.A(new_n24303_), .B(new_n23537_), .Y(new_n24304_));
  AOI21X1  g24112(.A0(new_n24302_), .A1(\asqrt[3] ), .B0(new_n24304_), .Y(new_n24305_));
  NOR3X1   g24113(.A(new_n24299_), .B(new_n24292_), .C(\asqrt[58] ), .Y(new_n24306_));
  OAI21X1  g24114(.A0(new_n24306_), .A1(new_n24305_), .B0(new_n24300_), .Y(new_n24307_));
  AND2X1   g24115(.A(new_n24307_), .B(\asqrt[59] ), .Y(new_n24308_));
  OR2X1    g24116(.A(new_n24306_), .B(new_n24305_), .Y(new_n24309_));
  AND2X1   g24117(.A(new_n23549_), .B(new_n23541_), .Y(new_n24310_));
  NOR3X1   g24118(.A(new_n24310_), .B(new_n23573_), .C(new_n23542_), .Y(new_n24311_));
  NOR3X1   g24119(.A(new_n23622_), .B(new_n24310_), .C(new_n23542_), .Y(new_n24312_));
  NOR2X1   g24120(.A(new_n24312_), .B(new_n23547_), .Y(new_n24313_));
  AOI21X1  g24121(.A0(new_n24311_), .A1(\asqrt[3] ), .B0(new_n24313_), .Y(new_n24314_));
  AND2X1   g24122(.A(new_n24300_), .B(new_n328_), .Y(new_n24315_));
  AOI21X1  g24123(.A0(new_n24315_), .A1(new_n24309_), .B0(new_n24314_), .Y(new_n24316_));
  OAI21X1  g24124(.A0(new_n24316_), .A1(new_n24308_), .B0(\asqrt[60] ), .Y(new_n24317_));
  OR4X1    g24125(.A(new_n23622_), .B(new_n23557_), .C(new_n23577_), .D(new_n23576_), .Y(new_n24318_));
  OR2X1    g24126(.A(new_n23557_), .B(new_n23576_), .Y(new_n24319_));
  OAI21X1  g24127(.A0(new_n24319_), .A1(new_n23622_), .B0(new_n23577_), .Y(new_n24320_));
  AND2X1   g24128(.A(new_n24320_), .B(new_n24318_), .Y(new_n24321_));
  INVX1    g24129(.A(new_n24321_), .Y(new_n24322_));
  AND2X1   g24130(.A(new_n24297_), .B(\asqrt[56] ), .Y(new_n24323_));
  OR2X1    g24131(.A(new_n24281_), .B(new_n24268_), .Y(new_n24324_));
  AND2X1   g24132(.A(new_n24289_), .B(new_n582_), .Y(new_n24325_));
  AOI21X1  g24133(.A0(new_n24325_), .A1(new_n24324_), .B0(new_n24287_), .Y(new_n24326_));
  OAI21X1  g24134(.A0(new_n24326_), .A1(new_n24323_), .B0(\asqrt[57] ), .Y(new_n24327_));
  INVX1    g24135(.A(new_n24296_), .Y(new_n24328_));
  OAI21X1  g24136(.A0(new_n24271_), .A1(new_n582_), .B0(new_n481_), .Y(new_n24329_));
  OAI21X1  g24137(.A0(new_n24329_), .A1(new_n24326_), .B0(new_n24328_), .Y(new_n24330_));
  AOI21X1  g24138(.A0(new_n24330_), .A1(new_n24327_), .B0(new_n399_), .Y(new_n24331_));
  INVX1    g24139(.A(new_n24305_), .Y(new_n24332_));
  NAND3X1  g24140(.A(new_n24330_), .B(new_n24327_), .C(new_n399_), .Y(new_n24333_));
  AOI21X1  g24141(.A0(new_n24333_), .A1(new_n24332_), .B0(new_n24331_), .Y(new_n24334_));
  OAI21X1  g24142(.A0(new_n24334_), .A1(new_n328_), .B0(new_n292_), .Y(new_n24335_));
  OAI21X1  g24143(.A0(new_n24335_), .A1(new_n24316_), .B0(new_n24322_), .Y(new_n24336_));
  AOI21X1  g24144(.A0(new_n24336_), .A1(new_n24317_), .B0(new_n217_), .Y(new_n24337_));
  AOI21X1  g24145(.A0(new_n23565_), .A1(new_n23560_), .B0(new_n23607_), .Y(new_n24338_));
  AND2X1   g24146(.A(new_n24338_), .B(new_n23605_), .Y(new_n24339_));
  AOI22X1  g24147(.A0(new_n23565_), .A1(new_n23560_), .B0(new_n23558_), .B1(\asqrt[60] ), .Y(new_n24340_));
  AOI21X1  g24148(.A0(new_n24340_), .A1(\asqrt[3] ), .B0(new_n23564_), .Y(new_n24341_));
  AOI21X1  g24149(.A0(new_n24339_), .A1(\asqrt[3] ), .B0(new_n24341_), .Y(new_n24342_));
  INVX1    g24150(.A(new_n24342_), .Y(new_n24343_));
  NAND3X1  g24151(.A(new_n24336_), .B(new_n24317_), .C(new_n217_), .Y(new_n24344_));
  AOI21X1  g24152(.A0(new_n24344_), .A1(new_n24343_), .B0(new_n24337_), .Y(new_n24345_));
  OR2X1    g24153(.A(new_n24345_), .B(new_n199_), .Y(new_n24346_));
  OR2X1    g24154(.A(new_n24334_), .B(new_n328_), .Y(new_n24347_));
  NOR2X1   g24155(.A(new_n24306_), .B(new_n24305_), .Y(new_n24348_));
  INVX1    g24156(.A(new_n24314_), .Y(new_n24349_));
  NAND2X1  g24157(.A(new_n24300_), .B(new_n328_), .Y(new_n24350_));
  OAI21X1  g24158(.A0(new_n24350_), .A1(new_n24348_), .B0(new_n24349_), .Y(new_n24351_));
  AOI21X1  g24159(.A0(new_n24351_), .A1(new_n24347_), .B0(new_n292_), .Y(new_n24352_));
  AOI21X1  g24160(.A0(new_n24307_), .A1(\asqrt[59] ), .B0(\asqrt[60] ), .Y(new_n24353_));
  AOI21X1  g24161(.A0(new_n24353_), .A1(new_n24351_), .B0(new_n24321_), .Y(new_n24354_));
  NOR3X1   g24162(.A(new_n24354_), .B(new_n24352_), .C(\asqrt[61] ), .Y(new_n24355_));
  NOR2X1   g24163(.A(new_n24355_), .B(new_n24342_), .Y(new_n24356_));
  OAI21X1  g24164(.A0(new_n24354_), .A1(new_n24352_), .B0(\asqrt[61] ), .Y(new_n24357_));
  NAND2X1  g24165(.A(new_n24357_), .B(new_n199_), .Y(new_n24358_));
  AND2X1   g24166(.A(new_n23611_), .B(new_n23609_), .Y(new_n24359_));
  NOR3X1   g24167(.A(new_n23586_), .B(new_n24359_), .C(new_n23610_), .Y(new_n24360_));
  NOR3X1   g24168(.A(new_n23622_), .B(new_n24359_), .C(new_n23610_), .Y(new_n24361_));
  NOR2X1   g24169(.A(new_n24361_), .B(new_n23585_), .Y(new_n24362_));
  AOI21X1  g24170(.A0(new_n24360_), .A1(\asqrt[3] ), .B0(new_n24362_), .Y(new_n24363_));
  INVX1    g24171(.A(new_n24363_), .Y(new_n24364_));
  OAI21X1  g24172(.A0(new_n24358_), .A1(new_n24356_), .B0(new_n24364_), .Y(new_n24365_));
  NAND4X1  g24173(.A(\asqrt[3] ), .B(new_n23595_), .C(new_n23593_), .D(new_n23615_), .Y(new_n24366_));
  NAND2X1  g24174(.A(new_n23595_), .B(new_n23615_), .Y(new_n24367_));
  OAI21X1  g24175(.A0(new_n24367_), .A1(new_n23622_), .B0(new_n23594_), .Y(new_n24368_));
  AND2X1   g24176(.A(new_n24368_), .B(new_n24366_), .Y(new_n24369_));
  NOR3X1   g24177(.A(new_n23622_), .B(new_n23600_), .C(new_n23596_), .Y(new_n24370_));
  NOR3X1   g24178(.A(new_n24370_), .B(new_n24369_), .C(new_n23647_), .Y(new_n24371_));
  INVX1    g24179(.A(new_n24371_), .Y(new_n24372_));
  AOI21X1  g24180(.A0(new_n24365_), .A1(new_n24346_), .B0(new_n24372_), .Y(new_n24373_));
  OAI21X1  g24181(.A0(new_n24355_), .A1(new_n24342_), .B0(new_n24357_), .Y(new_n24374_));
  INVX1    g24182(.A(new_n24369_), .Y(new_n24375_));
  AOI21X1  g24183(.A0(new_n24374_), .A1(\asqrt[62] ), .B0(new_n24375_), .Y(new_n24376_));
  INVX1    g24184(.A(new_n23600_), .Y(new_n24377_));
  AOI21X1  g24185(.A0(\asqrt[3] ), .A1(new_n24377_), .B0(new_n23630_), .Y(new_n24378_));
  OAI21X1  g24186(.A0(new_n23600_), .A1(new_n23596_), .B0(\asqrt[63] ), .Y(new_n24379_));
  NOR2X1   g24187(.A(new_n24379_), .B(new_n24378_), .Y(new_n24380_));
  AOI21X1  g24188(.A0(new_n24376_), .A1(new_n24365_), .B0(new_n24380_), .Y(new_n24381_));
  OAI21X1  g24189(.A0(new_n24373_), .A1(\asqrt[63] ), .B0(new_n24381_), .Y(\asqrt[2] ));
  MX2X1    g24190(.A(\asqrt[2] ), .B(new_n23625_), .S0(new_n23624_), .Y(new_n24383_));
  AND2X1   g24191(.A(new_n24383_), .B(\asqrt[3] ), .Y(new_n24384_));
  NOR3X1   g24192(.A(\a[4] ), .B(\a[3] ), .C(\a[2] ), .Y(new_n24385_));
  NOR4X1   g24193(.A(new_n24385_), .B(new_n23620_), .C(new_n23647_), .D(new_n23631_), .Y(new_n24386_));
  INVX1    g24194(.A(new_n24386_), .Y(new_n24387_));
  AOI21X1  g24195(.A0(\asqrt[2] ), .A1(\a[4] ), .B0(new_n24387_), .Y(new_n24388_));
  INVX1    g24196(.A(\a[5] ), .Y(new_n24389_));
  AOI21X1  g24197(.A0(\asqrt[2] ), .A1(new_n23624_), .B0(new_n24389_), .Y(new_n24390_));
  NOR2X1   g24198(.A(\a[5] ), .B(\a[4] ), .Y(new_n24391_));
  AND2X1   g24199(.A(\asqrt[2] ), .B(new_n24391_), .Y(new_n24392_));
  NOR3X1   g24200(.A(new_n24392_), .B(new_n24390_), .C(new_n24388_), .Y(new_n24393_));
  OAI21X1  g24201(.A0(new_n24393_), .A1(new_n24384_), .B0(\asqrt[4] ), .Y(new_n24394_));
  INVX1    g24202(.A(new_n23625_), .Y(new_n24395_));
  AND2X1   g24203(.A(new_n24374_), .B(\asqrt[62] ), .Y(new_n24396_));
  OR2X1    g24204(.A(new_n24355_), .B(new_n24342_), .Y(new_n24397_));
  AND2X1   g24205(.A(new_n24357_), .B(new_n199_), .Y(new_n24398_));
  AOI21X1  g24206(.A0(new_n24398_), .A1(new_n24397_), .B0(new_n24363_), .Y(new_n24399_));
  OAI21X1  g24207(.A0(new_n24399_), .A1(new_n24396_), .B0(new_n24371_), .Y(new_n24400_));
  OAI21X1  g24208(.A0(new_n24345_), .A1(new_n199_), .B0(new_n24369_), .Y(new_n24401_));
  OAI22X1  g24209(.A0(new_n24379_), .A1(new_n24378_), .B0(new_n24401_), .B1(new_n24399_), .Y(new_n24402_));
  AOI21X1  g24210(.A0(new_n24400_), .A1(new_n193_), .B0(new_n24402_), .Y(new_n24403_));
  MX2X1    g24211(.A(new_n24403_), .B(new_n24395_), .S0(new_n23624_), .Y(new_n24404_));
  OAI21X1  g24212(.A0(new_n24404_), .A1(new_n23622_), .B0(new_n22874_), .Y(new_n24405_));
  OR2X1    g24213(.A(new_n24373_), .B(\asqrt[63] ), .Y(new_n24406_));
  NOR2X1   g24214(.A(new_n24380_), .B(new_n23622_), .Y(new_n24407_));
  INVX1    g24215(.A(new_n24407_), .Y(new_n24408_));
  AOI21X1  g24216(.A0(new_n24376_), .A1(new_n24365_), .B0(new_n24408_), .Y(new_n24409_));
  AOI22X1  g24217(.A0(new_n24409_), .A1(new_n24406_), .B0(\asqrt[2] ), .B1(new_n24391_), .Y(new_n24410_));
  OAI21X1  g24218(.A0(new_n24373_), .A1(\asqrt[63] ), .B0(new_n24409_), .Y(new_n24411_));
  NAND2X1  g24219(.A(new_n24411_), .B(new_n23626_), .Y(new_n24412_));
  OAI22X1  g24220(.A0(new_n24412_), .A1(new_n24392_), .B0(new_n24410_), .B1(new_n23626_), .Y(new_n24413_));
  OAI21X1  g24221(.A0(new_n24405_), .A1(new_n24393_), .B0(new_n24413_), .Y(new_n24414_));
  AOI21X1  g24222(.A0(new_n24414_), .A1(new_n24394_), .B0(new_n22128_), .Y(new_n24415_));
  NOR2X1   g24223(.A(new_n23637_), .B(new_n23662_), .Y(new_n24416_));
  NAND3X1  g24224(.A(new_n24416_), .B(\asqrt[2] ), .C(new_n23642_), .Y(new_n24417_));
  INVX1    g24225(.A(new_n24416_), .Y(new_n24418_));
  OAI21X1  g24226(.A0(new_n24418_), .A1(new_n24403_), .B0(new_n23665_), .Y(new_n24419_));
  AND2X1   g24227(.A(new_n24419_), .B(new_n24417_), .Y(new_n24420_));
  INVX1    g24228(.A(new_n24420_), .Y(new_n24421_));
  NAND3X1  g24229(.A(new_n24414_), .B(new_n24394_), .C(new_n22128_), .Y(new_n24422_));
  AOI21X1  g24230(.A0(new_n24422_), .A1(new_n24421_), .B0(new_n24415_), .Y(new_n24423_));
  OR2X1    g24231(.A(new_n24423_), .B(new_n21393_), .Y(new_n24424_));
  AND2X1   g24232(.A(new_n24422_), .B(new_n24421_), .Y(new_n24425_));
  AOI21X1  g24233(.A0(new_n23646_), .A1(new_n23645_), .B0(new_n23691_), .Y(new_n24426_));
  NAND3X1  g24234(.A(new_n24426_), .B(\asqrt[2] ), .C(new_n23688_), .Y(new_n24427_));
  OAI22X1  g24235(.A0(new_n23690_), .A1(new_n23689_), .B0(new_n23666_), .B1(new_n22128_), .Y(new_n24428_));
  OAI21X1  g24236(.A0(new_n24428_), .A1(new_n24403_), .B0(new_n23691_), .Y(new_n24429_));
  AND2X1   g24237(.A(new_n24429_), .B(new_n24427_), .Y(new_n24430_));
  INVX1    g24238(.A(new_n24430_), .Y(new_n24431_));
  OR2X1    g24239(.A(new_n24415_), .B(\asqrt[6] ), .Y(new_n24432_));
  OAI21X1  g24240(.A0(new_n24432_), .A1(new_n24425_), .B0(new_n24431_), .Y(new_n24433_));
  AOI21X1  g24241(.A0(new_n24433_), .A1(new_n24424_), .B0(new_n20676_), .Y(new_n24434_));
  AND2X1   g24242(.A(new_n23694_), .B(new_n23692_), .Y(new_n24435_));
  OR4X1    g24243(.A(new_n24403_), .B(new_n24435_), .C(new_n23660_), .D(new_n23693_), .Y(new_n24436_));
  OR2X1    g24244(.A(new_n24435_), .B(new_n23693_), .Y(new_n24437_));
  OAI21X1  g24245(.A0(new_n24437_), .A1(new_n24403_), .B0(new_n23660_), .Y(new_n24438_));
  AND2X1   g24246(.A(new_n24438_), .B(new_n24436_), .Y(new_n24439_));
  OR2X1    g24247(.A(new_n24404_), .B(new_n23622_), .Y(new_n24440_));
  OAI21X1  g24248(.A0(new_n24403_), .A1(new_n23624_), .B0(new_n24386_), .Y(new_n24441_));
  OAI21X1  g24249(.A0(new_n24403_), .A1(\a[4] ), .B0(\a[5] ), .Y(new_n24442_));
  INVX1    g24250(.A(new_n24391_), .Y(new_n24443_));
  OR2X1    g24251(.A(new_n24403_), .B(new_n24443_), .Y(new_n24444_));
  NAND3X1  g24252(.A(new_n24444_), .B(new_n24442_), .C(new_n24441_), .Y(new_n24445_));
  AOI21X1  g24253(.A0(new_n24445_), .A1(new_n24440_), .B0(new_n22874_), .Y(new_n24446_));
  AOI21X1  g24254(.A0(new_n24383_), .A1(\asqrt[3] ), .B0(\asqrt[4] ), .Y(new_n24447_));
  OAI21X1  g24255(.A0(new_n24403_), .A1(new_n24443_), .B0(new_n24411_), .Y(new_n24448_));
  AND2X1   g24256(.A(new_n24411_), .B(new_n23626_), .Y(new_n24449_));
  AOI22X1  g24257(.A0(new_n24449_), .A1(new_n24444_), .B0(new_n24448_), .B1(\a[6] ), .Y(new_n24450_));
  AOI21X1  g24258(.A0(new_n24447_), .A1(new_n24445_), .B0(new_n24450_), .Y(new_n24451_));
  OAI21X1  g24259(.A0(new_n24451_), .A1(new_n24446_), .B0(\asqrt[5] ), .Y(new_n24452_));
  NOR3X1   g24260(.A(new_n24451_), .B(new_n24446_), .C(\asqrt[5] ), .Y(new_n24453_));
  OAI21X1  g24261(.A0(new_n24453_), .A1(new_n24420_), .B0(new_n24452_), .Y(new_n24454_));
  AOI21X1  g24262(.A0(new_n24454_), .A1(\asqrt[6] ), .B0(\asqrt[7] ), .Y(new_n24455_));
  AOI21X1  g24263(.A0(new_n24455_), .A1(new_n24433_), .B0(new_n24439_), .Y(new_n24456_));
  OAI21X1  g24264(.A0(new_n24456_), .A1(new_n24434_), .B0(\asqrt[8] ), .Y(new_n24457_));
  OR4X1    g24265(.A(new_n24403_), .B(new_n23704_), .C(new_n23677_), .D(new_n23669_), .Y(new_n24458_));
  NAND2X1  g24266(.A(new_n23678_), .B(new_n23696_), .Y(new_n24459_));
  OAI21X1  g24267(.A0(new_n24459_), .A1(new_n24403_), .B0(new_n23677_), .Y(new_n24460_));
  AND2X1   g24268(.A(new_n24460_), .B(new_n24458_), .Y(new_n24461_));
  NOR3X1   g24269(.A(new_n24456_), .B(new_n24434_), .C(\asqrt[8] ), .Y(new_n24462_));
  OAI21X1  g24270(.A0(new_n24462_), .A1(new_n24461_), .B0(new_n24457_), .Y(new_n24463_));
  AND2X1   g24271(.A(new_n24463_), .B(\asqrt[9] ), .Y(new_n24464_));
  INVX1    g24272(.A(new_n24461_), .Y(new_n24465_));
  AND2X1   g24273(.A(new_n24454_), .B(\asqrt[6] ), .Y(new_n24466_));
  NAND2X1  g24274(.A(new_n24422_), .B(new_n24421_), .Y(new_n24467_));
  NOR2X1   g24275(.A(new_n24415_), .B(\asqrt[6] ), .Y(new_n24468_));
  AOI21X1  g24276(.A0(new_n24468_), .A1(new_n24467_), .B0(new_n24430_), .Y(new_n24469_));
  OAI21X1  g24277(.A0(new_n24469_), .A1(new_n24466_), .B0(\asqrt[7] ), .Y(new_n24470_));
  INVX1    g24278(.A(new_n24439_), .Y(new_n24471_));
  OAI21X1  g24279(.A0(new_n24423_), .A1(new_n21393_), .B0(new_n20676_), .Y(new_n24472_));
  OAI21X1  g24280(.A0(new_n24472_), .A1(new_n24469_), .B0(new_n24471_), .Y(new_n24473_));
  NAND3X1  g24281(.A(new_n24473_), .B(new_n24470_), .C(new_n19976_), .Y(new_n24474_));
  NAND2X1  g24282(.A(new_n24474_), .B(new_n24465_), .Y(new_n24475_));
  AND2X1   g24283(.A(new_n23720_), .B(new_n23719_), .Y(new_n24476_));
  NOR4X1   g24284(.A(new_n24403_), .B(new_n24476_), .C(new_n23687_), .D(new_n23718_), .Y(new_n24477_));
  AOI22X1  g24285(.A0(new_n23720_), .A1(new_n23719_), .B0(new_n23705_), .B1(\asqrt[8] ), .Y(new_n24478_));
  AOI21X1  g24286(.A0(new_n24478_), .A1(\asqrt[2] ), .B0(new_n23686_), .Y(new_n24479_));
  NOR2X1   g24287(.A(new_n24479_), .B(new_n24477_), .Y(new_n24480_));
  AOI21X1  g24288(.A0(new_n24473_), .A1(new_n24470_), .B0(new_n19976_), .Y(new_n24481_));
  NOR2X1   g24289(.A(new_n24481_), .B(\asqrt[9] ), .Y(new_n24482_));
  AOI21X1  g24290(.A0(new_n24482_), .A1(new_n24475_), .B0(new_n24480_), .Y(new_n24483_));
  OAI21X1  g24291(.A0(new_n24483_), .A1(new_n24464_), .B0(\asqrt[10] ), .Y(new_n24484_));
  AND2X1   g24292(.A(new_n23706_), .B(new_n23698_), .Y(new_n24485_));
  OR4X1    g24293(.A(new_n24403_), .B(new_n24485_), .C(new_n23723_), .D(new_n23699_), .Y(new_n24486_));
  OR2X1    g24294(.A(new_n24485_), .B(new_n23699_), .Y(new_n24487_));
  OAI21X1  g24295(.A0(new_n24487_), .A1(new_n24403_), .B0(new_n23723_), .Y(new_n24488_));
  AND2X1   g24296(.A(new_n24488_), .B(new_n24486_), .Y(new_n24489_));
  INVX1    g24297(.A(new_n24489_), .Y(new_n24490_));
  AOI21X1  g24298(.A0(new_n24474_), .A1(new_n24465_), .B0(new_n24481_), .Y(new_n24491_));
  OAI21X1  g24299(.A0(new_n24491_), .A1(new_n19273_), .B0(new_n18591_), .Y(new_n24492_));
  OAI21X1  g24300(.A0(new_n24492_), .A1(new_n24483_), .B0(new_n24490_), .Y(new_n24493_));
  AOI21X1  g24301(.A0(new_n24493_), .A1(new_n24484_), .B0(new_n17927_), .Y(new_n24494_));
  NOR4X1   g24302(.A(new_n24403_), .B(new_n23714_), .C(new_n23717_), .D(new_n23733_), .Y(new_n24495_));
  AND2X1   g24303(.A(new_n23726_), .B(new_n23708_), .Y(new_n24496_));
  AOI21X1  g24304(.A0(new_n24496_), .A1(\asqrt[2] ), .B0(new_n23713_), .Y(new_n24497_));
  NOR2X1   g24305(.A(new_n24497_), .B(new_n24495_), .Y(new_n24498_));
  INVX1    g24306(.A(new_n24498_), .Y(new_n24499_));
  NAND3X1  g24307(.A(new_n24493_), .B(new_n24484_), .C(new_n17927_), .Y(new_n24500_));
  AOI21X1  g24308(.A0(new_n24500_), .A1(new_n24499_), .B0(new_n24494_), .Y(new_n24501_));
  OR2X1    g24309(.A(new_n24501_), .B(new_n17262_), .Y(new_n24502_));
  AND2X1   g24310(.A(new_n24500_), .B(new_n24499_), .Y(new_n24503_));
  OAI21X1  g24311(.A0(new_n23765_), .A1(new_n23763_), .B0(new_n23732_), .Y(new_n24504_));
  OR2X1    g24312(.A(new_n24504_), .B(new_n23716_), .Y(new_n24505_));
  AOI22X1  g24313(.A0(new_n23734_), .A1(new_n23727_), .B0(new_n23715_), .B1(\asqrt[11] ), .Y(new_n24506_));
  AND2X1   g24314(.A(new_n24506_), .B(\asqrt[2] ), .Y(new_n24507_));
  OAI22X1  g24315(.A0(new_n24507_), .A1(new_n23732_), .B0(new_n24505_), .B1(new_n24403_), .Y(new_n24508_));
  OR2X1    g24316(.A(new_n24494_), .B(\asqrt[12] ), .Y(new_n24509_));
  OAI21X1  g24317(.A0(new_n24509_), .A1(new_n24503_), .B0(new_n24508_), .Y(new_n24510_));
  AOI21X1  g24318(.A0(new_n24510_), .A1(new_n24502_), .B0(new_n16617_), .Y(new_n24511_));
  OR2X1    g24319(.A(new_n23743_), .B(new_n23735_), .Y(new_n24512_));
  NAND3X1  g24320(.A(new_n24512_), .B(new_n23740_), .C(new_n23736_), .Y(new_n24513_));
  NOR2X1   g24321(.A(new_n24513_), .B(new_n24403_), .Y(new_n24514_));
  AND2X1   g24322(.A(new_n24512_), .B(new_n23736_), .Y(new_n24515_));
  AOI21X1  g24323(.A0(new_n24515_), .A1(\asqrt[2] ), .B0(new_n23740_), .Y(new_n24516_));
  NOR2X1   g24324(.A(new_n24516_), .B(new_n24514_), .Y(new_n24517_));
  OR2X1    g24325(.A(new_n24491_), .B(new_n19273_), .Y(new_n24518_));
  AND2X1   g24326(.A(new_n24474_), .B(new_n24465_), .Y(new_n24519_));
  INVX1    g24327(.A(new_n24480_), .Y(new_n24520_));
  OR2X1    g24328(.A(new_n24481_), .B(\asqrt[9] ), .Y(new_n24521_));
  OAI21X1  g24329(.A0(new_n24521_), .A1(new_n24519_), .B0(new_n24520_), .Y(new_n24522_));
  AOI21X1  g24330(.A0(new_n24522_), .A1(new_n24518_), .B0(new_n18591_), .Y(new_n24523_));
  AOI21X1  g24331(.A0(new_n24463_), .A1(\asqrt[9] ), .B0(\asqrt[10] ), .Y(new_n24524_));
  AOI21X1  g24332(.A0(new_n24524_), .A1(new_n24522_), .B0(new_n24489_), .Y(new_n24525_));
  OAI21X1  g24333(.A0(new_n24525_), .A1(new_n24523_), .B0(\asqrt[11] ), .Y(new_n24526_));
  NOR3X1   g24334(.A(new_n24525_), .B(new_n24523_), .C(\asqrt[11] ), .Y(new_n24527_));
  OAI21X1  g24335(.A0(new_n24527_), .A1(new_n24498_), .B0(new_n24526_), .Y(new_n24528_));
  AOI21X1  g24336(.A0(new_n24528_), .A1(\asqrt[12] ), .B0(\asqrt[13] ), .Y(new_n24529_));
  AOI21X1  g24337(.A0(new_n24529_), .A1(new_n24510_), .B0(new_n24517_), .Y(new_n24530_));
  OAI21X1  g24338(.A0(new_n24530_), .A1(new_n24511_), .B0(\asqrt[14] ), .Y(new_n24531_));
  NOR4X1   g24339(.A(new_n24403_), .B(new_n23778_), .C(new_n23751_), .D(new_n23745_), .Y(new_n24532_));
  AND2X1   g24340(.A(new_n23752_), .B(new_n23770_), .Y(new_n24533_));
  AOI21X1  g24341(.A0(new_n24533_), .A1(\asqrt[2] ), .B0(new_n23750_), .Y(new_n24534_));
  NOR2X1   g24342(.A(new_n24534_), .B(new_n24532_), .Y(new_n24535_));
  NOR3X1   g24343(.A(new_n24530_), .B(new_n24511_), .C(\asqrt[14] ), .Y(new_n24536_));
  OAI21X1  g24344(.A0(new_n24536_), .A1(new_n24535_), .B0(new_n24531_), .Y(new_n24537_));
  AND2X1   g24345(.A(new_n24537_), .B(\asqrt[15] ), .Y(new_n24538_));
  INVX1    g24346(.A(new_n24535_), .Y(new_n24539_));
  AND2X1   g24347(.A(new_n24528_), .B(\asqrt[12] ), .Y(new_n24540_));
  NAND2X1  g24348(.A(new_n24500_), .B(new_n24499_), .Y(new_n24541_));
  INVX1    g24349(.A(new_n24508_), .Y(new_n24542_));
  NOR2X1   g24350(.A(new_n24494_), .B(\asqrt[12] ), .Y(new_n24543_));
  AOI21X1  g24351(.A0(new_n24543_), .A1(new_n24541_), .B0(new_n24542_), .Y(new_n24544_));
  OAI21X1  g24352(.A0(new_n24544_), .A1(new_n24540_), .B0(\asqrt[13] ), .Y(new_n24545_));
  INVX1    g24353(.A(new_n24517_), .Y(new_n24546_));
  OAI21X1  g24354(.A0(new_n24501_), .A1(new_n17262_), .B0(new_n16617_), .Y(new_n24547_));
  OAI21X1  g24355(.A0(new_n24547_), .A1(new_n24544_), .B0(new_n24546_), .Y(new_n24548_));
  NAND3X1  g24356(.A(new_n24548_), .B(new_n24545_), .C(new_n15990_), .Y(new_n24549_));
  NAND2X1  g24357(.A(new_n24549_), .B(new_n24539_), .Y(new_n24550_));
  AND2X1   g24358(.A(new_n23794_), .B(new_n23793_), .Y(new_n24551_));
  NOR4X1   g24359(.A(new_n24403_), .B(new_n24551_), .C(new_n23761_), .D(new_n23792_), .Y(new_n24552_));
  AOI22X1  g24360(.A0(new_n23794_), .A1(new_n23793_), .B0(new_n23779_), .B1(\asqrt[14] ), .Y(new_n24553_));
  AOI21X1  g24361(.A0(new_n24553_), .A1(\asqrt[2] ), .B0(new_n23760_), .Y(new_n24554_));
  NOR2X1   g24362(.A(new_n24554_), .B(new_n24552_), .Y(new_n24555_));
  AOI21X1  g24363(.A0(new_n24548_), .A1(new_n24545_), .B0(new_n15990_), .Y(new_n24556_));
  NOR2X1   g24364(.A(new_n24556_), .B(\asqrt[15] ), .Y(new_n24557_));
  AOI21X1  g24365(.A0(new_n24557_), .A1(new_n24550_), .B0(new_n24555_), .Y(new_n24558_));
  OAI21X1  g24366(.A0(new_n24558_), .A1(new_n24538_), .B0(\asqrt[16] ), .Y(new_n24559_));
  AND2X1   g24367(.A(new_n23780_), .B(new_n23772_), .Y(new_n24560_));
  OR4X1    g24368(.A(new_n24403_), .B(new_n24560_), .C(new_n23797_), .D(new_n23773_), .Y(new_n24561_));
  OR2X1    g24369(.A(new_n24560_), .B(new_n23773_), .Y(new_n24562_));
  OAI21X1  g24370(.A0(new_n24562_), .A1(new_n24403_), .B0(new_n23797_), .Y(new_n24563_));
  AND2X1   g24371(.A(new_n24563_), .B(new_n24561_), .Y(new_n24564_));
  INVX1    g24372(.A(new_n24564_), .Y(new_n24565_));
  AOI21X1  g24373(.A0(new_n24549_), .A1(new_n24539_), .B0(new_n24556_), .Y(new_n24566_));
  OAI21X1  g24374(.A0(new_n24566_), .A1(new_n15362_), .B0(new_n14754_), .Y(new_n24567_));
  OAI21X1  g24375(.A0(new_n24567_), .A1(new_n24558_), .B0(new_n24565_), .Y(new_n24568_));
  AOI21X1  g24376(.A0(new_n24568_), .A1(new_n24559_), .B0(new_n14165_), .Y(new_n24569_));
  OR4X1    g24377(.A(new_n24403_), .B(new_n23788_), .C(new_n23791_), .D(new_n23815_), .Y(new_n24570_));
  NAND2X1  g24378(.A(new_n23800_), .B(new_n23782_), .Y(new_n24571_));
  OAI21X1  g24379(.A0(new_n24571_), .A1(new_n24403_), .B0(new_n23791_), .Y(new_n24572_));
  AND2X1   g24380(.A(new_n24572_), .B(new_n24570_), .Y(new_n24573_));
  INVX1    g24381(.A(new_n24573_), .Y(new_n24574_));
  NAND3X1  g24382(.A(new_n24568_), .B(new_n24559_), .C(new_n14165_), .Y(new_n24575_));
  AOI21X1  g24383(.A0(new_n24575_), .A1(new_n24574_), .B0(new_n24569_), .Y(new_n24576_));
  OR2X1    g24384(.A(new_n24576_), .B(new_n13571_), .Y(new_n24577_));
  AND2X1   g24385(.A(new_n24575_), .B(new_n24574_), .Y(new_n24578_));
  OAI21X1  g24386(.A0(new_n23839_), .A1(new_n23837_), .B0(new_n23806_), .Y(new_n24579_));
  NOR3X1   g24387(.A(new_n24579_), .B(new_n24403_), .C(new_n23790_), .Y(new_n24580_));
  AOI22X1  g24388(.A0(new_n23807_), .A1(new_n23801_), .B0(new_n23789_), .B1(\asqrt[17] ), .Y(new_n24581_));
  AOI21X1  g24389(.A0(new_n24581_), .A1(\asqrt[2] ), .B0(new_n23806_), .Y(new_n24582_));
  NOR2X1   g24390(.A(new_n24582_), .B(new_n24580_), .Y(new_n24583_));
  INVX1    g24391(.A(new_n24583_), .Y(new_n24584_));
  OR2X1    g24392(.A(new_n24569_), .B(\asqrt[18] ), .Y(new_n24585_));
  OAI21X1  g24393(.A0(new_n24585_), .A1(new_n24578_), .B0(new_n24584_), .Y(new_n24586_));
  AOI21X1  g24394(.A0(new_n24586_), .A1(new_n24577_), .B0(new_n13000_), .Y(new_n24587_));
  AND2X1   g24395(.A(new_n23842_), .B(new_n23840_), .Y(new_n24588_));
  OR4X1    g24396(.A(new_n24403_), .B(new_n24588_), .C(new_n23814_), .D(new_n23841_), .Y(new_n24589_));
  OR2X1    g24397(.A(new_n24588_), .B(new_n23841_), .Y(new_n24590_));
  OAI21X1  g24398(.A0(new_n24590_), .A1(new_n24403_), .B0(new_n23814_), .Y(new_n24591_));
  AND2X1   g24399(.A(new_n24591_), .B(new_n24589_), .Y(new_n24592_));
  OR2X1    g24400(.A(new_n24566_), .B(new_n15362_), .Y(new_n24593_));
  AND2X1   g24401(.A(new_n24549_), .B(new_n24539_), .Y(new_n24594_));
  INVX1    g24402(.A(new_n24555_), .Y(new_n24595_));
  OR2X1    g24403(.A(new_n24556_), .B(\asqrt[15] ), .Y(new_n24596_));
  OAI21X1  g24404(.A0(new_n24596_), .A1(new_n24594_), .B0(new_n24595_), .Y(new_n24597_));
  AOI21X1  g24405(.A0(new_n24597_), .A1(new_n24593_), .B0(new_n14754_), .Y(new_n24598_));
  AOI21X1  g24406(.A0(new_n24537_), .A1(\asqrt[15] ), .B0(\asqrt[16] ), .Y(new_n24599_));
  AOI21X1  g24407(.A0(new_n24599_), .A1(new_n24597_), .B0(new_n24564_), .Y(new_n24600_));
  OAI21X1  g24408(.A0(new_n24600_), .A1(new_n24598_), .B0(\asqrt[17] ), .Y(new_n24601_));
  NOR3X1   g24409(.A(new_n24600_), .B(new_n24598_), .C(\asqrt[17] ), .Y(new_n24602_));
  OAI21X1  g24410(.A0(new_n24602_), .A1(new_n24573_), .B0(new_n24601_), .Y(new_n24603_));
  AOI21X1  g24411(.A0(new_n24603_), .A1(\asqrt[18] ), .B0(\asqrt[19] ), .Y(new_n24604_));
  AOI21X1  g24412(.A0(new_n24604_), .A1(new_n24586_), .B0(new_n24592_), .Y(new_n24605_));
  OAI21X1  g24413(.A0(new_n24605_), .A1(new_n24587_), .B0(\asqrt[20] ), .Y(new_n24606_));
  NAND3X1  g24414(.A(new_n23826_), .B(new_n23824_), .C(new_n23844_), .Y(new_n24607_));
  NOR3X1   g24415(.A(new_n24403_), .B(new_n23852_), .C(new_n23819_), .Y(new_n24608_));
  OAI22X1  g24416(.A0(new_n24608_), .A1(new_n23824_), .B0(new_n24607_), .B1(new_n24403_), .Y(new_n24609_));
  INVX1    g24417(.A(new_n24609_), .Y(new_n24610_));
  NOR3X1   g24418(.A(new_n24605_), .B(new_n24587_), .C(\asqrt[20] ), .Y(new_n24611_));
  OAI21X1  g24419(.A0(new_n24611_), .A1(new_n24610_), .B0(new_n24606_), .Y(new_n24612_));
  AND2X1   g24420(.A(new_n24612_), .B(\asqrt[21] ), .Y(new_n24613_));
  AND2X1   g24421(.A(new_n24603_), .B(\asqrt[18] ), .Y(new_n24614_));
  NAND2X1  g24422(.A(new_n24575_), .B(new_n24574_), .Y(new_n24615_));
  NOR2X1   g24423(.A(new_n24569_), .B(\asqrt[18] ), .Y(new_n24616_));
  AOI21X1  g24424(.A0(new_n24616_), .A1(new_n24615_), .B0(new_n24583_), .Y(new_n24617_));
  OAI21X1  g24425(.A0(new_n24617_), .A1(new_n24614_), .B0(\asqrt[19] ), .Y(new_n24618_));
  INVX1    g24426(.A(new_n24592_), .Y(new_n24619_));
  OAI21X1  g24427(.A0(new_n24576_), .A1(new_n13571_), .B0(new_n13000_), .Y(new_n24620_));
  OAI21X1  g24428(.A0(new_n24620_), .A1(new_n24617_), .B0(new_n24619_), .Y(new_n24621_));
  NAND3X1  g24429(.A(new_n24621_), .B(new_n24618_), .C(new_n12447_), .Y(new_n24622_));
  NAND2X1  g24430(.A(new_n24622_), .B(new_n24609_), .Y(new_n24623_));
  AND2X1   g24431(.A(new_n23868_), .B(new_n23867_), .Y(new_n24624_));
  NOR4X1   g24432(.A(new_n24403_), .B(new_n24624_), .C(new_n23835_), .D(new_n23866_), .Y(new_n24625_));
  AOI22X1  g24433(.A0(new_n23868_), .A1(new_n23867_), .B0(new_n23853_), .B1(\asqrt[20] ), .Y(new_n24626_));
  AOI21X1  g24434(.A0(new_n24626_), .A1(\asqrt[2] ), .B0(new_n23834_), .Y(new_n24627_));
  NOR2X1   g24435(.A(new_n24627_), .B(new_n24625_), .Y(new_n24628_));
  AOI21X1  g24436(.A0(new_n24621_), .A1(new_n24618_), .B0(new_n12447_), .Y(new_n24629_));
  NOR2X1   g24437(.A(new_n24629_), .B(\asqrt[21] ), .Y(new_n24630_));
  AOI21X1  g24438(.A0(new_n24630_), .A1(new_n24623_), .B0(new_n24628_), .Y(new_n24631_));
  OAI21X1  g24439(.A0(new_n24631_), .A1(new_n24613_), .B0(\asqrt[22] ), .Y(new_n24632_));
  AND2X1   g24440(.A(new_n23854_), .B(new_n23846_), .Y(new_n24633_));
  NOR4X1   g24441(.A(new_n24403_), .B(new_n24633_), .C(new_n23871_), .D(new_n23847_), .Y(new_n24634_));
  NOR2X1   g24442(.A(new_n24633_), .B(new_n23847_), .Y(new_n24635_));
  AOI21X1  g24443(.A0(new_n24635_), .A1(\asqrt[2] ), .B0(new_n23851_), .Y(new_n24636_));
  NOR2X1   g24444(.A(new_n24636_), .B(new_n24634_), .Y(new_n24637_));
  INVX1    g24445(.A(new_n24637_), .Y(new_n24638_));
  AOI21X1  g24446(.A0(new_n24622_), .A1(new_n24609_), .B0(new_n24629_), .Y(new_n24639_));
  OAI21X1  g24447(.A0(new_n24639_), .A1(new_n11896_), .B0(new_n11362_), .Y(new_n24640_));
  OAI21X1  g24448(.A0(new_n24640_), .A1(new_n24631_), .B0(new_n24638_), .Y(new_n24641_));
  AOI21X1  g24449(.A0(new_n24641_), .A1(new_n24632_), .B0(new_n10849_), .Y(new_n24642_));
  OR4X1    g24450(.A(new_n24403_), .B(new_n23862_), .C(new_n23865_), .D(new_n23889_), .Y(new_n24643_));
  NAND2X1  g24451(.A(new_n23874_), .B(new_n23856_), .Y(new_n24644_));
  OAI21X1  g24452(.A0(new_n24644_), .A1(new_n24403_), .B0(new_n23865_), .Y(new_n24645_));
  AND2X1   g24453(.A(new_n24645_), .B(new_n24643_), .Y(new_n24646_));
  INVX1    g24454(.A(new_n24646_), .Y(new_n24647_));
  NAND3X1  g24455(.A(new_n24641_), .B(new_n24632_), .C(new_n10849_), .Y(new_n24648_));
  AOI21X1  g24456(.A0(new_n24648_), .A1(new_n24647_), .B0(new_n24642_), .Y(new_n24649_));
  OR2X1    g24457(.A(new_n24649_), .B(new_n10332_), .Y(new_n24650_));
  AND2X1   g24458(.A(new_n24648_), .B(new_n24647_), .Y(new_n24651_));
  OAI21X1  g24459(.A0(new_n23913_), .A1(new_n23911_), .B0(new_n23880_), .Y(new_n24652_));
  NOR3X1   g24460(.A(new_n24652_), .B(new_n24403_), .C(new_n23864_), .Y(new_n24653_));
  AOI22X1  g24461(.A0(new_n23881_), .A1(new_n23875_), .B0(new_n23863_), .B1(\asqrt[23] ), .Y(new_n24654_));
  AOI21X1  g24462(.A0(new_n24654_), .A1(\asqrt[2] ), .B0(new_n23880_), .Y(new_n24655_));
  NOR2X1   g24463(.A(new_n24655_), .B(new_n24653_), .Y(new_n24656_));
  INVX1    g24464(.A(new_n24656_), .Y(new_n24657_));
  OR2X1    g24465(.A(new_n24642_), .B(\asqrt[24] ), .Y(new_n24658_));
  OAI21X1  g24466(.A0(new_n24658_), .A1(new_n24651_), .B0(new_n24657_), .Y(new_n24659_));
  AOI21X1  g24467(.A0(new_n24659_), .A1(new_n24650_), .B0(new_n9833_), .Y(new_n24660_));
  AND2X1   g24468(.A(new_n23916_), .B(new_n23914_), .Y(new_n24661_));
  NAND2X1  g24469(.A(new_n23887_), .B(new_n23883_), .Y(new_n24662_));
  OR2X1    g24470(.A(new_n24662_), .B(new_n24661_), .Y(new_n24663_));
  NOR3X1   g24471(.A(new_n24403_), .B(new_n24661_), .C(new_n23915_), .Y(new_n24664_));
  OAI22X1  g24472(.A0(new_n24664_), .A1(new_n23887_), .B0(new_n24663_), .B1(new_n24403_), .Y(new_n24665_));
  INVX1    g24473(.A(new_n24665_), .Y(new_n24666_));
  OR2X1    g24474(.A(new_n24639_), .B(new_n11896_), .Y(new_n24667_));
  AND2X1   g24475(.A(new_n24622_), .B(new_n24609_), .Y(new_n24668_));
  INVX1    g24476(.A(new_n24628_), .Y(new_n24669_));
  OR2X1    g24477(.A(new_n24629_), .B(\asqrt[21] ), .Y(new_n24670_));
  OAI21X1  g24478(.A0(new_n24670_), .A1(new_n24668_), .B0(new_n24669_), .Y(new_n24671_));
  AOI21X1  g24479(.A0(new_n24671_), .A1(new_n24667_), .B0(new_n11362_), .Y(new_n24672_));
  AOI21X1  g24480(.A0(new_n24612_), .A1(\asqrt[21] ), .B0(\asqrt[22] ), .Y(new_n24673_));
  AOI21X1  g24481(.A0(new_n24673_), .A1(new_n24671_), .B0(new_n24637_), .Y(new_n24674_));
  OAI21X1  g24482(.A0(new_n24674_), .A1(new_n24672_), .B0(\asqrt[23] ), .Y(new_n24675_));
  NOR3X1   g24483(.A(new_n24674_), .B(new_n24672_), .C(\asqrt[23] ), .Y(new_n24676_));
  OAI21X1  g24484(.A0(new_n24676_), .A1(new_n24646_), .B0(new_n24675_), .Y(new_n24677_));
  AOI21X1  g24485(.A0(new_n24677_), .A1(\asqrt[24] ), .B0(\asqrt[25] ), .Y(new_n24678_));
  AOI21X1  g24486(.A0(new_n24678_), .A1(new_n24659_), .B0(new_n24666_), .Y(new_n24679_));
  OAI21X1  g24487(.A0(new_n24679_), .A1(new_n24660_), .B0(\asqrt[26] ), .Y(new_n24680_));
  OR4X1    g24488(.A(new_n24403_), .B(new_n23926_), .C(new_n23899_), .D(new_n23893_), .Y(new_n24681_));
  NAND2X1  g24489(.A(new_n23900_), .B(new_n23918_), .Y(new_n24682_));
  OAI21X1  g24490(.A0(new_n24682_), .A1(new_n24403_), .B0(new_n23899_), .Y(new_n24683_));
  AND2X1   g24491(.A(new_n24683_), .B(new_n24681_), .Y(new_n24684_));
  NOR3X1   g24492(.A(new_n24679_), .B(new_n24660_), .C(\asqrt[26] ), .Y(new_n24685_));
  OAI21X1  g24493(.A0(new_n24685_), .A1(new_n24684_), .B0(new_n24680_), .Y(new_n24686_));
  AND2X1   g24494(.A(new_n24686_), .B(\asqrt[27] ), .Y(new_n24687_));
  INVX1    g24495(.A(new_n24684_), .Y(new_n24688_));
  AND2X1   g24496(.A(new_n24677_), .B(\asqrt[24] ), .Y(new_n24689_));
  NAND2X1  g24497(.A(new_n24648_), .B(new_n24647_), .Y(new_n24690_));
  NOR2X1   g24498(.A(new_n24642_), .B(\asqrt[24] ), .Y(new_n24691_));
  AOI21X1  g24499(.A0(new_n24691_), .A1(new_n24690_), .B0(new_n24656_), .Y(new_n24692_));
  OAI21X1  g24500(.A0(new_n24692_), .A1(new_n24689_), .B0(\asqrt[25] ), .Y(new_n24693_));
  OAI21X1  g24501(.A0(new_n24649_), .A1(new_n10332_), .B0(new_n9833_), .Y(new_n24694_));
  OAI21X1  g24502(.A0(new_n24694_), .A1(new_n24692_), .B0(new_n24665_), .Y(new_n24695_));
  NAND3X1  g24503(.A(new_n24695_), .B(new_n24693_), .C(new_n9353_), .Y(new_n24696_));
  NAND2X1  g24504(.A(new_n24696_), .B(new_n24688_), .Y(new_n24697_));
  AND2X1   g24505(.A(new_n23942_), .B(new_n23941_), .Y(new_n24698_));
  NOR4X1   g24506(.A(new_n24403_), .B(new_n24698_), .C(new_n23909_), .D(new_n23940_), .Y(new_n24699_));
  AOI22X1  g24507(.A0(new_n23942_), .A1(new_n23941_), .B0(new_n23927_), .B1(\asqrt[26] ), .Y(new_n24700_));
  AOI21X1  g24508(.A0(new_n24700_), .A1(\asqrt[2] ), .B0(new_n23908_), .Y(new_n24701_));
  NOR2X1   g24509(.A(new_n24701_), .B(new_n24699_), .Y(new_n24702_));
  AOI21X1  g24510(.A0(new_n24695_), .A1(new_n24693_), .B0(new_n9353_), .Y(new_n24703_));
  NOR2X1   g24511(.A(new_n24703_), .B(\asqrt[27] ), .Y(new_n24704_));
  AOI21X1  g24512(.A0(new_n24704_), .A1(new_n24697_), .B0(new_n24702_), .Y(new_n24705_));
  OAI21X1  g24513(.A0(new_n24705_), .A1(new_n24687_), .B0(\asqrt[28] ), .Y(new_n24706_));
  AND2X1   g24514(.A(new_n23928_), .B(new_n23920_), .Y(new_n24707_));
  OR4X1    g24515(.A(new_n24403_), .B(new_n24707_), .C(new_n23945_), .D(new_n23921_), .Y(new_n24708_));
  OR2X1    g24516(.A(new_n24707_), .B(new_n23921_), .Y(new_n24709_));
  OAI21X1  g24517(.A0(new_n24709_), .A1(new_n24403_), .B0(new_n23945_), .Y(new_n24710_));
  AND2X1   g24518(.A(new_n24710_), .B(new_n24708_), .Y(new_n24711_));
  INVX1    g24519(.A(new_n24711_), .Y(new_n24712_));
  AOI21X1  g24520(.A0(new_n24696_), .A1(new_n24688_), .B0(new_n24703_), .Y(new_n24713_));
  OAI21X1  g24521(.A0(new_n24713_), .A1(new_n8874_), .B0(new_n8412_), .Y(new_n24714_));
  OAI21X1  g24522(.A0(new_n24714_), .A1(new_n24705_), .B0(new_n24712_), .Y(new_n24715_));
  AOI21X1  g24523(.A0(new_n24715_), .A1(new_n24706_), .B0(new_n7970_), .Y(new_n24716_));
  NAND3X1  g24524(.A(new_n23948_), .B(new_n23935_), .C(new_n23930_), .Y(new_n24717_));
  NOR3X1   g24525(.A(new_n24403_), .B(new_n23936_), .C(new_n23963_), .Y(new_n24718_));
  OAI22X1  g24526(.A0(new_n24718_), .A1(new_n23935_), .B0(new_n24717_), .B1(new_n24403_), .Y(new_n24719_));
  NAND3X1  g24527(.A(new_n24715_), .B(new_n24706_), .C(new_n7970_), .Y(new_n24720_));
  AOI21X1  g24528(.A0(new_n24720_), .A1(new_n24719_), .B0(new_n24716_), .Y(new_n24721_));
  OR2X1    g24529(.A(new_n24721_), .B(new_n7527_), .Y(new_n24722_));
  AND2X1   g24530(.A(new_n24720_), .B(new_n24719_), .Y(new_n24723_));
  AOI21X1  g24531(.A0(new_n23955_), .A1(new_n23949_), .B0(new_n23986_), .Y(new_n24724_));
  AND2X1   g24532(.A(new_n24724_), .B(new_n23984_), .Y(new_n24725_));
  AOI22X1  g24533(.A0(new_n23955_), .A1(new_n23949_), .B0(new_n23937_), .B1(\asqrt[29] ), .Y(new_n24726_));
  AOI21X1  g24534(.A0(new_n24726_), .A1(\asqrt[2] ), .B0(new_n23954_), .Y(new_n24727_));
  AOI21X1  g24535(.A0(new_n24725_), .A1(\asqrt[2] ), .B0(new_n24727_), .Y(new_n24728_));
  INVX1    g24536(.A(new_n24728_), .Y(new_n24729_));
  OR2X1    g24537(.A(new_n24716_), .B(\asqrt[30] ), .Y(new_n24730_));
  OAI21X1  g24538(.A0(new_n24730_), .A1(new_n24723_), .B0(new_n24729_), .Y(new_n24731_));
  AOI21X1  g24539(.A0(new_n24731_), .A1(new_n24722_), .B0(new_n7103_), .Y(new_n24732_));
  AND2X1   g24540(.A(new_n23990_), .B(new_n23988_), .Y(new_n24733_));
  NOR4X1   g24541(.A(new_n24403_), .B(new_n24733_), .C(new_n23962_), .D(new_n23989_), .Y(new_n24734_));
  NOR2X1   g24542(.A(new_n24733_), .B(new_n23989_), .Y(new_n24735_));
  AOI21X1  g24543(.A0(new_n24735_), .A1(\asqrt[2] ), .B0(new_n23961_), .Y(new_n24736_));
  NOR2X1   g24544(.A(new_n24736_), .B(new_n24734_), .Y(new_n24737_));
  OR2X1    g24545(.A(new_n24713_), .B(new_n8874_), .Y(new_n24738_));
  AND2X1   g24546(.A(new_n24696_), .B(new_n24688_), .Y(new_n24739_));
  INVX1    g24547(.A(new_n24702_), .Y(new_n24740_));
  OR2X1    g24548(.A(new_n24703_), .B(\asqrt[27] ), .Y(new_n24741_));
  OAI21X1  g24549(.A0(new_n24741_), .A1(new_n24739_), .B0(new_n24740_), .Y(new_n24742_));
  AOI21X1  g24550(.A0(new_n24742_), .A1(new_n24738_), .B0(new_n8412_), .Y(new_n24743_));
  AOI21X1  g24551(.A0(new_n24686_), .A1(\asqrt[27] ), .B0(\asqrt[28] ), .Y(new_n24744_));
  AOI21X1  g24552(.A0(new_n24744_), .A1(new_n24742_), .B0(new_n24711_), .Y(new_n24745_));
  OAI21X1  g24553(.A0(new_n24745_), .A1(new_n24743_), .B0(\asqrt[29] ), .Y(new_n24746_));
  INVX1    g24554(.A(new_n24719_), .Y(new_n24747_));
  NOR3X1   g24555(.A(new_n24745_), .B(new_n24743_), .C(\asqrt[29] ), .Y(new_n24748_));
  OAI21X1  g24556(.A0(new_n24748_), .A1(new_n24747_), .B0(new_n24746_), .Y(new_n24749_));
  AOI21X1  g24557(.A0(new_n24749_), .A1(\asqrt[30] ), .B0(\asqrt[31] ), .Y(new_n24750_));
  AOI21X1  g24558(.A0(new_n24750_), .A1(new_n24731_), .B0(new_n24737_), .Y(new_n24751_));
  OAI21X1  g24559(.A0(new_n24751_), .A1(new_n24732_), .B0(\asqrt[32] ), .Y(new_n24752_));
  NOR3X1   g24560(.A(new_n24000_), .B(new_n23973_), .C(new_n23967_), .Y(new_n24753_));
  AND2X1   g24561(.A(new_n23974_), .B(new_n23992_), .Y(new_n24754_));
  AOI21X1  g24562(.A0(new_n24754_), .A1(\asqrt[2] ), .B0(new_n23972_), .Y(new_n24755_));
  AOI21X1  g24563(.A0(new_n24753_), .A1(\asqrt[2] ), .B0(new_n24755_), .Y(new_n24756_));
  NOR3X1   g24564(.A(new_n24751_), .B(new_n24732_), .C(\asqrt[32] ), .Y(new_n24757_));
  OAI21X1  g24565(.A0(new_n24757_), .A1(new_n24756_), .B0(new_n24752_), .Y(new_n24758_));
  AND2X1   g24566(.A(new_n24758_), .B(\asqrt[33] ), .Y(new_n24759_));
  INVX1    g24567(.A(new_n24756_), .Y(new_n24760_));
  AND2X1   g24568(.A(new_n24749_), .B(\asqrt[30] ), .Y(new_n24761_));
  NAND2X1  g24569(.A(new_n24720_), .B(new_n24719_), .Y(new_n24762_));
  NOR2X1   g24570(.A(new_n24716_), .B(\asqrt[30] ), .Y(new_n24763_));
  AOI21X1  g24571(.A0(new_n24763_), .A1(new_n24762_), .B0(new_n24728_), .Y(new_n24764_));
  OAI21X1  g24572(.A0(new_n24764_), .A1(new_n24761_), .B0(\asqrt[31] ), .Y(new_n24765_));
  INVX1    g24573(.A(new_n24737_), .Y(new_n24766_));
  OAI21X1  g24574(.A0(new_n24721_), .A1(new_n7527_), .B0(new_n7103_), .Y(new_n24767_));
  OAI21X1  g24575(.A0(new_n24767_), .A1(new_n24764_), .B0(new_n24766_), .Y(new_n24768_));
  NAND3X1  g24576(.A(new_n24768_), .B(new_n24765_), .C(new_n6699_), .Y(new_n24769_));
  NAND2X1  g24577(.A(new_n24769_), .B(new_n24760_), .Y(new_n24770_));
  AND2X1   g24578(.A(new_n24016_), .B(new_n24015_), .Y(new_n24771_));
  NOR3X1   g24579(.A(new_n24771_), .B(new_n23983_), .C(new_n24014_), .Y(new_n24772_));
  AOI22X1  g24580(.A0(new_n24016_), .A1(new_n24015_), .B0(new_n24001_), .B1(\asqrt[32] ), .Y(new_n24773_));
  AOI21X1  g24581(.A0(new_n24773_), .A1(\asqrt[2] ), .B0(new_n23982_), .Y(new_n24774_));
  AOI21X1  g24582(.A0(new_n24772_), .A1(\asqrt[2] ), .B0(new_n24774_), .Y(new_n24775_));
  AOI21X1  g24583(.A0(new_n24768_), .A1(new_n24765_), .B0(new_n6699_), .Y(new_n24776_));
  NOR2X1   g24584(.A(new_n24776_), .B(\asqrt[33] ), .Y(new_n24777_));
  AOI21X1  g24585(.A0(new_n24777_), .A1(new_n24770_), .B0(new_n24775_), .Y(new_n24778_));
  OAI21X1  g24586(.A0(new_n24778_), .A1(new_n24759_), .B0(\asqrt[34] ), .Y(new_n24779_));
  AND2X1   g24587(.A(new_n24002_), .B(new_n23994_), .Y(new_n24780_));
  OR4X1    g24588(.A(new_n24403_), .B(new_n24780_), .C(new_n24019_), .D(new_n23995_), .Y(new_n24781_));
  OR2X1    g24589(.A(new_n24780_), .B(new_n23995_), .Y(new_n24782_));
  OAI21X1  g24590(.A0(new_n24782_), .A1(new_n24403_), .B0(new_n24019_), .Y(new_n24783_));
  AND2X1   g24591(.A(new_n24783_), .B(new_n24781_), .Y(new_n24784_));
  INVX1    g24592(.A(new_n24784_), .Y(new_n24785_));
  AOI21X1  g24593(.A0(new_n24769_), .A1(new_n24760_), .B0(new_n24776_), .Y(new_n24786_));
  OAI21X1  g24594(.A0(new_n24786_), .A1(new_n6294_), .B0(new_n5941_), .Y(new_n24787_));
  OAI21X1  g24595(.A0(new_n24787_), .A1(new_n24778_), .B0(new_n24785_), .Y(new_n24788_));
  AOI21X1  g24596(.A0(new_n24788_), .A1(new_n24779_), .B0(new_n5541_), .Y(new_n24789_));
  OR4X1    g24597(.A(new_n24403_), .B(new_n24010_), .C(new_n24013_), .D(new_n24037_), .Y(new_n24790_));
  NAND2X1  g24598(.A(new_n24022_), .B(new_n24004_), .Y(new_n24791_));
  OAI21X1  g24599(.A0(new_n24791_), .A1(new_n24403_), .B0(new_n24013_), .Y(new_n24792_));
  AND2X1   g24600(.A(new_n24792_), .B(new_n24790_), .Y(new_n24793_));
  INVX1    g24601(.A(new_n24793_), .Y(new_n24794_));
  NAND3X1  g24602(.A(new_n24788_), .B(new_n24779_), .C(new_n5541_), .Y(new_n24795_));
  AOI21X1  g24603(.A0(new_n24795_), .A1(new_n24794_), .B0(new_n24789_), .Y(new_n24796_));
  OR2X1    g24604(.A(new_n24796_), .B(new_n5176_), .Y(new_n24797_));
  AND2X1   g24605(.A(new_n24795_), .B(new_n24794_), .Y(new_n24798_));
  OAI21X1  g24606(.A0(new_n24054_), .A1(new_n24052_), .B0(new_n24028_), .Y(new_n24799_));
  NOR3X1   g24607(.A(new_n24799_), .B(new_n24403_), .C(new_n24012_), .Y(new_n24800_));
  AOI22X1  g24608(.A0(new_n24029_), .A1(new_n24023_), .B0(new_n24011_), .B1(\asqrt[35] ), .Y(new_n24801_));
  AOI21X1  g24609(.A0(new_n24801_), .A1(\asqrt[2] ), .B0(new_n24028_), .Y(new_n24802_));
  NOR2X1   g24610(.A(new_n24802_), .B(new_n24800_), .Y(new_n24803_));
  INVX1    g24611(.A(new_n24803_), .Y(new_n24804_));
  OR2X1    g24612(.A(new_n24789_), .B(\asqrt[36] ), .Y(new_n24805_));
  OAI21X1  g24613(.A0(new_n24805_), .A1(new_n24798_), .B0(new_n24804_), .Y(new_n24806_));
  AOI21X1  g24614(.A0(new_n24806_), .A1(new_n24797_), .B0(new_n4826_), .Y(new_n24807_));
  AND2X1   g24615(.A(new_n24057_), .B(new_n24055_), .Y(new_n24808_));
  OR4X1    g24616(.A(new_n24403_), .B(new_n24808_), .C(new_n24036_), .D(new_n24056_), .Y(new_n24809_));
  OR2X1    g24617(.A(new_n24808_), .B(new_n24056_), .Y(new_n24810_));
  OAI21X1  g24618(.A0(new_n24810_), .A1(new_n24403_), .B0(new_n24036_), .Y(new_n24811_));
  AND2X1   g24619(.A(new_n24811_), .B(new_n24809_), .Y(new_n24812_));
  OR2X1    g24620(.A(new_n24786_), .B(new_n6294_), .Y(new_n24813_));
  AND2X1   g24621(.A(new_n24769_), .B(new_n24760_), .Y(new_n24814_));
  INVX1    g24622(.A(new_n24775_), .Y(new_n24815_));
  OR2X1    g24623(.A(new_n24776_), .B(\asqrt[33] ), .Y(new_n24816_));
  OAI21X1  g24624(.A0(new_n24816_), .A1(new_n24814_), .B0(new_n24815_), .Y(new_n24817_));
  AOI21X1  g24625(.A0(new_n24817_), .A1(new_n24813_), .B0(new_n5941_), .Y(new_n24818_));
  AOI21X1  g24626(.A0(new_n24758_), .A1(\asqrt[33] ), .B0(\asqrt[34] ), .Y(new_n24819_));
  AOI21X1  g24627(.A0(new_n24819_), .A1(new_n24817_), .B0(new_n24784_), .Y(new_n24820_));
  OAI21X1  g24628(.A0(new_n24820_), .A1(new_n24818_), .B0(\asqrt[35] ), .Y(new_n24821_));
  NOR3X1   g24629(.A(new_n24820_), .B(new_n24818_), .C(\asqrt[35] ), .Y(new_n24822_));
  OAI21X1  g24630(.A0(new_n24822_), .A1(new_n24793_), .B0(new_n24821_), .Y(new_n24823_));
  AOI21X1  g24631(.A0(new_n24823_), .A1(\asqrt[36] ), .B0(\asqrt[37] ), .Y(new_n24824_));
  AOI21X1  g24632(.A0(new_n24824_), .A1(new_n24806_), .B0(new_n24812_), .Y(new_n24825_));
  OAI21X1  g24633(.A0(new_n24825_), .A1(new_n24807_), .B0(\asqrt[38] ), .Y(new_n24826_));
  NAND3X1  g24634(.A(new_n24048_), .B(new_n24046_), .C(new_n24067_), .Y(new_n24827_));
  NOR3X1   g24635(.A(new_n24403_), .B(new_n24059_), .C(new_n24041_), .Y(new_n24828_));
  OAI22X1  g24636(.A0(new_n24828_), .A1(new_n24046_), .B0(new_n24827_), .B1(new_n24403_), .Y(new_n24829_));
  INVX1    g24637(.A(new_n24829_), .Y(new_n24830_));
  NOR3X1   g24638(.A(new_n24825_), .B(new_n24807_), .C(\asqrt[38] ), .Y(new_n24831_));
  OAI21X1  g24639(.A0(new_n24831_), .A1(new_n24830_), .B0(new_n24826_), .Y(new_n24832_));
  AND2X1   g24640(.A(new_n24832_), .B(\asqrt[39] ), .Y(new_n24833_));
  AND2X1   g24641(.A(new_n24823_), .B(\asqrt[36] ), .Y(new_n24834_));
  NAND2X1  g24642(.A(new_n24795_), .B(new_n24794_), .Y(new_n24835_));
  NOR2X1   g24643(.A(new_n24789_), .B(\asqrt[36] ), .Y(new_n24836_));
  AOI21X1  g24644(.A0(new_n24836_), .A1(new_n24835_), .B0(new_n24803_), .Y(new_n24837_));
  OAI21X1  g24645(.A0(new_n24837_), .A1(new_n24834_), .B0(\asqrt[37] ), .Y(new_n24838_));
  INVX1    g24646(.A(new_n24812_), .Y(new_n24839_));
  OAI21X1  g24647(.A0(new_n24796_), .A1(new_n5176_), .B0(new_n4826_), .Y(new_n24840_));
  OAI21X1  g24648(.A0(new_n24840_), .A1(new_n24837_), .B0(new_n24839_), .Y(new_n24841_));
  NAND3X1  g24649(.A(new_n24841_), .B(new_n24838_), .C(new_n4493_), .Y(new_n24842_));
  NAND2X1  g24650(.A(new_n24842_), .B(new_n24829_), .Y(new_n24843_));
  AND2X1   g24651(.A(new_n24103_), .B(new_n24102_), .Y(new_n24844_));
  NOR4X1   g24652(.A(new_n24403_), .B(new_n24844_), .C(new_n24066_), .D(new_n24101_), .Y(new_n24845_));
  AOI22X1  g24653(.A0(new_n24103_), .A1(new_n24102_), .B0(new_n24075_), .B1(\asqrt[38] ), .Y(new_n24846_));
  AOI21X1  g24654(.A0(new_n24846_), .A1(\asqrt[2] ), .B0(new_n24065_), .Y(new_n24847_));
  NOR2X1   g24655(.A(new_n24847_), .B(new_n24845_), .Y(new_n24848_));
  AOI21X1  g24656(.A0(new_n24841_), .A1(new_n24838_), .B0(new_n4493_), .Y(new_n24849_));
  NOR2X1   g24657(.A(new_n24849_), .B(\asqrt[39] ), .Y(new_n24850_));
  AOI21X1  g24658(.A0(new_n24850_), .A1(new_n24843_), .B0(new_n24848_), .Y(new_n24851_));
  OAI21X1  g24659(.A0(new_n24851_), .A1(new_n24833_), .B0(\asqrt[40] ), .Y(new_n24852_));
  AND2X1   g24660(.A(new_n24076_), .B(new_n24069_), .Y(new_n24853_));
  NOR3X1   g24661(.A(new_n24853_), .B(new_n24106_), .C(new_n24070_), .Y(new_n24854_));
  NOR2X1   g24662(.A(new_n24853_), .B(new_n24070_), .Y(new_n24855_));
  AOI21X1  g24663(.A0(new_n24855_), .A1(\asqrt[2] ), .B0(new_n24074_), .Y(new_n24856_));
  AOI21X1  g24664(.A0(new_n24854_), .A1(\asqrt[2] ), .B0(new_n24856_), .Y(new_n24857_));
  INVX1    g24665(.A(new_n24857_), .Y(new_n24858_));
  AOI21X1  g24666(.A0(new_n24842_), .A1(new_n24829_), .B0(new_n24849_), .Y(new_n24859_));
  OAI21X1  g24667(.A0(new_n24859_), .A1(new_n4165_), .B0(new_n3863_), .Y(new_n24860_));
  OAI21X1  g24668(.A0(new_n24860_), .A1(new_n24851_), .B0(new_n24858_), .Y(new_n24861_));
  AOI21X1  g24669(.A0(new_n24861_), .A1(new_n24852_), .B0(new_n3564_), .Y(new_n24862_));
  OR4X1    g24670(.A(new_n24403_), .B(new_n24084_), .C(new_n24110_), .D(new_n24109_), .Y(new_n24863_));
  OR2X1    g24671(.A(new_n24084_), .B(new_n24109_), .Y(new_n24864_));
  OAI21X1  g24672(.A0(new_n24864_), .A1(new_n24403_), .B0(new_n24110_), .Y(new_n24865_));
  AND2X1   g24673(.A(new_n24865_), .B(new_n24863_), .Y(new_n24866_));
  INVX1    g24674(.A(new_n24866_), .Y(new_n24867_));
  NAND3X1  g24675(.A(new_n24861_), .B(new_n24852_), .C(new_n3564_), .Y(new_n24868_));
  AOI21X1  g24676(.A0(new_n24868_), .A1(new_n24867_), .B0(new_n24862_), .Y(new_n24869_));
  OR2X1    g24677(.A(new_n24869_), .B(new_n3276_), .Y(new_n24870_));
  AND2X1   g24678(.A(new_n24868_), .B(new_n24867_), .Y(new_n24871_));
  OAI21X1  g24679(.A0(new_n24128_), .A1(new_n24126_), .B0(new_n24092_), .Y(new_n24872_));
  NOR3X1   g24680(.A(new_n24872_), .B(new_n24403_), .C(new_n24086_), .Y(new_n24873_));
  AOI22X1  g24681(.A0(new_n24093_), .A1(new_n24087_), .B0(new_n24085_), .B1(\asqrt[41] ), .Y(new_n24874_));
  AOI21X1  g24682(.A0(new_n24874_), .A1(\asqrt[2] ), .B0(new_n24092_), .Y(new_n24875_));
  NOR2X1   g24683(.A(new_n24875_), .B(new_n24873_), .Y(new_n24876_));
  INVX1    g24684(.A(new_n24876_), .Y(new_n24877_));
  OR2X1    g24685(.A(new_n24862_), .B(\asqrt[42] ), .Y(new_n24878_));
  OAI21X1  g24686(.A0(new_n24878_), .A1(new_n24871_), .B0(new_n24877_), .Y(new_n24879_));
  AOI21X1  g24687(.A0(new_n24879_), .A1(new_n24870_), .B0(new_n3008_), .Y(new_n24880_));
  AND2X1   g24688(.A(new_n24131_), .B(new_n24129_), .Y(new_n24881_));
  OR4X1    g24689(.A(new_n24403_), .B(new_n24881_), .C(new_n24100_), .D(new_n24130_), .Y(new_n24882_));
  OR2X1    g24690(.A(new_n24881_), .B(new_n24130_), .Y(new_n24883_));
  OAI21X1  g24691(.A0(new_n24883_), .A1(new_n24403_), .B0(new_n24100_), .Y(new_n24884_));
  AND2X1   g24692(.A(new_n24884_), .B(new_n24882_), .Y(new_n24885_));
  OR2X1    g24693(.A(new_n24859_), .B(new_n4165_), .Y(new_n24886_));
  AND2X1   g24694(.A(new_n24842_), .B(new_n24829_), .Y(new_n24887_));
  INVX1    g24695(.A(new_n24848_), .Y(new_n24888_));
  OR2X1    g24696(.A(new_n24849_), .B(\asqrt[39] ), .Y(new_n24889_));
  OAI21X1  g24697(.A0(new_n24889_), .A1(new_n24887_), .B0(new_n24888_), .Y(new_n24890_));
  AOI21X1  g24698(.A0(new_n24890_), .A1(new_n24886_), .B0(new_n3863_), .Y(new_n24891_));
  AOI21X1  g24699(.A0(new_n24832_), .A1(\asqrt[39] ), .B0(\asqrt[40] ), .Y(new_n24892_));
  AOI21X1  g24700(.A0(new_n24892_), .A1(new_n24890_), .B0(new_n24857_), .Y(new_n24893_));
  OAI21X1  g24701(.A0(new_n24893_), .A1(new_n24891_), .B0(\asqrt[41] ), .Y(new_n24894_));
  NOR3X1   g24702(.A(new_n24893_), .B(new_n24891_), .C(\asqrt[41] ), .Y(new_n24895_));
  OAI21X1  g24703(.A0(new_n24895_), .A1(new_n24866_), .B0(new_n24894_), .Y(new_n24896_));
  AOI21X1  g24704(.A0(new_n24896_), .A1(\asqrt[42] ), .B0(\asqrt[43] ), .Y(new_n24897_));
  AOI21X1  g24705(.A0(new_n24897_), .A1(new_n24879_), .B0(new_n24885_), .Y(new_n24898_));
  OAI21X1  g24706(.A0(new_n24898_), .A1(new_n24880_), .B0(\asqrt[44] ), .Y(new_n24899_));
  OR4X1    g24707(.A(new_n24403_), .B(new_n24133_), .C(new_n24121_), .D(new_n24115_), .Y(new_n24900_));
  OR2X1    g24708(.A(new_n24133_), .B(new_n24115_), .Y(new_n24901_));
  OAI21X1  g24709(.A0(new_n24901_), .A1(new_n24403_), .B0(new_n24121_), .Y(new_n24902_));
  AND2X1   g24710(.A(new_n24902_), .B(new_n24900_), .Y(new_n24903_));
  NOR3X1   g24711(.A(new_n24898_), .B(new_n24880_), .C(\asqrt[44] ), .Y(new_n24904_));
  OAI21X1  g24712(.A0(new_n24904_), .A1(new_n24903_), .B0(new_n24899_), .Y(new_n24905_));
  AND2X1   g24713(.A(new_n24905_), .B(\asqrt[45] ), .Y(new_n24906_));
  INVX1    g24714(.A(new_n24903_), .Y(new_n24907_));
  AND2X1   g24715(.A(new_n24896_), .B(\asqrt[42] ), .Y(new_n24908_));
  NAND2X1  g24716(.A(new_n24868_), .B(new_n24867_), .Y(new_n24909_));
  NOR2X1   g24717(.A(new_n24862_), .B(\asqrt[42] ), .Y(new_n24910_));
  AOI21X1  g24718(.A0(new_n24910_), .A1(new_n24909_), .B0(new_n24876_), .Y(new_n24911_));
  OAI21X1  g24719(.A0(new_n24911_), .A1(new_n24908_), .B0(\asqrt[43] ), .Y(new_n24912_));
  INVX1    g24720(.A(new_n24885_), .Y(new_n24913_));
  OAI21X1  g24721(.A0(new_n24869_), .A1(new_n3276_), .B0(new_n3008_), .Y(new_n24914_));
  OAI21X1  g24722(.A0(new_n24914_), .A1(new_n24911_), .B0(new_n24913_), .Y(new_n24915_));
  NAND3X1  g24723(.A(new_n24915_), .B(new_n24912_), .C(new_n2769_), .Y(new_n24916_));
  NAND2X1  g24724(.A(new_n24916_), .B(new_n24907_), .Y(new_n24917_));
  AND2X1   g24725(.A(new_n24177_), .B(new_n24176_), .Y(new_n24918_));
  NOR3X1   g24726(.A(new_n24918_), .B(new_n24140_), .C(new_n24175_), .Y(new_n24919_));
  AOI22X1  g24727(.A0(new_n24177_), .A1(new_n24176_), .B0(new_n24149_), .B1(\asqrt[44] ), .Y(new_n24920_));
  AOI21X1  g24728(.A0(new_n24920_), .A1(\asqrt[2] ), .B0(new_n24139_), .Y(new_n24921_));
  AOI21X1  g24729(.A0(new_n24919_), .A1(\asqrt[2] ), .B0(new_n24921_), .Y(new_n24922_));
  AOI21X1  g24730(.A0(new_n24915_), .A1(new_n24912_), .B0(new_n2769_), .Y(new_n24923_));
  NOR2X1   g24731(.A(new_n24923_), .B(\asqrt[45] ), .Y(new_n24924_));
  AOI21X1  g24732(.A0(new_n24924_), .A1(new_n24917_), .B0(new_n24922_), .Y(new_n24925_));
  OAI21X1  g24733(.A0(new_n24925_), .A1(new_n24906_), .B0(\asqrt[46] ), .Y(new_n24926_));
  AND2X1   g24734(.A(new_n24150_), .B(new_n24143_), .Y(new_n24927_));
  NOR3X1   g24735(.A(new_n24927_), .B(new_n24180_), .C(new_n24144_), .Y(new_n24928_));
  NOR2X1   g24736(.A(new_n24927_), .B(new_n24144_), .Y(new_n24929_));
  AOI21X1  g24737(.A0(new_n24929_), .A1(\asqrt[2] ), .B0(new_n24148_), .Y(new_n24930_));
  AOI21X1  g24738(.A0(new_n24928_), .A1(\asqrt[2] ), .B0(new_n24930_), .Y(new_n24931_));
  INVX1    g24739(.A(new_n24931_), .Y(new_n24932_));
  AOI21X1  g24740(.A0(new_n24916_), .A1(new_n24907_), .B0(new_n24923_), .Y(new_n24933_));
  OAI21X1  g24741(.A0(new_n24933_), .A1(new_n2570_), .B0(new_n2263_), .Y(new_n24934_));
  OAI21X1  g24742(.A0(new_n24934_), .A1(new_n24925_), .B0(new_n24932_), .Y(new_n24935_));
  AOI21X1  g24743(.A0(new_n24935_), .A1(new_n24926_), .B0(new_n2040_), .Y(new_n24936_));
  OR4X1    g24744(.A(new_n24403_), .B(new_n24158_), .C(new_n24184_), .D(new_n24183_), .Y(new_n24937_));
  OR2X1    g24745(.A(new_n24158_), .B(new_n24183_), .Y(new_n24938_));
  OAI21X1  g24746(.A0(new_n24938_), .A1(new_n24403_), .B0(new_n24184_), .Y(new_n24939_));
  AND2X1   g24747(.A(new_n24939_), .B(new_n24937_), .Y(new_n24940_));
  INVX1    g24748(.A(new_n24940_), .Y(new_n24941_));
  NAND3X1  g24749(.A(new_n24935_), .B(new_n24926_), .C(new_n2040_), .Y(new_n24942_));
  AOI21X1  g24750(.A0(new_n24942_), .A1(new_n24941_), .B0(new_n24936_), .Y(new_n24943_));
  OR2X1    g24751(.A(new_n24943_), .B(new_n1834_), .Y(new_n24944_));
  AND2X1   g24752(.A(new_n24942_), .B(new_n24941_), .Y(new_n24945_));
  OAI21X1  g24753(.A0(new_n24202_), .A1(new_n24200_), .B0(new_n24166_), .Y(new_n24946_));
  NOR3X1   g24754(.A(new_n24946_), .B(new_n24403_), .C(new_n24160_), .Y(new_n24947_));
  AOI22X1  g24755(.A0(new_n24167_), .A1(new_n24161_), .B0(new_n24159_), .B1(\asqrt[47] ), .Y(new_n24948_));
  AOI21X1  g24756(.A0(new_n24948_), .A1(\asqrt[2] ), .B0(new_n24166_), .Y(new_n24949_));
  NOR2X1   g24757(.A(new_n24949_), .B(new_n24947_), .Y(new_n24950_));
  INVX1    g24758(.A(new_n24950_), .Y(new_n24951_));
  OR2X1    g24759(.A(new_n24936_), .B(\asqrt[48] ), .Y(new_n24952_));
  OAI21X1  g24760(.A0(new_n24952_), .A1(new_n24945_), .B0(new_n24951_), .Y(new_n24953_));
  AOI21X1  g24761(.A0(new_n24953_), .A1(new_n24944_), .B0(new_n1632_), .Y(new_n24954_));
  AND2X1   g24762(.A(new_n24205_), .B(new_n24203_), .Y(new_n24955_));
  OR4X1    g24763(.A(new_n24403_), .B(new_n24955_), .C(new_n24174_), .D(new_n24204_), .Y(new_n24956_));
  OR2X1    g24764(.A(new_n24955_), .B(new_n24204_), .Y(new_n24957_));
  OAI21X1  g24765(.A0(new_n24957_), .A1(new_n24403_), .B0(new_n24174_), .Y(new_n24958_));
  AND2X1   g24766(.A(new_n24958_), .B(new_n24956_), .Y(new_n24959_));
  OR2X1    g24767(.A(new_n24933_), .B(new_n2570_), .Y(new_n24960_));
  AND2X1   g24768(.A(new_n24916_), .B(new_n24907_), .Y(new_n24961_));
  INVX1    g24769(.A(new_n24922_), .Y(new_n24962_));
  OR2X1    g24770(.A(new_n24923_), .B(\asqrt[45] ), .Y(new_n24963_));
  OAI21X1  g24771(.A0(new_n24963_), .A1(new_n24961_), .B0(new_n24962_), .Y(new_n24964_));
  AOI21X1  g24772(.A0(new_n24964_), .A1(new_n24960_), .B0(new_n2263_), .Y(new_n24965_));
  AOI21X1  g24773(.A0(new_n24905_), .A1(\asqrt[45] ), .B0(\asqrt[46] ), .Y(new_n24966_));
  AOI21X1  g24774(.A0(new_n24966_), .A1(new_n24964_), .B0(new_n24931_), .Y(new_n24967_));
  OAI21X1  g24775(.A0(new_n24967_), .A1(new_n24965_), .B0(\asqrt[47] ), .Y(new_n24968_));
  NOR3X1   g24776(.A(new_n24967_), .B(new_n24965_), .C(\asqrt[47] ), .Y(new_n24969_));
  OAI21X1  g24777(.A0(new_n24969_), .A1(new_n24940_), .B0(new_n24968_), .Y(new_n24970_));
  AOI21X1  g24778(.A0(new_n24970_), .A1(\asqrt[48] ), .B0(\asqrt[49] ), .Y(new_n24971_));
  AOI21X1  g24779(.A0(new_n24971_), .A1(new_n24953_), .B0(new_n24959_), .Y(new_n24972_));
  OAI21X1  g24780(.A0(new_n24972_), .A1(new_n24954_), .B0(\asqrt[50] ), .Y(new_n24973_));
  OR4X1    g24781(.A(new_n24403_), .B(new_n24207_), .C(new_n24195_), .D(new_n24189_), .Y(new_n24974_));
  OR2X1    g24782(.A(new_n24207_), .B(new_n24189_), .Y(new_n24975_));
  OAI21X1  g24783(.A0(new_n24975_), .A1(new_n24403_), .B0(new_n24195_), .Y(new_n24976_));
  AND2X1   g24784(.A(new_n24976_), .B(new_n24974_), .Y(new_n24977_));
  NOR3X1   g24785(.A(new_n24972_), .B(new_n24954_), .C(\asqrt[50] ), .Y(new_n24978_));
  OAI21X1  g24786(.A0(new_n24978_), .A1(new_n24977_), .B0(new_n24973_), .Y(new_n24979_));
  AND2X1   g24787(.A(new_n24979_), .B(\asqrt[51] ), .Y(new_n24980_));
  INVX1    g24788(.A(new_n24977_), .Y(new_n24981_));
  AND2X1   g24789(.A(new_n24970_), .B(\asqrt[48] ), .Y(new_n24982_));
  NAND2X1  g24790(.A(new_n24942_), .B(new_n24941_), .Y(new_n24983_));
  NOR2X1   g24791(.A(new_n24936_), .B(\asqrt[48] ), .Y(new_n24984_));
  AOI21X1  g24792(.A0(new_n24984_), .A1(new_n24983_), .B0(new_n24950_), .Y(new_n24985_));
  OAI21X1  g24793(.A0(new_n24985_), .A1(new_n24982_), .B0(\asqrt[49] ), .Y(new_n24986_));
  INVX1    g24794(.A(new_n24959_), .Y(new_n24987_));
  OAI21X1  g24795(.A0(new_n24943_), .A1(new_n1834_), .B0(new_n1632_), .Y(new_n24988_));
  OAI21X1  g24796(.A0(new_n24988_), .A1(new_n24985_), .B0(new_n24987_), .Y(new_n24989_));
  NAND3X1  g24797(.A(new_n24989_), .B(new_n24986_), .C(new_n1469_), .Y(new_n24990_));
  NAND2X1  g24798(.A(new_n24990_), .B(new_n24981_), .Y(new_n24991_));
  AND2X1   g24799(.A(new_n24251_), .B(new_n24250_), .Y(new_n24992_));
  NOR4X1   g24800(.A(new_n24403_), .B(new_n24992_), .C(new_n24214_), .D(new_n24249_), .Y(new_n24993_));
  AOI22X1  g24801(.A0(new_n24251_), .A1(new_n24250_), .B0(new_n24223_), .B1(\asqrt[50] ), .Y(new_n24994_));
  AOI21X1  g24802(.A0(new_n24994_), .A1(\asqrt[2] ), .B0(new_n24213_), .Y(new_n24995_));
  NOR2X1   g24803(.A(new_n24995_), .B(new_n24993_), .Y(new_n24996_));
  AOI21X1  g24804(.A0(new_n24989_), .A1(new_n24986_), .B0(new_n1469_), .Y(new_n24997_));
  NOR2X1   g24805(.A(new_n24997_), .B(\asqrt[51] ), .Y(new_n24998_));
  AOI21X1  g24806(.A0(new_n24998_), .A1(new_n24991_), .B0(new_n24996_), .Y(new_n24999_));
  OAI21X1  g24807(.A0(new_n24999_), .A1(new_n24980_), .B0(\asqrt[52] ), .Y(new_n25000_));
  AND2X1   g24808(.A(new_n24224_), .B(new_n24217_), .Y(new_n25001_));
  OR4X1    g24809(.A(new_n24403_), .B(new_n25001_), .C(new_n24254_), .D(new_n24218_), .Y(new_n25002_));
  OR2X1    g24810(.A(new_n25001_), .B(new_n24218_), .Y(new_n25003_));
  OAI21X1  g24811(.A0(new_n25003_), .A1(new_n24403_), .B0(new_n24254_), .Y(new_n25004_));
  AND2X1   g24812(.A(new_n25004_), .B(new_n25002_), .Y(new_n25005_));
  INVX1    g24813(.A(new_n25005_), .Y(new_n25006_));
  AOI21X1  g24814(.A0(new_n24990_), .A1(new_n24981_), .B0(new_n24997_), .Y(new_n25007_));
  OAI21X1  g24815(.A0(new_n25007_), .A1(new_n1277_), .B0(new_n1111_), .Y(new_n25008_));
  OAI21X1  g24816(.A0(new_n25008_), .A1(new_n24999_), .B0(new_n25006_), .Y(new_n25009_));
  AOI21X1  g24817(.A0(new_n25009_), .A1(new_n25000_), .B0(new_n968_), .Y(new_n25010_));
  OR4X1    g24818(.A(new_n24403_), .B(new_n24232_), .C(new_n24258_), .D(new_n24257_), .Y(new_n25011_));
  OR2X1    g24819(.A(new_n24232_), .B(new_n24257_), .Y(new_n25012_));
  OAI21X1  g24820(.A0(new_n25012_), .A1(new_n24403_), .B0(new_n24258_), .Y(new_n25013_));
  AND2X1   g24821(.A(new_n25013_), .B(new_n25011_), .Y(new_n25014_));
  INVX1    g24822(.A(new_n25014_), .Y(new_n25015_));
  NAND3X1  g24823(.A(new_n25009_), .B(new_n25000_), .C(new_n968_), .Y(new_n25016_));
  AOI21X1  g24824(.A0(new_n25016_), .A1(new_n25015_), .B0(new_n25010_), .Y(new_n25017_));
  OR2X1    g24825(.A(new_n25017_), .B(new_n902_), .Y(new_n25018_));
  AND2X1   g24826(.A(new_n25016_), .B(new_n25015_), .Y(new_n25019_));
  OAI21X1  g24827(.A0(new_n24276_), .A1(new_n24274_), .B0(new_n24240_), .Y(new_n25020_));
  NOR3X1   g24828(.A(new_n25020_), .B(new_n24403_), .C(new_n24234_), .Y(new_n25021_));
  AOI22X1  g24829(.A0(new_n24241_), .A1(new_n24235_), .B0(new_n24233_), .B1(\asqrt[53] ), .Y(new_n25022_));
  AOI21X1  g24830(.A0(new_n25022_), .A1(\asqrt[2] ), .B0(new_n24240_), .Y(new_n25023_));
  NOR2X1   g24831(.A(new_n25023_), .B(new_n25021_), .Y(new_n25024_));
  INVX1    g24832(.A(new_n25024_), .Y(new_n25025_));
  OR2X1    g24833(.A(new_n25010_), .B(\asqrt[54] ), .Y(new_n25026_));
  OAI21X1  g24834(.A0(new_n25026_), .A1(new_n25019_), .B0(new_n25025_), .Y(new_n25027_));
  AOI21X1  g24835(.A0(new_n25027_), .A1(new_n25018_), .B0(new_n697_), .Y(new_n25028_));
  AND2X1   g24836(.A(new_n24279_), .B(new_n24277_), .Y(new_n25029_));
  NOR4X1   g24837(.A(new_n24403_), .B(new_n25029_), .C(new_n24248_), .D(new_n24278_), .Y(new_n25030_));
  NOR2X1   g24838(.A(new_n25029_), .B(new_n24278_), .Y(new_n25031_));
  AOI21X1  g24839(.A0(new_n25031_), .A1(\asqrt[2] ), .B0(new_n24247_), .Y(new_n25032_));
  NOR2X1   g24840(.A(new_n25032_), .B(new_n25030_), .Y(new_n25033_));
  OR2X1    g24841(.A(new_n25007_), .B(new_n1277_), .Y(new_n25034_));
  AND2X1   g24842(.A(new_n24990_), .B(new_n24981_), .Y(new_n25035_));
  INVX1    g24843(.A(new_n24996_), .Y(new_n25036_));
  OR2X1    g24844(.A(new_n24997_), .B(\asqrt[51] ), .Y(new_n25037_));
  OAI21X1  g24845(.A0(new_n25037_), .A1(new_n25035_), .B0(new_n25036_), .Y(new_n25038_));
  AOI21X1  g24846(.A0(new_n25038_), .A1(new_n25034_), .B0(new_n1111_), .Y(new_n25039_));
  AOI21X1  g24847(.A0(new_n24979_), .A1(\asqrt[51] ), .B0(\asqrt[52] ), .Y(new_n25040_));
  AOI21X1  g24848(.A0(new_n25040_), .A1(new_n25038_), .B0(new_n25005_), .Y(new_n25041_));
  OAI21X1  g24849(.A0(new_n25041_), .A1(new_n25039_), .B0(\asqrt[53] ), .Y(new_n25042_));
  NOR3X1   g24850(.A(new_n25041_), .B(new_n25039_), .C(\asqrt[53] ), .Y(new_n25043_));
  OAI21X1  g24851(.A0(new_n25043_), .A1(new_n25014_), .B0(new_n25042_), .Y(new_n25044_));
  AOI21X1  g24852(.A0(new_n25044_), .A1(\asqrt[54] ), .B0(\asqrt[55] ), .Y(new_n25045_));
  AOI21X1  g24853(.A0(new_n25045_), .A1(new_n25027_), .B0(new_n25033_), .Y(new_n25046_));
  OAI21X1  g24854(.A0(new_n25046_), .A1(new_n25028_), .B0(\asqrt[56] ), .Y(new_n25047_));
  NAND3X1  g24855(.A(new_n24270_), .B(new_n24268_), .C(new_n24289_), .Y(new_n25048_));
  NOR3X1   g24856(.A(new_n24403_), .B(new_n24281_), .C(new_n24263_), .Y(new_n25049_));
  OAI22X1  g24857(.A0(new_n25049_), .A1(new_n24268_), .B0(new_n25048_), .B1(new_n24403_), .Y(new_n25050_));
  INVX1    g24858(.A(new_n25050_), .Y(new_n25051_));
  NOR3X1   g24859(.A(new_n25046_), .B(new_n25028_), .C(\asqrt[56] ), .Y(new_n25052_));
  OAI21X1  g24860(.A0(new_n25052_), .A1(new_n25051_), .B0(new_n25047_), .Y(new_n25053_));
  AND2X1   g24861(.A(new_n25053_), .B(\asqrt[57] ), .Y(new_n25054_));
  AND2X1   g24862(.A(new_n25044_), .B(\asqrt[54] ), .Y(new_n25055_));
  NAND2X1  g24863(.A(new_n25016_), .B(new_n25015_), .Y(new_n25056_));
  NOR2X1   g24864(.A(new_n25010_), .B(\asqrt[54] ), .Y(new_n25057_));
  AOI21X1  g24865(.A0(new_n25057_), .A1(new_n25056_), .B0(new_n25024_), .Y(new_n25058_));
  OAI21X1  g24866(.A0(new_n25058_), .A1(new_n25055_), .B0(\asqrt[55] ), .Y(new_n25059_));
  INVX1    g24867(.A(new_n25033_), .Y(new_n25060_));
  OAI21X1  g24868(.A0(new_n25017_), .A1(new_n902_), .B0(new_n697_), .Y(new_n25061_));
  OAI21X1  g24869(.A0(new_n25061_), .A1(new_n25058_), .B0(new_n25060_), .Y(new_n25062_));
  NAND3X1  g24870(.A(new_n25062_), .B(new_n25059_), .C(new_n582_), .Y(new_n25063_));
  NAND2X1  g24871(.A(new_n25063_), .B(new_n25050_), .Y(new_n25064_));
  AND2X1   g24872(.A(new_n24325_), .B(new_n24324_), .Y(new_n25065_));
  NOR4X1   g24873(.A(new_n24403_), .B(new_n25065_), .C(new_n24288_), .D(new_n24323_), .Y(new_n25066_));
  AOI22X1  g24874(.A0(new_n24325_), .A1(new_n24324_), .B0(new_n24297_), .B1(\asqrt[56] ), .Y(new_n25067_));
  AOI21X1  g24875(.A0(new_n25067_), .A1(\asqrt[2] ), .B0(new_n24287_), .Y(new_n25068_));
  NOR2X1   g24876(.A(new_n25068_), .B(new_n25066_), .Y(new_n25069_));
  AOI21X1  g24877(.A0(new_n25062_), .A1(new_n25059_), .B0(new_n582_), .Y(new_n25070_));
  NOR2X1   g24878(.A(new_n25070_), .B(\asqrt[57] ), .Y(new_n25071_));
  AOI21X1  g24879(.A0(new_n25071_), .A1(new_n25064_), .B0(new_n25069_), .Y(new_n25072_));
  OAI21X1  g24880(.A0(new_n25072_), .A1(new_n25054_), .B0(\asqrt[58] ), .Y(new_n25073_));
  AND2X1   g24881(.A(new_n24298_), .B(new_n24291_), .Y(new_n25074_));
  OR4X1    g24882(.A(new_n24403_), .B(new_n25074_), .C(new_n24328_), .D(new_n24292_), .Y(new_n25075_));
  OR2X1    g24883(.A(new_n25074_), .B(new_n24292_), .Y(new_n25076_));
  OAI21X1  g24884(.A0(new_n25076_), .A1(new_n24403_), .B0(new_n24328_), .Y(new_n25077_));
  AND2X1   g24885(.A(new_n25077_), .B(new_n25075_), .Y(new_n25078_));
  INVX1    g24886(.A(new_n25078_), .Y(new_n25079_));
  AOI21X1  g24887(.A0(new_n25063_), .A1(new_n25050_), .B0(new_n25070_), .Y(new_n25080_));
  OAI21X1  g24888(.A0(new_n25080_), .A1(new_n481_), .B0(new_n399_), .Y(new_n25081_));
  OAI21X1  g24889(.A0(new_n25081_), .A1(new_n25072_), .B0(new_n25079_), .Y(new_n25082_));
  AOI21X1  g24890(.A0(new_n25082_), .A1(new_n25073_), .B0(new_n328_), .Y(new_n25083_));
  OR4X1    g24891(.A(new_n24403_), .B(new_n24306_), .C(new_n24332_), .D(new_n24331_), .Y(new_n25084_));
  OR2X1    g24892(.A(new_n24306_), .B(new_n24331_), .Y(new_n25085_));
  OAI21X1  g24893(.A0(new_n25085_), .A1(new_n24403_), .B0(new_n24332_), .Y(new_n25086_));
  AND2X1   g24894(.A(new_n25086_), .B(new_n25084_), .Y(new_n25087_));
  INVX1    g24895(.A(new_n25087_), .Y(new_n25088_));
  NAND3X1  g24896(.A(new_n25082_), .B(new_n25073_), .C(new_n328_), .Y(new_n25089_));
  AOI21X1  g24897(.A0(new_n25089_), .A1(new_n25088_), .B0(new_n25083_), .Y(new_n25090_));
  OR2X1    g24898(.A(new_n25090_), .B(new_n292_), .Y(new_n25091_));
  AND2X1   g24899(.A(new_n25089_), .B(new_n25088_), .Y(new_n25092_));
  OAI21X1  g24900(.A0(new_n24350_), .A1(new_n24348_), .B0(new_n24314_), .Y(new_n25093_));
  NOR3X1   g24901(.A(new_n25093_), .B(new_n24403_), .C(new_n24308_), .Y(new_n25094_));
  AOI22X1  g24902(.A0(new_n24315_), .A1(new_n24309_), .B0(new_n24307_), .B1(\asqrt[59] ), .Y(new_n25095_));
  AOI21X1  g24903(.A0(new_n25095_), .A1(\asqrt[2] ), .B0(new_n24314_), .Y(new_n25096_));
  NOR2X1   g24904(.A(new_n25096_), .B(new_n25094_), .Y(new_n25097_));
  INVX1    g24905(.A(new_n25097_), .Y(new_n25098_));
  OR2X1    g24906(.A(new_n25083_), .B(\asqrt[60] ), .Y(new_n25099_));
  OAI21X1  g24907(.A0(new_n25099_), .A1(new_n25092_), .B0(new_n25098_), .Y(new_n25100_));
  AOI21X1  g24908(.A0(new_n25100_), .A1(new_n25091_), .B0(new_n217_), .Y(new_n25101_));
  AND2X1   g24909(.A(new_n24353_), .B(new_n24351_), .Y(new_n25102_));
  OR4X1    g24910(.A(new_n24403_), .B(new_n25102_), .C(new_n24322_), .D(new_n24352_), .Y(new_n25103_));
  OR2X1    g24911(.A(new_n25102_), .B(new_n24352_), .Y(new_n25104_));
  OAI21X1  g24912(.A0(new_n25104_), .A1(new_n24403_), .B0(new_n24322_), .Y(new_n25105_));
  AND2X1   g24913(.A(new_n25105_), .B(new_n25103_), .Y(new_n25106_));
  OR2X1    g24914(.A(new_n25080_), .B(new_n481_), .Y(new_n25107_));
  AND2X1   g24915(.A(new_n25063_), .B(new_n25050_), .Y(new_n25108_));
  INVX1    g24916(.A(new_n25069_), .Y(new_n25109_));
  OR2X1    g24917(.A(new_n25070_), .B(\asqrt[57] ), .Y(new_n25110_));
  OAI21X1  g24918(.A0(new_n25110_), .A1(new_n25108_), .B0(new_n25109_), .Y(new_n25111_));
  AOI21X1  g24919(.A0(new_n25111_), .A1(new_n25107_), .B0(new_n399_), .Y(new_n25112_));
  AOI21X1  g24920(.A0(new_n25053_), .A1(\asqrt[57] ), .B0(\asqrt[58] ), .Y(new_n25113_));
  AOI21X1  g24921(.A0(new_n25113_), .A1(new_n25111_), .B0(new_n25078_), .Y(new_n25114_));
  OAI21X1  g24922(.A0(new_n25114_), .A1(new_n25112_), .B0(\asqrt[59] ), .Y(new_n25115_));
  NOR3X1   g24923(.A(new_n25114_), .B(new_n25112_), .C(\asqrt[59] ), .Y(new_n25116_));
  OAI21X1  g24924(.A0(new_n25116_), .A1(new_n25087_), .B0(new_n25115_), .Y(new_n25117_));
  AOI21X1  g24925(.A0(new_n25117_), .A1(\asqrt[60] ), .B0(\asqrt[61] ), .Y(new_n25118_));
  AOI21X1  g24926(.A0(new_n25118_), .A1(new_n25100_), .B0(new_n25106_), .Y(new_n25119_));
  OAI21X1  g24927(.A0(new_n25119_), .A1(new_n25101_), .B0(\asqrt[62] ), .Y(new_n25120_));
  NAND3X1  g24928(.A(new_n24344_), .B(new_n24342_), .C(new_n24357_), .Y(new_n25121_));
  NOR3X1   g24929(.A(new_n24403_), .B(new_n24355_), .C(new_n24337_), .Y(new_n25122_));
  OAI22X1  g24930(.A0(new_n25122_), .A1(new_n24342_), .B0(new_n25121_), .B1(new_n24403_), .Y(new_n25123_));
  INVX1    g24931(.A(new_n25123_), .Y(new_n25124_));
  NOR3X1   g24932(.A(new_n25119_), .B(new_n25101_), .C(\asqrt[62] ), .Y(new_n25125_));
  OAI21X1  g24933(.A0(new_n25125_), .A1(new_n25124_), .B0(new_n25120_), .Y(new_n25126_));
  AND2X1   g24934(.A(new_n24398_), .B(new_n24397_), .Y(new_n25127_));
  OR4X1    g24935(.A(new_n24403_), .B(new_n24364_), .C(new_n25127_), .D(new_n24396_), .Y(new_n25128_));
  OAI22X1  g24936(.A0(new_n24358_), .A1(new_n24356_), .B0(new_n24345_), .B1(new_n199_), .Y(new_n25129_));
  OAI21X1  g24937(.A0(new_n25129_), .A1(new_n24403_), .B0(new_n24364_), .Y(new_n25130_));
  NAND2X1  g24938(.A(new_n25130_), .B(new_n25128_), .Y(new_n25131_));
  AOI21X1  g24939(.A0(new_n24365_), .A1(new_n24346_), .B0(new_n24369_), .Y(new_n25132_));
  AOI22X1  g24940(.A0(new_n25132_), .A1(\asqrt[2] ), .B0(new_n24376_), .B1(new_n24365_), .Y(new_n25133_));
  AND2X1   g24941(.A(new_n25133_), .B(new_n25131_), .Y(new_n25134_));
  AOI21X1  g24942(.A0(new_n25134_), .A1(new_n25126_), .B0(\asqrt[63] ), .Y(new_n25135_));
  AND2X1   g24943(.A(new_n25117_), .B(\asqrt[60] ), .Y(new_n25136_));
  NAND2X1  g24944(.A(new_n25089_), .B(new_n25088_), .Y(new_n25137_));
  NOR2X1   g24945(.A(new_n25083_), .B(\asqrt[60] ), .Y(new_n25138_));
  AOI21X1  g24946(.A0(new_n25138_), .A1(new_n25137_), .B0(new_n25097_), .Y(new_n25139_));
  OAI21X1  g24947(.A0(new_n25139_), .A1(new_n25136_), .B0(\asqrt[61] ), .Y(new_n25140_));
  INVX1    g24948(.A(new_n25106_), .Y(new_n25141_));
  OAI21X1  g24949(.A0(new_n25090_), .A1(new_n292_), .B0(new_n217_), .Y(new_n25142_));
  OAI21X1  g24950(.A0(new_n25142_), .A1(new_n25139_), .B0(new_n25141_), .Y(new_n25143_));
  NAND3X1  g24951(.A(new_n25143_), .B(new_n25140_), .C(new_n199_), .Y(new_n25144_));
  AND2X1   g24952(.A(new_n25144_), .B(new_n25123_), .Y(new_n25145_));
  AOI21X1  g24953(.A0(new_n25143_), .A1(new_n25140_), .B0(new_n199_), .Y(new_n25146_));
  OR2X1    g24954(.A(new_n25131_), .B(new_n25146_), .Y(new_n25147_));
  AND2X1   g24955(.A(new_n24365_), .B(new_n24346_), .Y(new_n25148_));
  OAI21X1  g24956(.A0(new_n24403_), .A1(new_n24369_), .B0(new_n25148_), .Y(new_n25149_));
  NOR2X1   g24957(.A(new_n25132_), .B(new_n193_), .Y(new_n25150_));
  AND2X1   g24958(.A(new_n25150_), .B(new_n25149_), .Y(new_n25151_));
  INVX1    g24959(.A(new_n25151_), .Y(new_n25152_));
  OAI21X1  g24960(.A0(new_n25147_), .A1(new_n25145_), .B0(new_n25152_), .Y(new_n25153_));
  OAI21X1  g24961(.A0(new_n25153_), .A1(new_n25135_), .B0(new_n23625_), .Y(new_n25154_));
  NAND2X1  g24962(.A(new_n25144_), .B(new_n25123_), .Y(new_n25155_));
  NOR2X1   g24963(.A(new_n25131_), .B(new_n25146_), .Y(new_n25156_));
  AND2X1   g24964(.A(new_n25156_), .B(new_n25155_), .Y(new_n25157_));
  OR4X1    g24965(.A(new_n25151_), .B(new_n25157_), .C(new_n25135_), .D(new_n24403_), .Y(new_n25158_));
  AOI21X1  g24966(.A0(new_n25158_), .A1(new_n25154_), .B0(new_n23624_), .Y(new_n25159_));
  AOI21X1  g24967(.A0(new_n25144_), .A1(new_n25123_), .B0(new_n25146_), .Y(new_n25160_));
  INVX1    g24968(.A(new_n25134_), .Y(new_n25161_));
  OAI21X1  g24969(.A0(new_n25161_), .A1(new_n25160_), .B0(new_n193_), .Y(new_n25162_));
  AOI21X1  g24970(.A0(new_n25156_), .A1(new_n25155_), .B0(new_n25151_), .Y(new_n25163_));
  AOI21X1  g24971(.A0(new_n25163_), .A1(new_n25162_), .B0(new_n24395_), .Y(new_n25164_));
  NOR4X1   g24972(.A(new_n25151_), .B(new_n25157_), .C(new_n25135_), .D(new_n24403_), .Y(new_n25165_));
  NOR3X1   g24973(.A(new_n25165_), .B(new_n25164_), .C(\a[4] ), .Y(new_n25166_));
  NOR2X1   g24974(.A(new_n25166_), .B(new_n25159_), .Y(new_n25167_));
  INVX1    g24975(.A(\a[2] ), .Y(new_n25168_));
  OAI21X1  g24976(.A0(new_n25153_), .A1(new_n25135_), .B0(new_n25168_), .Y(new_n25169_));
  NAND2X1  g24977(.A(new_n25169_), .B(\a[3] ), .Y(new_n25170_));
  OAI21X1  g24978(.A0(\a[1] ), .A1(\a[0] ), .B0(new_n25168_), .Y(new_n25171_));
  INVX1    g24979(.A(new_n25171_), .Y(new_n25172_));
  AOI21X1  g24980(.A0(new_n25150_), .A1(new_n25149_), .B0(new_n25168_), .Y(new_n25173_));
  INVX1    g24981(.A(new_n25173_), .Y(new_n25174_));
  AOI21X1  g24982(.A0(new_n25156_), .A1(new_n25155_), .B0(new_n25174_), .Y(new_n25175_));
  AOI21X1  g24983(.A0(new_n25175_), .A1(new_n25162_), .B0(new_n25172_), .Y(new_n25176_));
  AND2X1   g24984(.A(new_n25176_), .B(new_n25154_), .Y(new_n25177_));
  AOI21X1  g24985(.A0(new_n25177_), .A1(new_n25170_), .B0(\asqrt[2] ), .Y(new_n25178_));
  AOI21X1  g24986(.A0(new_n25170_), .A1(new_n25154_), .B0(new_n25176_), .Y(new_n25179_));
  NOR3X1   g24987(.A(new_n25179_), .B(new_n25178_), .C(new_n25167_), .Y(new_n25180_));
  OR2X1    g24988(.A(new_n25180_), .B(\asqrt[3] ), .Y(new_n25181_));
  AND2X1   g24989(.A(new_n24444_), .B(new_n24442_), .Y(new_n25182_));
  NOR3X1   g24990(.A(new_n25182_), .B(new_n24388_), .C(new_n24384_), .Y(new_n25183_));
  OAI21X1  g24991(.A0(new_n25153_), .A1(new_n25135_), .B0(new_n25183_), .Y(new_n25184_));
  AOI21X1  g24992(.A0(new_n24383_), .A1(\asqrt[3] ), .B0(new_n24388_), .Y(new_n25185_));
  OAI21X1  g24993(.A0(new_n25153_), .A1(new_n25135_), .B0(new_n25185_), .Y(new_n25186_));
  NAND2X1  g24994(.A(new_n25186_), .B(new_n25182_), .Y(new_n25187_));
  NAND2X1  g24995(.A(new_n25187_), .B(new_n25184_), .Y(new_n25188_));
  OAI21X1  g24996(.A0(new_n25179_), .A1(new_n25178_), .B0(new_n25167_), .Y(new_n25189_));
  AND2X1   g24997(.A(new_n25189_), .B(new_n25188_), .Y(new_n25190_));
  AOI21X1  g24998(.A0(new_n25190_), .A1(new_n25181_), .B0(\asqrt[4] ), .Y(new_n25191_));
  OR2X1    g24999(.A(new_n25166_), .B(new_n25159_), .Y(new_n25192_));
  AND2X1   g25000(.A(new_n25169_), .B(\a[3] ), .Y(new_n25193_));
  OAI21X1  g25001(.A0(new_n25147_), .A1(new_n25145_), .B0(new_n25173_), .Y(new_n25194_));
  OAI21X1  g25002(.A0(new_n25194_), .A1(new_n25135_), .B0(new_n25171_), .Y(new_n25195_));
  OR2X1    g25003(.A(new_n25195_), .B(new_n25164_), .Y(new_n25196_));
  OAI21X1  g25004(.A0(new_n25196_), .A1(new_n25193_), .B0(new_n24403_), .Y(new_n25197_));
  OAI21X1  g25005(.A0(new_n25193_), .A1(new_n25164_), .B0(new_n25195_), .Y(new_n25198_));
  NAND3X1  g25006(.A(new_n25198_), .B(new_n25197_), .C(new_n25192_), .Y(new_n25199_));
  AOI21X1  g25007(.A0(new_n25198_), .A1(new_n25197_), .B0(new_n25192_), .Y(new_n25200_));
  AOI21X1  g25008(.A0(new_n25199_), .A1(new_n23622_), .B0(new_n25200_), .Y(new_n25201_));
  AND2X1   g25009(.A(new_n24447_), .B(new_n24445_), .Y(new_n25202_));
  NOR2X1   g25010(.A(new_n25153_), .B(new_n25135_), .Y(new_n25203_));
  NOR3X1   g25011(.A(new_n25203_), .B(new_n25202_), .C(new_n24446_), .Y(new_n25204_));
  NOR3X1   g25012(.A(new_n24413_), .B(new_n25202_), .C(new_n24446_), .Y(new_n25205_));
  OAI21X1  g25013(.A0(new_n25153_), .A1(new_n25135_), .B0(new_n25205_), .Y(new_n25206_));
  OAI21X1  g25014(.A0(new_n25204_), .A1(new_n24450_), .B0(new_n25206_), .Y(new_n25207_));
  OAI21X1  g25015(.A0(new_n25201_), .A1(new_n25188_), .B0(new_n25207_), .Y(new_n25208_));
  OAI21X1  g25016(.A0(new_n25208_), .A1(new_n25191_), .B0(new_n22128_), .Y(new_n25209_));
  INVX1    g25017(.A(new_n25203_), .Y(\asqrt[1] ));
  NOR3X1   g25018(.A(new_n24453_), .B(new_n24421_), .C(new_n24415_), .Y(new_n25211_));
  NAND3X1  g25019(.A(\asqrt[1] ), .B(new_n24422_), .C(new_n24452_), .Y(new_n25212_));
  AOI22X1  g25020(.A0(new_n25212_), .A1(new_n24421_), .B0(new_n25211_), .B1(\asqrt[1] ), .Y(new_n25213_));
  INVX1    g25021(.A(new_n25213_), .Y(new_n25214_));
  INVX1    g25022(.A(new_n25188_), .Y(new_n25215_));
  OAI21X1  g25023(.A0(new_n25180_), .A1(\asqrt[3] ), .B0(new_n25189_), .Y(new_n25216_));
  AND2X1   g25024(.A(new_n25216_), .B(new_n25215_), .Y(new_n25217_));
  INVX1    g25025(.A(new_n25207_), .Y(new_n25218_));
  OAI21X1  g25026(.A0(new_n25217_), .A1(new_n25191_), .B0(new_n25218_), .Y(new_n25219_));
  NAND3X1  g25027(.A(new_n25219_), .B(new_n25214_), .C(new_n25209_), .Y(new_n25220_));
  NAND2X1  g25028(.A(new_n25220_), .B(new_n21393_), .Y(new_n25221_));
  AOI21X1  g25029(.A0(new_n25219_), .A1(new_n25209_), .B0(new_n25214_), .Y(new_n25222_));
  AOI22X1  g25030(.A0(new_n24468_), .A1(new_n24467_), .B0(new_n24454_), .B1(\asqrt[6] ), .Y(new_n25223_));
  AOI21X1  g25031(.A0(new_n25223_), .A1(\asqrt[1] ), .B0(new_n24430_), .Y(new_n25224_));
  OAI21X1  g25032(.A0(new_n24432_), .A1(new_n24425_), .B0(new_n24430_), .Y(new_n25225_));
  NOR2X1   g25033(.A(new_n25225_), .B(new_n24466_), .Y(new_n25226_));
  AOI21X1  g25034(.A0(new_n25226_), .A1(\asqrt[1] ), .B0(new_n25224_), .Y(new_n25227_));
  NOR2X1   g25035(.A(new_n25227_), .B(new_n25222_), .Y(new_n25228_));
  AOI21X1  g25036(.A0(new_n25228_), .A1(new_n25221_), .B0(\asqrt[7] ), .Y(new_n25229_));
  INVX1    g25037(.A(new_n25227_), .Y(new_n25230_));
  AND2X1   g25038(.A(new_n24455_), .B(new_n24433_), .Y(new_n25231_));
  OR2X1    g25039(.A(new_n25231_), .B(new_n24434_), .Y(new_n25232_));
  OAI21X1  g25040(.A0(new_n25232_), .A1(new_n25203_), .B0(new_n24471_), .Y(new_n25233_));
  OR4X1    g25041(.A(new_n25203_), .B(new_n25231_), .C(new_n24471_), .D(new_n24434_), .Y(new_n25234_));
  AND2X1   g25042(.A(new_n25234_), .B(new_n25233_), .Y(new_n25235_));
  INVX1    g25043(.A(new_n25235_), .Y(new_n25236_));
  AOI21X1  g25044(.A0(new_n25220_), .A1(new_n21393_), .B0(new_n25222_), .Y(new_n25237_));
  OAI21X1  g25045(.A0(new_n25237_), .A1(new_n25230_), .B0(new_n25236_), .Y(new_n25238_));
  OAI21X1  g25046(.A0(new_n25238_), .A1(new_n25229_), .B0(new_n19976_), .Y(new_n25239_));
  AND2X1   g25047(.A(new_n25199_), .B(new_n23622_), .Y(new_n25240_));
  NAND2X1  g25048(.A(new_n25189_), .B(new_n25188_), .Y(new_n25241_));
  OAI21X1  g25049(.A0(new_n25241_), .A1(new_n25240_), .B0(new_n22874_), .Y(new_n25242_));
  AOI21X1  g25050(.A0(new_n25216_), .A1(new_n25215_), .B0(new_n25218_), .Y(new_n25243_));
  AOI21X1  g25051(.A0(new_n25243_), .A1(new_n25242_), .B0(\asqrt[5] ), .Y(new_n25244_));
  OR2X1    g25052(.A(new_n25201_), .B(new_n25188_), .Y(new_n25245_));
  AOI21X1  g25053(.A0(new_n25245_), .A1(new_n25242_), .B0(new_n25207_), .Y(new_n25246_));
  NOR3X1   g25054(.A(new_n25246_), .B(new_n25213_), .C(new_n25244_), .Y(new_n25247_));
  OAI21X1  g25055(.A0(new_n25246_), .A1(new_n25244_), .B0(new_n25213_), .Y(new_n25248_));
  OAI21X1  g25056(.A0(new_n25247_), .A1(\asqrt[6] ), .B0(new_n25248_), .Y(new_n25249_));
  AND2X1   g25057(.A(new_n25249_), .B(new_n25227_), .Y(new_n25250_));
  OAI21X1  g25058(.A0(new_n25250_), .A1(new_n25229_), .B0(new_n25235_), .Y(new_n25251_));
  NOR3X1   g25059(.A(new_n25203_), .B(new_n24462_), .C(new_n24481_), .Y(new_n25252_));
  NOR2X1   g25060(.A(new_n25252_), .B(new_n24461_), .Y(new_n25253_));
  NOR3X1   g25061(.A(new_n24462_), .B(new_n24465_), .C(new_n24481_), .Y(new_n25254_));
  AOI21X1  g25062(.A0(new_n25254_), .A1(\asqrt[1] ), .B0(new_n25253_), .Y(new_n25255_));
  INVX1    g25063(.A(new_n25255_), .Y(new_n25256_));
  NAND3X1  g25064(.A(new_n25256_), .B(new_n25251_), .C(new_n25239_), .Y(new_n25257_));
  NAND2X1  g25065(.A(new_n25257_), .B(new_n19273_), .Y(new_n25258_));
  AND2X1   g25066(.A(new_n24482_), .B(new_n24475_), .Y(new_n25259_));
  NOR3X1   g25067(.A(new_n25203_), .B(new_n25259_), .C(new_n24464_), .Y(new_n25260_));
  NOR2X1   g25068(.A(new_n25260_), .B(new_n24480_), .Y(new_n25261_));
  NOR3X1   g25069(.A(new_n25259_), .B(new_n24520_), .C(new_n24464_), .Y(new_n25262_));
  AOI21X1  g25070(.A0(new_n25262_), .A1(\asqrt[1] ), .B0(new_n25261_), .Y(new_n25263_));
  AOI21X1  g25071(.A0(new_n25251_), .A1(new_n25239_), .B0(new_n25256_), .Y(new_n25264_));
  NOR2X1   g25072(.A(new_n25264_), .B(new_n25263_), .Y(new_n25265_));
  AOI21X1  g25073(.A0(new_n25265_), .A1(new_n25258_), .B0(\asqrt[10] ), .Y(new_n25266_));
  INVX1    g25074(.A(new_n25263_), .Y(new_n25267_));
  AOI21X1  g25075(.A0(new_n25257_), .A1(new_n19273_), .B0(new_n25264_), .Y(new_n25268_));
  AND2X1   g25076(.A(new_n24524_), .B(new_n24522_), .Y(new_n25269_));
  OR2X1    g25077(.A(new_n25269_), .B(new_n24523_), .Y(new_n25270_));
  OAI21X1  g25078(.A0(new_n25270_), .A1(new_n25203_), .B0(new_n24490_), .Y(new_n25271_));
  OR4X1    g25079(.A(new_n25203_), .B(new_n25269_), .C(new_n24490_), .D(new_n24523_), .Y(new_n25272_));
  AND2X1   g25080(.A(new_n25272_), .B(new_n25271_), .Y(new_n25273_));
  INVX1    g25081(.A(new_n25273_), .Y(new_n25274_));
  OAI21X1  g25082(.A0(new_n25268_), .A1(new_n25267_), .B0(new_n25274_), .Y(new_n25275_));
  OAI21X1  g25083(.A0(new_n25275_), .A1(new_n25266_), .B0(new_n17927_), .Y(new_n25276_));
  NOR3X1   g25084(.A(new_n25203_), .B(new_n24527_), .C(new_n24494_), .Y(new_n25277_));
  NOR2X1   g25085(.A(new_n25277_), .B(new_n24498_), .Y(new_n25278_));
  NOR3X1   g25086(.A(new_n24527_), .B(new_n24499_), .C(new_n24494_), .Y(new_n25279_));
  AOI21X1  g25087(.A0(new_n25279_), .A1(\asqrt[1] ), .B0(new_n25278_), .Y(new_n25280_));
  INVX1    g25088(.A(new_n25280_), .Y(new_n25281_));
  AND2X1   g25089(.A(new_n25220_), .B(new_n21393_), .Y(new_n25282_));
  OR2X1    g25090(.A(new_n25227_), .B(new_n25222_), .Y(new_n25283_));
  OAI21X1  g25091(.A0(new_n25283_), .A1(new_n25282_), .B0(new_n20676_), .Y(new_n25284_));
  AOI21X1  g25092(.A0(new_n25249_), .A1(new_n25227_), .B0(new_n25235_), .Y(new_n25285_));
  AOI21X1  g25093(.A0(new_n25285_), .A1(new_n25284_), .B0(\asqrt[8] ), .Y(new_n25286_));
  OR2X1    g25094(.A(new_n25237_), .B(new_n25230_), .Y(new_n25287_));
  AOI21X1  g25095(.A0(new_n25287_), .A1(new_n25284_), .B0(new_n25236_), .Y(new_n25288_));
  NOR3X1   g25096(.A(new_n25255_), .B(new_n25288_), .C(new_n25286_), .Y(new_n25289_));
  OAI21X1  g25097(.A0(new_n25288_), .A1(new_n25286_), .B0(new_n25255_), .Y(new_n25290_));
  OAI21X1  g25098(.A0(new_n25289_), .A1(\asqrt[9] ), .B0(new_n25290_), .Y(new_n25291_));
  AND2X1   g25099(.A(new_n25291_), .B(new_n25263_), .Y(new_n25292_));
  OAI21X1  g25100(.A0(new_n25292_), .A1(new_n25266_), .B0(new_n25273_), .Y(new_n25293_));
  NAND3X1  g25101(.A(new_n25293_), .B(new_n25281_), .C(new_n25276_), .Y(new_n25294_));
  NAND2X1  g25102(.A(new_n25294_), .B(new_n17262_), .Y(new_n25295_));
  AOI21X1  g25103(.A0(new_n25293_), .A1(new_n25276_), .B0(new_n25281_), .Y(new_n25296_));
  AOI22X1  g25104(.A0(new_n24543_), .A1(new_n24541_), .B0(new_n24528_), .B1(\asqrt[12] ), .Y(new_n25297_));
  AOI21X1  g25105(.A0(new_n25297_), .A1(\asqrt[1] ), .B0(new_n24542_), .Y(new_n25298_));
  OAI21X1  g25106(.A0(new_n24509_), .A1(new_n24503_), .B0(new_n24542_), .Y(new_n25299_));
  NOR2X1   g25107(.A(new_n25299_), .B(new_n24540_), .Y(new_n25300_));
  AOI21X1  g25108(.A0(new_n25300_), .A1(\asqrt[1] ), .B0(new_n25298_), .Y(new_n25301_));
  NOR2X1   g25109(.A(new_n25301_), .B(new_n25296_), .Y(new_n25302_));
  AOI21X1  g25110(.A0(new_n25302_), .A1(new_n25295_), .B0(\asqrt[13] ), .Y(new_n25303_));
  INVX1    g25111(.A(new_n25301_), .Y(new_n25304_));
  AND2X1   g25112(.A(new_n24529_), .B(new_n24510_), .Y(new_n25305_));
  OR2X1    g25113(.A(new_n25305_), .B(new_n24511_), .Y(new_n25306_));
  OAI21X1  g25114(.A0(new_n25306_), .A1(new_n25203_), .B0(new_n24546_), .Y(new_n25307_));
  OR4X1    g25115(.A(new_n25203_), .B(new_n25305_), .C(new_n24546_), .D(new_n24511_), .Y(new_n25308_));
  AND2X1   g25116(.A(new_n25308_), .B(new_n25307_), .Y(new_n25309_));
  INVX1    g25117(.A(new_n25309_), .Y(new_n25310_));
  AOI21X1  g25118(.A0(new_n25294_), .A1(new_n17262_), .B0(new_n25296_), .Y(new_n25311_));
  OAI21X1  g25119(.A0(new_n25311_), .A1(new_n25304_), .B0(new_n25310_), .Y(new_n25312_));
  OAI21X1  g25120(.A0(new_n25312_), .A1(new_n25303_), .B0(new_n15990_), .Y(new_n25313_));
  AND2X1   g25121(.A(new_n25257_), .B(new_n19273_), .Y(new_n25314_));
  OR2X1    g25122(.A(new_n25264_), .B(new_n25263_), .Y(new_n25315_));
  OAI21X1  g25123(.A0(new_n25315_), .A1(new_n25314_), .B0(new_n18591_), .Y(new_n25316_));
  AOI21X1  g25124(.A0(new_n25291_), .A1(new_n25263_), .B0(new_n25273_), .Y(new_n25317_));
  AOI21X1  g25125(.A0(new_n25317_), .A1(new_n25316_), .B0(\asqrt[11] ), .Y(new_n25318_));
  OR2X1    g25126(.A(new_n25268_), .B(new_n25267_), .Y(new_n25319_));
  AOI21X1  g25127(.A0(new_n25319_), .A1(new_n25316_), .B0(new_n25274_), .Y(new_n25320_));
  NOR3X1   g25128(.A(new_n25320_), .B(new_n25280_), .C(new_n25318_), .Y(new_n25321_));
  OAI21X1  g25129(.A0(new_n25320_), .A1(new_n25318_), .B0(new_n25280_), .Y(new_n25322_));
  OAI21X1  g25130(.A0(new_n25321_), .A1(\asqrt[12] ), .B0(new_n25322_), .Y(new_n25323_));
  AND2X1   g25131(.A(new_n25323_), .B(new_n25301_), .Y(new_n25324_));
  OAI21X1  g25132(.A0(new_n25324_), .A1(new_n25303_), .B0(new_n25309_), .Y(new_n25325_));
  NOR3X1   g25133(.A(new_n25203_), .B(new_n24536_), .C(new_n24556_), .Y(new_n25326_));
  NOR2X1   g25134(.A(new_n25326_), .B(new_n24535_), .Y(new_n25327_));
  NOR3X1   g25135(.A(new_n24536_), .B(new_n24539_), .C(new_n24556_), .Y(new_n25328_));
  AOI21X1  g25136(.A0(new_n25328_), .A1(\asqrt[1] ), .B0(new_n25327_), .Y(new_n25329_));
  INVX1    g25137(.A(new_n25329_), .Y(new_n25330_));
  NAND3X1  g25138(.A(new_n25330_), .B(new_n25325_), .C(new_n25313_), .Y(new_n25331_));
  NAND2X1  g25139(.A(new_n25331_), .B(new_n15362_), .Y(new_n25332_));
  AND2X1   g25140(.A(new_n24557_), .B(new_n24550_), .Y(new_n25333_));
  NOR3X1   g25141(.A(new_n25203_), .B(new_n25333_), .C(new_n24538_), .Y(new_n25334_));
  NOR2X1   g25142(.A(new_n25334_), .B(new_n24555_), .Y(new_n25335_));
  NOR3X1   g25143(.A(new_n25333_), .B(new_n24595_), .C(new_n24538_), .Y(new_n25336_));
  AOI21X1  g25144(.A0(new_n25336_), .A1(\asqrt[1] ), .B0(new_n25335_), .Y(new_n25337_));
  AOI21X1  g25145(.A0(new_n25325_), .A1(new_n25313_), .B0(new_n25330_), .Y(new_n25338_));
  NOR2X1   g25146(.A(new_n25338_), .B(new_n25337_), .Y(new_n25339_));
  AOI21X1  g25147(.A0(new_n25339_), .A1(new_n25332_), .B0(\asqrt[16] ), .Y(new_n25340_));
  INVX1    g25148(.A(new_n25337_), .Y(new_n25341_));
  AOI21X1  g25149(.A0(new_n25331_), .A1(new_n15362_), .B0(new_n25338_), .Y(new_n25342_));
  AND2X1   g25150(.A(new_n24599_), .B(new_n24597_), .Y(new_n25343_));
  OR2X1    g25151(.A(new_n25343_), .B(new_n24598_), .Y(new_n25344_));
  OAI21X1  g25152(.A0(new_n25344_), .A1(new_n25203_), .B0(new_n24565_), .Y(new_n25345_));
  OR4X1    g25153(.A(new_n25203_), .B(new_n25343_), .C(new_n24565_), .D(new_n24598_), .Y(new_n25346_));
  AND2X1   g25154(.A(new_n25346_), .B(new_n25345_), .Y(new_n25347_));
  INVX1    g25155(.A(new_n25347_), .Y(new_n25348_));
  OAI21X1  g25156(.A0(new_n25342_), .A1(new_n25341_), .B0(new_n25348_), .Y(new_n25349_));
  OAI21X1  g25157(.A0(new_n25349_), .A1(new_n25340_), .B0(new_n14165_), .Y(new_n25350_));
  NOR3X1   g25158(.A(new_n25203_), .B(new_n24602_), .C(new_n24569_), .Y(new_n25351_));
  NOR2X1   g25159(.A(new_n25351_), .B(new_n24573_), .Y(new_n25352_));
  NOR3X1   g25160(.A(new_n24602_), .B(new_n24574_), .C(new_n24569_), .Y(new_n25353_));
  AOI21X1  g25161(.A0(new_n25353_), .A1(\asqrt[1] ), .B0(new_n25352_), .Y(new_n25354_));
  INVX1    g25162(.A(new_n25354_), .Y(new_n25355_));
  AND2X1   g25163(.A(new_n25294_), .B(new_n17262_), .Y(new_n25356_));
  OR2X1    g25164(.A(new_n25301_), .B(new_n25296_), .Y(new_n25357_));
  OAI21X1  g25165(.A0(new_n25357_), .A1(new_n25356_), .B0(new_n16617_), .Y(new_n25358_));
  AOI21X1  g25166(.A0(new_n25323_), .A1(new_n25301_), .B0(new_n25309_), .Y(new_n25359_));
  AOI21X1  g25167(.A0(new_n25359_), .A1(new_n25358_), .B0(\asqrt[14] ), .Y(new_n25360_));
  OR2X1    g25168(.A(new_n25311_), .B(new_n25304_), .Y(new_n25361_));
  AOI21X1  g25169(.A0(new_n25361_), .A1(new_n25358_), .B0(new_n25310_), .Y(new_n25362_));
  NOR3X1   g25170(.A(new_n25329_), .B(new_n25362_), .C(new_n25360_), .Y(new_n25363_));
  OAI21X1  g25171(.A0(new_n25362_), .A1(new_n25360_), .B0(new_n25329_), .Y(new_n25364_));
  OAI21X1  g25172(.A0(new_n25363_), .A1(\asqrt[15] ), .B0(new_n25364_), .Y(new_n25365_));
  AND2X1   g25173(.A(new_n25365_), .B(new_n25337_), .Y(new_n25366_));
  OAI21X1  g25174(.A0(new_n25366_), .A1(new_n25340_), .B0(new_n25347_), .Y(new_n25367_));
  NAND3X1  g25175(.A(new_n25367_), .B(new_n25355_), .C(new_n25350_), .Y(new_n25368_));
  NAND2X1  g25176(.A(new_n25368_), .B(new_n13571_), .Y(new_n25369_));
  AOI21X1  g25177(.A0(new_n25367_), .A1(new_n25350_), .B0(new_n25355_), .Y(new_n25370_));
  AND2X1   g25178(.A(new_n24616_), .B(new_n24615_), .Y(new_n25371_));
  NOR3X1   g25179(.A(new_n25203_), .B(new_n25371_), .C(new_n24614_), .Y(new_n25372_));
  NOR2X1   g25180(.A(new_n25372_), .B(new_n24583_), .Y(new_n25373_));
  NOR3X1   g25181(.A(new_n25371_), .B(new_n24584_), .C(new_n24614_), .Y(new_n25374_));
  AOI21X1  g25182(.A0(new_n25374_), .A1(\asqrt[1] ), .B0(new_n25373_), .Y(new_n25375_));
  NOR2X1   g25183(.A(new_n25375_), .B(new_n25370_), .Y(new_n25376_));
  AOI21X1  g25184(.A0(new_n25376_), .A1(new_n25369_), .B0(\asqrt[19] ), .Y(new_n25377_));
  INVX1    g25185(.A(new_n25375_), .Y(new_n25378_));
  AND2X1   g25186(.A(new_n24604_), .B(new_n24586_), .Y(new_n25379_));
  OR2X1    g25187(.A(new_n25379_), .B(new_n24587_), .Y(new_n25380_));
  OAI21X1  g25188(.A0(new_n25380_), .A1(new_n25203_), .B0(new_n24619_), .Y(new_n25381_));
  OR4X1    g25189(.A(new_n25203_), .B(new_n25379_), .C(new_n24619_), .D(new_n24587_), .Y(new_n25382_));
  AND2X1   g25190(.A(new_n25382_), .B(new_n25381_), .Y(new_n25383_));
  INVX1    g25191(.A(new_n25383_), .Y(new_n25384_));
  AOI21X1  g25192(.A0(new_n25368_), .A1(new_n13571_), .B0(new_n25370_), .Y(new_n25385_));
  OAI21X1  g25193(.A0(new_n25385_), .A1(new_n25378_), .B0(new_n25384_), .Y(new_n25386_));
  OAI21X1  g25194(.A0(new_n25386_), .A1(new_n25377_), .B0(new_n12447_), .Y(new_n25387_));
  AND2X1   g25195(.A(new_n25331_), .B(new_n15362_), .Y(new_n25388_));
  OR2X1    g25196(.A(new_n25338_), .B(new_n25337_), .Y(new_n25389_));
  OAI21X1  g25197(.A0(new_n25389_), .A1(new_n25388_), .B0(new_n14754_), .Y(new_n25390_));
  AOI21X1  g25198(.A0(new_n25365_), .A1(new_n25337_), .B0(new_n25347_), .Y(new_n25391_));
  AOI21X1  g25199(.A0(new_n25391_), .A1(new_n25390_), .B0(\asqrt[17] ), .Y(new_n25392_));
  OR2X1    g25200(.A(new_n25342_), .B(new_n25341_), .Y(new_n25393_));
  AOI21X1  g25201(.A0(new_n25393_), .A1(new_n25390_), .B0(new_n25348_), .Y(new_n25394_));
  NOR3X1   g25202(.A(new_n25394_), .B(new_n25354_), .C(new_n25392_), .Y(new_n25395_));
  OAI21X1  g25203(.A0(new_n25394_), .A1(new_n25392_), .B0(new_n25354_), .Y(new_n25396_));
  OAI21X1  g25204(.A0(new_n25395_), .A1(\asqrt[18] ), .B0(new_n25396_), .Y(new_n25397_));
  AND2X1   g25205(.A(new_n25397_), .B(new_n25375_), .Y(new_n25398_));
  OAI21X1  g25206(.A0(new_n25398_), .A1(new_n25377_), .B0(new_n25383_), .Y(new_n25399_));
  NOR3X1   g25207(.A(new_n25203_), .B(new_n24611_), .C(new_n24629_), .Y(new_n25400_));
  NOR2X1   g25208(.A(new_n25400_), .B(new_n24610_), .Y(new_n25401_));
  NOR3X1   g25209(.A(new_n24611_), .B(new_n24609_), .C(new_n24629_), .Y(new_n25402_));
  AOI21X1  g25210(.A0(new_n25402_), .A1(\asqrt[1] ), .B0(new_n25401_), .Y(new_n25403_));
  INVX1    g25211(.A(new_n25403_), .Y(new_n25404_));
  NAND3X1  g25212(.A(new_n25404_), .B(new_n25399_), .C(new_n25387_), .Y(new_n25405_));
  NAND2X1  g25213(.A(new_n25405_), .B(new_n11896_), .Y(new_n25406_));
  OAI22X1  g25214(.A0(new_n24670_), .A1(new_n24668_), .B0(new_n24639_), .B1(new_n11896_), .Y(new_n25407_));
  OAI21X1  g25215(.A0(new_n25407_), .A1(new_n25203_), .B0(new_n24669_), .Y(new_n25408_));
  AND2X1   g25216(.A(new_n24630_), .B(new_n24623_), .Y(new_n25409_));
  OR4X1    g25217(.A(new_n25203_), .B(new_n25409_), .C(new_n24669_), .D(new_n24613_), .Y(new_n25410_));
  AND2X1   g25218(.A(new_n25410_), .B(new_n25408_), .Y(new_n25411_));
  AOI21X1  g25219(.A0(new_n25399_), .A1(new_n25387_), .B0(new_n25404_), .Y(new_n25412_));
  NOR2X1   g25220(.A(new_n25412_), .B(new_n25411_), .Y(new_n25413_));
  AOI21X1  g25221(.A0(new_n25413_), .A1(new_n25406_), .B0(\asqrt[22] ), .Y(new_n25414_));
  INVX1    g25222(.A(new_n25411_), .Y(new_n25415_));
  AOI21X1  g25223(.A0(new_n25405_), .A1(new_n11896_), .B0(new_n25412_), .Y(new_n25416_));
  AND2X1   g25224(.A(new_n24673_), .B(new_n24671_), .Y(new_n25417_));
  OR2X1    g25225(.A(new_n25417_), .B(new_n24672_), .Y(new_n25418_));
  OAI21X1  g25226(.A0(new_n25418_), .A1(new_n25203_), .B0(new_n24638_), .Y(new_n25419_));
  OR4X1    g25227(.A(new_n25203_), .B(new_n25417_), .C(new_n24638_), .D(new_n24672_), .Y(new_n25420_));
  AND2X1   g25228(.A(new_n25420_), .B(new_n25419_), .Y(new_n25421_));
  INVX1    g25229(.A(new_n25421_), .Y(new_n25422_));
  OAI21X1  g25230(.A0(new_n25416_), .A1(new_n25415_), .B0(new_n25422_), .Y(new_n25423_));
  OAI21X1  g25231(.A0(new_n25423_), .A1(new_n25414_), .B0(new_n10849_), .Y(new_n25424_));
  NAND2X1  g25232(.A(new_n24648_), .B(new_n24675_), .Y(new_n25425_));
  OAI21X1  g25233(.A0(new_n25425_), .A1(new_n25203_), .B0(new_n24647_), .Y(new_n25426_));
  NAND4X1  g25234(.A(\asqrt[1] ), .B(new_n24648_), .C(new_n24646_), .D(new_n24675_), .Y(new_n25427_));
  AND2X1   g25235(.A(new_n25427_), .B(new_n25426_), .Y(new_n25428_));
  INVX1    g25236(.A(new_n25428_), .Y(new_n25429_));
  AND2X1   g25237(.A(new_n25368_), .B(new_n13571_), .Y(new_n25430_));
  OR2X1    g25238(.A(new_n25375_), .B(new_n25370_), .Y(new_n25431_));
  OAI21X1  g25239(.A0(new_n25431_), .A1(new_n25430_), .B0(new_n13000_), .Y(new_n25432_));
  AOI21X1  g25240(.A0(new_n25397_), .A1(new_n25375_), .B0(new_n25383_), .Y(new_n25433_));
  AOI21X1  g25241(.A0(new_n25433_), .A1(new_n25432_), .B0(\asqrt[20] ), .Y(new_n25434_));
  OR2X1    g25242(.A(new_n25385_), .B(new_n25378_), .Y(new_n25435_));
  AOI21X1  g25243(.A0(new_n25435_), .A1(new_n25432_), .B0(new_n25384_), .Y(new_n25436_));
  NOR3X1   g25244(.A(new_n25403_), .B(new_n25436_), .C(new_n25434_), .Y(new_n25437_));
  OAI21X1  g25245(.A0(new_n25436_), .A1(new_n25434_), .B0(new_n25403_), .Y(new_n25438_));
  OAI21X1  g25246(.A0(new_n25437_), .A1(\asqrt[21] ), .B0(new_n25438_), .Y(new_n25439_));
  AND2X1   g25247(.A(new_n25439_), .B(new_n25411_), .Y(new_n25440_));
  OAI21X1  g25248(.A0(new_n25440_), .A1(new_n25414_), .B0(new_n25421_), .Y(new_n25441_));
  NAND3X1  g25249(.A(new_n25441_), .B(new_n25429_), .C(new_n25424_), .Y(new_n25442_));
  NAND2X1  g25250(.A(new_n25442_), .B(new_n10332_), .Y(new_n25443_));
  AOI21X1  g25251(.A0(new_n25441_), .A1(new_n25424_), .B0(new_n25429_), .Y(new_n25444_));
  OAI22X1  g25252(.A0(new_n24658_), .A1(new_n24651_), .B0(new_n24649_), .B1(new_n10332_), .Y(new_n25445_));
  OAI21X1  g25253(.A0(new_n25445_), .A1(new_n25203_), .B0(new_n24657_), .Y(new_n25446_));
  AND2X1   g25254(.A(new_n24691_), .B(new_n24690_), .Y(new_n25447_));
  OR4X1    g25255(.A(new_n25203_), .B(new_n25447_), .C(new_n24657_), .D(new_n24689_), .Y(new_n25448_));
  AND2X1   g25256(.A(new_n25448_), .B(new_n25446_), .Y(new_n25449_));
  NOR2X1   g25257(.A(new_n25449_), .B(new_n25444_), .Y(new_n25450_));
  AOI21X1  g25258(.A0(new_n25450_), .A1(new_n25443_), .B0(\asqrt[25] ), .Y(new_n25451_));
  INVX1    g25259(.A(new_n25449_), .Y(new_n25452_));
  AND2X1   g25260(.A(new_n24678_), .B(new_n24659_), .Y(new_n25453_));
  OR2X1    g25261(.A(new_n25453_), .B(new_n24660_), .Y(new_n25454_));
  OAI21X1  g25262(.A0(new_n25454_), .A1(new_n25203_), .B0(new_n24665_), .Y(new_n25455_));
  OR4X1    g25263(.A(new_n25203_), .B(new_n25453_), .C(new_n24665_), .D(new_n24660_), .Y(new_n25456_));
  AND2X1   g25264(.A(new_n25456_), .B(new_n25455_), .Y(new_n25457_));
  INVX1    g25265(.A(new_n25457_), .Y(new_n25458_));
  AOI21X1  g25266(.A0(new_n25442_), .A1(new_n10332_), .B0(new_n25444_), .Y(new_n25459_));
  OAI21X1  g25267(.A0(new_n25459_), .A1(new_n25452_), .B0(new_n25458_), .Y(new_n25460_));
  OAI21X1  g25268(.A0(new_n25460_), .A1(new_n25451_), .B0(new_n9353_), .Y(new_n25461_));
  AND2X1   g25269(.A(new_n25405_), .B(new_n11896_), .Y(new_n25462_));
  OR2X1    g25270(.A(new_n25412_), .B(new_n25411_), .Y(new_n25463_));
  OAI21X1  g25271(.A0(new_n25463_), .A1(new_n25462_), .B0(new_n11362_), .Y(new_n25464_));
  AOI21X1  g25272(.A0(new_n25439_), .A1(new_n25411_), .B0(new_n25421_), .Y(new_n25465_));
  AOI21X1  g25273(.A0(new_n25465_), .A1(new_n25464_), .B0(\asqrt[23] ), .Y(new_n25466_));
  OR2X1    g25274(.A(new_n25416_), .B(new_n25415_), .Y(new_n25467_));
  AOI21X1  g25275(.A0(new_n25467_), .A1(new_n25464_), .B0(new_n25422_), .Y(new_n25468_));
  NOR3X1   g25276(.A(new_n25468_), .B(new_n25428_), .C(new_n25466_), .Y(new_n25469_));
  OAI21X1  g25277(.A0(new_n25468_), .A1(new_n25466_), .B0(new_n25428_), .Y(new_n25470_));
  OAI21X1  g25278(.A0(new_n25469_), .A1(\asqrt[24] ), .B0(new_n25470_), .Y(new_n25471_));
  AND2X1   g25279(.A(new_n25471_), .B(new_n25449_), .Y(new_n25472_));
  OAI21X1  g25280(.A0(new_n25472_), .A1(new_n25451_), .B0(new_n25457_), .Y(new_n25473_));
  NAND2X1  g25281(.A(new_n24696_), .B(new_n24680_), .Y(new_n25474_));
  OAI21X1  g25282(.A0(new_n25474_), .A1(new_n25203_), .B0(new_n24688_), .Y(new_n25475_));
  NAND4X1  g25283(.A(\asqrt[1] ), .B(new_n24696_), .C(new_n24684_), .D(new_n24680_), .Y(new_n25476_));
  AND2X1   g25284(.A(new_n25476_), .B(new_n25475_), .Y(new_n25477_));
  INVX1    g25285(.A(new_n25477_), .Y(new_n25478_));
  NAND3X1  g25286(.A(new_n25478_), .B(new_n25473_), .C(new_n25461_), .Y(new_n25479_));
  NAND2X1  g25287(.A(new_n25479_), .B(new_n8874_), .Y(new_n25480_));
  OAI22X1  g25288(.A0(new_n24741_), .A1(new_n24739_), .B0(new_n24713_), .B1(new_n8874_), .Y(new_n25481_));
  OAI21X1  g25289(.A0(new_n25481_), .A1(new_n25203_), .B0(new_n24740_), .Y(new_n25482_));
  AND2X1   g25290(.A(new_n24704_), .B(new_n24697_), .Y(new_n25483_));
  OR4X1    g25291(.A(new_n25203_), .B(new_n25483_), .C(new_n24740_), .D(new_n24687_), .Y(new_n25484_));
  AND2X1   g25292(.A(new_n25484_), .B(new_n25482_), .Y(new_n25485_));
  AOI21X1  g25293(.A0(new_n25473_), .A1(new_n25461_), .B0(new_n25478_), .Y(new_n25486_));
  NOR2X1   g25294(.A(new_n25486_), .B(new_n25485_), .Y(new_n25487_));
  AOI21X1  g25295(.A0(new_n25487_), .A1(new_n25480_), .B0(\asqrt[28] ), .Y(new_n25488_));
  INVX1    g25296(.A(new_n25485_), .Y(new_n25489_));
  AOI21X1  g25297(.A0(new_n25479_), .A1(new_n8874_), .B0(new_n25486_), .Y(new_n25490_));
  AND2X1   g25298(.A(new_n24744_), .B(new_n24742_), .Y(new_n25491_));
  OR2X1    g25299(.A(new_n25491_), .B(new_n24743_), .Y(new_n25492_));
  OAI21X1  g25300(.A0(new_n25492_), .A1(new_n25203_), .B0(new_n24712_), .Y(new_n25493_));
  OR4X1    g25301(.A(new_n25203_), .B(new_n25491_), .C(new_n24712_), .D(new_n24743_), .Y(new_n25494_));
  AND2X1   g25302(.A(new_n25494_), .B(new_n25493_), .Y(new_n25495_));
  INVX1    g25303(.A(new_n25495_), .Y(new_n25496_));
  OAI21X1  g25304(.A0(new_n25490_), .A1(new_n25489_), .B0(new_n25496_), .Y(new_n25497_));
  OAI21X1  g25305(.A0(new_n25497_), .A1(new_n25488_), .B0(new_n7970_), .Y(new_n25498_));
  NAND2X1  g25306(.A(new_n24720_), .B(new_n24746_), .Y(new_n25499_));
  OAI21X1  g25307(.A0(new_n25499_), .A1(new_n25203_), .B0(new_n24719_), .Y(new_n25500_));
  NAND4X1  g25308(.A(\asqrt[1] ), .B(new_n24720_), .C(new_n24747_), .D(new_n24746_), .Y(new_n25501_));
  AND2X1   g25309(.A(new_n25501_), .B(new_n25500_), .Y(new_n25502_));
  INVX1    g25310(.A(new_n25502_), .Y(new_n25503_));
  AND2X1   g25311(.A(new_n25442_), .B(new_n10332_), .Y(new_n25504_));
  OR2X1    g25312(.A(new_n25449_), .B(new_n25444_), .Y(new_n25505_));
  OAI21X1  g25313(.A0(new_n25505_), .A1(new_n25504_), .B0(new_n9833_), .Y(new_n25506_));
  AOI21X1  g25314(.A0(new_n25471_), .A1(new_n25449_), .B0(new_n25457_), .Y(new_n25507_));
  AOI21X1  g25315(.A0(new_n25507_), .A1(new_n25506_), .B0(\asqrt[26] ), .Y(new_n25508_));
  OR2X1    g25316(.A(new_n25459_), .B(new_n25452_), .Y(new_n25509_));
  AOI21X1  g25317(.A0(new_n25509_), .A1(new_n25506_), .B0(new_n25458_), .Y(new_n25510_));
  NOR3X1   g25318(.A(new_n25477_), .B(new_n25510_), .C(new_n25508_), .Y(new_n25511_));
  OAI21X1  g25319(.A0(new_n25510_), .A1(new_n25508_), .B0(new_n25477_), .Y(new_n25512_));
  OAI21X1  g25320(.A0(new_n25511_), .A1(\asqrt[27] ), .B0(new_n25512_), .Y(new_n25513_));
  AND2X1   g25321(.A(new_n25513_), .B(new_n25485_), .Y(new_n25514_));
  OAI21X1  g25322(.A0(new_n25514_), .A1(new_n25488_), .B0(new_n25495_), .Y(new_n25515_));
  NAND3X1  g25323(.A(new_n25515_), .B(new_n25503_), .C(new_n25498_), .Y(new_n25516_));
  NAND2X1  g25324(.A(new_n25516_), .B(new_n7527_), .Y(new_n25517_));
  AOI21X1  g25325(.A0(new_n25515_), .A1(new_n25498_), .B0(new_n25503_), .Y(new_n25518_));
  OAI22X1  g25326(.A0(new_n24730_), .A1(new_n24723_), .B0(new_n24721_), .B1(new_n7527_), .Y(new_n25519_));
  OAI21X1  g25327(.A0(new_n25519_), .A1(new_n25203_), .B0(new_n24729_), .Y(new_n25520_));
  AND2X1   g25328(.A(new_n24763_), .B(new_n24762_), .Y(new_n25521_));
  OR4X1    g25329(.A(new_n25203_), .B(new_n25521_), .C(new_n24729_), .D(new_n24761_), .Y(new_n25522_));
  AND2X1   g25330(.A(new_n25522_), .B(new_n25520_), .Y(new_n25523_));
  NOR2X1   g25331(.A(new_n25523_), .B(new_n25518_), .Y(new_n25524_));
  AOI21X1  g25332(.A0(new_n25524_), .A1(new_n25517_), .B0(\asqrt[31] ), .Y(new_n25525_));
  INVX1    g25333(.A(new_n25523_), .Y(new_n25526_));
  AND2X1   g25334(.A(new_n24750_), .B(new_n24731_), .Y(new_n25527_));
  OR2X1    g25335(.A(new_n25527_), .B(new_n24732_), .Y(new_n25528_));
  OAI21X1  g25336(.A0(new_n25528_), .A1(new_n25203_), .B0(new_n24766_), .Y(new_n25529_));
  OR4X1    g25337(.A(new_n25203_), .B(new_n25527_), .C(new_n24766_), .D(new_n24732_), .Y(new_n25530_));
  AND2X1   g25338(.A(new_n25530_), .B(new_n25529_), .Y(new_n25531_));
  INVX1    g25339(.A(new_n25531_), .Y(new_n25532_));
  AOI21X1  g25340(.A0(new_n25516_), .A1(new_n7527_), .B0(new_n25518_), .Y(new_n25533_));
  OAI21X1  g25341(.A0(new_n25533_), .A1(new_n25526_), .B0(new_n25532_), .Y(new_n25534_));
  OAI21X1  g25342(.A0(new_n25534_), .A1(new_n25525_), .B0(new_n6699_), .Y(new_n25535_));
  AND2X1   g25343(.A(new_n25479_), .B(new_n8874_), .Y(new_n25536_));
  OR2X1    g25344(.A(new_n25486_), .B(new_n25485_), .Y(new_n25537_));
  OAI21X1  g25345(.A0(new_n25537_), .A1(new_n25536_), .B0(new_n8412_), .Y(new_n25538_));
  AOI21X1  g25346(.A0(new_n25513_), .A1(new_n25485_), .B0(new_n25495_), .Y(new_n25539_));
  AOI21X1  g25347(.A0(new_n25539_), .A1(new_n25538_), .B0(\asqrt[29] ), .Y(new_n25540_));
  OR2X1    g25348(.A(new_n25490_), .B(new_n25489_), .Y(new_n25541_));
  AOI21X1  g25349(.A0(new_n25541_), .A1(new_n25538_), .B0(new_n25496_), .Y(new_n25542_));
  NOR3X1   g25350(.A(new_n25542_), .B(new_n25502_), .C(new_n25540_), .Y(new_n25543_));
  OAI21X1  g25351(.A0(new_n25542_), .A1(new_n25540_), .B0(new_n25502_), .Y(new_n25544_));
  OAI21X1  g25352(.A0(new_n25543_), .A1(\asqrt[30] ), .B0(new_n25544_), .Y(new_n25545_));
  AND2X1   g25353(.A(new_n25545_), .B(new_n25523_), .Y(new_n25546_));
  OAI21X1  g25354(.A0(new_n25546_), .A1(new_n25525_), .B0(new_n25531_), .Y(new_n25547_));
  NAND2X1  g25355(.A(new_n24769_), .B(new_n24752_), .Y(new_n25548_));
  OAI21X1  g25356(.A0(new_n25548_), .A1(new_n25203_), .B0(new_n24760_), .Y(new_n25549_));
  OR4X1    g25357(.A(new_n25203_), .B(new_n24757_), .C(new_n24760_), .D(new_n24776_), .Y(new_n25550_));
  AND2X1   g25358(.A(new_n25550_), .B(new_n25549_), .Y(new_n25551_));
  INVX1    g25359(.A(new_n25551_), .Y(new_n25552_));
  NAND3X1  g25360(.A(new_n25552_), .B(new_n25547_), .C(new_n25535_), .Y(new_n25553_));
  NAND2X1  g25361(.A(new_n25553_), .B(new_n6294_), .Y(new_n25554_));
  OAI22X1  g25362(.A0(new_n24816_), .A1(new_n24814_), .B0(new_n24786_), .B1(new_n6294_), .Y(new_n25555_));
  OAI21X1  g25363(.A0(new_n25555_), .A1(new_n25203_), .B0(new_n24815_), .Y(new_n25556_));
  AND2X1   g25364(.A(new_n24777_), .B(new_n24770_), .Y(new_n25557_));
  OR4X1    g25365(.A(new_n25203_), .B(new_n25557_), .C(new_n24815_), .D(new_n24759_), .Y(new_n25558_));
  AND2X1   g25366(.A(new_n25558_), .B(new_n25556_), .Y(new_n25559_));
  AOI21X1  g25367(.A0(new_n25547_), .A1(new_n25535_), .B0(new_n25552_), .Y(new_n25560_));
  NOR2X1   g25368(.A(new_n25560_), .B(new_n25559_), .Y(new_n25561_));
  AOI21X1  g25369(.A0(new_n25561_), .A1(new_n25554_), .B0(\asqrt[34] ), .Y(new_n25562_));
  INVX1    g25370(.A(new_n25559_), .Y(new_n25563_));
  AOI21X1  g25371(.A0(new_n25553_), .A1(new_n6294_), .B0(new_n25560_), .Y(new_n25564_));
  AND2X1   g25372(.A(new_n24819_), .B(new_n24817_), .Y(new_n25565_));
  OR2X1    g25373(.A(new_n25565_), .B(new_n24818_), .Y(new_n25566_));
  OAI21X1  g25374(.A0(new_n25566_), .A1(new_n25203_), .B0(new_n24785_), .Y(new_n25567_));
  OR4X1    g25375(.A(new_n25203_), .B(new_n25565_), .C(new_n24785_), .D(new_n24818_), .Y(new_n25568_));
  AND2X1   g25376(.A(new_n25568_), .B(new_n25567_), .Y(new_n25569_));
  INVX1    g25377(.A(new_n25569_), .Y(new_n25570_));
  OAI21X1  g25378(.A0(new_n25564_), .A1(new_n25563_), .B0(new_n25570_), .Y(new_n25571_));
  OAI21X1  g25379(.A0(new_n25571_), .A1(new_n25562_), .B0(new_n5541_), .Y(new_n25572_));
  NAND2X1  g25380(.A(new_n24795_), .B(new_n24821_), .Y(new_n25573_));
  OAI21X1  g25381(.A0(new_n25573_), .A1(new_n25203_), .B0(new_n24794_), .Y(new_n25574_));
  NAND4X1  g25382(.A(\asqrt[1] ), .B(new_n24795_), .C(new_n24793_), .D(new_n24821_), .Y(new_n25575_));
  AND2X1   g25383(.A(new_n25575_), .B(new_n25574_), .Y(new_n25576_));
  INVX1    g25384(.A(new_n25576_), .Y(new_n25577_));
  AND2X1   g25385(.A(new_n25516_), .B(new_n7527_), .Y(new_n25578_));
  OR2X1    g25386(.A(new_n25523_), .B(new_n25518_), .Y(new_n25579_));
  OAI21X1  g25387(.A0(new_n25579_), .A1(new_n25578_), .B0(new_n7103_), .Y(new_n25580_));
  AOI21X1  g25388(.A0(new_n25545_), .A1(new_n25523_), .B0(new_n25531_), .Y(new_n25581_));
  AOI21X1  g25389(.A0(new_n25581_), .A1(new_n25580_), .B0(\asqrt[32] ), .Y(new_n25582_));
  OR2X1    g25390(.A(new_n25533_), .B(new_n25526_), .Y(new_n25583_));
  AOI21X1  g25391(.A0(new_n25583_), .A1(new_n25580_), .B0(new_n25532_), .Y(new_n25584_));
  NOR3X1   g25392(.A(new_n25551_), .B(new_n25584_), .C(new_n25582_), .Y(new_n25585_));
  OAI21X1  g25393(.A0(new_n25584_), .A1(new_n25582_), .B0(new_n25551_), .Y(new_n25586_));
  OAI21X1  g25394(.A0(new_n25585_), .A1(\asqrt[33] ), .B0(new_n25586_), .Y(new_n25587_));
  AND2X1   g25395(.A(new_n25587_), .B(new_n25559_), .Y(new_n25588_));
  OAI21X1  g25396(.A0(new_n25588_), .A1(new_n25562_), .B0(new_n25569_), .Y(new_n25589_));
  NAND3X1  g25397(.A(new_n25589_), .B(new_n25577_), .C(new_n25572_), .Y(new_n25590_));
  NAND2X1  g25398(.A(new_n25590_), .B(new_n5176_), .Y(new_n25591_));
  AOI21X1  g25399(.A0(new_n25589_), .A1(new_n25572_), .B0(new_n25577_), .Y(new_n25592_));
  OAI22X1  g25400(.A0(new_n24805_), .A1(new_n24798_), .B0(new_n24796_), .B1(new_n5176_), .Y(new_n25593_));
  OAI21X1  g25401(.A0(new_n25593_), .A1(new_n25203_), .B0(new_n24804_), .Y(new_n25594_));
  AND2X1   g25402(.A(new_n24836_), .B(new_n24835_), .Y(new_n25595_));
  OR4X1    g25403(.A(new_n25203_), .B(new_n25595_), .C(new_n24804_), .D(new_n24834_), .Y(new_n25596_));
  AND2X1   g25404(.A(new_n25596_), .B(new_n25594_), .Y(new_n25597_));
  NOR2X1   g25405(.A(new_n25597_), .B(new_n25592_), .Y(new_n25598_));
  AOI21X1  g25406(.A0(new_n25598_), .A1(new_n25591_), .B0(\asqrt[37] ), .Y(new_n25599_));
  INVX1    g25407(.A(new_n25597_), .Y(new_n25600_));
  AND2X1   g25408(.A(new_n24824_), .B(new_n24806_), .Y(new_n25601_));
  OR2X1    g25409(.A(new_n25601_), .B(new_n24807_), .Y(new_n25602_));
  OAI21X1  g25410(.A0(new_n25602_), .A1(new_n25203_), .B0(new_n24839_), .Y(new_n25603_));
  OR4X1    g25411(.A(new_n25203_), .B(new_n25601_), .C(new_n24839_), .D(new_n24807_), .Y(new_n25604_));
  AND2X1   g25412(.A(new_n25604_), .B(new_n25603_), .Y(new_n25605_));
  INVX1    g25413(.A(new_n25605_), .Y(new_n25606_));
  AOI21X1  g25414(.A0(new_n25590_), .A1(new_n5176_), .B0(new_n25592_), .Y(new_n25607_));
  OAI21X1  g25415(.A0(new_n25607_), .A1(new_n25600_), .B0(new_n25606_), .Y(new_n25608_));
  OAI21X1  g25416(.A0(new_n25608_), .A1(new_n25599_), .B0(new_n4493_), .Y(new_n25609_));
  AND2X1   g25417(.A(new_n25553_), .B(new_n6294_), .Y(new_n25610_));
  OR2X1    g25418(.A(new_n25560_), .B(new_n25559_), .Y(new_n25611_));
  OAI21X1  g25419(.A0(new_n25611_), .A1(new_n25610_), .B0(new_n5941_), .Y(new_n25612_));
  AOI21X1  g25420(.A0(new_n25587_), .A1(new_n25559_), .B0(new_n25569_), .Y(new_n25613_));
  AOI21X1  g25421(.A0(new_n25613_), .A1(new_n25612_), .B0(\asqrt[35] ), .Y(new_n25614_));
  OR2X1    g25422(.A(new_n25564_), .B(new_n25563_), .Y(new_n25615_));
  AOI21X1  g25423(.A0(new_n25615_), .A1(new_n25612_), .B0(new_n25570_), .Y(new_n25616_));
  NOR3X1   g25424(.A(new_n25616_), .B(new_n25576_), .C(new_n25614_), .Y(new_n25617_));
  OAI21X1  g25425(.A0(new_n25616_), .A1(new_n25614_), .B0(new_n25576_), .Y(new_n25618_));
  OAI21X1  g25426(.A0(new_n25617_), .A1(\asqrt[36] ), .B0(new_n25618_), .Y(new_n25619_));
  AND2X1   g25427(.A(new_n25619_), .B(new_n25597_), .Y(new_n25620_));
  OAI21X1  g25428(.A0(new_n25620_), .A1(new_n25599_), .B0(new_n25605_), .Y(new_n25621_));
  NAND2X1  g25429(.A(new_n24842_), .B(new_n24826_), .Y(new_n25622_));
  OAI21X1  g25430(.A0(new_n25622_), .A1(new_n25203_), .B0(new_n24829_), .Y(new_n25623_));
  NAND4X1  g25431(.A(\asqrt[1] ), .B(new_n24842_), .C(new_n24830_), .D(new_n24826_), .Y(new_n25624_));
  AND2X1   g25432(.A(new_n25624_), .B(new_n25623_), .Y(new_n25625_));
  INVX1    g25433(.A(new_n25625_), .Y(new_n25626_));
  NAND3X1  g25434(.A(new_n25626_), .B(new_n25621_), .C(new_n25609_), .Y(new_n25627_));
  NAND2X1  g25435(.A(new_n25627_), .B(new_n4165_), .Y(new_n25628_));
  OAI22X1  g25436(.A0(new_n24889_), .A1(new_n24887_), .B0(new_n24859_), .B1(new_n4165_), .Y(new_n25629_));
  OAI21X1  g25437(.A0(new_n25629_), .A1(new_n25203_), .B0(new_n24888_), .Y(new_n25630_));
  AND2X1   g25438(.A(new_n24850_), .B(new_n24843_), .Y(new_n25631_));
  OR4X1    g25439(.A(new_n25203_), .B(new_n25631_), .C(new_n24888_), .D(new_n24833_), .Y(new_n25632_));
  AND2X1   g25440(.A(new_n25632_), .B(new_n25630_), .Y(new_n25633_));
  AOI21X1  g25441(.A0(new_n25621_), .A1(new_n25609_), .B0(new_n25626_), .Y(new_n25634_));
  NOR2X1   g25442(.A(new_n25634_), .B(new_n25633_), .Y(new_n25635_));
  AOI21X1  g25443(.A0(new_n25635_), .A1(new_n25628_), .B0(\asqrt[40] ), .Y(new_n25636_));
  INVX1    g25444(.A(new_n25633_), .Y(new_n25637_));
  AOI21X1  g25445(.A0(new_n25627_), .A1(new_n4165_), .B0(new_n25634_), .Y(new_n25638_));
  AND2X1   g25446(.A(new_n24892_), .B(new_n24890_), .Y(new_n25639_));
  OR2X1    g25447(.A(new_n25639_), .B(new_n24891_), .Y(new_n25640_));
  OAI21X1  g25448(.A0(new_n25640_), .A1(new_n25203_), .B0(new_n24858_), .Y(new_n25641_));
  OR4X1    g25449(.A(new_n25203_), .B(new_n25639_), .C(new_n24858_), .D(new_n24891_), .Y(new_n25642_));
  AND2X1   g25450(.A(new_n25642_), .B(new_n25641_), .Y(new_n25643_));
  INVX1    g25451(.A(new_n25643_), .Y(new_n25644_));
  OAI21X1  g25452(.A0(new_n25638_), .A1(new_n25637_), .B0(new_n25644_), .Y(new_n25645_));
  OAI21X1  g25453(.A0(new_n25645_), .A1(new_n25636_), .B0(new_n3564_), .Y(new_n25646_));
  NAND2X1  g25454(.A(new_n24868_), .B(new_n24894_), .Y(new_n25647_));
  OAI21X1  g25455(.A0(new_n25647_), .A1(new_n25203_), .B0(new_n24867_), .Y(new_n25648_));
  NAND4X1  g25456(.A(\asqrt[1] ), .B(new_n24868_), .C(new_n24866_), .D(new_n24894_), .Y(new_n25649_));
  AND2X1   g25457(.A(new_n25649_), .B(new_n25648_), .Y(new_n25650_));
  INVX1    g25458(.A(new_n25650_), .Y(new_n25651_));
  AND2X1   g25459(.A(new_n25590_), .B(new_n5176_), .Y(new_n25652_));
  OR2X1    g25460(.A(new_n25597_), .B(new_n25592_), .Y(new_n25653_));
  OAI21X1  g25461(.A0(new_n25653_), .A1(new_n25652_), .B0(new_n4826_), .Y(new_n25654_));
  AOI21X1  g25462(.A0(new_n25619_), .A1(new_n25597_), .B0(new_n25605_), .Y(new_n25655_));
  AOI21X1  g25463(.A0(new_n25655_), .A1(new_n25654_), .B0(\asqrt[38] ), .Y(new_n25656_));
  OR2X1    g25464(.A(new_n25607_), .B(new_n25600_), .Y(new_n25657_));
  AOI21X1  g25465(.A0(new_n25657_), .A1(new_n25654_), .B0(new_n25606_), .Y(new_n25658_));
  NOR3X1   g25466(.A(new_n25625_), .B(new_n25658_), .C(new_n25656_), .Y(new_n25659_));
  OAI21X1  g25467(.A0(new_n25658_), .A1(new_n25656_), .B0(new_n25625_), .Y(new_n25660_));
  OAI21X1  g25468(.A0(new_n25659_), .A1(\asqrt[39] ), .B0(new_n25660_), .Y(new_n25661_));
  AND2X1   g25469(.A(new_n25661_), .B(new_n25633_), .Y(new_n25662_));
  OAI21X1  g25470(.A0(new_n25662_), .A1(new_n25636_), .B0(new_n25643_), .Y(new_n25663_));
  NAND3X1  g25471(.A(new_n25663_), .B(new_n25651_), .C(new_n25646_), .Y(new_n25664_));
  AND2X1   g25472(.A(new_n25664_), .B(new_n3276_), .Y(new_n25665_));
  AOI21X1  g25473(.A0(new_n25663_), .A1(new_n25646_), .B0(new_n25651_), .Y(new_n25666_));
  OAI22X1  g25474(.A0(new_n24878_), .A1(new_n24871_), .B0(new_n24869_), .B1(new_n3276_), .Y(new_n25667_));
  OAI21X1  g25475(.A0(new_n25667_), .A1(new_n25203_), .B0(new_n24877_), .Y(new_n25668_));
  AND2X1   g25476(.A(new_n24910_), .B(new_n24909_), .Y(new_n25669_));
  OR4X1    g25477(.A(new_n25203_), .B(new_n25669_), .C(new_n24877_), .D(new_n24908_), .Y(new_n25670_));
  AND2X1   g25478(.A(new_n25670_), .B(new_n25668_), .Y(new_n25671_));
  OR2X1    g25479(.A(new_n25671_), .B(new_n25666_), .Y(new_n25672_));
  OAI21X1  g25480(.A0(new_n25672_), .A1(new_n25665_), .B0(new_n3008_), .Y(new_n25673_));
  AND2X1   g25481(.A(new_n24897_), .B(new_n24879_), .Y(new_n25674_));
  OR2X1    g25482(.A(new_n25674_), .B(new_n24880_), .Y(new_n25675_));
  OAI21X1  g25483(.A0(new_n25675_), .A1(new_n25203_), .B0(new_n24913_), .Y(new_n25676_));
  OR4X1    g25484(.A(new_n25203_), .B(new_n25674_), .C(new_n24913_), .D(new_n24880_), .Y(new_n25677_));
  AND2X1   g25485(.A(new_n25677_), .B(new_n25676_), .Y(new_n25678_));
  AND2X1   g25486(.A(new_n25627_), .B(new_n4165_), .Y(new_n25679_));
  OR2X1    g25487(.A(new_n25634_), .B(new_n25633_), .Y(new_n25680_));
  OAI21X1  g25488(.A0(new_n25680_), .A1(new_n25679_), .B0(new_n3863_), .Y(new_n25681_));
  AOI21X1  g25489(.A0(new_n25661_), .A1(new_n25633_), .B0(new_n25643_), .Y(new_n25682_));
  AOI21X1  g25490(.A0(new_n25682_), .A1(new_n25681_), .B0(\asqrt[41] ), .Y(new_n25683_));
  OR2X1    g25491(.A(new_n25638_), .B(new_n25637_), .Y(new_n25684_));
  AOI21X1  g25492(.A0(new_n25684_), .A1(new_n25681_), .B0(new_n25644_), .Y(new_n25685_));
  NOR3X1   g25493(.A(new_n25685_), .B(new_n25650_), .C(new_n25683_), .Y(new_n25686_));
  OAI21X1  g25494(.A0(new_n25685_), .A1(new_n25683_), .B0(new_n25650_), .Y(new_n25687_));
  OAI21X1  g25495(.A0(new_n25686_), .A1(\asqrt[42] ), .B0(new_n25687_), .Y(new_n25688_));
  AOI21X1  g25496(.A0(new_n25688_), .A1(new_n25671_), .B0(new_n25678_), .Y(new_n25689_));
  AOI21X1  g25497(.A0(new_n25689_), .A1(new_n25673_), .B0(\asqrt[44] ), .Y(new_n25690_));
  INVX1    g25498(.A(new_n25678_), .Y(new_n25691_));
  INVX1    g25499(.A(new_n25671_), .Y(new_n25692_));
  AOI21X1  g25500(.A0(new_n25664_), .A1(new_n3276_), .B0(new_n25666_), .Y(new_n25693_));
  OR2X1    g25501(.A(new_n25693_), .B(new_n25692_), .Y(new_n25694_));
  AOI21X1  g25502(.A0(new_n25694_), .A1(new_n25673_), .B0(new_n25691_), .Y(new_n25695_));
  NAND2X1  g25503(.A(new_n24916_), .B(new_n24899_), .Y(new_n25696_));
  OAI21X1  g25504(.A0(new_n25696_), .A1(new_n25203_), .B0(new_n24907_), .Y(new_n25697_));
  NAND4X1  g25505(.A(\asqrt[1] ), .B(new_n24916_), .C(new_n24903_), .D(new_n24899_), .Y(new_n25698_));
  AND2X1   g25506(.A(new_n25698_), .B(new_n25697_), .Y(new_n25699_));
  NOR3X1   g25507(.A(new_n25699_), .B(new_n25695_), .C(new_n25690_), .Y(new_n25700_));
  OR2X1    g25508(.A(new_n25700_), .B(\asqrt[45] ), .Y(new_n25701_));
  OAI22X1  g25509(.A0(new_n24963_), .A1(new_n24961_), .B0(new_n24933_), .B1(new_n2570_), .Y(new_n25702_));
  OAI21X1  g25510(.A0(new_n25702_), .A1(new_n25203_), .B0(new_n24962_), .Y(new_n25703_));
  AND2X1   g25511(.A(new_n24924_), .B(new_n24917_), .Y(new_n25704_));
  OR4X1    g25512(.A(new_n25203_), .B(new_n25704_), .C(new_n24962_), .D(new_n24906_), .Y(new_n25705_));
  AND2X1   g25513(.A(new_n25705_), .B(new_n25703_), .Y(new_n25706_));
  INVX1    g25514(.A(new_n25706_), .Y(new_n25707_));
  OAI21X1  g25515(.A0(new_n25695_), .A1(new_n25690_), .B0(new_n25699_), .Y(new_n25708_));
  AND2X1   g25516(.A(new_n25708_), .B(new_n25707_), .Y(new_n25709_));
  AOI21X1  g25517(.A0(new_n25709_), .A1(new_n25701_), .B0(\asqrt[46] ), .Y(new_n25710_));
  OR2X1    g25518(.A(new_n25686_), .B(\asqrt[42] ), .Y(new_n25711_));
  AND2X1   g25519(.A(new_n25692_), .B(new_n25687_), .Y(new_n25712_));
  AOI21X1  g25520(.A0(new_n25712_), .A1(new_n25711_), .B0(\asqrt[43] ), .Y(new_n25713_));
  OAI21X1  g25521(.A0(new_n25693_), .A1(new_n25692_), .B0(new_n25691_), .Y(new_n25714_));
  OAI21X1  g25522(.A0(new_n25714_), .A1(new_n25713_), .B0(new_n2769_), .Y(new_n25715_));
  AND2X1   g25523(.A(new_n25688_), .B(new_n25671_), .Y(new_n25716_));
  OAI21X1  g25524(.A0(new_n25716_), .A1(new_n25713_), .B0(new_n25678_), .Y(new_n25717_));
  INVX1    g25525(.A(new_n25699_), .Y(new_n25718_));
  NAND3X1  g25526(.A(new_n25718_), .B(new_n25717_), .C(new_n25715_), .Y(new_n25719_));
  AOI21X1  g25527(.A0(new_n25717_), .A1(new_n25715_), .B0(new_n25718_), .Y(new_n25720_));
  AOI21X1  g25528(.A0(new_n25719_), .A1(new_n2570_), .B0(new_n25720_), .Y(new_n25721_));
  AND2X1   g25529(.A(new_n24966_), .B(new_n24964_), .Y(new_n25722_));
  OR2X1    g25530(.A(new_n25722_), .B(new_n24965_), .Y(new_n25723_));
  OAI21X1  g25531(.A0(new_n25723_), .A1(new_n25203_), .B0(new_n24932_), .Y(new_n25724_));
  OR4X1    g25532(.A(new_n25203_), .B(new_n25722_), .C(new_n24932_), .D(new_n24965_), .Y(new_n25725_));
  AND2X1   g25533(.A(new_n25725_), .B(new_n25724_), .Y(new_n25726_));
  INVX1    g25534(.A(new_n25726_), .Y(new_n25727_));
  OAI21X1  g25535(.A0(new_n25721_), .A1(new_n25707_), .B0(new_n25727_), .Y(new_n25728_));
  OAI21X1  g25536(.A0(new_n25728_), .A1(new_n25710_), .B0(new_n2040_), .Y(new_n25729_));
  NAND2X1  g25537(.A(new_n24942_), .B(new_n24968_), .Y(new_n25730_));
  OAI21X1  g25538(.A0(new_n25730_), .A1(new_n25203_), .B0(new_n24941_), .Y(new_n25731_));
  NAND4X1  g25539(.A(\asqrt[1] ), .B(new_n24942_), .C(new_n24940_), .D(new_n24968_), .Y(new_n25732_));
  AND2X1   g25540(.A(new_n25732_), .B(new_n25731_), .Y(new_n25733_));
  INVX1    g25541(.A(new_n25733_), .Y(new_n25734_));
  OAI21X1  g25542(.A0(new_n25700_), .A1(\asqrt[45] ), .B0(new_n25708_), .Y(new_n25735_));
  AND2X1   g25543(.A(new_n25735_), .B(new_n25706_), .Y(new_n25736_));
  OAI21X1  g25544(.A0(new_n25736_), .A1(new_n25710_), .B0(new_n25726_), .Y(new_n25737_));
  NAND3X1  g25545(.A(new_n25737_), .B(new_n25734_), .C(new_n25729_), .Y(new_n25738_));
  AND2X1   g25546(.A(new_n25738_), .B(new_n1834_), .Y(new_n25739_));
  AOI21X1  g25547(.A0(new_n25737_), .A1(new_n25729_), .B0(new_n25734_), .Y(new_n25740_));
  OAI22X1  g25548(.A0(new_n24952_), .A1(new_n24945_), .B0(new_n24943_), .B1(new_n1834_), .Y(new_n25741_));
  OAI21X1  g25549(.A0(new_n25741_), .A1(new_n25203_), .B0(new_n24951_), .Y(new_n25742_));
  AND2X1   g25550(.A(new_n24984_), .B(new_n24983_), .Y(new_n25743_));
  OR4X1    g25551(.A(new_n25203_), .B(new_n25743_), .C(new_n24951_), .D(new_n24982_), .Y(new_n25744_));
  AND2X1   g25552(.A(new_n25744_), .B(new_n25742_), .Y(new_n25745_));
  OR2X1    g25553(.A(new_n25745_), .B(new_n25740_), .Y(new_n25746_));
  OAI21X1  g25554(.A0(new_n25746_), .A1(new_n25739_), .B0(new_n1632_), .Y(new_n25747_));
  AND2X1   g25555(.A(new_n24971_), .B(new_n24953_), .Y(new_n25748_));
  OR2X1    g25556(.A(new_n25748_), .B(new_n24954_), .Y(new_n25749_));
  OAI21X1  g25557(.A0(new_n25749_), .A1(new_n25203_), .B0(new_n24987_), .Y(new_n25750_));
  OR4X1    g25558(.A(new_n25203_), .B(new_n25748_), .C(new_n24987_), .D(new_n24954_), .Y(new_n25751_));
  AND2X1   g25559(.A(new_n25751_), .B(new_n25750_), .Y(new_n25752_));
  NOR2X1   g25560(.A(new_n25700_), .B(\asqrt[45] ), .Y(new_n25753_));
  NAND2X1  g25561(.A(new_n25708_), .B(new_n25707_), .Y(new_n25754_));
  OAI21X1  g25562(.A0(new_n25754_), .A1(new_n25753_), .B0(new_n2263_), .Y(new_n25755_));
  AOI21X1  g25563(.A0(new_n25735_), .A1(new_n25706_), .B0(new_n25726_), .Y(new_n25756_));
  AOI21X1  g25564(.A0(new_n25756_), .A1(new_n25755_), .B0(\asqrt[47] ), .Y(new_n25757_));
  OR2X1    g25565(.A(new_n25721_), .B(new_n25707_), .Y(new_n25758_));
  AOI21X1  g25566(.A0(new_n25758_), .A1(new_n25755_), .B0(new_n25727_), .Y(new_n25759_));
  NOR3X1   g25567(.A(new_n25759_), .B(new_n25733_), .C(new_n25757_), .Y(new_n25760_));
  OAI21X1  g25568(.A0(new_n25759_), .A1(new_n25757_), .B0(new_n25733_), .Y(new_n25761_));
  OAI21X1  g25569(.A0(new_n25760_), .A1(\asqrt[48] ), .B0(new_n25761_), .Y(new_n25762_));
  AOI21X1  g25570(.A0(new_n25762_), .A1(new_n25745_), .B0(new_n25752_), .Y(new_n25763_));
  AOI21X1  g25571(.A0(new_n25763_), .A1(new_n25747_), .B0(\asqrt[50] ), .Y(new_n25764_));
  INVX1    g25572(.A(new_n25752_), .Y(new_n25765_));
  INVX1    g25573(.A(new_n25745_), .Y(new_n25766_));
  AOI21X1  g25574(.A0(new_n25738_), .A1(new_n1834_), .B0(new_n25740_), .Y(new_n25767_));
  OR2X1    g25575(.A(new_n25767_), .B(new_n25766_), .Y(new_n25768_));
  AOI21X1  g25576(.A0(new_n25768_), .A1(new_n25747_), .B0(new_n25765_), .Y(new_n25769_));
  NAND2X1  g25577(.A(new_n24990_), .B(new_n24973_), .Y(new_n25770_));
  OAI21X1  g25578(.A0(new_n25770_), .A1(new_n25203_), .B0(new_n24981_), .Y(new_n25771_));
  NAND4X1  g25579(.A(\asqrt[1] ), .B(new_n24990_), .C(new_n24977_), .D(new_n24973_), .Y(new_n25772_));
  AND2X1   g25580(.A(new_n25772_), .B(new_n25771_), .Y(new_n25773_));
  NOR3X1   g25581(.A(new_n25773_), .B(new_n25769_), .C(new_n25764_), .Y(new_n25774_));
  NOR2X1   g25582(.A(new_n25774_), .B(\asqrt[51] ), .Y(new_n25775_));
  OAI22X1  g25583(.A0(new_n25037_), .A1(new_n25035_), .B0(new_n25007_), .B1(new_n1277_), .Y(new_n25776_));
  OAI21X1  g25584(.A0(new_n25776_), .A1(new_n25203_), .B0(new_n25036_), .Y(new_n25777_));
  AND2X1   g25585(.A(new_n24998_), .B(new_n24991_), .Y(new_n25778_));
  OR4X1    g25586(.A(new_n25203_), .B(new_n25778_), .C(new_n25036_), .D(new_n24980_), .Y(new_n25779_));
  AND2X1   g25587(.A(new_n25779_), .B(new_n25777_), .Y(new_n25780_));
  OR2X1    g25588(.A(new_n25760_), .B(\asqrt[48] ), .Y(new_n25781_));
  AND2X1   g25589(.A(new_n25766_), .B(new_n25761_), .Y(new_n25782_));
  AOI21X1  g25590(.A0(new_n25782_), .A1(new_n25781_), .B0(\asqrt[49] ), .Y(new_n25783_));
  OAI21X1  g25591(.A0(new_n25767_), .A1(new_n25766_), .B0(new_n25765_), .Y(new_n25784_));
  OAI21X1  g25592(.A0(new_n25784_), .A1(new_n25783_), .B0(new_n1469_), .Y(new_n25785_));
  AND2X1   g25593(.A(new_n25762_), .B(new_n25745_), .Y(new_n25786_));
  OAI21X1  g25594(.A0(new_n25786_), .A1(new_n25783_), .B0(new_n25752_), .Y(new_n25787_));
  INVX1    g25595(.A(new_n25773_), .Y(new_n25788_));
  AOI21X1  g25596(.A0(new_n25787_), .A1(new_n25785_), .B0(new_n25788_), .Y(new_n25789_));
  OR2X1    g25597(.A(new_n25789_), .B(new_n25780_), .Y(new_n25790_));
  OAI21X1  g25598(.A0(new_n25790_), .A1(new_n25775_), .B0(new_n1111_), .Y(new_n25791_));
  OAI21X1  g25599(.A0(new_n25769_), .A1(new_n25764_), .B0(new_n25773_), .Y(new_n25792_));
  OAI21X1  g25600(.A0(new_n25774_), .A1(\asqrt[51] ), .B0(new_n25792_), .Y(new_n25793_));
  AND2X1   g25601(.A(new_n25040_), .B(new_n25038_), .Y(new_n25794_));
  OR2X1    g25602(.A(new_n25794_), .B(new_n25039_), .Y(new_n25795_));
  OAI21X1  g25603(.A0(new_n25795_), .A1(new_n25203_), .B0(new_n25006_), .Y(new_n25796_));
  OR4X1    g25604(.A(new_n25203_), .B(new_n25794_), .C(new_n25006_), .D(new_n25039_), .Y(new_n25797_));
  AND2X1   g25605(.A(new_n25797_), .B(new_n25796_), .Y(new_n25798_));
  AOI21X1  g25606(.A0(new_n25793_), .A1(new_n25780_), .B0(new_n25798_), .Y(new_n25799_));
  AOI21X1  g25607(.A0(new_n25799_), .A1(new_n25791_), .B0(\asqrt[53] ), .Y(new_n25800_));
  NAND2X1  g25608(.A(new_n25016_), .B(new_n25042_), .Y(new_n25801_));
  OAI21X1  g25609(.A0(new_n25801_), .A1(new_n25203_), .B0(new_n25015_), .Y(new_n25802_));
  NAND4X1  g25610(.A(\asqrt[1] ), .B(new_n25016_), .C(new_n25014_), .D(new_n25042_), .Y(new_n25803_));
  AND2X1   g25611(.A(new_n25803_), .B(new_n25802_), .Y(new_n25804_));
  INVX1    g25612(.A(new_n25780_), .Y(new_n25805_));
  NAND3X1  g25613(.A(new_n25788_), .B(new_n25787_), .C(new_n25785_), .Y(new_n25806_));
  AOI21X1  g25614(.A0(new_n25806_), .A1(new_n1277_), .B0(new_n25789_), .Y(new_n25807_));
  OR2X1    g25615(.A(new_n25807_), .B(new_n25805_), .Y(new_n25808_));
  INVX1    g25616(.A(new_n25798_), .Y(new_n25809_));
  AOI21X1  g25617(.A0(new_n25808_), .A1(new_n25791_), .B0(new_n25809_), .Y(new_n25810_));
  NOR3X1   g25618(.A(new_n25810_), .B(new_n25804_), .C(new_n25800_), .Y(new_n25811_));
  OR2X1    g25619(.A(new_n25811_), .B(\asqrt[54] ), .Y(new_n25812_));
  OAI21X1  g25620(.A0(new_n25810_), .A1(new_n25800_), .B0(new_n25804_), .Y(new_n25813_));
  OAI22X1  g25621(.A0(new_n25026_), .A1(new_n25019_), .B0(new_n25017_), .B1(new_n902_), .Y(new_n25814_));
  OAI21X1  g25622(.A0(new_n25814_), .A1(new_n25203_), .B0(new_n25025_), .Y(new_n25815_));
  AND2X1   g25623(.A(new_n25057_), .B(new_n25056_), .Y(new_n25816_));
  OR4X1    g25624(.A(new_n25203_), .B(new_n25816_), .C(new_n25025_), .D(new_n25055_), .Y(new_n25817_));
  AND2X1   g25625(.A(new_n25817_), .B(new_n25815_), .Y(new_n25818_));
  INVX1    g25626(.A(new_n25818_), .Y(new_n25819_));
  AND2X1   g25627(.A(new_n25819_), .B(new_n25813_), .Y(new_n25820_));
  AOI21X1  g25628(.A0(new_n25820_), .A1(new_n25812_), .B0(\asqrt[55] ), .Y(new_n25821_));
  AND2X1   g25629(.A(new_n25045_), .B(new_n25027_), .Y(new_n25822_));
  OR2X1    g25630(.A(new_n25822_), .B(new_n25028_), .Y(new_n25823_));
  OAI21X1  g25631(.A0(new_n25823_), .A1(new_n25203_), .B0(new_n25060_), .Y(new_n25824_));
  OR4X1    g25632(.A(new_n25203_), .B(new_n25822_), .C(new_n25060_), .D(new_n25028_), .Y(new_n25825_));
  AND2X1   g25633(.A(new_n25825_), .B(new_n25824_), .Y(new_n25826_));
  INVX1    g25634(.A(new_n25826_), .Y(new_n25827_));
  OR2X1    g25635(.A(new_n25774_), .B(\asqrt[51] ), .Y(new_n25828_));
  AND2X1   g25636(.A(new_n25792_), .B(new_n25805_), .Y(new_n25829_));
  AOI21X1  g25637(.A0(new_n25829_), .A1(new_n25828_), .B0(\asqrt[52] ), .Y(new_n25830_));
  OAI21X1  g25638(.A0(new_n25807_), .A1(new_n25805_), .B0(new_n25809_), .Y(new_n25831_));
  OAI21X1  g25639(.A0(new_n25831_), .A1(new_n25830_), .B0(new_n968_), .Y(new_n25832_));
  INVX1    g25640(.A(new_n25804_), .Y(new_n25833_));
  AND2X1   g25641(.A(new_n25793_), .B(new_n25780_), .Y(new_n25834_));
  OAI21X1  g25642(.A0(new_n25834_), .A1(new_n25830_), .B0(new_n25798_), .Y(new_n25835_));
  NAND3X1  g25643(.A(new_n25835_), .B(new_n25833_), .C(new_n25832_), .Y(new_n25836_));
  AOI21X1  g25644(.A0(new_n25835_), .A1(new_n25832_), .B0(new_n25833_), .Y(new_n25837_));
  AOI21X1  g25645(.A0(new_n25836_), .A1(new_n902_), .B0(new_n25837_), .Y(new_n25838_));
  OAI21X1  g25646(.A0(new_n25838_), .A1(new_n25819_), .B0(new_n25827_), .Y(new_n25839_));
  OAI21X1  g25647(.A0(new_n25839_), .A1(new_n25821_), .B0(new_n582_), .Y(new_n25840_));
  OAI21X1  g25648(.A0(new_n25811_), .A1(\asqrt[54] ), .B0(new_n25813_), .Y(new_n25841_));
  AND2X1   g25649(.A(new_n25841_), .B(new_n25818_), .Y(new_n25842_));
  OAI21X1  g25650(.A0(new_n25842_), .A1(new_n25821_), .B0(new_n25826_), .Y(new_n25843_));
  NAND2X1  g25651(.A(new_n25063_), .B(new_n25047_), .Y(new_n25844_));
  OAI21X1  g25652(.A0(new_n25844_), .A1(new_n25203_), .B0(new_n25050_), .Y(new_n25845_));
  OR4X1    g25653(.A(new_n25203_), .B(new_n25052_), .C(new_n25050_), .D(new_n25070_), .Y(new_n25846_));
  AND2X1   g25654(.A(new_n25846_), .B(new_n25845_), .Y(new_n25847_));
  INVX1    g25655(.A(new_n25847_), .Y(new_n25848_));
  NAND3X1  g25656(.A(new_n25848_), .B(new_n25843_), .C(new_n25840_), .Y(new_n25849_));
  AND2X1   g25657(.A(new_n25849_), .B(new_n481_), .Y(new_n25850_));
  OAI22X1  g25658(.A0(new_n25110_), .A1(new_n25108_), .B0(new_n25080_), .B1(new_n481_), .Y(new_n25851_));
  OAI21X1  g25659(.A0(new_n25851_), .A1(new_n25203_), .B0(new_n25109_), .Y(new_n25852_));
  AND2X1   g25660(.A(new_n25071_), .B(new_n25064_), .Y(new_n25853_));
  OR4X1    g25661(.A(new_n25203_), .B(new_n25853_), .C(new_n25109_), .D(new_n25054_), .Y(new_n25854_));
  AND2X1   g25662(.A(new_n25854_), .B(new_n25852_), .Y(new_n25855_));
  AOI21X1  g25663(.A0(new_n25843_), .A1(new_n25840_), .B0(new_n25848_), .Y(new_n25856_));
  OR2X1    g25664(.A(new_n25856_), .B(new_n25855_), .Y(new_n25857_));
  OAI21X1  g25665(.A0(new_n25857_), .A1(new_n25850_), .B0(new_n399_), .Y(new_n25858_));
  AND2X1   g25666(.A(new_n25836_), .B(new_n902_), .Y(new_n25859_));
  OR2X1    g25667(.A(new_n25818_), .B(new_n25837_), .Y(new_n25860_));
  OAI21X1  g25668(.A0(new_n25860_), .A1(new_n25859_), .B0(new_n697_), .Y(new_n25861_));
  AOI21X1  g25669(.A0(new_n25841_), .A1(new_n25818_), .B0(new_n25826_), .Y(new_n25862_));
  AOI21X1  g25670(.A0(new_n25862_), .A1(new_n25861_), .B0(\asqrt[56] ), .Y(new_n25863_));
  OR2X1    g25671(.A(new_n25838_), .B(new_n25819_), .Y(new_n25864_));
  AOI21X1  g25672(.A0(new_n25864_), .A1(new_n25861_), .B0(new_n25827_), .Y(new_n25865_));
  NOR3X1   g25673(.A(new_n25847_), .B(new_n25865_), .C(new_n25863_), .Y(new_n25866_));
  OAI21X1  g25674(.A0(new_n25865_), .A1(new_n25863_), .B0(new_n25847_), .Y(new_n25867_));
  OAI21X1  g25675(.A0(new_n25866_), .A1(\asqrt[57] ), .B0(new_n25867_), .Y(new_n25868_));
  AND2X1   g25676(.A(new_n25113_), .B(new_n25111_), .Y(new_n25869_));
  OR2X1    g25677(.A(new_n25869_), .B(new_n25112_), .Y(new_n25870_));
  OAI21X1  g25678(.A0(new_n25870_), .A1(new_n25203_), .B0(new_n25079_), .Y(new_n25871_));
  OR4X1    g25679(.A(new_n25203_), .B(new_n25869_), .C(new_n25079_), .D(new_n25112_), .Y(new_n25872_));
  AND2X1   g25680(.A(new_n25872_), .B(new_n25871_), .Y(new_n25873_));
  AOI21X1  g25681(.A0(new_n25868_), .A1(new_n25855_), .B0(new_n25873_), .Y(new_n25874_));
  AOI21X1  g25682(.A0(new_n25874_), .A1(new_n25858_), .B0(\asqrt[59] ), .Y(new_n25875_));
  NAND2X1  g25683(.A(new_n25089_), .B(new_n25115_), .Y(new_n25876_));
  OAI21X1  g25684(.A0(new_n25876_), .A1(new_n25203_), .B0(new_n25088_), .Y(new_n25877_));
  NAND4X1  g25685(.A(\asqrt[1] ), .B(new_n25089_), .C(new_n25087_), .D(new_n25115_), .Y(new_n25878_));
  AND2X1   g25686(.A(new_n25878_), .B(new_n25877_), .Y(new_n25879_));
  INVX1    g25687(.A(new_n25855_), .Y(new_n25880_));
  AOI21X1  g25688(.A0(new_n25849_), .A1(new_n481_), .B0(new_n25856_), .Y(new_n25881_));
  OR2X1    g25689(.A(new_n25881_), .B(new_n25880_), .Y(new_n25882_));
  INVX1    g25690(.A(new_n25873_), .Y(new_n25883_));
  AOI21X1  g25691(.A0(new_n25882_), .A1(new_n25858_), .B0(new_n25883_), .Y(new_n25884_));
  NOR3X1   g25692(.A(new_n25884_), .B(new_n25879_), .C(new_n25875_), .Y(new_n25885_));
  NOR2X1   g25693(.A(new_n25885_), .B(\asqrt[60] ), .Y(new_n25886_));
  OAI21X1  g25694(.A0(new_n25884_), .A1(new_n25875_), .B0(new_n25879_), .Y(new_n25887_));
  OAI22X1  g25695(.A0(new_n25099_), .A1(new_n25092_), .B0(new_n25090_), .B1(new_n292_), .Y(new_n25888_));
  OAI21X1  g25696(.A0(new_n25888_), .A1(new_n25203_), .B0(new_n25098_), .Y(new_n25889_));
  AND2X1   g25697(.A(new_n25138_), .B(new_n25137_), .Y(new_n25890_));
  OR4X1    g25698(.A(new_n25203_), .B(new_n25890_), .C(new_n25098_), .D(new_n25136_), .Y(new_n25891_));
  AND2X1   g25699(.A(new_n25891_), .B(new_n25889_), .Y(new_n25892_));
  INVX1    g25700(.A(new_n25892_), .Y(new_n25893_));
  NAND2X1  g25701(.A(new_n25893_), .B(new_n25887_), .Y(new_n25894_));
  OAI21X1  g25702(.A0(new_n25894_), .A1(new_n25886_), .B0(new_n217_), .Y(new_n25895_));
  AND2X1   g25703(.A(new_n25118_), .B(new_n25100_), .Y(new_n25896_));
  OR2X1    g25704(.A(new_n25896_), .B(new_n25101_), .Y(new_n25897_));
  OAI21X1  g25705(.A0(new_n25897_), .A1(new_n25203_), .B0(new_n25141_), .Y(new_n25898_));
  OR4X1    g25706(.A(new_n25203_), .B(new_n25896_), .C(new_n25141_), .D(new_n25101_), .Y(new_n25899_));
  AND2X1   g25707(.A(new_n25899_), .B(new_n25898_), .Y(new_n25900_));
  OAI21X1  g25708(.A0(new_n25885_), .A1(\asqrt[60] ), .B0(new_n25887_), .Y(new_n25901_));
  AOI21X1  g25709(.A0(new_n25901_), .A1(new_n25892_), .B0(new_n25900_), .Y(new_n25902_));
  AOI21X1  g25710(.A0(new_n25902_), .A1(new_n25895_), .B0(\asqrt[62] ), .Y(new_n25903_));
  INVX1    g25711(.A(new_n25900_), .Y(new_n25904_));
  NAND2X1  g25712(.A(new_n25901_), .B(new_n25892_), .Y(new_n25905_));
  AOI21X1  g25713(.A0(new_n25905_), .A1(new_n25895_), .B0(new_n25904_), .Y(new_n25906_));
  NAND2X1  g25714(.A(new_n25144_), .B(new_n25120_), .Y(new_n25907_));
  OAI21X1  g25715(.A0(new_n25907_), .A1(new_n25203_), .B0(new_n25123_), .Y(new_n25908_));
  OR4X1    g25716(.A(new_n25203_), .B(new_n25125_), .C(new_n25123_), .D(new_n25146_), .Y(new_n25909_));
  AND2X1   g25717(.A(new_n25909_), .B(new_n25908_), .Y(new_n25910_));
  AND2X1   g25718(.A(new_n25131_), .B(new_n25126_), .Y(new_n25911_));
  AND2X1   g25719(.A(new_n25911_), .B(\asqrt[1] ), .Y(new_n25912_));
  OR4X1    g25720(.A(new_n25912_), .B(new_n25910_), .C(new_n25906_), .D(new_n25157_), .Y(new_n25913_));
  OAI21X1  g25721(.A0(new_n25913_), .A1(new_n25903_), .B0(new_n193_), .Y(new_n25914_));
  OAI21X1  g25722(.A0(new_n25906_), .A1(new_n25903_), .B0(new_n25910_), .Y(new_n25915_));
  AOI21X1  g25723(.A0(\asqrt[1] ), .A1(new_n25131_), .B0(new_n25126_), .Y(new_n25916_));
  OR2X1    g25724(.A(new_n25911_), .B(new_n193_), .Y(new_n25917_));
  OR2X1    g25725(.A(new_n25917_), .B(new_n25916_), .Y(new_n25918_));
  NAND3X1  g25726(.A(new_n25918_), .B(new_n25915_), .C(new_n25914_), .Y(\asqrt[0] ));
endmodule


