//Converted to Combinational (Partial output: n70) , Module name: s1494_n70
module s1494_n70 ( v1, CLR, v7, v10, v9, v12, v2, v8, v11, v5, v4, v3, v6, v0, n70 );
input v1, CLR, v7, v10, v9, v12, v2, v8, v11, v5, v4, v3, v6, v0;
output n70;
wire n267, n365, n374, n68, n346, n364, n373, n116, n369, n62, n341, n345, n363, n349, n372, n93, n139, n160, n368, n244, n70_1, n67, n84, n45, n343, n344, n362, n354, n348, n174, n124, n272, n371, n87, n119, n366, n367, n94, n137, n342, n357, n360, n361, n350, n353, n304, n347, n107, n74, n370, n111, n136, n100, n355, n356, n358, n359, n123, n86, n352, n351, n53, n54, n64, n140, n254, n83;
AOI21X1  g329(.A0(n374), .A1(n365), .B0(n267), .Y(n70));
INVX1    g221(.A(CLR), .Y(n267));
OAI21X1  g319(.A0(n364), .A1(n346), .B0(n68), .Y(n365));
AOI22X1  g328(.A0(n369), .A1(n116), .B0(v7), .B1(n373), .Y(n374));
INVX1    g023(.A(v7), .Y(n68));
AOI21X1  g300(.A0(n345), .A1(n341), .B0(n62), .Y(n346));
OAI21X1  g318(.A0(n349), .A1(v10), .B0(n363), .Y(n364));
OAI22X1  g327(.A0(n160), .A1(n139), .B0(n93), .B1(n372), .Y(n373));
NOR2X1   g071(.A(v9), .B(v10), .Y(n116));
OAI21X1  g323(.A0(n244), .A1(v12), .B0(n368), .Y(n369));
INVX1    g017(.A(v2), .Y(n62));
NAND4X1  g295(.A(v10), .B(n84), .C(n67), .D(n70_1), .Y(n341));
OAI21X1  g299(.A0(n344), .A1(n343), .B0(n45), .Y(n345));
AOI21X1  g317(.A0(n354), .A1(n93), .B0(n362), .Y(n363));
AOI22X1  g303(.A0(n272), .A1(n124), .B0(n174), .B1(n348), .Y(n349));
AOI22X1  g326(.A0(n87), .A1(n67), .B0(n70_1), .B1(n371), .Y(n372));
INVX1    g048(.A(v8), .Y(n93));
NAND2X1  g093(.A(v11), .B(n67), .Y(n139));
NOR2X1   g114(.A(v9), .B(n45), .Y(n160));
OAI21X1  g322(.A0(n367), .A1(n366), .B0(n119), .Y(n368));
INVX1    g198(.A(n94), .Y(n244));
INVX1    g025(.A(v9), .Y(n70_1));
INVX1    g022(.A(v12), .Y(n67));
INVX1    g039(.A(v11), .Y(n84));
INVX1    g000(.A(v10), .Y(n45));
AOI21X1  g297(.A0(n342), .A1(n70_1), .B0(n137), .Y(n343));
NOR4X1   g298(.A(n70_1), .B(v11), .C(v12), .D(v8), .Y(n344));
NAND3X1  g316(.A(n361), .B(n360), .C(n357), .Y(n362));
OAI21X1  g308(.A0(n353), .A1(v9), .B0(n350), .Y(n354));
OAI22X1  g302(.A0(n74), .A1(n107), .B0(n347), .B1(n304), .Y(n348));
INVX1    g128(.A(v1), .Y(n174));
AND2X1   g078(.A(v4), .B(v5), .Y(n124));
NOR3X1   g226(.A(v9), .B(v11), .C(v12), .Y(n272));
OAI21X1  g325(.A0(n111), .A1(n84), .B0(n370), .Y(n371));
OR2X1    g042(.A(v10), .B(v11), .Y(n87));
INVX1    g073(.A(v3), .Y(n119));
NOR4X1   g320(.A(v8), .B(n67), .C(v6), .D(v7), .Y(n366));
NOR2X1   g321(.A(n93), .B(v12), .Y(n367));
NOR2X1   g049(.A(n93), .B(v11), .Y(n94));
INVX1    g091(.A(n136), .Y(n137));
NAND2X1  g296(.A(v12), .B(v1), .Y(n342));
OAI21X1  g311(.A0(n356), .A1(n355), .B0(n100), .Y(n357));
OAI21X1  g314(.A0(n359), .A1(n358), .B0(v8), .Y(n360));
NAND4X1  g315(.A(v10), .B(n84), .C(v12), .D(v9), .Y(n361));
NAND4X1  g304(.A(v9), .B(n67), .C(n86), .D(n123), .Y(n350));
AOI22X1  g307(.A0(n53), .A1(n45), .B0(n351), .B1(n352), .Y(n353));
NAND2X1  g258(.A(n93), .B(v9), .Y(n304));
INVX1    g301(.A(n54), .Y(n347));
NAND2X1  g062(.A(v11), .B(v12), .Y(n107));
NAND2X1  g029(.A(v8), .B(n62), .Y(n74));
AOI21X1  g324(.A0(v10), .A1(n84), .B0(n67), .Y(n370));
AND2X1   g066(.A(v10), .B(v2), .Y(n111));
AND2X1   g090(.A(v8), .B(v11), .Y(n136));
NAND2X1  g055(.A(v4), .B(v5), .Y(n100));
NOR3X1   g309(.A(n64), .B(v8), .C(n45), .Y(n355));
NOR4X1   g310(.A(n70_1), .B(v10), .C(n84), .D(n93), .Y(n356));
NOR3X1   g312(.A(n87), .B(v12), .C(n119), .Y(n358));
AND2X1   g313(.A(n254), .B(n140), .Y(n359));
NOR2X1   g077(.A(v10), .B(v11), .Y(n123));
INVX1    g041(.A(v6), .Y(n86));
NAND2X1  g306(.A(v11), .B(n83), .Y(n352));
NOR2X1   g305(.A(n45), .B(v12), .Y(n351));
AND2X1   g008(.A(v11), .B(v12), .Y(n53));
NOR2X1   g009(.A(v11), .B(v12), .Y(n54));
OR2X1    g019(.A(v9), .B(v12), .Y(n64));
NAND2X1  g094(.A(v10), .B(v11), .Y(n140));
AND2X1   g208(.A(v9), .B(v12), .Y(n254));
INVX1    g038(.A(v0), .Y(n83));

endmodule
