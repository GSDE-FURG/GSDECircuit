//Converted to Combinational (Partial output: n2727) , Module name: s35932_n2727 , Timestamp: 2018-12-03T15:51:09.032984 
module s35932_n2727 ( RESET, TM1, TM0, WX3071, WX3295, WX3423, WX4588, WX4716, WX3231, WX3359, WX4524, WX4652, WX3425, WX3427, WX3429, WX3431, WX3433, WX3435, WX3437, WX3439, WX3441, WX3443, WX3445, WX3447, WX3449, WX3451, WX3453, WX3455, WX3457, WX3459, WX3461, WX3463, WX3465, WX3467, WX3469, WX3471, WX3473, WX3475, WX3477, WX3479, WX3481, WX3483, WX3485, n2727 );
input RESET, TM1, TM0, WX3071, WX3295, WX3423, WX4588, WX4716, WX3231, WX3359, WX4524, WX4652, WX3425, WX3427, WX3429, WX3431, WX3433, WX3435, WX3437, WX3439, WX3441, WX3443, WX3445, WX3447, WX3449, WX3451, WX3453, WX3455, WX3457, WX3459, WX3461, WX3463, WX3465, WX3467, WX3469, WX3471, WX3473, WX3475, WX3477, WX3479, WX3481, WX3483, WX3485;
output n2727;
wire n5827, n6997, n6996, n6994_1, n5539, n6413, n6995, n6992, n6987, n6410, n6412, n6989_1, n6991, CRC_OUT_7_31, n6409_1, n6411, n6988, n6990, n7532_1, CRC_OUT_7_30, n7530, CRC_OUT_7_29, n7528, CRC_OUT_7_28, n7526, CRC_OUT_7_27, n7524, CRC_OUT_7_26, n7522_1, CRC_OUT_7_25, n7520, CRC_OUT_7_24, n7518, CRC_OUT_7_23, n7516, CRC_OUT_7_22, n7514, CRC_OUT_7_21, n7512_1, CRC_OUT_7_20, n7510, CRC_OUT_7_19, n7508, CRC_OUT_7_18, n7506, CRC_OUT_7_17, n7504, CRC_OUT_7_16, n7502_1, CRC_OUT_7_15, n7501, n7499, CRC_OUT_7_14, n7497_1, CRC_OUT_7_13, n7495, CRC_OUT_7_12, n7493, CRC_OUT_7_11, n7491, CRC_OUT_7_10, n7490, n7488, CRC_OUT_7_9, n7486, CRC_OUT_7_8, n7484, CRC_OUT_7_7, n7482_1, CRC_OUT_7_6, n7480, CRC_OUT_7_5, n7478, CRC_OUT_7_4, n7476, CRC_OUT_7_3, n7475, n7473, CRC_OUT_7_2, n7471, CRC_OUT_7_1, n7469, CRC_OUT_7_0, n7467_1;
NOR2X1   g1394(.A(n6997), .B(n5827), .Y(n2727));
INVX1    g0288(.A(RESET), .Y(n5827));
MX2X1    g1393(.A(n6994_1), .B(n6996), .S0(TM1), .Y(n6997));
MX2X1    g1392(.A(n6995), .B(n6413), .S0(n5539), .Y(n6996));
MX2X1    g1390(.A(n6987), .B(n6992), .S0(n5539), .Y(n6994_1));
INVX1    g0000(.A(TM0), .Y(n5539));
XOR2X1   g0842(.A(n6412), .B(n6410), .Y(n6413));
INVX1    g1391(.A(WX3071), .Y(n6995));
XOR2X1   g1389(.A(n6991), .B(n6989_1), .Y(n6992));
INVX1    g1384(.A(CRC_OUT_7_31), .Y(n6987));
XOR2X1   g0839(.A(n6409_1), .B(WX3295), .Y(n6410));
XOR2X1   g0841(.A(WX3423), .B(n6411), .Y(n6412));
XOR2X1   g1386(.A(n6988), .B(WX4588), .Y(n6989_1));
XOR2X1   g1388(.A(WX4716), .B(n6990), .Y(n6991));
NOR2X1   g1898(.A(n7532_1), .B(n5827), .Y(CRC_OUT_7_31));
XOR2X1   g0838(.A(WX3231), .B(TM1), .Y(n6409_1));
INVX1    g0840(.A(WX3359), .Y(n6411));
XOR2X1   g1385(.A(WX4524), .B(TM1), .Y(n6988));
INVX1    g1387(.A(WX4652), .Y(n6990));
XOR2X1   g1897(.A(CRC_OUT_7_30), .B(WX3423), .Y(n7532_1));
NOR2X1   g1896(.A(n7530), .B(n5827), .Y(CRC_OUT_7_30));
XOR2X1   g1895(.A(CRC_OUT_7_29), .B(WX3425), .Y(n7530));
NOR2X1   g1894(.A(n7528), .B(n5827), .Y(CRC_OUT_7_29));
XOR2X1   g1893(.A(CRC_OUT_7_28), .B(WX3427), .Y(n7528));
NOR2X1   g1892(.A(n7526), .B(n5827), .Y(CRC_OUT_7_28));
XOR2X1   g1891(.A(CRC_OUT_7_27), .B(WX3429), .Y(n7526));
NOR2X1   g1890(.A(n7524), .B(n5827), .Y(CRC_OUT_7_27));
XOR2X1   g1889(.A(CRC_OUT_7_26), .B(WX3431), .Y(n7524));
NOR2X1   g1888(.A(n7522_1), .B(n5827), .Y(CRC_OUT_7_26));
XOR2X1   g1887(.A(CRC_OUT_7_25), .B(WX3433), .Y(n7522_1));
NOR2X1   g1886(.A(n7520), .B(n5827), .Y(CRC_OUT_7_25));
XOR2X1   g1885(.A(CRC_OUT_7_24), .B(WX3435), .Y(n7520));
NOR2X1   g1884(.A(n7518), .B(n5827), .Y(CRC_OUT_7_24));
XOR2X1   g1883(.A(CRC_OUT_7_23), .B(WX3437), .Y(n7518));
NOR2X1   g1882(.A(n7516), .B(n5827), .Y(CRC_OUT_7_23));
XOR2X1   g1881(.A(CRC_OUT_7_22), .B(WX3439), .Y(n7516));
NOR2X1   g1880(.A(n7514), .B(n5827), .Y(CRC_OUT_7_22));
XOR2X1   g1879(.A(CRC_OUT_7_21), .B(WX3441), .Y(n7514));
NOR2X1   g1878(.A(n7512_1), .B(n5827), .Y(CRC_OUT_7_21));
XOR2X1   g1877(.A(CRC_OUT_7_20), .B(WX3443), .Y(n7512_1));
NOR2X1   g1876(.A(n7510), .B(n5827), .Y(CRC_OUT_7_20));
XOR2X1   g1875(.A(CRC_OUT_7_19), .B(WX3445), .Y(n7510));
NOR2X1   g1874(.A(n7508), .B(n5827), .Y(CRC_OUT_7_19));
XOR2X1   g1873(.A(CRC_OUT_7_18), .B(WX3447), .Y(n7508));
NOR2X1   g1872(.A(n7506), .B(n5827), .Y(CRC_OUT_7_18));
XOR2X1   g1871(.A(CRC_OUT_7_17), .B(WX3449), .Y(n7506));
NOR2X1   g1870(.A(n7504), .B(n5827), .Y(CRC_OUT_7_17));
XOR2X1   g1869(.A(CRC_OUT_7_16), .B(WX3451), .Y(n7504));
NOR2X1   g1868(.A(n7502_1), .B(n5827), .Y(CRC_OUT_7_16));
XOR2X1   g1867(.A(n7501), .B(CRC_OUT_7_15), .Y(n7502_1));
NOR2X1   g1865(.A(n7499), .B(n5827), .Y(CRC_OUT_7_15));
XOR2X1   g1866(.A(CRC_OUT_7_31), .B(WX3453), .Y(n7501));
XOR2X1   g1864(.A(CRC_OUT_7_14), .B(WX3455), .Y(n7499));
NOR2X1   g1863(.A(n7497_1), .B(n5827), .Y(CRC_OUT_7_14));
XOR2X1   g1862(.A(CRC_OUT_7_13), .B(WX3457), .Y(n7497_1));
NOR2X1   g1861(.A(n7495), .B(n5827), .Y(CRC_OUT_7_13));
XOR2X1   g1860(.A(CRC_OUT_7_12), .B(WX3459), .Y(n7495));
NOR2X1   g1859(.A(n7493), .B(n5827), .Y(CRC_OUT_7_12));
XOR2X1   g1858(.A(CRC_OUT_7_11), .B(WX3461), .Y(n7493));
NOR2X1   g1857(.A(n7491), .B(n5827), .Y(CRC_OUT_7_11));
XOR2X1   g1856(.A(n7490), .B(CRC_OUT_7_10), .Y(n7491));
NOR2X1   g1854(.A(n7488), .B(n5827), .Y(CRC_OUT_7_10));
XOR2X1   g1855(.A(CRC_OUT_7_31), .B(WX3463), .Y(n7490));
XOR2X1   g1853(.A(CRC_OUT_7_9), .B(WX3465), .Y(n7488));
NOR2X1   g1852(.A(n7486), .B(n5827), .Y(CRC_OUT_7_9));
XOR2X1   g1851(.A(CRC_OUT_7_8), .B(WX3467), .Y(n7486));
NOR2X1   g1850(.A(n7484), .B(n5827), .Y(CRC_OUT_7_8));
XOR2X1   g1849(.A(CRC_OUT_7_7), .B(WX3469), .Y(n7484));
NOR2X1   g1848(.A(n7482_1), .B(n5827), .Y(CRC_OUT_7_7));
XOR2X1   g1847(.A(CRC_OUT_7_6), .B(WX3471), .Y(n7482_1));
NOR2X1   g1846(.A(n7480), .B(n5827), .Y(CRC_OUT_7_6));
XOR2X1   g1845(.A(CRC_OUT_7_5), .B(WX3473), .Y(n7480));
NOR2X1   g1844(.A(n7478), .B(n5827), .Y(CRC_OUT_7_5));
XOR2X1   g1843(.A(CRC_OUT_7_4), .B(WX3475), .Y(n7478));
NOR2X1   g1842(.A(n7476), .B(n5827), .Y(CRC_OUT_7_4));
XOR2X1   g1841(.A(n7475), .B(CRC_OUT_7_3), .Y(n7476));
NOR2X1   g1839(.A(n7473), .B(n5827), .Y(CRC_OUT_7_3));
XOR2X1   g1840(.A(CRC_OUT_7_31), .B(WX3477), .Y(n7475));
XOR2X1   g1838(.A(CRC_OUT_7_2), .B(WX3479), .Y(n7473));
NOR2X1   g1837(.A(n7471), .B(n5827), .Y(CRC_OUT_7_2));
XOR2X1   g1836(.A(CRC_OUT_7_1), .B(WX3481), .Y(n7471));
NOR2X1   g1835(.A(n7469), .B(n5827), .Y(CRC_OUT_7_1));
XOR2X1   g1834(.A(CRC_OUT_7_0), .B(WX3483), .Y(n7469));
NOR2X1   g1833(.A(n7467_1), .B(n5827), .Y(CRC_OUT_7_0));
XOR2X1   g1832(.A(CRC_OUT_7_31), .B(WX3485), .Y(n7467_1));

endmodule
