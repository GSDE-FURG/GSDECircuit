//Converted to Combinational (Partial output: g10379) , Module name: s15850_g10379 , Timestamp: 2018-12-03T15:51:07.632441 
module s15850_g10379 ( g30, g41, g31, g48, g1191, g1311, g284, g919, g947, g1741, g40, g1589, g1546, g46, g43, g45, g47, g44, g42, g10379 );
input g30, g41, g31, g48, g1191, g1311, g284, g919, g947, g1741, g40, g1589, g1546, g46, g43, g45, g47, g44, g42;
output g10379;
wire n1892, n2004, n1887, n2003, n1994, n1997_1, n2000, n1959, n2001, n2002_1, n1993, n1987_1, n1989, n1990, n1996, n1903, n1909_1, n1995, n1931, n1943, n1999, n1944, n1902, n1908, n1938_1, n1900_1, n1992_1, n1927, n1986, n1950, n1915, n1910, n1897, n1905_1, n1911, n1930, n1923, n1925, n1934, n1939, n1942_1, n1998, n1899, n1940, n1885_1, n1896, n1901, n1907, n1937, n1895_1, n1991, n1894, n1906, n1926, n1919_1, n1924_1, n1949, n1913, n1914_1, n1893, n1904, n1928_1, n1929, n1922, n1933_1, n1936, n1941, n1884, n1898, n1918, n1920, n1921, n1932, n1935;
NAND2X1  g0174(.A(n2004), .B(n1892), .Y(g10379));
NOR4X1   g0063(.A(g31), .B(g41), .C(n1887), .D(g30), .Y(n1892));
NOR4X1   g0173(.A(n2000), .B(n1997_1), .C(n1994), .D(n2003), .Y(n2004));
INVX1    g0058(.A(g48), .Y(n1887));
AOI21X1  g0172(.A0(n2002_1), .A1(n2001), .B0(n1959), .Y(n2003));
NAND4X1  g0163(.A(n1990), .B(n1989), .C(n1987_1), .D(n1993), .Y(n1994));
OAI22X1  g0166(.A0(n1995), .A1(n1909_1), .B0(n1903), .B1(n1996), .Y(n1997_1));
NOR3X1   g0169(.A(n1999), .B(n1943), .C(n1931), .Y(n2000));
OAI21X1  g0130(.A0(n1908), .A1(n1902), .B0(n1944), .Y(n1959));
NAND3X1  g0170(.A(n1944), .B(n1908), .C(g1191), .Y(n2001));
NAND3X1  g0171(.A(n1944), .B(n1902), .C(g1311), .Y(n2002_1));
NAND4X1  g0162(.A(n1992_1), .B(n1900_1), .C(g284), .D(n1938_1), .Y(n1993));
AOI22X1  g0157(.A0(n1986), .A1(g947), .B0(g919), .B1(n1927), .Y(n1987_1));
NAND3X1  g0158(.A(n1950), .B(n1944), .C(g1741), .Y(n1989));
OAI21X1  g0159(.A0(g31), .A1(n1887), .B0(g40), .Y(n1990));
OAI21X1  g0165(.A0(n1910), .A1(n1915), .B0(g1589), .Y(n1996));
OAI21X1  g0074(.A0(n1902), .A1(n1897), .B0(n1900_1), .Y(n1903));
OAI21X1  g0080(.A0(n1908), .A1(n1905_1), .B0(n1900_1), .Y(n1909_1));
OAI21X1  g0164(.A0(n1911), .A1(n1910), .B0(g1546), .Y(n1995));
OR4X1    g0102(.A(n1927), .B(n1925), .C(n1923), .D(n1930), .Y(n1931));
NAND3X1  g0114(.A(n1942_1), .B(n1939), .C(n1934), .Y(n1943));
NAND4X1  g0168(.A(n1998), .B(n1909_1), .C(n1903), .D(n1959), .Y(n1999));
NOR4X1   g0115(.A(n1885_1), .B(n1940), .C(g46), .D(n1899), .Y(n1944));
NOR4X1   g0073(.A(g41), .B(n1887), .C(n1901), .D(n1896), .Y(n1902));
NOR4X1   g0079(.A(g41), .B(n1887), .C(n1901), .D(n1907), .Y(n1908));
NOR4X1   g0109(.A(n1895_1), .B(g45), .C(g43), .D(n1937), .Y(n1938_1));
NOR4X1   g0071(.A(n1885_1), .B(g47), .C(g46), .D(n1899), .Y(n1900_1));
NAND4X1  g0161(.A(g44), .B(n1906), .C(n1894), .D(n1991), .Y(n1992_1));
NOR2X1   g0098(.A(n1919_1), .B(n1926), .Y(n1927));
NOR2X1   g0156(.A(n1919_1), .B(n1924_1), .Y(n1986));
NOR4X1   g0121(.A(g41), .B(n1887), .C(n1901), .D(n1949), .Y(n1950));
NAND3X1  g0086(.A(n1914_1), .B(n1913), .C(g48), .Y(n1915));
OR4X1    g0081(.A(n1885_1), .B(g47), .C(g46), .D(n1899), .Y(n1910));
NOR3X1   g0068(.A(n1896), .B(n1893), .C(n1887), .Y(n1897));
AND2X1   g0076(.A(n1904), .B(g48), .Y(n1905_1));
NAND2X1  g0082(.A(n1904), .B(g48), .Y(n1911));
NOR3X1   g0101(.A(n1929), .B(n1919_1), .C(n1928_1), .Y(n1930));
AOI21X1  g0094(.A0(n1922), .A1(n1911), .B0(n1919_1), .Y(n1923));
AOI21X1  g0096(.A0(n1924_1), .A1(n1915), .B0(n1919_1), .Y(n1925));
INVX1    g0105(.A(n1933_1), .Y(n1934));
OAI21X1  g0110(.A0(n1938_1), .A1(n1936), .B0(n1900_1), .Y(n1939));
OR4X1    g0113(.A(n1899), .B(n1885_1), .C(n1940), .D(n1941), .Y(n1942_1));
NAND2X1  g0167(.A(n1950), .B(n1944), .Y(n1998));
OAI21X1  g0070(.A0(n1898), .A1(g48), .B0(n1884), .Y(n1899));
INVX1    g0111(.A(g47), .Y(n1940));
AND2X1   g0056(.A(g31), .B(g48), .Y(n1885_1));
NAND3X1  g0067(.A(n1895_1), .B(g45), .C(n1894), .Y(n1896));
INVX1    g0072(.A(g42), .Y(n1901));
NAND3X1  g0078(.A(g44), .B(n1906), .C(g43), .Y(n1907));
NAND3X1  g0108(.A(n1884), .B(g48), .C(g42), .Y(n1937));
INVX1    g0066(.A(g44), .Y(n1895_1));
NOR3X1   g0160(.A(g41), .B(n1887), .C(g42), .Y(n1991));
INVX1    g0065(.A(g43), .Y(n1894));
INVX1    g0077(.A(g45), .Y(n1906));
OR4X1    g0097(.A(g41), .B(n1887), .C(n1901), .D(n1907), .Y(n1926));
OR4X1    g0090(.A(n1885_1), .B(g47), .C(n1918), .D(n1899), .Y(n1919_1));
NAND4X1  g0095(.A(n1884), .B(g48), .C(g42), .D(n1914_1), .Y(n1924_1));
NAND3X1  g0120(.A(g44), .B(g45), .C(g43), .Y(n1949));
NOR2X1   g0084(.A(g41), .B(g42), .Y(n1913));
NOR3X1   g0085(.A(g44), .B(n1906), .C(g43), .Y(n1914_1));
OR2X1    g0064(.A(g41), .B(g42), .Y(n1893));
NOR4X1   g0075(.A(n1895_1), .B(g45), .C(n1894), .D(n1893), .Y(n1904));
NAND2X1  g0099(.A(n1895_1), .B(g45), .Y(n1928_1));
NAND4X1  g0100(.A(n1884), .B(g48), .C(g42), .D(g43), .Y(n1929));
OR2X1    g0093(.A(n1921), .B(n1920), .Y(n1922));
NAND2X1  g0104(.A(n1932), .B(g48), .Y(n1933_1));
NOR4X1   g0107(.A(n1895_1), .B(g45), .C(g43), .D(n1935), .Y(n1936));
NAND3X1  g0112(.A(n1904), .B(g46), .C(g48), .Y(n1941));
INVX1    g0055(.A(g41), .Y(n1884));
INVX1    g0069(.A(g30), .Y(n1898));
INVX1    g0089(.A(g46), .Y(n1918));
NAND2X1  g0091(.A(g44), .B(g45), .Y(n1920));
NAND4X1  g0092(.A(n1884), .B(g48), .C(g42), .D(n1894), .Y(n1921));
INVX1    g0103(.A(g31), .Y(n1932));
NAND3X1  g0106(.A(n1884), .B(g48), .C(n1901), .Y(n1935));

endmodule
