//Converted to Combinational , Module name: s1238 , Timestamp: 2018-12-03T15:51:02.329060 
module s1238 ( G0, G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G40, G41, G42, G43, G44, G46, G549, G550, G551, G552, G542, G546, G547, G548, G530, G532, G535, G537, G45, G539, n57, n62, n67, n72, n77, n82, n87, n92, n97, n102, n107, n112, n117, n122, n127, n132, n141 );
input G0, G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G40, G41, G42, G43, G44, G46;
output G549, G550, G551, G552, G542, G546, G547, G548, G530, G532, G535, G537, G45, G539, n57, n62, n67, n72, n77, n82, n87, n92, n97, n102, n107, n112, n117, n122, n127, n132, n141;
wire n82_1, n83, n84, n85, n86, n87_1, n88, n89, n90, n91, n92_1, n93, n94, n95, n96, n97_1, n98, n99, n100, n101, n102_1, n103, n104, n105, n106, n107_1, n108, n109, n110, n111, n112_1, n113, n114, n115, n116, n117_1, n118, n119, n120, n121, n122_1, n123, n124, n125, n126, n127_1, n128, n129, n130, n131, n132_1, n133, n134, n135, n136, n137_1, n138, n139, n140, n141_1, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n230, n231, n232, n233, n234, n235, n236, n237, n239, n240, n241, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n364, n365, n366, n368, n372, n373, n375, n376, n378, n380, n382, n387, n388, n389, n390, n392, n393, n394, n396, n397, n398, n399, n401, n402, n403, n404, n406, n407, n408, n410, n411, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424;
INVX1    g000(.A(G12), .Y(n82_1));
INVX1    g001(.A(G4), .Y(n83));
NOR2X1   g002(.A(G5), .B(n83), .Y(n84));
INVX1    g003(.A(G0), .Y(n85));
NAND3X1  g004(.A(n83), .B(G3), .C(n85), .Y(n86));
INVX1    g005(.A(G5), .Y(n87_1));
NOR3X1   g006(.A(G3), .B(G2), .C(n85), .Y(n88));
INVX1    g007(.A(G2), .Y(n89));
INVX1    g008(.A(G3), .Y(n90));
INVX1    g009(.A(G1), .Y(n91));
NAND2X1  g010(.A(G5), .B(G3), .Y(n92_1));
AOI22X1  g011(.A0(G5), .A1(n91), .B0(G4), .B1(n92_1), .Y(n93));
OAI21X1  g012(.A0(n93), .A1(n89), .B0(n90), .Y(n94));
AOI21X1  g013(.A0(n94), .A1(G0), .B0(G4), .Y(n95));
OAI21X1  g014(.A0(n95), .A1(n88), .B0(n87_1), .Y(n96));
AOI21X1  g015(.A0(n96), .A1(n86), .B0(n84), .Y(n97_1));
INVX1    g016(.A(G46), .Y(n98));
INVX1    g017(.A(G11), .Y(n99));
INVX1    g018(.A(G8), .Y(n100));
INVX1    g019(.A(G7), .Y(n101));
INVX1    g020(.A(G30), .Y(n102_1));
NOR3X1   g021(.A(n102_1), .B(n101), .C(G6), .Y(n103));
INVX1    g022(.A(G9), .Y(n104));
AND2X1   g023(.A(G10), .B(G8), .Y(n105));
NOR2X1   g024(.A(n105), .B(n104), .Y(n106));
OR4X1    g025(.A(n103), .B(G31), .C(n100), .D(n106), .Y(n107_1));
NOR3X1   g026(.A(G9), .B(G8), .C(G7), .Y(n108));
NOR2X1   g027(.A(G30), .B(G6), .Y(n109));
NOR2X1   g028(.A(n109), .B(n108), .Y(n110));
AOI21X1  g029(.A0(n110), .A1(n107_1), .B0(n99), .Y(n111));
NOR2X1   g030(.A(G11), .B(G10), .Y(n112_1));
NAND2X1  g031(.A(n112_1), .B(n104), .Y(n113));
AND2X1   g032(.A(G31), .B(G8), .Y(n114));
NOR3X1   g033(.A(n114), .B(n113), .C(n103), .Y(n115));
INVX1    g034(.A(G10), .Y(n116));
MX2X1    g035(.A(n116), .B(G31), .S0(G8), .Y(n117_1));
NOR4X1   g036(.A(G11), .B(n104), .C(G7), .D(n117_1), .Y(n118));
OR4X1    g037(.A(n115), .B(n111), .C(n98), .D(n118), .Y(n119));
OR4X1    g038(.A(n97_1), .B(G13), .C(n82_1), .D(n119), .Y(n120));
AND2X1   g039(.A(G4), .B(G1), .Y(n121));
NAND2X1  g040(.A(G3), .B(G0), .Y(n122_1));
NAND2X1  g041(.A(n122_1), .B(n121), .Y(n123));
AND2X1   g042(.A(G11), .B(G9), .Y(n124));
NAND2X1  g043(.A(G10), .B(G7), .Y(n125));
AOI21X1  g044(.A0(n124), .A1(G8), .B0(n125), .Y(n126));
NAND2X1  g045(.A(n116), .B(G9), .Y(n127_1));
NAND2X1  g046(.A(G8), .B(n101), .Y(n128));
OAI22X1  g047(.A0(n127_1), .A1(n101), .B0(n102_1), .B1(n128), .Y(n129));
INVX1    g048(.A(G6), .Y(n130));
XOR2X1   g049(.A(G3), .B(G2), .Y(n131));
AOI21X1  g050(.A0(n92_1), .A1(G4), .B0(n131), .Y(n132_1));
OR2X1    g051(.A(n132_1), .B(n130), .Y(n133));
AND2X1   g052(.A(G6), .B(G4), .Y(n134));
OR2X1    g053(.A(G6), .B(G4), .Y(n135));
OAI21X1  g054(.A0(n134), .A1(n90), .B0(n135), .Y(n136));
AOI22X1  g055(.A0(n84), .A1(n90), .B0(G5), .B1(n136), .Y(n137_1));
AOI21X1  g056(.A0(n137_1), .A1(n133), .B0(n91), .Y(n138));
OAI21X1  g057(.A0(n130), .A1(G4), .B0(n87_1), .Y(n139));
NOR2X1   g058(.A(n89), .B(G1), .Y(n140));
NAND2X1  g059(.A(n140), .B(n139), .Y(n141_1));
AOI21X1  g060(.A0(G4), .A1(G1), .B0(G5), .Y(n142));
NAND2X1  g061(.A(n130), .B(G2), .Y(n143));
OAI21X1  g062(.A0(n143), .A1(n142), .B0(n141_1), .Y(n144));
OAI22X1  g063(.A0(n138), .A1(n144), .B0(n129), .B1(n126), .Y(n145));
NOR2X1   g064(.A(n145), .B(n91), .Y(n146));
MX2X1    g065(.A(n89), .B(n134), .S0(n90), .Y(n147));
NAND2X1  g066(.A(n147), .B(G5), .Y(n148));
NAND3X1  g067(.A(G6), .B(n90), .C(G2), .Y(n149));
OAI21X1  g068(.A0(n130), .A1(G3), .B0(G5), .Y(n150));
AOI21X1  g069(.A0(n150), .A1(n149), .B0(G4), .Y(n151));
NOR3X1   g070(.A(G5), .B(n83), .C(n89), .Y(n152));
NOR2X1   g071(.A(n152), .B(n151), .Y(n153));
INVX1    g072(.A(G13), .Y(n154));
NOR2X1   g073(.A(n154), .B(G12), .Y(n155));
INVX1    g074(.A(n155), .Y(n156));
AOI21X1  g075(.A0(n153), .A1(n148), .B0(n156), .Y(n157));
NOR2X1   g076(.A(G33), .B(G13), .Y(n158));
NAND2X1  g077(.A(n158), .B(G3), .Y(n159));
INVX1    g078(.A(G32), .Y(n160));
NOR2X1   g079(.A(n129), .B(n126), .Y(n161));
NOR4X1   g080(.A(n160), .B(G13), .C(G12), .D(n161), .Y(n162));
INVX1    g081(.A(n162), .Y(n163));
AND2X1   g082(.A(G5), .B(G2), .Y(n164));
OAI21X1  g083(.A0(n83), .A1(n90), .B0(n164), .Y(n165));
OAI21X1  g084(.A0(n165), .A1(n163), .B0(n159), .Y(n166));
AOI21X1  g085(.A0(n157), .A1(n146), .B0(n166), .Y(n167));
OAI21X1  g086(.A0(n123), .A1(n120), .B0(n167), .Y(G549));
NOR4X1   g087(.A(n90), .B(n91), .C(G0), .D(n83), .Y(n169));
NOR2X1   g088(.A(G29), .B(n85), .Y(n170));
NOR2X1   g089(.A(n170), .B(n169), .Y(n171));
OR2X1    g090(.A(n121), .B(n87_1), .Y(n172));
OR4X1    g091(.A(G5), .B(n83), .C(n91), .D(n145), .Y(n173));
OAI21X1  g092(.A0(n172), .A1(n145), .B0(n173), .Y(n174));
NOR3X1   g093(.A(n154), .B(G12), .C(n89), .Y(n175));
INVX1    g094(.A(n92_1), .Y(n176));
OAI21X1  g095(.A0(n83), .A1(n89), .B0(n176), .Y(n177));
OAI21X1  g096(.A0(n177), .A1(n163), .B0(n159), .Y(n178));
AOI21X1  g097(.A0(n175), .A1(n174), .B0(n178), .Y(n179));
OAI21X1  g098(.A0(n171), .A1(n120), .B0(n179), .Y(G550));
NOR3X1   g099(.A(n119), .B(n97_1), .C(n82_1), .Y(n181));
AND2X1   g100(.A(G2), .B(G0), .Y(n182));
MX2X1    g101(.A(n91), .B(n83), .S0(n182), .Y(n183));
MX2X1    g102(.A(n122_1), .B(G0), .S0(n121), .Y(n184));
OAI21X1  g103(.A0(n183), .A1(G3), .B0(n184), .Y(n185));
NAND4X1  g104(.A(n181), .B(n154), .C(G5), .D(n185), .Y(n186));
OR4X1    g105(.A(n83), .B(n89), .C(G1), .D(n145), .Y(n187));
NOR2X1   g106(.A(n90), .B(G2), .Y(n188));
NOR2X1   g107(.A(n144), .B(n138), .Y(n189));
NOR2X1   g108(.A(n189), .B(n161), .Y(n190));
NAND3X1  g109(.A(n190), .B(n188), .C(n121), .Y(n191));
AOI21X1  g110(.A0(n191), .A1(n187), .B0(n87_1), .Y(n192));
NOR3X1   g111(.A(n130), .B(n90), .C(G2), .Y(n193));
INVX1    g112(.A(n84), .Y(n194));
NAND2X1  g113(.A(G6), .B(G4), .Y(n195));
OAI22X1  g114(.A0(n188), .A1(n194), .B0(G3), .B1(n195), .Y(n196));
AOI21X1  g115(.A0(n193), .A1(n87_1), .B0(n196), .Y(n197));
NOR3X1   g116(.A(n197), .B(n145), .C(n91), .Y(n198));
OAI21X1  g117(.A0(n198), .A1(n192), .B0(n155), .Y(n199));
NAND3X1  g118(.A(n162), .B(G39), .C(G4), .Y(n200));
NAND3X1  g119(.A(n200), .B(n199), .C(n186), .Y(G551));
INVX1    g120(.A(n193), .Y(n202));
XOR2X1   g121(.A(G5), .B(G4), .Y(n203));
AOI22X1  g122(.A0(n134), .A1(n90), .B0(G6), .B1(n203), .Y(n204));
OAI22X1  g123(.A0(n202), .A1(n84), .B0(n89), .B1(n204), .Y(n205));
OR4X1    g124(.A(n130), .B(n83), .C(n91), .D(n164), .Y(n206));
OAI22X1  g125(.A0(G4), .A1(G3), .B0(G1), .B1(n84), .Y(n207));
NOR3X1   g126(.A(n92_1), .B(G4), .C(n91), .Y(n208));
AOI21X1  g127(.A0(n207), .A1(G2), .B0(n208), .Y(n209));
OAI21X1  g128(.A0(n209), .A1(n130), .B0(n206), .Y(n210));
AND2X1   g129(.A(n210), .B(n155), .Y(n211));
AOI22X1  g130(.A0(n205), .A1(n162), .B0(n190), .B1(n211), .Y(n212));
OAI21X1  g131(.A0(n120), .A1(G40), .B0(n212), .Y(G552));
NOR3X1   g132(.A(G10), .B(n104), .C(n101), .Y(n214));
INVX1    g133(.A(G34), .Y(n215));
OAI22X1  g134(.A0(n215), .A1(n100), .B0(n130), .B1(n120), .Y(n216));
NAND2X1  g135(.A(n216), .B(n214), .Y(n217));
INVX1    g136(.A(n125), .Y(n218));
NOR2X1   g137(.A(n120), .B(n130), .Y(n219));
AOI21X1  g138(.A0(G9), .A1(G8), .B0(n215), .Y(n220));
NAND2X1  g139(.A(n100), .B(G7), .Y(n221));
MX2X1    g140(.A(n116), .B(n221), .S0(G11), .Y(n222));
NAND2X1  g141(.A(G9), .B(G7), .Y(n223));
NOR4X1   g142(.A(n116), .B(n104), .C(G8), .D(n99), .Y(n224));
AOI21X1  g143(.A0(n223), .A1(n105), .B0(n224), .Y(n225));
OAI21X1  g144(.A0(n222), .A1(G9), .B0(n225), .Y(n226));
AOI22X1  g145(.A0(n220), .A1(n218), .B0(n219), .B1(n226), .Y(n227));
NAND2X1  g146(.A(n227), .B(n217), .Y(G542));
INVX1    g147(.A(G41), .Y(G546));
XOR2X1   g148(.A(n105), .B(G7), .Y(n230));
NAND3X1  g149(.A(n230), .B(G34), .C(G9), .Y(n231));
NOR3X1   g150(.A(n125), .B(n104), .C(G6), .Y(n232));
MX2X1    g151(.A(n104), .B(n99), .S0(n116), .Y(n233));
INVX1    g152(.A(n127_1), .Y(n234));
AOI22X1  g153(.A0(n234), .A1(n128), .B0(n124), .B1(n100), .Y(n235));
OAI21X1  g154(.A0(n233), .A1(n128), .B0(n235), .Y(n236));
AOI21X1  g155(.A0(n236), .A1(G6), .B0(n232), .Y(n237));
OAI21X1  g156(.A0(n237), .A1(n120), .B0(n231), .Y(G547));
NOR4X1   g157(.A(n99), .B(n104), .C(n101), .D(n105), .Y(n239));
OAI22X1  g158(.A0(n234), .A1(n128), .B0(n125), .B1(G9), .Y(n240));
AOI21X1  g159(.A0(n240), .A1(G11), .B0(n239), .Y(n241));
OAI22X1  g160(.A0(n120), .A1(G42), .B0(n215), .B1(n241), .Y(G548));
AOI21X1  g161(.A0(G5), .A1(n90), .B0(G4), .Y(n243));
NOR3X1   g162(.A(n243), .B(n91), .C(G0), .Y(n244));
AND2X1   g163(.A(G3), .B(G1), .Y(n245));
AOI22X1  g164(.A0(n176), .A1(n83), .B0(n87_1), .B1(n245), .Y(n246));
AOI21X1  g165(.A0(n246), .A1(n93), .B0(n85), .Y(n247));
OAI21X1  g166(.A0(n247), .A1(n244), .B0(G2), .Y(n248));
INVX1    g167(.A(G36), .Y(n249));
NOR4X1   g168(.A(n104), .B(G8), .C(G7), .D(n116), .Y(n250));
NOR4X1   g169(.A(G9), .B(n100), .C(n101), .D(G10), .Y(n251));
NOR2X1   g170(.A(n251), .B(n250), .Y(n252));
NAND4X1  g171(.A(G6), .B(G5), .C(G4), .D(G11), .Y(n253));
OAI22X1  g172(.A0(n252), .A1(n253), .B0(n249), .B1(G6), .Y(n254));
AND2X1   g173(.A(n254), .B(n90), .Y(n255));
INVX1    g174(.A(n255), .Y(n256));
OR2X1    g175(.A(n251), .B(n250), .Y(n257));
NOR4X1   g176(.A(n104), .B(n100), .C(G7), .D(G10), .Y(n258));
NAND3X1  g177(.A(G6), .B(G4), .C(G3), .Y(n259));
NOR4X1   g178(.A(n99), .B(G5), .C(G2), .D(n259), .Y(n260));
OAI21X1  g179(.A0(n258), .A1(n257), .B0(n260), .Y(n261));
NOR3X1   g180(.A(G11), .B(G8), .C(G7), .Y(n262));
NAND4X1  g181(.A(n116), .B(G9), .C(G5), .D(n262), .Y(n263));
NOR2X1   g182(.A(n263), .B(n259), .Y(n264));
NAND3X1  g183(.A(G11), .B(G9), .C(G8), .Y(n265));
NOR4X1   g184(.A(n125), .B(n265), .C(n92_1), .D(n195), .Y(n266));
NAND3X1  g185(.A(G35), .B(G11), .C(G3), .Y(n267));
NOR3X1   g186(.A(n267), .B(G5), .C(G4), .Y(n268));
NOR3X1   g187(.A(n268), .B(n266), .C(n264), .Y(n269));
OAI21X1  g188(.A0(n269), .A1(n89), .B0(n261), .Y(n270));
AOI21X1  g189(.A0(n255), .A1(n89), .B0(n270), .Y(n271));
OAI21X1  g190(.A0(n161), .A1(n160), .B0(n154), .Y(n272));
OR4X1    g191(.A(n271), .B(G12), .C(G2), .D(n272), .Y(n273));
OAI22X1  g192(.A0(n256), .A1(n273), .B0(n248), .B1(n120), .Y(G530));
OR2X1    g193(.A(n245), .B(n89), .Y(n275));
NOR2X1   g194(.A(G5), .B(G3), .Y(n276));
AOI21X1  g195(.A0(n176), .A1(n89), .B0(n276), .Y(n277));
AOI21X1  g196(.A0(n277), .A1(n275), .B0(n83), .Y(n278));
NAND4X1  g197(.A(n90), .B(n89), .C(G1), .D(G5), .Y(n279));
NAND2X1  g198(.A(n245), .B(n83), .Y(n280));
NAND2X1  g199(.A(n280), .B(n279), .Y(n281));
OAI21X1  g200(.A0(n281), .A1(n278), .B0(G0), .Y(n282));
NOR2X1   g201(.A(n259), .B(G1), .Y(n283));
NOR4X1   g202(.A(G4), .B(n90), .C(n91), .D(n130), .Y(n284));
OR2X1    g203(.A(n283), .B(n284), .Y(n285));
NOR2X1   g204(.A(n265), .B(G10), .Y(n286));
AOI22X1  g205(.A0(n285), .A1(n224), .B0(n283), .B1(n286), .Y(n287));
NAND4X1  g206(.A(n116), .B(n104), .C(G7), .D(G11), .Y(n288));
NOR4X1   g207(.A(G8), .B(n90), .C(G1), .D(n135), .Y(n289));
AOI21X1  g208(.A0(n285), .A1(G8), .B0(n289), .Y(n290));
OAI22X1  g209(.A0(n288), .A1(n290), .B0(n287), .B1(G7), .Y(n291));
NOR2X1   g210(.A(G5), .B(n89), .Y(n292));
NAND3X1  g211(.A(n262), .B(n116), .C(G9), .Y(n293));
OR2X1    g212(.A(n125), .B(n265), .Y(n294));
NAND2X1  g213(.A(n294), .B(n293), .Y(n295));
NAND3X1  g214(.A(G5), .B(G3), .C(G1), .Y(n296));
NOR3X1   g215(.A(n296), .B(n195), .C(n89), .Y(n297));
AOI22X1  g216(.A0(n295), .A1(n297), .B0(n292), .B1(n291), .Y(n298));
OR4X1    g217(.A(n190), .B(n154), .C(G1), .D(n298), .Y(n299));
OR4X1    g218(.A(n195), .B(n90), .C(n89), .D(n299), .Y(n300));
OR4X1    g219(.A(n271), .B(n259), .C(G2), .D(n272), .Y(n301));
NAND3X1  g220(.A(n224), .B(n101), .C(n87_1), .Y(n302));
AOI21X1  g221(.A0(n301), .A1(n300), .B0(n302), .Y(n303));
NOR2X1   g222(.A(n272), .B(n271), .Y(n304));
NOR4X1   g223(.A(n190), .B(n154), .C(n91), .D(n298), .Y(n305));
NOR2X1   g224(.A(n305), .B(n304), .Y(n306));
NOR4X1   g225(.A(n99), .B(G5), .C(G4), .D(n252), .Y(n307));
NOR2X1   g226(.A(n263), .B(n83), .Y(n308));
NOR3X1   g227(.A(n130), .B(n90), .C(n89), .Y(n309));
OAI21X1  g228(.A0(n308), .A1(n307), .B0(n309), .Y(n310));
NOR2X1   g229(.A(n310), .B(n306), .Y(n311));
NOR4X1   g230(.A(n195), .B(n100), .C(n87_1), .D(n288), .Y(n312));
NOR2X1   g231(.A(n135), .B(n249), .Y(n313));
OAI21X1  g232(.A0(n313), .A1(n312), .B0(n90), .Y(n314));
NOR4X1   g233(.A(n272), .B(n271), .C(G2), .D(n314), .Y(n315));
NOR3X1   g234(.A(n145), .B(G43), .C(n154), .Y(n316));
NOR4X1   g235(.A(n315), .B(n311), .C(n303), .D(n316), .Y(n317));
OAI22X1  g236(.A0(n282), .A1(n120), .B0(G12), .B1(n317), .Y(G532));
NOR4X1   g237(.A(G8), .B(G7), .C(G5), .D(n116), .Y(n319));
NAND4X1  g238(.A(n104), .B(G6), .C(n90), .D(n319), .Y(n320));
NAND2X1  g239(.A(G37), .B(G8), .Y(n321));
OR4X1    g240(.A(n92_1), .B(G10), .C(n101), .D(n321), .Y(n322));
NAND3X1  g241(.A(G11), .B(n83), .C(n85), .Y(n323));
AOI21X1  g242(.A0(n322), .A1(n320), .B0(n323), .Y(n324));
AOI21X1  g243(.A0(n266), .A1(G0), .B0(n324), .Y(n325));
NAND2X1  g244(.A(G2), .B(G1), .Y(n326));
NOR2X1   g245(.A(n326), .B(n325), .Y(n327));
INVX1    g246(.A(n327), .Y(n328));
NOR2X1   g247(.A(G13), .B(n82_1), .Y(n329));
OAI21X1  g248(.A0(n119), .A1(n97_1), .B0(n329), .Y(n330));
NOR4X1   g249(.A(n328), .B(n296), .C(n100), .D(n330), .Y(n331));
AND2X1   g250(.A(G38), .B(G37), .Y(n332));
NAND3X1  g251(.A(n257), .B(n87_1), .C(n83), .Y(n333));
NAND3X1  g252(.A(n116), .B(n104), .C(G7), .Y(n334));
NAND3X1  g253(.A(n116), .B(G9), .C(n101), .Y(n335));
AOI21X1  g254(.A0(n335), .A1(n334), .B0(n100), .Y(n336));
NAND2X1  g255(.A(n336), .B(n84), .Y(n337));
OAI22X1  g256(.A0(n333), .A1(n306), .B0(n299), .B1(n337), .Y(n338));
NOR3X1   g257(.A(G12), .B(n130), .C(n90), .Y(n339));
AOI22X1  g258(.A0(n338), .A1(n339), .B0(n332), .B1(n331), .Y(n340));
NAND2X1  g259(.A(G11), .B(G2), .Y(n341));
NOR3X1   g260(.A(n259), .B(n99), .C(G5), .Y(n342));
NOR2X1   g261(.A(G44), .B(G3), .Y(n343));
AOI21X1  g262(.A0(n336), .A1(n342), .B0(n343), .Y(n344));
OAI22X1  g263(.A0(n341), .A1(n340), .B0(n273), .B1(n344), .Y(G535));
NAND4X1  g264(.A(n87_1), .B(n83), .C(G3), .D(G6), .Y(n346));
NAND4X1  g265(.A(G10), .B(G9), .C(G7), .D(n134), .Y(n347));
OAI22X1  g266(.A0(n346), .A1(n334), .B0(n92_1), .B1(n347), .Y(n348));
NAND2X1  g267(.A(n348), .B(G8), .Y(n349));
OR4X1    g268(.A(n195), .B(G5), .C(n90), .D(n252), .Y(n350));
OAI22X1  g269(.A0(n349), .A1(n306), .B0(n299), .B1(n350), .Y(n351));
NAND3X1  g270(.A(G38), .B(n104), .C(G6), .Y(n352));
OAI21X1  g271(.A0(n347), .A1(n85), .B0(n352), .Y(n353));
AOI22X1  g272(.A0(n351), .A1(n82_1), .B0(n331), .B1(n353), .Y(n354));
OR2X1    g273(.A(G8), .B(G7), .Y(n355));
OR4X1    g274(.A(G6), .B(G5), .C(n83), .D(n125), .Y(n356));
OR4X1    g275(.A(G11), .B(G10), .C(G5), .D(n135), .Y(n357));
NAND4X1  g276(.A(n124), .B(G10), .C(G5), .D(n134), .Y(n358));
AND2X1   g277(.A(n358), .B(n357), .Y(n359));
OAI22X1  g278(.A0(n356), .A1(n265), .B0(n355), .B1(n359), .Y(n360));
NOR4X1   g279(.A(n252), .B(n99), .C(G5), .D(n259), .Y(n361));
AOI21X1  g280(.A0(n360), .A1(n90), .B0(n361), .Y(n362));
OAI22X1  g281(.A0(n354), .A1(n341), .B0(n273), .B1(n362), .Y(G537));
AND2X1   g282(.A(n155), .B(n145), .Y(n364));
NOR2X1   g283(.A(n272), .B(G12), .Y(n365));
AOI22X1  g284(.A0(n364), .A1(n298), .B0(n271), .B1(n365), .Y(n366));
OAI21X1  g285(.A0(n330), .A1(n327), .B0(n366), .Y(G539));
MX2X1    g286(.A(G5), .B(G3), .S0(G4), .Y(n368));
AOI22X1  g287(.A0(n140), .A1(n368), .B0(n188), .B1(n194), .Y(n57));
OAI21X1  g288(.A0(n99), .A1(G9), .B0(n116), .Y(n62));
OAI22X1  g289(.A0(n99), .A1(G7), .B0(n116), .B1(n124), .Y(n67));
NAND2X1  g290(.A(n259), .B(n164), .Y(n372));
AOI21X1  g291(.A0(n139), .A1(n188), .B0(n152), .Y(n373));
NAND2X1  g292(.A(n373), .B(n372), .Y(n72));
NOR3X1   g293(.A(n161), .B(n160), .C(G12), .Y(n375));
NOR3X1   g294(.A(G4), .B(n91), .C(n85), .Y(n376));
AOI22X1  g295(.A0(n375), .A1(n152), .B0(n181), .B1(n376), .Y(n77));
MX2X1    g296(.A(n160), .B(n189), .S0(G13), .Y(n378));
NOR3X1   g297(.A(n378), .B(n161), .C(G12), .Y(n82));
OR2X1    g298(.A(G8), .B(G6), .Y(n380));
OAI22X1  g299(.A0(n252), .A1(n130), .B0(n334), .B1(n380), .Y(n87));
OR4X1    g300(.A(G10), .B(G8), .C(G7), .D(G11), .Y(n382));
AOI21X1  g301(.A0(n382), .A1(n294), .B0(G5), .Y(n92));
XOR2X1   g302(.A(G9), .B(G6), .Y(n97));
NOR4X1   g303(.A(n101), .B(G4), .C(G0), .D(G10), .Y(n102));
XOR2X1   g304(.A(n92_1), .B(n89), .Y(n107));
AND2X1   g305(.A(G9), .B(G6), .Y(n387));
AOI22X1  g306(.A0(G30), .A1(n130), .B0(n99), .B1(n387), .Y(n388));
NAND2X1  g307(.A(G31), .B(G6), .Y(n389));
OAI21X1  g308(.A0(n388), .A1(n101), .B0(n389), .Y(n390));
AOI22X1  g309(.A0(n286), .A1(G6), .B0(G8), .B1(n390), .Y(n112));
OR2X1    g310(.A(n387), .B(n125), .Y(n392));
NAND3X1  g311(.A(n223), .B(n105), .C(G34), .Y(n393));
OAI21X1  g312(.A0(n392), .A1(n120), .B0(n393), .Y(n394));
AOI21X1  g313(.A0(n216), .A1(n214), .B0(n394), .Y(n117));
NOR4X1   g314(.A(n99), .B(n104), .C(n130), .D(n218), .Y(n396));
NAND3X1  g315(.A(n127_1), .B(G7), .C(n130), .Y(n397));
AOI22X1  g316(.A0(n100), .A1(G7), .B0(G6), .B1(n105), .Y(n398));
OAI21X1  g317(.A0(n398), .A1(G9), .B0(n397), .Y(n399));
AOI21X1  g318(.A0(n399), .A1(G11), .B0(n396), .Y(n122));
NAND3X1  g319(.A(n130), .B(G4), .C(G2), .Y(n401));
AOI22X1  g320(.A0(n84), .A1(G6), .B0(G5), .B1(n195), .Y(n402));
NAND2X1  g321(.A(n402), .B(n401), .Y(n403));
OAI22X1  g322(.A0(n141_1), .A1(n90), .B0(n91), .B1(n202), .Y(n404));
AOI21X1  g323(.A0(n403), .A1(n245), .B0(n404), .Y(n127));
NOR4X1   g324(.A(n125), .B(n265), .C(G5), .D(n135), .Y(n406));
NAND4X1  g325(.A(n104), .B(n130), .C(n87_1), .D(n112_1), .Y(n407));
AOI21X1  g326(.A0(n407), .A1(n358), .B0(n355), .Y(n408));
NOR2X1   g327(.A(n408), .B(n406), .Y(n132));
NOR3X1   g328(.A(n298), .B(n156), .C(n190), .Y(n410));
AOI21X1  g329(.A0(n304), .A1(n82_1), .B0(n410), .Y(n411));
OAI21X1  g330(.A0(n330), .A1(n328), .B0(n411), .Y(G45));
NOR4X1   g331(.A(n83), .B(n90), .C(G2), .D(G5), .Y(n413));
NOR2X1   g332(.A(n413), .B(n85), .Y(n414));
OAI21X1  g333(.A0(n94), .A1(n84), .B0(n414), .Y(n415));
OAI21X1  g334(.A0(n84), .A1(n85), .B0(G1), .Y(n416));
NOR2X1   g335(.A(n92_1), .B(n83), .Y(n417));
NAND2X1  g336(.A(n90), .B(G0), .Y(n418));
NAND3X1  g337(.A(n87_1), .B(G3), .C(n91), .Y(n419));
OAI21X1  g338(.A0(n418), .A1(n84), .B0(n419), .Y(n420));
AOI21X1  g339(.A0(n417), .A1(n416), .B0(n420), .Y(n421));
NAND2X1  g340(.A(n93), .B(G2), .Y(n422));
AOI22X1  g341(.A0(n116), .A1(n109), .B0(n101), .B1(n130), .Y(n423));
OAI21X1  g342(.A0(n422), .A1(n421), .B0(n423), .Y(n424));
AOI21X1  g343(.A0(n415), .A1(n91), .B0(n424), .Y(n141));
endmodule
