// Benchmark "top" written by ABC on Mon Sep 21 04:00:31 2020

module top ( 
    \priority[0] , \priority[1] , \priority[2] , \priority[3] ,
    \priority[4] , \priority[5] , \priority[6] , \priority[7] ,
    \priority[8] , \priority[9] , \priority[10] , \priority[11] ,
    \priority[12] , \priority[13] , \priority[14] , \priority[15] ,
    \priority[16] , \priority[17] , \priority[18] , \priority[19] ,
    \priority[20] , \priority[21] , \priority[22] , \priority[23] ,
    \priority[24] , \priority[25] , \priority[26] , \priority[27] ,
    \priority[28] , \priority[29] , \priority[30] , \priority[31] ,
    \priority[32] , \priority[33] , \priority[34] , \priority[35] ,
    \priority[36] , \priority[37] , \priority[38] , \priority[39] ,
    \priority[40] , \priority[41] , \priority[42] , \priority[43] ,
    \priority[44] , \priority[45] , \priority[46] , \priority[47] ,
    \priority[48] , \priority[49] , \priority[50] , \priority[51] ,
    \priority[52] , \priority[53] , \priority[54] , \priority[55] ,
    \priority[56] , \priority[57] , \priority[58] , \priority[59] ,
    \priority[60] , \priority[61] , \priority[62] , \priority[63] ,
    \priority[64] , \priority[65] , \priority[66] , \priority[67] ,
    \priority[68] , \priority[69] , \priority[70] , \priority[71] ,
    \priority[72] , \priority[73] , \priority[74] , \priority[75] ,
    \priority[76] , \priority[77] , \priority[78] , \priority[79] ,
    \priority[80] , \priority[81] , \priority[82] , \priority[83] ,
    \priority[84] , \priority[85] , \priority[86] , \priority[87] ,
    \priority[88] , \priority[89] , \priority[90] , \priority[91] ,
    \priority[92] , \priority[93] , \priority[94] , \priority[95] ,
    \priority[96] , \priority[97] , \priority[98] , \priority[99] ,
    \priority[100] , \priority[101] , \priority[102] , \priority[103] ,
    \priority[104] , \priority[105] , \priority[106] , \priority[107] ,
    \priority[108] , \priority[109] , \priority[110] , \priority[111] ,
    \priority[112] , \priority[113] , \priority[114] , \priority[115] ,
    \priority[116] , \priority[117] , \priority[118] , \priority[119] ,
    \priority[120] , \priority[121] , \priority[122] , \priority[123] ,
    \priority[124] , \priority[125] , \priority[126] , \priority[127] ,
    \req[0] , \req[1] , \req[2] , \req[3] , \req[4] , \req[5] , \req[6] ,
    \req[7] , \req[8] , \req[9] , \req[10] , \req[11] , \req[12] ,
    \req[13] , \req[14] , \req[15] , \req[16] , \req[17] , \req[18] ,
    \req[19] , \req[20] , \req[21] , \req[22] , \req[23] , \req[24] ,
    \req[25] , \req[26] , \req[27] , \req[28] , \req[29] , \req[30] ,
    \req[31] , \req[32] , \req[33] , \req[34] , \req[35] , \req[36] ,
    \req[37] , \req[38] , \req[39] , \req[40] , \req[41] , \req[42] ,
    \req[43] , \req[44] , \req[45] , \req[46] , \req[47] , \req[48] ,
    \req[49] , \req[50] , \req[51] , \req[52] , \req[53] , \req[54] ,
    \req[55] , \req[56] , \req[57] , \req[58] , \req[59] , \req[60] ,
    \req[61] , \req[62] , \req[63] , \req[64] , \req[65] , \req[66] ,
    \req[67] , \req[68] , \req[69] , \req[70] , \req[71] , \req[72] ,
    \req[73] , \req[74] , \req[75] , \req[76] , \req[77] , \req[78] ,
    \req[79] , \req[80] , \req[81] , \req[82] , \req[83] , \req[84] ,
    \req[85] , \req[86] , \req[87] , \req[88] , \req[89] , \req[90] ,
    \req[91] , \req[92] , \req[93] , \req[94] , \req[95] , \req[96] ,
    \req[97] , \req[98] , \req[99] , \req[100] , \req[101] , \req[102] ,
    \req[103] , \req[104] , \req[105] , \req[106] , \req[107] , \req[108] ,
    \req[109] , \req[110] , \req[111] , \req[112] , \req[113] , \req[114] ,
    \req[115] , \req[116] , \req[117] , \req[118] , \req[119] , \req[120] ,
    \req[121] , \req[122] , \req[123] , \req[124] , \req[125] , \req[126] ,
    \req[127] ,
    \grant[0] , \grant[1] , \grant[2] , \grant[3] , \grant[4] , \grant[5] ,
    \grant[6] , \grant[7] , \grant[8] , \grant[9] , \grant[10] ,
    \grant[11] , \grant[12] , \grant[13] , \grant[14] , \grant[15] ,
    \grant[16] , \grant[17] , \grant[18] , \grant[19] , \grant[20] ,
    \grant[21] , \grant[22] , \grant[23] , \grant[24] , \grant[25] ,
    \grant[26] , \grant[27] , \grant[28] , \grant[29] , \grant[30] ,
    \grant[31] , \grant[32] , \grant[33] , \grant[34] , \grant[35] ,
    \grant[36] , \grant[37] , \grant[38] , \grant[39] , \grant[40] ,
    \grant[41] , \grant[42] , \grant[43] , \grant[44] , \grant[45] ,
    \grant[46] , \grant[47] , \grant[48] , \grant[49] , \grant[50] ,
    \grant[51] , \grant[52] , \grant[53] , \grant[54] , \grant[55] ,
    \grant[56] , \grant[57] , \grant[58] , \grant[59] , \grant[60] ,
    \grant[61] , \grant[62] , \grant[63] , \grant[64] , \grant[65] ,
    \grant[66] , \grant[67] , \grant[68] , \grant[69] , \grant[70] ,
    \grant[71] , \grant[72] , \grant[73] , \grant[74] , \grant[75] ,
    \grant[76] , \grant[77] , \grant[78] , \grant[79] , \grant[80] ,
    \grant[81] , \grant[82] , \grant[83] , \grant[84] , \grant[85] ,
    \grant[86] , \grant[87] , \grant[88] , \grant[89] , \grant[90] ,
    \grant[91] , \grant[92] , \grant[93] , \grant[94] , \grant[95] ,
    \grant[96] , \grant[97] , \grant[98] , \grant[99] , \grant[100] ,
    \grant[101] , \grant[102] , \grant[103] , \grant[104] , \grant[105] ,
    \grant[106] , \grant[107] , \grant[108] , \grant[109] , \grant[110] ,
    \grant[111] , \grant[112] , \grant[113] , \grant[114] , \grant[115] ,
    \grant[116] , \grant[117] , \grant[118] , \grant[119] , \grant[120] ,
    \grant[121] , \grant[122] , \grant[123] , \grant[124] , \grant[125] ,
    \grant[126] , \grant[127] , anyGrant  );
  input  \priority[0] , \priority[1] , \priority[2] , \priority[3] ,
    \priority[4] , \priority[5] , \priority[6] , \priority[7] ,
    \priority[8] , \priority[9] , \priority[10] , \priority[11] ,
    \priority[12] , \priority[13] , \priority[14] , \priority[15] ,
    \priority[16] , \priority[17] , \priority[18] , \priority[19] ,
    \priority[20] , \priority[21] , \priority[22] , \priority[23] ,
    \priority[24] , \priority[25] , \priority[26] , \priority[27] ,
    \priority[28] , \priority[29] , \priority[30] , \priority[31] ,
    \priority[32] , \priority[33] , \priority[34] , \priority[35] ,
    \priority[36] , \priority[37] , \priority[38] , \priority[39] ,
    \priority[40] , \priority[41] , \priority[42] , \priority[43] ,
    \priority[44] , \priority[45] , \priority[46] , \priority[47] ,
    \priority[48] , \priority[49] , \priority[50] , \priority[51] ,
    \priority[52] , \priority[53] , \priority[54] , \priority[55] ,
    \priority[56] , \priority[57] , \priority[58] , \priority[59] ,
    \priority[60] , \priority[61] , \priority[62] , \priority[63] ,
    \priority[64] , \priority[65] , \priority[66] , \priority[67] ,
    \priority[68] , \priority[69] , \priority[70] , \priority[71] ,
    \priority[72] , \priority[73] , \priority[74] , \priority[75] ,
    \priority[76] , \priority[77] , \priority[78] , \priority[79] ,
    \priority[80] , \priority[81] , \priority[82] , \priority[83] ,
    \priority[84] , \priority[85] , \priority[86] , \priority[87] ,
    \priority[88] , \priority[89] , \priority[90] , \priority[91] ,
    \priority[92] , \priority[93] , \priority[94] , \priority[95] ,
    \priority[96] , \priority[97] , \priority[98] , \priority[99] ,
    \priority[100] , \priority[101] , \priority[102] , \priority[103] ,
    \priority[104] , \priority[105] , \priority[106] , \priority[107] ,
    \priority[108] , \priority[109] , \priority[110] , \priority[111] ,
    \priority[112] , \priority[113] , \priority[114] , \priority[115] ,
    \priority[116] , \priority[117] , \priority[118] , \priority[119] ,
    \priority[120] , \priority[121] , \priority[122] , \priority[123] ,
    \priority[124] , \priority[125] , \priority[126] , \priority[127] ,
    \req[0] , \req[1] , \req[2] , \req[3] , \req[4] , \req[5] , \req[6] ,
    \req[7] , \req[8] , \req[9] , \req[10] , \req[11] , \req[12] ,
    \req[13] , \req[14] , \req[15] , \req[16] , \req[17] , \req[18] ,
    \req[19] , \req[20] , \req[21] , \req[22] , \req[23] , \req[24] ,
    \req[25] , \req[26] , \req[27] , \req[28] , \req[29] , \req[30] ,
    \req[31] , \req[32] , \req[33] , \req[34] , \req[35] , \req[36] ,
    \req[37] , \req[38] , \req[39] , \req[40] , \req[41] , \req[42] ,
    \req[43] , \req[44] , \req[45] , \req[46] , \req[47] , \req[48] ,
    \req[49] , \req[50] , \req[51] , \req[52] , \req[53] , \req[54] ,
    \req[55] , \req[56] , \req[57] , \req[58] , \req[59] , \req[60] ,
    \req[61] , \req[62] , \req[63] , \req[64] , \req[65] , \req[66] ,
    \req[67] , \req[68] , \req[69] , \req[70] , \req[71] , \req[72] ,
    \req[73] , \req[74] , \req[75] , \req[76] , \req[77] , \req[78] ,
    \req[79] , \req[80] , \req[81] , \req[82] , \req[83] , \req[84] ,
    \req[85] , \req[86] , \req[87] , \req[88] , \req[89] , \req[90] ,
    \req[91] , \req[92] , \req[93] , \req[94] , \req[95] , \req[96] ,
    \req[97] , \req[98] , \req[99] , \req[100] , \req[101] , \req[102] ,
    \req[103] , \req[104] , \req[105] , \req[106] , \req[107] , \req[108] ,
    \req[109] , \req[110] , \req[111] , \req[112] , \req[113] , \req[114] ,
    \req[115] , \req[116] , \req[117] , \req[118] , \req[119] , \req[120] ,
    \req[121] , \req[122] , \req[123] , \req[124] , \req[125] , \req[126] ,
    \req[127] ;
  output \grant[0] , \grant[1] , \grant[2] , \grant[3] , \grant[4] ,
    \grant[5] , \grant[6] , \grant[7] , \grant[8] , \grant[9] ,
    \grant[10] , \grant[11] , \grant[12] , \grant[13] , \grant[14] ,
    \grant[15] , \grant[16] , \grant[17] , \grant[18] , \grant[19] ,
    \grant[20] , \grant[21] , \grant[22] , \grant[23] , \grant[24] ,
    \grant[25] , \grant[26] , \grant[27] , \grant[28] , \grant[29] ,
    \grant[30] , \grant[31] , \grant[32] , \grant[33] , \grant[34] ,
    \grant[35] , \grant[36] , \grant[37] , \grant[38] , \grant[39] ,
    \grant[40] , \grant[41] , \grant[42] , \grant[43] , \grant[44] ,
    \grant[45] , \grant[46] , \grant[47] , \grant[48] , \grant[49] ,
    \grant[50] , \grant[51] , \grant[52] , \grant[53] , \grant[54] ,
    \grant[55] , \grant[56] , \grant[57] , \grant[58] , \grant[59] ,
    \grant[60] , \grant[61] , \grant[62] , \grant[63] , \grant[64] ,
    \grant[65] , \grant[66] , \grant[67] , \grant[68] , \grant[69] ,
    \grant[70] , \grant[71] , \grant[72] , \grant[73] , \grant[74] ,
    \grant[75] , \grant[76] , \grant[77] , \grant[78] , \grant[79] ,
    \grant[80] , \grant[81] , \grant[82] , \grant[83] , \grant[84] ,
    \grant[85] , \grant[86] , \grant[87] , \grant[88] , \grant[89] ,
    \grant[90] , \grant[91] , \grant[92] , \grant[93] , \grant[94] ,
    \grant[95] , \grant[96] , \grant[97] , \grant[98] , \grant[99] ,
    \grant[100] , \grant[101] , \grant[102] , \grant[103] , \grant[104] ,
    \grant[105] , \grant[106] , \grant[107] , \grant[108] , \grant[109] ,
    \grant[110] , \grant[111] , \grant[112] , \grant[113] , \grant[114] ,
    \grant[115] , \grant[116] , \grant[117] , \grant[118] , \grant[119] ,
    \grant[120] , \grant[121] , \grant[122] , \grant[123] , \grant[124] ,
    \grant[125] , \grant[126] , \grant[127] , anyGrant;
  wire new_n386_, new_n387_, new_n388_, new_n389_, new_n390_, new_n391_,
    new_n392_, new_n393_, new_n394_, new_n395_, new_n396_, new_n397_,
    new_n398_, new_n399_, new_n400_, new_n401_, new_n402_, new_n403_,
    new_n404_, new_n405_, new_n406_, new_n407_, new_n408_, new_n409_,
    new_n410_, new_n411_, new_n412_, new_n413_, new_n414_, new_n415_,
    new_n416_, new_n417_, new_n418_, new_n419_, new_n420_, new_n421_,
    new_n422_, new_n423_, new_n424_, new_n425_, new_n426_, new_n427_,
    new_n428_, new_n429_, new_n430_, new_n431_, new_n432_, new_n433_,
    new_n434_, new_n435_, new_n436_, new_n437_, new_n438_, new_n439_,
    new_n440_, new_n441_, new_n442_, new_n443_, new_n444_, new_n445_,
    new_n446_, new_n447_, new_n448_, new_n449_, new_n450_, new_n451_,
    new_n452_, new_n453_, new_n454_, new_n455_, new_n456_, new_n457_,
    new_n458_, new_n459_, new_n460_, new_n461_, new_n462_, new_n463_,
    new_n464_, new_n465_, new_n466_, new_n467_, new_n468_, new_n469_,
    new_n470_, new_n471_, new_n472_, new_n473_, new_n474_, new_n475_,
    new_n476_, new_n477_, new_n478_, new_n479_, new_n480_, new_n481_,
    new_n482_, new_n483_, new_n484_, new_n485_, new_n486_, new_n487_,
    new_n488_, new_n489_, new_n490_, new_n491_, new_n492_, new_n493_,
    new_n494_, new_n495_, new_n496_, new_n497_, new_n498_, new_n499_,
    new_n500_, new_n501_, new_n502_, new_n503_, new_n504_, new_n505_,
    new_n506_, new_n507_, new_n508_, new_n509_, new_n510_, new_n511_,
    new_n512_, new_n513_, new_n514_, new_n515_, new_n516_, new_n517_,
    new_n518_, new_n519_, new_n520_, new_n521_, new_n522_, new_n523_,
    new_n524_, new_n525_, new_n526_, new_n527_, new_n528_, new_n529_,
    new_n530_, new_n531_, new_n532_, new_n533_, new_n534_, new_n535_,
    new_n536_, new_n537_, new_n538_, new_n539_, new_n540_, new_n541_,
    new_n542_, new_n543_, new_n544_, new_n545_, new_n546_, new_n547_,
    new_n548_, new_n549_, new_n550_, new_n551_, new_n552_, new_n553_,
    new_n554_, new_n555_, new_n556_, new_n557_, new_n558_, new_n559_,
    new_n560_, new_n561_, new_n562_, new_n563_, new_n564_, new_n565_,
    new_n566_, new_n567_, new_n568_, new_n569_, new_n570_, new_n571_,
    new_n572_, new_n573_, new_n574_, new_n575_, new_n576_, new_n577_,
    new_n578_, new_n579_, new_n580_, new_n581_, new_n582_, new_n583_,
    new_n584_, new_n585_, new_n586_, new_n587_, new_n588_, new_n589_,
    new_n590_, new_n591_, new_n592_, new_n593_, new_n594_, new_n595_,
    new_n596_, new_n597_, new_n598_, new_n599_, new_n600_, new_n601_,
    new_n602_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n759_, new_n760_, new_n761_, new_n762_, new_n763_, new_n764_,
    new_n765_, new_n766_, new_n767_, new_n768_, new_n769_, new_n770_,
    new_n771_, new_n772_, new_n773_, new_n774_, new_n775_, new_n776_,
    new_n777_, new_n778_, new_n779_, new_n780_, new_n781_, new_n782_,
    new_n783_, new_n784_, new_n785_, new_n786_, new_n787_, new_n788_,
    new_n789_, new_n790_, new_n791_, new_n792_, new_n793_, new_n794_,
    new_n795_, new_n796_, new_n797_, new_n798_, new_n799_, new_n800_,
    new_n801_, new_n802_, new_n803_, new_n804_, new_n805_, new_n806_,
    new_n807_, new_n808_, new_n809_, new_n810_, new_n811_, new_n812_,
    new_n813_, new_n814_, new_n815_, new_n816_, new_n817_, new_n818_,
    new_n819_, new_n820_, new_n821_, new_n822_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n846_, new_n847_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n870_, new_n871_, new_n872_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n877_, new_n878_,
    new_n879_, new_n880_, new_n881_, new_n882_, new_n883_, new_n884_,
    new_n885_, new_n886_, new_n887_, new_n888_, new_n889_, new_n890_,
    new_n891_, new_n892_, new_n893_, new_n894_, new_n895_, new_n896_,
    new_n897_, new_n898_, new_n899_, new_n900_, new_n901_, new_n902_,
    new_n903_, new_n904_, new_n905_, new_n906_, new_n907_, new_n908_,
    new_n909_, new_n910_, new_n911_, new_n912_, new_n913_, new_n914_,
    new_n915_, new_n916_, new_n917_, new_n918_, new_n919_, new_n920_,
    new_n921_, new_n922_, new_n923_, new_n924_, new_n925_, new_n926_,
    new_n927_, new_n928_, new_n929_, new_n930_, new_n931_, new_n932_,
    new_n933_, new_n934_, new_n935_, new_n936_, new_n937_, new_n938_,
    new_n939_, new_n940_, new_n941_, new_n942_, new_n943_, new_n944_,
    new_n945_, new_n946_, new_n947_, new_n948_, new_n949_, new_n950_,
    new_n951_, new_n952_, new_n953_, new_n954_, new_n955_, new_n956_,
    new_n957_, new_n958_, new_n959_, new_n960_, new_n961_, new_n962_,
    new_n963_, new_n964_, new_n965_, new_n966_, new_n967_, new_n968_,
    new_n969_, new_n970_, new_n971_, new_n972_, new_n973_, new_n974_,
    new_n975_, new_n976_, new_n977_, new_n978_, new_n979_, new_n980_,
    new_n981_, new_n982_, new_n983_, new_n984_, new_n985_, new_n986_,
    new_n987_, new_n988_, new_n989_, new_n990_, new_n991_, new_n992_,
    new_n993_, new_n994_, new_n995_, new_n996_, new_n997_, new_n998_,
    new_n999_, new_n1000_, new_n1001_, new_n1002_, new_n1003_, new_n1004_,
    new_n1005_, new_n1006_, new_n1007_, new_n1008_, new_n1009_, new_n1010_,
    new_n1011_, new_n1012_, new_n1013_, new_n1014_, new_n1015_, new_n1016_,
    new_n1017_, new_n1018_, new_n1019_, new_n1021_, new_n1022_, new_n1023_,
    new_n1024_, new_n1025_, new_n1026_, new_n1027_, new_n1028_, new_n1029_,
    new_n1030_, new_n1031_, new_n1032_, new_n1033_, new_n1034_, new_n1035_,
    new_n1036_, new_n1037_, new_n1038_, new_n1039_, new_n1040_, new_n1041_,
    new_n1042_, new_n1043_, new_n1044_, new_n1045_, new_n1046_, new_n1047_,
    new_n1048_, new_n1049_, new_n1050_, new_n1051_, new_n1052_, new_n1053_,
    new_n1054_, new_n1055_, new_n1056_, new_n1057_, new_n1058_, new_n1059_,
    new_n1060_, new_n1061_, new_n1062_, new_n1063_, new_n1064_, new_n1065_,
    new_n1066_, new_n1067_, new_n1068_, new_n1069_, new_n1070_, new_n1071_,
    new_n1072_, new_n1073_, new_n1074_, new_n1075_, new_n1076_, new_n1077_,
    new_n1078_, new_n1079_, new_n1080_, new_n1081_, new_n1082_, new_n1083_,
    new_n1084_, new_n1085_, new_n1086_, new_n1087_, new_n1088_, new_n1089_,
    new_n1090_, new_n1091_, new_n1092_, new_n1093_, new_n1094_, new_n1095_,
    new_n1096_, new_n1097_, new_n1098_, new_n1099_, new_n1100_, new_n1101_,
    new_n1102_, new_n1103_, new_n1104_, new_n1105_, new_n1106_, new_n1107_,
    new_n1108_, new_n1109_, new_n1110_, new_n1111_, new_n1112_, new_n1113_,
    new_n1114_, new_n1115_, new_n1116_, new_n1117_, new_n1118_, new_n1119_,
    new_n1120_, new_n1121_, new_n1122_, new_n1123_, new_n1124_, new_n1125_,
    new_n1126_, new_n1127_, new_n1128_, new_n1129_, new_n1130_, new_n1131_,
    new_n1132_, new_n1133_, new_n1134_, new_n1135_, new_n1136_, new_n1137_,
    new_n1138_, new_n1139_, new_n1140_, new_n1141_, new_n1142_, new_n1143_,
    new_n1144_, new_n1145_, new_n1146_, new_n1147_, new_n1148_, new_n1149_,
    new_n1150_, new_n1151_, new_n1152_, new_n1153_, new_n1154_, new_n1155_,
    new_n1156_, new_n1157_, new_n1158_, new_n1159_, new_n1160_, new_n1161_,
    new_n1162_, new_n1163_, new_n1164_, new_n1165_, new_n1166_, new_n1167_,
    new_n1168_, new_n1169_, new_n1170_, new_n1171_, new_n1172_, new_n1173_,
    new_n1174_, new_n1175_, new_n1176_, new_n1177_, new_n1178_, new_n1179_,
    new_n1180_, new_n1181_, new_n1182_, new_n1183_, new_n1184_, new_n1185_,
    new_n1186_, new_n1187_, new_n1188_, new_n1189_, new_n1190_, new_n1191_,
    new_n1192_, new_n1193_, new_n1194_, new_n1195_, new_n1196_, new_n1197_,
    new_n1198_, new_n1199_, new_n1200_, new_n1201_, new_n1202_, new_n1203_,
    new_n1204_, new_n1205_, new_n1206_, new_n1207_, new_n1208_, new_n1209_,
    new_n1210_, new_n1211_, new_n1212_, new_n1213_, new_n1214_, new_n1215_,
    new_n1216_, new_n1217_, new_n1218_, new_n1219_, new_n1220_, new_n1221_,
    new_n1222_, new_n1223_, new_n1224_, new_n1225_, new_n1226_, new_n1227_,
    new_n1228_, new_n1229_, new_n1230_, new_n1231_, new_n1232_, new_n1233_,
    new_n1234_, new_n1235_, new_n1236_, new_n1237_, new_n1238_, new_n1239_,
    new_n1240_, new_n1241_, new_n1242_, new_n1243_, new_n1244_, new_n1245_,
    new_n1246_, new_n1247_, new_n1248_, new_n1249_, new_n1250_, new_n1251_,
    new_n1252_, new_n1253_, new_n1254_, new_n1255_, new_n1256_, new_n1257_,
    new_n1258_, new_n1259_, new_n1260_, new_n1261_, new_n1262_, new_n1263_,
    new_n1264_, new_n1265_, new_n1266_, new_n1267_, new_n1268_, new_n1269_,
    new_n1270_, new_n1271_, new_n1272_, new_n1273_, new_n1274_, new_n1275_,
    new_n1276_, new_n1277_, new_n1278_, new_n1279_, new_n1280_, new_n1281_,
    new_n1282_, new_n1283_, new_n1284_, new_n1285_, new_n1286_, new_n1287_,
    new_n1288_, new_n1289_, new_n1290_, new_n1291_, new_n1292_, new_n1293_,
    new_n1294_, new_n1295_, new_n1296_, new_n1297_, new_n1298_, new_n1299_,
    new_n1300_, new_n1301_, new_n1302_, new_n1303_, new_n1304_, new_n1305_,
    new_n1306_, new_n1307_, new_n1308_, new_n1309_, new_n1310_, new_n1311_,
    new_n1312_, new_n1313_, new_n1314_, new_n1315_, new_n1316_, new_n1317_,
    new_n1318_, new_n1319_, new_n1320_, new_n1321_, new_n1322_, new_n1323_,
    new_n1324_, new_n1325_, new_n1326_, new_n1327_, new_n1328_, new_n1329_,
    new_n1330_, new_n1331_, new_n1332_, new_n1333_, new_n1335_, new_n1336_,
    new_n1337_, new_n1338_, new_n1339_, new_n1340_, new_n1341_, new_n1342_,
    new_n1343_, new_n1344_, new_n1345_, new_n1346_, new_n1347_, new_n1348_,
    new_n1349_, new_n1350_, new_n1351_, new_n1352_, new_n1353_, new_n1354_,
    new_n1355_, new_n1356_, new_n1357_, new_n1358_, new_n1359_, new_n1360_,
    new_n1361_, new_n1362_, new_n1363_, new_n1364_, new_n1365_, new_n1366_,
    new_n1367_, new_n1368_, new_n1369_, new_n1370_, new_n1371_, new_n1372_,
    new_n1373_, new_n1374_, new_n1375_, new_n1376_, new_n1377_, new_n1378_,
    new_n1379_, new_n1380_, new_n1381_, new_n1382_, new_n1383_, new_n1384_,
    new_n1385_, new_n1386_, new_n1387_, new_n1388_, new_n1389_, new_n1390_,
    new_n1391_, new_n1392_, new_n1393_, new_n1394_, new_n1395_, new_n1396_,
    new_n1397_, new_n1398_, new_n1399_, new_n1400_, new_n1401_, new_n1402_,
    new_n1403_, new_n1404_, new_n1405_, new_n1406_, new_n1407_, new_n1408_,
    new_n1409_, new_n1410_, new_n1411_, new_n1412_, new_n1413_, new_n1414_,
    new_n1415_, new_n1416_, new_n1417_, new_n1418_, new_n1419_, new_n1420_,
    new_n1421_, new_n1422_, new_n1423_, new_n1424_, new_n1425_, new_n1426_,
    new_n1427_, new_n1428_, new_n1429_, new_n1430_, new_n1431_, new_n1432_,
    new_n1433_, new_n1434_, new_n1435_, new_n1436_, new_n1437_, new_n1438_,
    new_n1439_, new_n1440_, new_n1441_, new_n1442_, new_n1444_, new_n1445_,
    new_n1446_, new_n1447_, new_n1448_, new_n1449_, new_n1450_, new_n1451_,
    new_n1452_, new_n1453_, new_n1454_, new_n1455_, new_n1456_, new_n1457_,
    new_n1458_, new_n1459_, new_n1460_, new_n1461_, new_n1462_, new_n1463_,
    new_n1464_, new_n1465_, new_n1466_, new_n1467_, new_n1468_, new_n1469_,
    new_n1470_, new_n1471_, new_n1472_, new_n1473_, new_n1474_, new_n1475_,
    new_n1476_, new_n1477_, new_n1478_, new_n1479_, new_n1480_, new_n1481_,
    new_n1482_, new_n1483_, new_n1484_, new_n1485_, new_n1486_, new_n1487_,
    new_n1488_, new_n1489_, new_n1490_, new_n1491_, new_n1492_, new_n1493_,
    new_n1494_, new_n1495_, new_n1496_, new_n1497_, new_n1498_, new_n1499_,
    new_n1500_, new_n1501_, new_n1502_, new_n1503_, new_n1504_, new_n1505_,
    new_n1506_, new_n1507_, new_n1508_, new_n1509_, new_n1510_, new_n1511_,
    new_n1512_, new_n1513_, new_n1514_, new_n1515_, new_n1516_, new_n1517_,
    new_n1518_, new_n1519_, new_n1520_, new_n1521_, new_n1522_, new_n1523_,
    new_n1524_, new_n1525_, new_n1526_, new_n1527_, new_n1528_, new_n1529_,
    new_n1530_, new_n1531_, new_n1532_, new_n1533_, new_n1534_, new_n1535_,
    new_n1536_, new_n1537_, new_n1538_, new_n1539_, new_n1540_, new_n1541_,
    new_n1542_, new_n1543_, new_n1544_, new_n1545_, new_n1546_, new_n1547_,
    new_n1548_, new_n1549_, new_n1550_, new_n1552_, new_n1553_, new_n1554_,
    new_n1555_, new_n1556_, new_n1557_, new_n1558_, new_n1559_, new_n1560_,
    new_n1561_, new_n1562_, new_n1563_, new_n1564_, new_n1565_, new_n1566_,
    new_n1567_, new_n1568_, new_n1569_, new_n1570_, new_n1571_, new_n1572_,
    new_n1573_, new_n1574_, new_n1575_, new_n1576_, new_n1577_, new_n1578_,
    new_n1579_, new_n1580_, new_n1581_, new_n1582_, new_n1583_, new_n1584_,
    new_n1585_, new_n1586_, new_n1587_, new_n1588_, new_n1589_, new_n1590_,
    new_n1591_, new_n1592_, new_n1593_, new_n1594_, new_n1595_, new_n1596_,
    new_n1597_, new_n1598_, new_n1599_, new_n1600_, new_n1601_, new_n1602_,
    new_n1603_, new_n1604_, new_n1605_, new_n1606_, new_n1607_, new_n1608_,
    new_n1609_, new_n1610_, new_n1611_, new_n1612_, new_n1613_, new_n1614_,
    new_n1615_, new_n1616_, new_n1617_, new_n1618_, new_n1619_, new_n1620_,
    new_n1621_, new_n1622_, new_n1623_, new_n1624_, new_n1625_, new_n1626_,
    new_n1627_, new_n1628_, new_n1629_, new_n1630_, new_n1631_, new_n1632_,
    new_n1633_, new_n1634_, new_n1635_, new_n1636_, new_n1637_, new_n1638_,
    new_n1639_, new_n1640_, new_n1641_, new_n1642_, new_n1643_, new_n1644_,
    new_n1645_, new_n1646_, new_n1647_, new_n1648_, new_n1649_, new_n1650_,
    new_n1651_, new_n1652_, new_n1653_, new_n1654_, new_n1655_, new_n1656_,
    new_n1657_, new_n1658_, new_n1660_, new_n1661_, new_n1662_, new_n1663_,
    new_n1664_, new_n1665_, new_n1666_, new_n1667_, new_n1668_, new_n1669_,
    new_n1670_, new_n1671_, new_n1672_, new_n1673_, new_n1674_, new_n1675_,
    new_n1676_, new_n1677_, new_n1678_, new_n1679_, new_n1680_, new_n1681_,
    new_n1682_, new_n1683_, new_n1684_, new_n1685_, new_n1686_, new_n1687_,
    new_n1688_, new_n1689_, new_n1690_, new_n1691_, new_n1692_, new_n1693_,
    new_n1694_, new_n1695_, new_n1696_, new_n1697_, new_n1698_, new_n1699_,
    new_n1700_, new_n1701_, new_n1702_, new_n1703_, new_n1704_, new_n1705_,
    new_n1706_, new_n1707_, new_n1709_, new_n1710_, new_n1711_, new_n1712_,
    new_n1713_, new_n1714_, new_n1715_, new_n1716_, new_n1717_, new_n1718_,
    new_n1719_, new_n1720_, new_n1721_, new_n1722_, new_n1723_, new_n1724_,
    new_n1725_, new_n1726_, new_n1727_, new_n1728_, new_n1729_, new_n1730_,
    new_n1731_, new_n1732_, new_n1733_, new_n1734_, new_n1735_, new_n1736_,
    new_n1737_, new_n1738_, new_n1739_, new_n1740_, new_n1741_, new_n1742_,
    new_n1743_, new_n1744_, new_n1745_, new_n1746_, new_n1747_, new_n1748_,
    new_n1749_, new_n1750_, new_n1751_, new_n1752_, new_n1753_, new_n1754_,
    new_n1755_, new_n1756_, new_n1758_, new_n1759_, new_n1760_, new_n1761_,
    new_n1762_, new_n1763_, new_n1764_, new_n1765_, new_n1766_, new_n1767_,
    new_n1768_, new_n1769_, new_n1770_, new_n1771_, new_n1772_, new_n1773_,
    new_n1774_, new_n1775_, new_n1776_, new_n1777_, new_n1778_, new_n1779_,
    new_n1780_, new_n1781_, new_n1782_, new_n1783_, new_n1784_, new_n1785_,
    new_n1786_, new_n1787_, new_n1788_, new_n1789_, new_n1790_, new_n1791_,
    new_n1792_, new_n1793_, new_n1794_, new_n1795_, new_n1796_, new_n1797_,
    new_n1798_, new_n1799_, new_n1800_, new_n1801_, new_n1803_, new_n1804_,
    new_n1805_, new_n1806_, new_n1807_, new_n1808_, new_n1809_, new_n1810_,
    new_n1811_, new_n1812_, new_n1813_, new_n1814_, new_n1815_, new_n1816_,
    new_n1817_, new_n1818_, new_n1819_, new_n1820_, new_n1821_, new_n1822_,
    new_n1823_, new_n1824_, new_n1825_, new_n1826_, new_n1827_, new_n1828_,
    new_n1829_, new_n1830_, new_n1831_, new_n1832_, new_n1833_, new_n1834_,
    new_n1835_, new_n1836_, new_n1837_, new_n1838_, new_n1839_, new_n1840_,
    new_n1841_, new_n1842_, new_n1843_, new_n1844_, new_n1845_, new_n1846_,
    new_n1848_, new_n1849_, new_n1850_, new_n1851_, new_n1852_, new_n1853_,
    new_n1854_, new_n1855_, new_n1856_, new_n1857_, new_n1858_, new_n1859_,
    new_n1860_, new_n1861_, new_n1862_, new_n1863_, new_n1864_, new_n1865_,
    new_n1866_, new_n1867_, new_n1868_, new_n1869_, new_n1870_, new_n1871_,
    new_n1872_, new_n1873_, new_n1874_, new_n1875_, new_n1876_, new_n1877_,
    new_n1878_, new_n1879_, new_n1880_, new_n1881_, new_n1882_, new_n1883_,
    new_n1884_, new_n1885_, new_n1886_, new_n1887_, new_n1888_, new_n1889_,
    new_n1890_, new_n1891_, new_n1893_, new_n1894_, new_n1895_, new_n1896_,
    new_n1897_, new_n1898_, new_n1899_, new_n1900_, new_n1901_, new_n1902_,
    new_n1903_, new_n1904_, new_n1905_, new_n1906_, new_n1907_, new_n1908_,
    new_n1909_, new_n1910_, new_n1911_, new_n1912_, new_n1913_, new_n1914_,
    new_n1915_, new_n1916_, new_n1917_, new_n1918_, new_n1919_, new_n1920_,
    new_n1921_, new_n1922_, new_n1923_, new_n1924_, new_n1925_, new_n1926_,
    new_n1927_, new_n1928_, new_n1929_, new_n1930_, new_n1931_, new_n1932_,
    new_n1933_, new_n1934_, new_n1935_, new_n1936_, new_n1938_, new_n1939_,
    new_n1940_, new_n1941_, new_n1942_, new_n1943_, new_n1944_, new_n1945_,
    new_n1946_, new_n1947_, new_n1948_, new_n1949_, new_n1950_, new_n1951_,
    new_n1952_, new_n1953_, new_n1954_, new_n1955_, new_n1956_, new_n1957_,
    new_n1958_, new_n1959_, new_n1960_, new_n1961_, new_n1962_, new_n1963_,
    new_n1964_, new_n1965_, new_n1966_, new_n1967_, new_n1968_, new_n1969_,
    new_n1970_, new_n1971_, new_n1972_, new_n1973_, new_n1974_, new_n1975_,
    new_n1976_, new_n1977_, new_n1978_, new_n1979_, new_n1980_, new_n1981_,
    new_n1983_, new_n1984_, new_n1985_, new_n1986_, new_n1987_, new_n1988_,
    new_n1989_, new_n1990_, new_n1991_, new_n1992_, new_n1993_, new_n1994_,
    new_n1995_, new_n1996_, new_n1997_, new_n1998_, new_n1999_, new_n2000_,
    new_n2001_, new_n2002_, new_n2003_, new_n2004_, new_n2005_, new_n2006_,
    new_n2007_, new_n2008_, new_n2009_, new_n2010_, new_n2011_, new_n2012_,
    new_n2013_, new_n2014_, new_n2015_, new_n2016_, new_n2017_, new_n2018_,
    new_n2019_, new_n2020_, new_n2021_, new_n2022_, new_n2023_, new_n2024_,
    new_n2025_, new_n2026_, new_n2028_, new_n2029_, new_n2030_, new_n2031_,
    new_n2032_, new_n2033_, new_n2034_, new_n2035_, new_n2036_, new_n2037_,
    new_n2038_, new_n2039_, new_n2040_, new_n2041_, new_n2042_, new_n2043_,
    new_n2044_, new_n2045_, new_n2046_, new_n2047_, new_n2048_, new_n2049_,
    new_n2050_, new_n2051_, new_n2052_, new_n2053_, new_n2054_, new_n2055_,
    new_n2056_, new_n2057_, new_n2058_, new_n2059_, new_n2060_, new_n2061_,
    new_n2062_, new_n2063_, new_n2064_, new_n2065_, new_n2066_, new_n2067_,
    new_n2068_, new_n2069_, new_n2070_, new_n2072_, new_n2073_, new_n2074_,
    new_n2075_, new_n2076_, new_n2077_, new_n2078_, new_n2079_, new_n2080_,
    new_n2081_, new_n2082_, new_n2083_, new_n2084_, new_n2085_, new_n2086_,
    new_n2087_, new_n2088_, new_n2089_, new_n2090_, new_n2091_, new_n2092_,
    new_n2093_, new_n2094_, new_n2095_, new_n2096_, new_n2097_, new_n2098_,
    new_n2099_, new_n2100_, new_n2101_, new_n2102_, new_n2103_, new_n2104_,
    new_n2105_, new_n2106_, new_n2107_, new_n2108_, new_n2109_, new_n2110_,
    new_n2111_, new_n2112_, new_n2113_, new_n2114_, new_n2116_, new_n2117_,
    new_n2118_, new_n2119_, new_n2120_, new_n2121_, new_n2122_, new_n2123_,
    new_n2124_, new_n2125_, new_n2126_, new_n2127_, new_n2128_, new_n2129_,
    new_n2130_, new_n2131_, new_n2132_, new_n2133_, new_n2134_, new_n2135_,
    new_n2136_, new_n2137_, new_n2138_, new_n2139_, new_n2140_, new_n2141_,
    new_n2142_, new_n2143_, new_n2144_, new_n2145_, new_n2146_, new_n2147_,
    new_n2148_, new_n2149_, new_n2150_, new_n2151_, new_n2152_, new_n2153_,
    new_n2154_, new_n2155_, new_n2156_, new_n2157_, new_n2158_, new_n2160_,
    new_n2161_, new_n2162_, new_n2163_, new_n2164_, new_n2165_, new_n2166_,
    new_n2167_, new_n2168_, new_n2169_, new_n2170_, new_n2171_, new_n2172_,
    new_n2173_, new_n2174_, new_n2175_, new_n2176_, new_n2177_, new_n2178_,
    new_n2179_, new_n2180_, new_n2181_, new_n2182_, new_n2183_, new_n2184_,
    new_n2185_, new_n2186_, new_n2187_, new_n2188_, new_n2189_, new_n2190_,
    new_n2191_, new_n2192_, new_n2193_, new_n2194_, new_n2195_, new_n2196_,
    new_n2197_, new_n2198_, new_n2199_, new_n2200_, new_n2201_, new_n2202_,
    new_n2204_, new_n2205_, new_n2206_, new_n2207_, new_n2208_, new_n2209_,
    new_n2210_, new_n2211_, new_n2212_, new_n2213_, new_n2214_, new_n2215_,
    new_n2216_, new_n2217_, new_n2218_, new_n2219_, new_n2220_, new_n2221_,
    new_n2222_, new_n2223_, new_n2224_, new_n2225_, new_n2226_, new_n2227_,
    new_n2228_, new_n2229_, new_n2230_, new_n2231_, new_n2232_, new_n2233_,
    new_n2234_, new_n2235_, new_n2236_, new_n2237_, new_n2238_, new_n2239_,
    new_n2240_, new_n2241_, new_n2242_, new_n2243_, new_n2244_, new_n2245_,
    new_n2246_, new_n2248_, new_n2249_, new_n2250_, new_n2251_, new_n2252_,
    new_n2253_, new_n2254_, new_n2255_, new_n2256_, new_n2257_, new_n2258_,
    new_n2259_, new_n2260_, new_n2261_, new_n2262_, new_n2263_, new_n2264_,
    new_n2265_, new_n2266_, new_n2267_, new_n2268_, new_n2269_, new_n2270_,
    new_n2271_, new_n2272_, new_n2273_, new_n2274_, new_n2275_, new_n2276_,
    new_n2277_, new_n2278_, new_n2279_, new_n2280_, new_n2281_, new_n2282_,
    new_n2283_, new_n2284_, new_n2285_, new_n2286_, new_n2287_, new_n2288_,
    new_n2289_, new_n2290_, new_n2292_, new_n2293_, new_n2294_, new_n2295_,
    new_n2296_, new_n2297_, new_n2298_, new_n2299_, new_n2300_, new_n2301_,
    new_n2302_, new_n2303_, new_n2304_, new_n2305_, new_n2306_, new_n2307_,
    new_n2308_, new_n2309_, new_n2310_, new_n2311_, new_n2312_, new_n2313_,
    new_n2314_, new_n2315_, new_n2316_, new_n2317_, new_n2318_, new_n2319_,
    new_n2320_, new_n2321_, new_n2322_, new_n2323_, new_n2324_, new_n2325_,
    new_n2326_, new_n2327_, new_n2328_, new_n2329_, new_n2330_, new_n2331_,
    new_n2332_, new_n2333_, new_n2334_, new_n2336_, new_n2337_, new_n2338_,
    new_n2339_, new_n2340_, new_n2341_, new_n2342_, new_n2343_, new_n2344_,
    new_n2345_, new_n2346_, new_n2347_, new_n2348_, new_n2349_, new_n2350_,
    new_n2351_, new_n2352_, new_n2353_, new_n2354_, new_n2355_, new_n2356_,
    new_n2357_, new_n2358_, new_n2359_, new_n2360_, new_n2361_, new_n2362_,
    new_n2363_, new_n2364_, new_n2365_, new_n2366_, new_n2367_, new_n2368_,
    new_n2369_, new_n2370_, new_n2371_, new_n2372_, new_n2373_, new_n2374_,
    new_n2375_, new_n2376_, new_n2377_, new_n2378_, new_n2380_, new_n2381_,
    new_n2382_, new_n2383_, new_n2384_, new_n2385_, new_n2386_, new_n2387_,
    new_n2388_, new_n2389_, new_n2390_, new_n2391_, new_n2392_, new_n2393_,
    new_n2394_, new_n2395_, new_n2396_, new_n2397_, new_n2398_, new_n2399_,
    new_n2400_, new_n2401_, new_n2402_, new_n2403_, new_n2404_, new_n2405_,
    new_n2406_, new_n2407_, new_n2408_, new_n2409_, new_n2410_, new_n2411_,
    new_n2412_, new_n2413_, new_n2414_, new_n2415_, new_n2416_, new_n2417_,
    new_n2418_, new_n2419_, new_n2420_, new_n2421_, new_n2422_, new_n2424_,
    new_n2425_, new_n2426_, new_n2427_, new_n2428_, new_n2429_, new_n2430_,
    new_n2431_, new_n2432_, new_n2433_, new_n2434_, new_n2435_, new_n2436_,
    new_n2437_, new_n2438_, new_n2439_, new_n2440_, new_n2441_, new_n2442_,
    new_n2443_, new_n2444_, new_n2445_, new_n2446_, new_n2447_, new_n2448_,
    new_n2449_, new_n2450_, new_n2451_, new_n2452_, new_n2453_, new_n2454_,
    new_n2455_, new_n2456_, new_n2457_, new_n2458_, new_n2459_, new_n2460_,
    new_n2461_, new_n2462_, new_n2463_, new_n2464_, new_n2465_, new_n2466_,
    new_n2468_, new_n2469_, new_n2470_, new_n2471_, new_n2472_, new_n2473_,
    new_n2474_, new_n2475_, new_n2476_, new_n2477_, new_n2478_, new_n2479_,
    new_n2480_, new_n2481_, new_n2482_, new_n2483_, new_n2484_, new_n2485_,
    new_n2486_, new_n2487_, new_n2488_, new_n2489_, new_n2490_, new_n2491_,
    new_n2492_, new_n2493_, new_n2494_, new_n2495_, new_n2496_, new_n2497_,
    new_n2498_, new_n2499_, new_n2500_, new_n2501_, new_n2502_, new_n2503_,
    new_n2504_, new_n2505_, new_n2506_, new_n2507_, new_n2508_, new_n2509_,
    new_n2510_, new_n2512_, new_n2513_, new_n2514_, new_n2515_, new_n2516_,
    new_n2517_, new_n2518_, new_n2519_, new_n2520_, new_n2521_, new_n2522_,
    new_n2523_, new_n2524_, new_n2525_, new_n2526_, new_n2527_, new_n2528_,
    new_n2529_, new_n2530_, new_n2531_, new_n2532_, new_n2533_, new_n2534_,
    new_n2535_, new_n2536_, new_n2537_, new_n2538_, new_n2539_, new_n2540_,
    new_n2541_, new_n2542_, new_n2543_, new_n2544_, new_n2545_, new_n2546_,
    new_n2547_, new_n2548_, new_n2549_, new_n2550_, new_n2551_, new_n2552_,
    new_n2553_, new_n2554_, new_n2556_, new_n2557_, new_n2558_, new_n2559_,
    new_n2560_, new_n2561_, new_n2562_, new_n2563_, new_n2564_, new_n2565_,
    new_n2566_, new_n2567_, new_n2568_, new_n2569_, new_n2570_, new_n2571_,
    new_n2572_, new_n2573_, new_n2574_, new_n2575_, new_n2576_, new_n2577_,
    new_n2578_, new_n2579_, new_n2580_, new_n2581_, new_n2582_, new_n2583_,
    new_n2584_, new_n2585_, new_n2586_, new_n2587_, new_n2588_, new_n2589_,
    new_n2590_, new_n2591_, new_n2592_, new_n2593_, new_n2594_, new_n2595_,
    new_n2596_, new_n2597_, new_n2598_, new_n2600_, new_n2601_, new_n2602_,
    new_n2603_, new_n2604_, new_n2605_, new_n2606_, new_n2607_, new_n2608_,
    new_n2609_, new_n2610_, new_n2611_, new_n2612_, new_n2613_, new_n2614_,
    new_n2615_, new_n2616_, new_n2617_, new_n2618_, new_n2619_, new_n2620_,
    new_n2621_, new_n2622_, new_n2623_, new_n2624_, new_n2625_, new_n2626_,
    new_n2627_, new_n2628_, new_n2629_, new_n2630_, new_n2631_, new_n2632_,
    new_n2633_, new_n2634_, new_n2635_, new_n2636_, new_n2637_, new_n2638_,
    new_n2639_, new_n2640_, new_n2641_, new_n2642_, new_n2644_, new_n2645_,
    new_n2646_, new_n2647_, new_n2648_, new_n2649_, new_n2650_, new_n2651_,
    new_n2652_, new_n2653_, new_n2654_, new_n2655_, new_n2656_, new_n2657_,
    new_n2658_, new_n2659_, new_n2660_, new_n2661_, new_n2662_, new_n2663_,
    new_n2664_, new_n2665_, new_n2666_, new_n2667_, new_n2668_, new_n2669_,
    new_n2670_, new_n2671_, new_n2672_, new_n2673_, new_n2674_, new_n2675_,
    new_n2676_, new_n2677_, new_n2678_, new_n2679_, new_n2680_, new_n2681_,
    new_n2682_, new_n2683_, new_n2684_, new_n2685_, new_n2686_, new_n2688_,
    new_n2689_, new_n2690_, new_n2691_, new_n2692_, new_n2693_, new_n2694_,
    new_n2695_, new_n2696_, new_n2697_, new_n2698_, new_n2699_, new_n2700_,
    new_n2701_, new_n2702_, new_n2703_, new_n2704_, new_n2705_, new_n2706_,
    new_n2707_, new_n2708_, new_n2709_, new_n2710_, new_n2711_, new_n2712_,
    new_n2713_, new_n2714_, new_n2715_, new_n2716_, new_n2717_, new_n2718_,
    new_n2719_, new_n2720_, new_n2721_, new_n2722_, new_n2723_, new_n2724_,
    new_n2725_, new_n2726_, new_n2727_, new_n2728_, new_n2729_, new_n2730_,
    new_n2732_, new_n2733_, new_n2734_, new_n2735_, new_n2736_, new_n2737_,
    new_n2738_, new_n2739_, new_n2740_, new_n2741_, new_n2742_, new_n2743_,
    new_n2744_, new_n2745_, new_n2746_, new_n2747_, new_n2748_, new_n2749_,
    new_n2750_, new_n2751_, new_n2752_, new_n2753_, new_n2754_, new_n2755_,
    new_n2756_, new_n2757_, new_n2758_, new_n2759_, new_n2760_, new_n2761_,
    new_n2762_, new_n2763_, new_n2764_, new_n2765_, new_n2766_, new_n2767_,
    new_n2768_, new_n2769_, new_n2770_, new_n2771_, new_n2772_, new_n2773_,
    new_n2774_, new_n2776_, new_n2777_, new_n2778_, new_n2779_, new_n2780_,
    new_n2781_, new_n2782_, new_n2783_, new_n2784_, new_n2785_, new_n2786_,
    new_n2787_, new_n2788_, new_n2789_, new_n2790_, new_n2791_, new_n2792_,
    new_n2793_, new_n2794_, new_n2795_, new_n2796_, new_n2797_, new_n2798_,
    new_n2799_, new_n2800_, new_n2801_, new_n2802_, new_n2803_, new_n2804_,
    new_n2805_, new_n2806_, new_n2807_, new_n2808_, new_n2809_, new_n2810_,
    new_n2811_, new_n2812_, new_n2813_, new_n2814_, new_n2815_, new_n2816_,
    new_n2817_, new_n2818_, new_n2820_, new_n2821_, new_n2822_, new_n2823_,
    new_n2824_, new_n2825_, new_n2826_, new_n2827_, new_n2828_, new_n2829_,
    new_n2830_, new_n2831_, new_n2832_, new_n2833_, new_n2834_, new_n2835_,
    new_n2836_, new_n2837_, new_n2838_, new_n2839_, new_n2840_, new_n2841_,
    new_n2842_, new_n2843_, new_n2844_, new_n2845_, new_n2846_, new_n2847_,
    new_n2848_, new_n2849_, new_n2850_, new_n2851_, new_n2852_, new_n2853_,
    new_n2854_, new_n2855_, new_n2856_, new_n2857_, new_n2858_, new_n2859_,
    new_n2860_, new_n2861_, new_n2862_, new_n2864_, new_n2865_, new_n2866_,
    new_n2867_, new_n2868_, new_n2869_, new_n2870_, new_n2871_, new_n2872_,
    new_n2873_, new_n2874_, new_n2875_, new_n2876_, new_n2877_, new_n2878_,
    new_n2879_, new_n2880_, new_n2881_, new_n2882_, new_n2883_, new_n2884_,
    new_n2885_, new_n2886_, new_n2887_, new_n2888_, new_n2889_, new_n2890_,
    new_n2891_, new_n2892_, new_n2893_, new_n2894_, new_n2895_, new_n2896_,
    new_n2897_, new_n2898_, new_n2899_, new_n2900_, new_n2901_, new_n2902_,
    new_n2903_, new_n2904_, new_n2905_, new_n2906_, new_n2908_, new_n2909_,
    new_n2910_, new_n2911_, new_n2912_, new_n2913_, new_n2914_, new_n2915_,
    new_n2916_, new_n2917_, new_n2918_, new_n2919_, new_n2920_, new_n2921_,
    new_n2922_, new_n2923_, new_n2924_, new_n2925_, new_n2926_, new_n2927_,
    new_n2928_, new_n2929_, new_n2930_, new_n2931_, new_n2932_, new_n2933_,
    new_n2934_, new_n2935_, new_n2936_, new_n2937_, new_n2938_, new_n2939_,
    new_n2940_, new_n2941_, new_n2942_, new_n2943_, new_n2944_, new_n2945_,
    new_n2946_, new_n2947_, new_n2948_, new_n2949_, new_n2950_, new_n2952_,
    new_n2953_, new_n2954_, new_n2955_, new_n2956_, new_n2957_, new_n2958_,
    new_n2959_, new_n2960_, new_n2961_, new_n2962_, new_n2963_, new_n2964_,
    new_n2965_, new_n2966_, new_n2967_, new_n2968_, new_n2969_, new_n2970_,
    new_n2971_, new_n2972_, new_n2973_, new_n2974_, new_n2975_, new_n2976_,
    new_n2977_, new_n2978_, new_n2979_, new_n2980_, new_n2981_, new_n2982_,
    new_n2983_, new_n2984_, new_n2985_, new_n2986_, new_n2987_, new_n2988_,
    new_n2989_, new_n2990_, new_n2991_, new_n2992_, new_n2993_, new_n2994_,
    new_n2996_, new_n2997_, new_n2998_, new_n2999_, new_n3000_, new_n3001_,
    new_n3002_, new_n3003_, new_n3004_, new_n3005_, new_n3006_, new_n3007_,
    new_n3008_, new_n3009_, new_n3010_, new_n3011_, new_n3012_, new_n3013_,
    new_n3014_, new_n3015_, new_n3016_, new_n3017_, new_n3018_, new_n3019_,
    new_n3020_, new_n3021_, new_n3022_, new_n3023_, new_n3024_, new_n3025_,
    new_n3026_, new_n3027_, new_n3028_, new_n3029_, new_n3030_, new_n3031_,
    new_n3032_, new_n3033_, new_n3034_, new_n3035_, new_n3036_, new_n3037_,
    new_n3038_, new_n3040_, new_n3041_, new_n3042_, new_n3043_, new_n3044_,
    new_n3045_, new_n3046_, new_n3047_, new_n3048_, new_n3049_, new_n3050_,
    new_n3051_, new_n3052_, new_n3053_, new_n3054_, new_n3055_, new_n3056_,
    new_n3057_, new_n3058_, new_n3059_, new_n3060_, new_n3061_, new_n3062_,
    new_n3063_, new_n3064_, new_n3065_, new_n3066_, new_n3067_, new_n3068_,
    new_n3069_, new_n3070_, new_n3071_, new_n3072_, new_n3073_, new_n3074_,
    new_n3075_, new_n3076_, new_n3077_, new_n3078_, new_n3079_, new_n3080_,
    new_n3081_, new_n3082_, new_n3084_, new_n3085_, new_n3086_, new_n3087_,
    new_n3088_, new_n3089_, new_n3090_, new_n3091_, new_n3092_, new_n3093_,
    new_n3094_, new_n3095_, new_n3096_, new_n3097_, new_n3098_, new_n3099_,
    new_n3100_, new_n3101_, new_n3102_, new_n3103_, new_n3104_, new_n3105_,
    new_n3106_, new_n3107_, new_n3108_, new_n3109_, new_n3110_, new_n3111_,
    new_n3112_, new_n3113_, new_n3114_, new_n3115_, new_n3116_, new_n3117_,
    new_n3118_, new_n3119_, new_n3120_, new_n3121_, new_n3122_, new_n3123_,
    new_n3124_, new_n3125_, new_n3126_, new_n3128_, new_n3129_, new_n3130_,
    new_n3131_, new_n3132_, new_n3133_, new_n3134_, new_n3135_, new_n3136_,
    new_n3137_, new_n3138_, new_n3139_, new_n3140_, new_n3141_, new_n3142_,
    new_n3143_, new_n3144_, new_n3145_, new_n3146_, new_n3147_, new_n3148_,
    new_n3149_, new_n3150_, new_n3151_, new_n3152_, new_n3153_, new_n3154_,
    new_n3155_, new_n3156_, new_n3157_, new_n3158_, new_n3159_, new_n3160_,
    new_n3161_, new_n3162_, new_n3163_, new_n3164_, new_n3165_, new_n3166_,
    new_n3167_, new_n3168_, new_n3169_, new_n3170_, new_n3172_, new_n3173_,
    new_n3174_, new_n3175_, new_n3176_, new_n3177_, new_n3178_, new_n3179_,
    new_n3180_, new_n3181_, new_n3182_, new_n3183_, new_n3184_, new_n3185_,
    new_n3186_, new_n3187_, new_n3188_, new_n3189_, new_n3190_, new_n3191_,
    new_n3192_, new_n3193_, new_n3194_, new_n3195_, new_n3196_, new_n3197_,
    new_n3198_, new_n3199_, new_n3200_, new_n3201_, new_n3202_, new_n3203_,
    new_n3204_, new_n3205_, new_n3206_, new_n3207_, new_n3208_, new_n3209_,
    new_n3210_, new_n3211_, new_n3212_, new_n3213_, new_n3214_, new_n3216_,
    new_n3217_, new_n3218_, new_n3219_, new_n3220_, new_n3221_, new_n3222_,
    new_n3223_, new_n3224_, new_n3225_, new_n3226_, new_n3227_, new_n3228_,
    new_n3229_, new_n3230_, new_n3231_, new_n3232_, new_n3233_, new_n3234_,
    new_n3235_, new_n3236_, new_n3237_, new_n3238_, new_n3239_, new_n3240_,
    new_n3241_, new_n3242_, new_n3243_, new_n3244_, new_n3245_, new_n3246_,
    new_n3247_, new_n3248_, new_n3249_, new_n3250_, new_n3251_, new_n3252_,
    new_n3253_, new_n3254_, new_n3255_, new_n3256_, new_n3257_, new_n3258_,
    new_n3260_, new_n3261_, new_n3262_, new_n3263_, new_n3264_, new_n3265_,
    new_n3266_, new_n3267_, new_n3268_, new_n3269_, new_n3270_, new_n3271_,
    new_n3272_, new_n3273_, new_n3274_, new_n3275_, new_n3276_, new_n3277_,
    new_n3278_, new_n3279_, new_n3280_, new_n3281_, new_n3282_, new_n3283_,
    new_n3284_, new_n3285_, new_n3286_, new_n3287_, new_n3288_, new_n3289_,
    new_n3290_, new_n3291_, new_n3292_, new_n3293_, new_n3294_, new_n3295_,
    new_n3296_, new_n3297_, new_n3298_, new_n3299_, new_n3300_, new_n3301_,
    new_n3302_, new_n3304_, new_n3305_, new_n3306_, new_n3307_, new_n3308_,
    new_n3309_, new_n3310_, new_n3311_, new_n3312_, new_n3313_, new_n3314_,
    new_n3315_, new_n3316_, new_n3317_, new_n3318_, new_n3319_, new_n3320_,
    new_n3321_, new_n3322_, new_n3323_, new_n3324_, new_n3325_, new_n3326_,
    new_n3327_, new_n3328_, new_n3329_, new_n3330_, new_n3331_, new_n3332_,
    new_n3333_, new_n3334_, new_n3335_, new_n3336_, new_n3337_, new_n3338_,
    new_n3339_, new_n3340_, new_n3341_, new_n3342_, new_n3343_, new_n3344_,
    new_n3345_, new_n3346_, new_n3348_, new_n3349_, new_n3350_, new_n3351_,
    new_n3352_, new_n3353_, new_n3354_, new_n3355_, new_n3356_, new_n3357_,
    new_n3358_, new_n3359_, new_n3360_, new_n3361_, new_n3362_, new_n3363_,
    new_n3364_, new_n3365_, new_n3366_, new_n3367_, new_n3368_, new_n3369_,
    new_n3370_, new_n3371_, new_n3372_, new_n3373_, new_n3374_, new_n3375_,
    new_n3376_, new_n3377_, new_n3378_, new_n3379_, new_n3380_, new_n3381_,
    new_n3382_, new_n3383_, new_n3384_, new_n3385_, new_n3386_, new_n3387_,
    new_n3388_, new_n3389_, new_n3390_, new_n3392_, new_n3393_, new_n3394_,
    new_n3395_, new_n3396_, new_n3397_, new_n3398_, new_n3399_, new_n3400_,
    new_n3401_, new_n3402_, new_n3403_, new_n3404_, new_n3405_, new_n3406_,
    new_n3407_, new_n3408_, new_n3409_, new_n3410_, new_n3411_, new_n3412_,
    new_n3413_, new_n3414_, new_n3415_, new_n3416_, new_n3417_, new_n3418_,
    new_n3419_, new_n3420_, new_n3421_, new_n3422_, new_n3423_, new_n3424_,
    new_n3425_, new_n3426_, new_n3427_, new_n3428_, new_n3429_, new_n3430_,
    new_n3431_, new_n3432_, new_n3433_, new_n3434_, new_n3436_, new_n3437_,
    new_n3438_, new_n3439_, new_n3440_, new_n3441_, new_n3442_, new_n3443_,
    new_n3444_, new_n3445_, new_n3446_, new_n3447_, new_n3448_, new_n3449_,
    new_n3450_, new_n3451_, new_n3452_, new_n3453_, new_n3454_, new_n3455_,
    new_n3456_, new_n3457_, new_n3458_, new_n3459_, new_n3460_, new_n3461_,
    new_n3462_, new_n3463_, new_n3464_, new_n3465_, new_n3466_, new_n3467_,
    new_n3468_, new_n3469_, new_n3470_, new_n3471_, new_n3472_, new_n3473_,
    new_n3474_, new_n3475_, new_n3476_, new_n3477_, new_n3478_, new_n3480_,
    new_n3481_, new_n3482_, new_n3483_, new_n3484_, new_n3485_, new_n3486_,
    new_n3487_, new_n3488_, new_n3489_, new_n3490_, new_n3491_, new_n3492_,
    new_n3493_, new_n3494_, new_n3495_, new_n3496_, new_n3497_, new_n3498_,
    new_n3499_, new_n3500_, new_n3501_, new_n3502_, new_n3503_, new_n3504_,
    new_n3505_, new_n3506_, new_n3507_, new_n3508_, new_n3509_, new_n3510_,
    new_n3511_, new_n3512_, new_n3513_, new_n3514_, new_n3515_, new_n3516_,
    new_n3517_, new_n3518_, new_n3519_, new_n3520_, new_n3521_, new_n3522_,
    new_n3524_, new_n3525_, new_n3526_, new_n3527_, new_n3528_, new_n3529_,
    new_n3530_, new_n3531_, new_n3532_, new_n3533_, new_n3534_, new_n3535_,
    new_n3536_, new_n3537_, new_n3538_, new_n3539_, new_n3540_, new_n3541_,
    new_n3542_, new_n3543_, new_n3544_, new_n3545_, new_n3546_, new_n3547_,
    new_n3548_, new_n3549_, new_n3550_, new_n3551_, new_n3552_, new_n3553_,
    new_n3554_, new_n3555_, new_n3556_, new_n3557_, new_n3558_, new_n3559_,
    new_n3560_, new_n3561_, new_n3562_, new_n3563_, new_n3564_, new_n3565_,
    new_n3566_, new_n3568_, new_n3569_, new_n3570_, new_n3571_, new_n3572_,
    new_n3573_, new_n3574_, new_n3575_, new_n3576_, new_n3577_, new_n3578_,
    new_n3579_, new_n3580_, new_n3581_, new_n3582_, new_n3583_, new_n3584_,
    new_n3585_, new_n3586_, new_n3587_, new_n3588_, new_n3589_, new_n3590_,
    new_n3591_, new_n3592_, new_n3593_, new_n3594_, new_n3595_, new_n3596_,
    new_n3597_, new_n3598_, new_n3599_, new_n3600_, new_n3601_, new_n3602_,
    new_n3603_, new_n3604_, new_n3605_, new_n3606_, new_n3607_, new_n3608_,
    new_n3609_, new_n3610_, new_n3612_, new_n3613_, new_n3614_, new_n3615_,
    new_n3616_, new_n3617_, new_n3618_, new_n3619_, new_n3620_, new_n3621_,
    new_n3622_, new_n3623_, new_n3624_, new_n3625_, new_n3626_, new_n3627_,
    new_n3628_, new_n3629_, new_n3630_, new_n3631_, new_n3632_, new_n3633_,
    new_n3634_, new_n3635_, new_n3636_, new_n3637_, new_n3638_, new_n3639_,
    new_n3640_, new_n3641_, new_n3642_, new_n3643_, new_n3644_, new_n3645_,
    new_n3646_, new_n3647_, new_n3648_, new_n3649_, new_n3650_, new_n3651_,
    new_n3652_, new_n3653_, new_n3654_, new_n3656_, new_n3657_, new_n3658_,
    new_n3659_, new_n3660_, new_n3661_, new_n3662_, new_n3663_, new_n3664_,
    new_n3665_, new_n3666_, new_n3667_, new_n3668_, new_n3669_, new_n3670_,
    new_n3671_, new_n3672_, new_n3673_, new_n3674_, new_n3675_, new_n3676_,
    new_n3677_, new_n3678_, new_n3679_, new_n3680_, new_n3681_, new_n3682_,
    new_n3683_, new_n3684_, new_n3685_, new_n3686_, new_n3687_, new_n3688_,
    new_n3689_, new_n3690_, new_n3691_, new_n3692_, new_n3693_, new_n3694_,
    new_n3695_, new_n3696_, new_n3697_, new_n3698_, new_n3700_, new_n3701_,
    new_n3702_, new_n3703_, new_n3704_, new_n3705_, new_n3706_, new_n3707_,
    new_n3708_, new_n3709_, new_n3710_, new_n3711_, new_n3712_, new_n3713_,
    new_n3714_, new_n3715_, new_n3716_, new_n3717_, new_n3718_, new_n3719_,
    new_n3720_, new_n3721_, new_n3722_, new_n3723_, new_n3724_, new_n3725_,
    new_n3726_, new_n3727_, new_n3728_, new_n3729_, new_n3730_, new_n3731_,
    new_n3732_, new_n3733_, new_n3734_, new_n3735_, new_n3736_, new_n3737_,
    new_n3738_, new_n3739_, new_n3740_, new_n3741_, new_n3742_, new_n3744_,
    new_n3745_, new_n3746_, new_n3747_, new_n3748_, new_n3749_, new_n3750_,
    new_n3751_, new_n3752_, new_n3753_, new_n3754_, new_n3755_, new_n3756_,
    new_n3757_, new_n3758_, new_n3759_, new_n3760_, new_n3761_, new_n3762_,
    new_n3763_, new_n3764_, new_n3765_, new_n3766_, new_n3767_, new_n3768_,
    new_n3769_, new_n3770_, new_n3771_, new_n3772_, new_n3773_, new_n3774_,
    new_n3775_, new_n3776_, new_n3777_, new_n3778_, new_n3779_, new_n3780_,
    new_n3781_, new_n3782_, new_n3783_, new_n3784_, new_n3785_, new_n3786_,
    new_n3788_, new_n3789_, new_n3790_, new_n3791_, new_n3792_, new_n3793_,
    new_n3794_, new_n3795_, new_n3796_, new_n3797_, new_n3798_, new_n3799_,
    new_n3800_, new_n3801_, new_n3802_, new_n3803_, new_n3804_, new_n3805_,
    new_n3806_, new_n3807_, new_n3808_, new_n3809_, new_n3810_, new_n3811_,
    new_n3812_, new_n3813_, new_n3814_, new_n3815_, new_n3816_, new_n3817_,
    new_n3818_, new_n3819_, new_n3820_, new_n3821_, new_n3822_, new_n3823_,
    new_n3824_, new_n3825_, new_n3826_, new_n3827_, new_n3828_, new_n3829_,
    new_n3830_, new_n3832_, new_n3833_, new_n3834_, new_n3835_, new_n3836_,
    new_n3837_, new_n3838_, new_n3839_, new_n3840_, new_n3841_, new_n3842_,
    new_n3843_, new_n3844_, new_n3845_, new_n3846_, new_n3847_, new_n3848_,
    new_n3849_, new_n3850_, new_n3851_, new_n3852_, new_n3853_, new_n3854_,
    new_n3855_, new_n3856_, new_n3857_, new_n3858_, new_n3859_, new_n3860_,
    new_n3861_, new_n3862_, new_n3863_, new_n3864_, new_n3865_, new_n3866_,
    new_n3867_, new_n3868_, new_n3869_, new_n3870_, new_n3871_, new_n3872_,
    new_n3873_, new_n3874_, new_n3876_, new_n3877_, new_n3878_, new_n3879_,
    new_n3880_, new_n3881_, new_n3882_, new_n3883_, new_n3884_, new_n3885_,
    new_n3886_, new_n3887_, new_n3888_, new_n3889_, new_n3890_, new_n3891_,
    new_n3892_, new_n3893_, new_n3894_, new_n3895_, new_n3896_, new_n3897_,
    new_n3898_, new_n3899_, new_n3900_, new_n3901_, new_n3902_, new_n3903_,
    new_n3904_, new_n3905_, new_n3906_, new_n3907_, new_n3908_, new_n3909_,
    new_n3910_, new_n3911_, new_n3912_, new_n3913_, new_n3914_, new_n3915_,
    new_n3916_, new_n3917_, new_n3918_, new_n3920_, new_n3921_, new_n3922_,
    new_n3923_, new_n3924_, new_n3925_, new_n3926_, new_n3927_, new_n3928_,
    new_n3929_, new_n3930_, new_n3931_, new_n3932_, new_n3933_, new_n3934_,
    new_n3935_, new_n3936_, new_n3937_, new_n3938_, new_n3939_, new_n3940_,
    new_n3941_, new_n3942_, new_n3943_, new_n3944_, new_n3945_, new_n3946_,
    new_n3947_, new_n3948_, new_n3949_, new_n3950_, new_n3951_, new_n3952_,
    new_n3953_, new_n3954_, new_n3955_, new_n3956_, new_n3957_, new_n3958_,
    new_n3959_, new_n3960_, new_n3961_, new_n3962_, new_n3964_, new_n3965_,
    new_n3966_, new_n3967_, new_n3968_, new_n3969_, new_n3970_, new_n3971_,
    new_n3972_, new_n3973_, new_n3974_, new_n3975_, new_n3976_, new_n3977_,
    new_n3978_, new_n3979_, new_n3980_, new_n3981_, new_n3982_, new_n3983_,
    new_n3984_, new_n3985_, new_n3986_, new_n3987_, new_n3988_, new_n3989_,
    new_n3990_, new_n3991_, new_n3992_, new_n3993_, new_n3994_, new_n3995_,
    new_n3996_, new_n3997_, new_n3998_, new_n3999_, new_n4000_, new_n4001_,
    new_n4002_, new_n4003_, new_n4004_, new_n4005_, new_n4006_, new_n4008_,
    new_n4009_, new_n4010_, new_n4011_, new_n4012_, new_n4013_, new_n4014_,
    new_n4015_, new_n4016_, new_n4017_, new_n4018_, new_n4019_, new_n4020_,
    new_n4021_, new_n4022_, new_n4023_, new_n4024_, new_n4025_, new_n4026_,
    new_n4027_, new_n4028_, new_n4029_, new_n4030_, new_n4031_, new_n4032_,
    new_n4033_, new_n4034_, new_n4035_, new_n4036_, new_n4037_, new_n4038_,
    new_n4039_, new_n4040_, new_n4041_, new_n4042_, new_n4043_, new_n4044_,
    new_n4045_, new_n4046_, new_n4047_, new_n4048_, new_n4049_, new_n4050_,
    new_n4052_, new_n4053_, new_n4054_, new_n4055_, new_n4056_, new_n4057_,
    new_n4058_, new_n4059_, new_n4060_, new_n4061_, new_n4062_, new_n4063_,
    new_n4064_, new_n4065_, new_n4066_, new_n4067_, new_n4068_, new_n4069_,
    new_n4070_, new_n4071_, new_n4072_, new_n4073_, new_n4074_, new_n4075_,
    new_n4076_, new_n4077_, new_n4078_, new_n4079_, new_n4080_, new_n4081_,
    new_n4082_, new_n4083_, new_n4084_, new_n4085_, new_n4086_, new_n4087_,
    new_n4088_, new_n4089_, new_n4090_, new_n4091_, new_n4092_, new_n4093_,
    new_n4094_, new_n4096_, new_n4097_, new_n4098_, new_n4099_, new_n4100_,
    new_n4101_, new_n4102_, new_n4103_, new_n4104_, new_n4105_, new_n4106_,
    new_n4107_, new_n4108_, new_n4109_, new_n4110_, new_n4111_, new_n4112_,
    new_n4113_, new_n4114_, new_n4115_, new_n4116_, new_n4117_, new_n4118_,
    new_n4119_, new_n4120_, new_n4121_, new_n4122_, new_n4123_, new_n4124_,
    new_n4125_, new_n4126_, new_n4127_, new_n4128_, new_n4129_, new_n4130_,
    new_n4131_, new_n4132_, new_n4133_, new_n4134_, new_n4135_, new_n4136_,
    new_n4137_, new_n4138_, new_n4140_, new_n4141_, new_n4142_, new_n4143_,
    new_n4144_, new_n4145_, new_n4146_, new_n4147_, new_n4148_, new_n4149_,
    new_n4150_, new_n4151_, new_n4152_, new_n4153_, new_n4154_, new_n4155_,
    new_n4156_, new_n4157_, new_n4158_, new_n4159_, new_n4160_, new_n4161_,
    new_n4162_, new_n4163_, new_n4164_, new_n4165_, new_n4166_, new_n4167_,
    new_n4168_, new_n4169_, new_n4170_, new_n4171_, new_n4172_, new_n4173_,
    new_n4174_, new_n4175_, new_n4176_, new_n4177_, new_n4178_, new_n4179_,
    new_n4180_, new_n4181_, new_n4182_, new_n4184_, new_n4185_, new_n4186_,
    new_n4187_, new_n4188_, new_n4189_, new_n4190_, new_n4191_, new_n4192_,
    new_n4193_, new_n4194_, new_n4195_, new_n4196_, new_n4197_, new_n4198_,
    new_n4199_, new_n4200_, new_n4201_, new_n4202_, new_n4203_, new_n4204_,
    new_n4205_, new_n4206_, new_n4207_, new_n4208_, new_n4209_, new_n4210_,
    new_n4211_, new_n4212_, new_n4213_, new_n4214_, new_n4215_, new_n4216_,
    new_n4217_, new_n4218_, new_n4219_, new_n4220_, new_n4221_, new_n4222_,
    new_n4223_, new_n4224_, new_n4225_, new_n4226_, new_n4228_, new_n4229_,
    new_n4230_, new_n4231_, new_n4232_, new_n4233_, new_n4234_, new_n4235_,
    new_n4236_, new_n4237_, new_n4238_, new_n4239_, new_n4240_, new_n4241_,
    new_n4242_, new_n4243_, new_n4244_, new_n4245_, new_n4246_, new_n4247_,
    new_n4248_, new_n4249_, new_n4250_, new_n4251_, new_n4252_, new_n4253_,
    new_n4254_, new_n4255_, new_n4256_, new_n4257_, new_n4258_, new_n4259_,
    new_n4260_, new_n4261_, new_n4262_, new_n4263_, new_n4264_, new_n4265_,
    new_n4266_, new_n4267_, new_n4268_, new_n4269_, new_n4270_, new_n4272_,
    new_n4273_, new_n4274_, new_n4275_, new_n4276_, new_n4277_, new_n4278_,
    new_n4279_, new_n4280_, new_n4281_, new_n4282_, new_n4283_, new_n4284_,
    new_n4285_, new_n4286_, new_n4287_, new_n4288_, new_n4289_, new_n4290_,
    new_n4291_, new_n4292_, new_n4293_, new_n4294_, new_n4295_, new_n4296_,
    new_n4297_, new_n4298_, new_n4299_, new_n4300_, new_n4301_, new_n4302_,
    new_n4303_, new_n4304_, new_n4305_, new_n4306_, new_n4307_, new_n4308_,
    new_n4309_, new_n4310_, new_n4311_, new_n4312_, new_n4313_, new_n4314_,
    new_n4316_, new_n4317_, new_n4318_, new_n4319_, new_n4320_, new_n4321_,
    new_n4322_, new_n4323_, new_n4324_, new_n4325_, new_n4326_, new_n4327_,
    new_n4328_, new_n4329_, new_n4330_, new_n4331_, new_n4332_, new_n4333_,
    new_n4334_, new_n4335_, new_n4336_, new_n4337_, new_n4338_, new_n4339_,
    new_n4340_, new_n4341_, new_n4342_, new_n4343_, new_n4344_, new_n4345_,
    new_n4346_, new_n4347_, new_n4348_, new_n4349_, new_n4350_, new_n4351_,
    new_n4352_, new_n4353_, new_n4354_, new_n4355_, new_n4356_, new_n4357_,
    new_n4358_, new_n4360_, new_n4361_, new_n4362_, new_n4363_, new_n4364_,
    new_n4365_, new_n4366_, new_n4367_, new_n4368_, new_n4369_, new_n4370_,
    new_n4371_, new_n4372_, new_n4373_, new_n4374_, new_n4375_, new_n4376_,
    new_n4377_, new_n4378_, new_n4379_, new_n4380_, new_n4381_, new_n4382_,
    new_n4383_, new_n4384_, new_n4385_, new_n4386_, new_n4387_, new_n4388_,
    new_n4389_, new_n4390_, new_n4391_, new_n4392_, new_n4393_, new_n4394_,
    new_n4395_, new_n4396_, new_n4397_, new_n4398_, new_n4399_, new_n4400_,
    new_n4401_, new_n4402_, new_n4404_, new_n4405_, new_n4406_, new_n4407_,
    new_n4408_, new_n4409_, new_n4410_, new_n4411_, new_n4412_, new_n4413_,
    new_n4414_, new_n4415_, new_n4416_, new_n4417_, new_n4418_, new_n4419_,
    new_n4420_, new_n4421_, new_n4422_, new_n4423_, new_n4424_, new_n4425_,
    new_n4426_, new_n4427_, new_n4428_, new_n4429_, new_n4430_, new_n4431_,
    new_n4432_, new_n4433_, new_n4434_, new_n4435_, new_n4436_, new_n4437_,
    new_n4438_, new_n4439_, new_n4440_, new_n4441_, new_n4442_, new_n4443_,
    new_n4444_, new_n4445_, new_n4446_, new_n4448_, new_n4449_, new_n4450_,
    new_n4451_, new_n4452_, new_n4453_, new_n4454_, new_n4455_, new_n4456_,
    new_n4457_, new_n4458_, new_n4459_, new_n4460_, new_n4461_, new_n4462_,
    new_n4463_, new_n4464_, new_n4465_, new_n4466_, new_n4467_, new_n4468_,
    new_n4469_, new_n4470_, new_n4471_, new_n4472_, new_n4473_, new_n4474_,
    new_n4475_, new_n4476_, new_n4477_, new_n4478_, new_n4479_, new_n4480_,
    new_n4481_, new_n4482_, new_n4483_, new_n4484_, new_n4485_, new_n4486_,
    new_n4487_, new_n4488_, new_n4489_, new_n4490_, new_n4492_, new_n4493_,
    new_n4494_, new_n4495_, new_n4496_, new_n4497_, new_n4498_, new_n4499_,
    new_n4500_, new_n4501_, new_n4502_, new_n4503_, new_n4504_, new_n4505_,
    new_n4506_, new_n4507_, new_n4508_, new_n4509_, new_n4510_, new_n4511_,
    new_n4512_, new_n4513_, new_n4514_, new_n4515_, new_n4516_, new_n4517_,
    new_n4518_, new_n4519_, new_n4520_, new_n4521_, new_n4522_, new_n4523_,
    new_n4524_, new_n4525_, new_n4526_, new_n4527_, new_n4528_, new_n4529_,
    new_n4530_, new_n4531_, new_n4532_, new_n4533_, new_n4534_, new_n4536_,
    new_n4537_, new_n4538_, new_n4539_, new_n4540_, new_n4541_, new_n4542_,
    new_n4543_, new_n4544_, new_n4545_, new_n4546_, new_n4547_, new_n4548_,
    new_n4549_, new_n4550_, new_n4551_, new_n4552_, new_n4553_, new_n4554_,
    new_n4555_, new_n4556_, new_n4557_, new_n4558_, new_n4559_, new_n4560_,
    new_n4561_, new_n4562_, new_n4563_, new_n4564_, new_n4565_, new_n4566_,
    new_n4567_, new_n4568_, new_n4569_, new_n4570_, new_n4571_, new_n4572_,
    new_n4573_, new_n4574_, new_n4575_, new_n4576_, new_n4577_, new_n4578_,
    new_n4580_, new_n4581_, new_n4582_, new_n4583_, new_n4584_, new_n4585_,
    new_n4586_, new_n4587_, new_n4588_, new_n4589_, new_n4590_, new_n4591_,
    new_n4592_, new_n4593_, new_n4594_, new_n4595_, new_n4596_, new_n4597_,
    new_n4598_, new_n4599_, new_n4600_, new_n4601_, new_n4602_, new_n4603_,
    new_n4604_, new_n4605_, new_n4606_, new_n4607_, new_n4608_, new_n4609_,
    new_n4610_, new_n4611_, new_n4612_, new_n4613_, new_n4614_, new_n4615_,
    new_n4616_, new_n4617_, new_n4618_, new_n4619_, new_n4620_, new_n4621_,
    new_n4622_, new_n4624_, new_n4625_, new_n4626_, new_n4627_, new_n4628_,
    new_n4629_, new_n4630_, new_n4631_, new_n4632_, new_n4633_, new_n4634_,
    new_n4635_, new_n4636_, new_n4637_, new_n4638_, new_n4639_, new_n4640_,
    new_n4641_, new_n4642_, new_n4643_, new_n4644_, new_n4645_, new_n4646_,
    new_n4647_, new_n4648_, new_n4649_, new_n4650_, new_n4651_, new_n4652_,
    new_n4653_, new_n4654_, new_n4655_, new_n4656_, new_n4657_, new_n4658_,
    new_n4659_, new_n4660_, new_n4661_, new_n4662_, new_n4663_, new_n4664_,
    new_n4665_, new_n4666_, new_n4668_, new_n4669_, new_n4670_, new_n4671_,
    new_n4672_, new_n4673_, new_n4674_, new_n4675_, new_n4676_, new_n4677_,
    new_n4678_, new_n4679_, new_n4680_, new_n4681_, new_n4682_, new_n4683_,
    new_n4684_, new_n4685_, new_n4686_, new_n4687_, new_n4688_, new_n4689_,
    new_n4690_, new_n4691_, new_n4692_, new_n4693_, new_n4694_, new_n4695_,
    new_n4696_, new_n4697_, new_n4698_, new_n4699_, new_n4700_, new_n4701_,
    new_n4702_, new_n4703_, new_n4704_, new_n4705_, new_n4706_, new_n4707_,
    new_n4708_, new_n4709_, new_n4710_, new_n4712_, new_n4713_, new_n4714_,
    new_n4715_, new_n4716_, new_n4717_, new_n4718_, new_n4719_, new_n4720_,
    new_n4721_, new_n4722_, new_n4723_, new_n4724_, new_n4725_, new_n4726_,
    new_n4727_, new_n4728_, new_n4729_, new_n4730_, new_n4731_, new_n4732_,
    new_n4733_, new_n4734_, new_n4735_, new_n4736_, new_n4737_, new_n4738_,
    new_n4739_, new_n4740_, new_n4741_, new_n4742_, new_n4743_, new_n4744_,
    new_n4745_, new_n4746_, new_n4747_, new_n4748_, new_n4749_, new_n4750_,
    new_n4751_, new_n4752_, new_n4753_, new_n4754_, new_n4756_, new_n4757_,
    new_n4758_, new_n4759_, new_n4760_, new_n4761_, new_n4762_, new_n4763_,
    new_n4764_, new_n4765_, new_n4766_, new_n4767_, new_n4768_, new_n4769_,
    new_n4770_, new_n4771_, new_n4772_, new_n4773_, new_n4774_, new_n4775_,
    new_n4776_, new_n4777_, new_n4778_, new_n4779_, new_n4780_, new_n4781_,
    new_n4782_, new_n4783_, new_n4784_, new_n4785_, new_n4786_, new_n4787_,
    new_n4788_, new_n4789_, new_n4790_, new_n4791_, new_n4792_, new_n4793_,
    new_n4794_, new_n4795_, new_n4796_, new_n4797_, new_n4798_, new_n4800_,
    new_n4801_, new_n4802_, new_n4803_, new_n4804_, new_n4805_, new_n4806_,
    new_n4807_, new_n4808_, new_n4809_, new_n4810_, new_n4811_, new_n4812_,
    new_n4813_, new_n4814_, new_n4815_, new_n4816_, new_n4817_, new_n4818_,
    new_n4819_, new_n4820_, new_n4821_, new_n4822_, new_n4823_, new_n4824_,
    new_n4825_, new_n4826_, new_n4827_, new_n4828_, new_n4829_, new_n4830_,
    new_n4831_, new_n4832_, new_n4833_, new_n4834_, new_n4835_, new_n4836_,
    new_n4837_, new_n4838_, new_n4839_, new_n4840_, new_n4841_, new_n4842_,
    new_n4844_, new_n4845_, new_n4846_, new_n4847_, new_n4848_, new_n4849_,
    new_n4850_, new_n4851_, new_n4852_, new_n4853_, new_n4854_, new_n4855_,
    new_n4856_, new_n4857_, new_n4858_, new_n4859_, new_n4860_, new_n4861_,
    new_n4862_, new_n4863_, new_n4864_, new_n4865_, new_n4866_, new_n4867_,
    new_n4868_, new_n4869_, new_n4870_, new_n4871_, new_n4872_, new_n4873_,
    new_n4874_, new_n4875_, new_n4876_, new_n4877_, new_n4878_, new_n4879_,
    new_n4880_, new_n4881_, new_n4882_, new_n4883_, new_n4884_, new_n4885_,
    new_n4886_, new_n4888_, new_n4889_, new_n4890_, new_n4891_, new_n4892_,
    new_n4893_, new_n4894_, new_n4895_, new_n4896_, new_n4897_, new_n4898_,
    new_n4899_, new_n4900_, new_n4901_, new_n4902_, new_n4903_, new_n4904_,
    new_n4905_, new_n4906_, new_n4907_, new_n4908_, new_n4909_, new_n4910_,
    new_n4911_, new_n4912_, new_n4913_, new_n4914_, new_n4915_, new_n4916_,
    new_n4917_, new_n4918_, new_n4919_, new_n4920_, new_n4921_, new_n4922_,
    new_n4923_, new_n4924_, new_n4925_, new_n4926_, new_n4927_, new_n4928_,
    new_n4929_, new_n4930_, new_n4932_, new_n4933_, new_n4934_, new_n4935_,
    new_n4936_, new_n4937_, new_n4938_, new_n4939_, new_n4940_, new_n4941_,
    new_n4942_, new_n4943_, new_n4944_, new_n4945_, new_n4946_, new_n4947_,
    new_n4948_, new_n4949_, new_n4950_, new_n4951_, new_n4952_, new_n4953_,
    new_n4954_, new_n4955_, new_n4956_, new_n4957_, new_n4958_, new_n4959_,
    new_n4960_, new_n4961_, new_n4962_, new_n4963_, new_n4964_, new_n4965_,
    new_n4966_, new_n4967_, new_n4968_, new_n4969_, new_n4970_, new_n4971_,
    new_n4972_, new_n4973_, new_n4974_, new_n4976_, new_n4977_, new_n4978_,
    new_n4979_, new_n4980_, new_n4981_, new_n4982_, new_n4983_, new_n4984_,
    new_n4985_, new_n4986_, new_n4987_, new_n4988_, new_n4989_, new_n4990_,
    new_n4991_, new_n4992_, new_n4993_, new_n4994_, new_n4995_, new_n4996_,
    new_n4997_, new_n4998_, new_n4999_, new_n5000_, new_n5001_, new_n5002_,
    new_n5003_, new_n5004_, new_n5005_, new_n5006_, new_n5007_, new_n5008_,
    new_n5009_, new_n5010_, new_n5011_, new_n5012_, new_n5013_, new_n5014_,
    new_n5015_, new_n5016_, new_n5017_, new_n5018_, new_n5020_, new_n5021_,
    new_n5022_, new_n5023_, new_n5024_, new_n5025_, new_n5026_, new_n5027_,
    new_n5028_, new_n5029_, new_n5030_, new_n5031_, new_n5032_, new_n5033_,
    new_n5034_, new_n5035_, new_n5036_, new_n5037_, new_n5038_, new_n5039_,
    new_n5040_, new_n5041_, new_n5042_, new_n5043_, new_n5044_, new_n5045_,
    new_n5046_, new_n5047_, new_n5048_, new_n5049_, new_n5050_, new_n5051_,
    new_n5052_, new_n5053_, new_n5054_, new_n5055_, new_n5056_, new_n5057_,
    new_n5058_, new_n5059_, new_n5060_, new_n5061_, new_n5062_, new_n5064_,
    new_n5065_, new_n5066_, new_n5067_, new_n5068_, new_n5069_, new_n5070_,
    new_n5071_, new_n5072_, new_n5073_, new_n5074_, new_n5075_, new_n5076_,
    new_n5077_, new_n5078_, new_n5079_, new_n5080_, new_n5081_, new_n5082_,
    new_n5083_, new_n5084_, new_n5085_, new_n5086_, new_n5087_, new_n5088_,
    new_n5089_, new_n5090_, new_n5091_, new_n5092_, new_n5093_, new_n5094_,
    new_n5095_, new_n5096_, new_n5097_, new_n5098_, new_n5099_, new_n5100_,
    new_n5101_, new_n5102_, new_n5103_, new_n5104_, new_n5105_, new_n5106_,
    new_n5108_, new_n5109_, new_n5110_, new_n5111_, new_n5112_, new_n5113_,
    new_n5114_, new_n5115_, new_n5116_, new_n5117_, new_n5118_, new_n5119_,
    new_n5120_, new_n5121_, new_n5122_, new_n5123_, new_n5124_, new_n5125_,
    new_n5126_, new_n5127_, new_n5128_, new_n5129_, new_n5130_, new_n5131_,
    new_n5132_, new_n5133_, new_n5134_, new_n5135_, new_n5136_, new_n5137_,
    new_n5138_, new_n5139_, new_n5140_, new_n5141_, new_n5142_, new_n5143_,
    new_n5144_, new_n5145_, new_n5146_, new_n5147_, new_n5148_, new_n5149_,
    new_n5150_, new_n5152_, new_n5153_, new_n5154_, new_n5155_, new_n5156_,
    new_n5157_, new_n5158_, new_n5159_, new_n5160_, new_n5161_, new_n5162_,
    new_n5163_, new_n5164_, new_n5165_, new_n5166_, new_n5167_, new_n5168_,
    new_n5169_, new_n5170_, new_n5171_, new_n5172_, new_n5173_, new_n5174_,
    new_n5175_, new_n5176_, new_n5177_, new_n5178_, new_n5179_, new_n5180_,
    new_n5181_, new_n5182_, new_n5183_, new_n5184_, new_n5185_, new_n5186_,
    new_n5187_, new_n5188_, new_n5189_, new_n5190_, new_n5191_, new_n5192_,
    new_n5193_, new_n5194_, new_n5196_, new_n5197_, new_n5198_, new_n5199_,
    new_n5200_, new_n5201_, new_n5202_, new_n5203_, new_n5204_, new_n5205_,
    new_n5206_, new_n5207_, new_n5208_, new_n5209_, new_n5210_, new_n5211_,
    new_n5212_, new_n5213_, new_n5214_, new_n5215_, new_n5216_, new_n5217_,
    new_n5218_, new_n5219_, new_n5220_, new_n5221_, new_n5222_, new_n5223_,
    new_n5224_, new_n5225_, new_n5226_, new_n5227_, new_n5228_, new_n5229_,
    new_n5230_, new_n5231_, new_n5232_, new_n5233_, new_n5234_, new_n5235_,
    new_n5236_, new_n5237_, new_n5238_, new_n5240_, new_n5241_, new_n5242_,
    new_n5243_, new_n5244_, new_n5245_, new_n5246_, new_n5247_, new_n5248_,
    new_n5249_, new_n5250_, new_n5251_, new_n5252_, new_n5253_, new_n5254_,
    new_n5255_, new_n5256_, new_n5257_, new_n5258_, new_n5259_, new_n5260_,
    new_n5261_, new_n5262_, new_n5263_, new_n5264_, new_n5265_, new_n5266_,
    new_n5267_, new_n5268_, new_n5269_, new_n5270_, new_n5271_, new_n5272_,
    new_n5273_, new_n5274_, new_n5275_, new_n5276_, new_n5277_, new_n5278_,
    new_n5279_, new_n5280_, new_n5281_, new_n5282_, new_n5284_, new_n5285_,
    new_n5286_, new_n5287_, new_n5288_, new_n5289_, new_n5290_, new_n5291_,
    new_n5292_, new_n5293_, new_n5294_, new_n5295_, new_n5296_, new_n5297_,
    new_n5298_, new_n5299_, new_n5300_, new_n5301_, new_n5302_, new_n5303_,
    new_n5304_, new_n5305_, new_n5306_, new_n5307_, new_n5308_, new_n5309_,
    new_n5310_, new_n5311_, new_n5312_, new_n5313_, new_n5314_, new_n5315_,
    new_n5316_, new_n5317_, new_n5318_, new_n5319_, new_n5320_, new_n5321_,
    new_n5322_, new_n5323_, new_n5324_, new_n5325_, new_n5326_, new_n5328_,
    new_n5329_, new_n5330_, new_n5331_, new_n5332_, new_n5333_, new_n5334_,
    new_n5335_, new_n5336_, new_n5337_, new_n5338_, new_n5339_, new_n5340_,
    new_n5341_, new_n5342_, new_n5343_, new_n5344_, new_n5345_, new_n5346_,
    new_n5347_, new_n5348_, new_n5349_, new_n5350_, new_n5351_, new_n5352_,
    new_n5353_, new_n5354_, new_n5355_, new_n5356_, new_n5357_, new_n5358_,
    new_n5359_, new_n5360_, new_n5361_, new_n5362_, new_n5363_, new_n5364_,
    new_n5365_, new_n5366_, new_n5367_, new_n5368_, new_n5369_, new_n5370_,
    new_n5372_, new_n5373_, new_n5374_, new_n5375_, new_n5376_, new_n5377_,
    new_n5378_, new_n5379_, new_n5380_, new_n5381_, new_n5382_, new_n5383_,
    new_n5384_, new_n5385_, new_n5386_, new_n5387_, new_n5388_, new_n5389_,
    new_n5390_, new_n5391_, new_n5392_, new_n5393_, new_n5394_, new_n5395_,
    new_n5396_, new_n5397_, new_n5398_, new_n5399_, new_n5400_, new_n5401_,
    new_n5402_, new_n5403_, new_n5404_, new_n5405_, new_n5406_, new_n5407_,
    new_n5408_, new_n5409_, new_n5410_, new_n5411_, new_n5412_, new_n5413_,
    new_n5414_, new_n5416_, new_n5417_, new_n5418_, new_n5419_, new_n5420_,
    new_n5421_, new_n5422_, new_n5423_, new_n5424_, new_n5425_, new_n5426_,
    new_n5427_, new_n5428_, new_n5429_, new_n5430_, new_n5431_, new_n5432_,
    new_n5433_, new_n5434_, new_n5435_, new_n5436_, new_n5437_, new_n5438_,
    new_n5439_, new_n5440_, new_n5441_, new_n5442_, new_n5443_, new_n5444_,
    new_n5445_, new_n5446_, new_n5447_, new_n5448_, new_n5449_, new_n5450_,
    new_n5451_, new_n5452_, new_n5453_, new_n5454_, new_n5455_, new_n5456_,
    new_n5457_, new_n5458_, new_n5460_, new_n5461_, new_n5462_, new_n5463_,
    new_n5464_, new_n5465_, new_n5466_, new_n5467_, new_n5468_, new_n5469_,
    new_n5470_, new_n5471_, new_n5472_, new_n5473_, new_n5474_, new_n5475_,
    new_n5476_, new_n5477_, new_n5478_, new_n5479_, new_n5480_, new_n5481_,
    new_n5482_, new_n5483_, new_n5484_, new_n5485_, new_n5486_, new_n5487_,
    new_n5488_, new_n5489_, new_n5490_, new_n5491_, new_n5492_, new_n5493_,
    new_n5494_, new_n5495_, new_n5496_, new_n5497_, new_n5498_, new_n5499_,
    new_n5500_, new_n5501_, new_n5502_, new_n5504_, new_n5505_, new_n5506_,
    new_n5507_, new_n5508_, new_n5509_, new_n5510_, new_n5511_, new_n5512_,
    new_n5513_, new_n5514_, new_n5515_, new_n5516_, new_n5517_, new_n5518_,
    new_n5519_, new_n5520_, new_n5521_, new_n5522_, new_n5523_, new_n5524_,
    new_n5525_, new_n5526_, new_n5527_, new_n5528_, new_n5529_, new_n5530_,
    new_n5531_, new_n5532_, new_n5533_, new_n5534_, new_n5535_, new_n5536_,
    new_n5537_, new_n5538_, new_n5539_, new_n5540_, new_n5541_, new_n5542_,
    new_n5543_, new_n5544_, new_n5545_, new_n5546_, new_n5548_, new_n5549_,
    new_n5550_, new_n5551_, new_n5552_, new_n5553_, new_n5554_, new_n5555_,
    new_n5556_, new_n5557_, new_n5558_, new_n5559_, new_n5560_, new_n5561_,
    new_n5562_, new_n5563_, new_n5564_, new_n5565_, new_n5566_, new_n5567_,
    new_n5568_, new_n5569_, new_n5570_, new_n5571_, new_n5572_, new_n5573_,
    new_n5574_, new_n5575_, new_n5576_, new_n5577_, new_n5578_, new_n5579_,
    new_n5580_, new_n5581_, new_n5582_, new_n5583_, new_n5584_, new_n5585_,
    new_n5586_, new_n5587_, new_n5588_, new_n5589_, new_n5590_, new_n5592_,
    new_n5593_, new_n5594_, new_n5595_, new_n5596_, new_n5597_, new_n5598_,
    new_n5599_, new_n5600_, new_n5601_, new_n5602_, new_n5603_, new_n5604_,
    new_n5605_, new_n5606_, new_n5607_, new_n5608_, new_n5609_, new_n5610_,
    new_n5611_, new_n5612_, new_n5613_, new_n5614_, new_n5615_, new_n5616_,
    new_n5617_, new_n5618_, new_n5619_, new_n5620_, new_n5621_, new_n5622_,
    new_n5623_, new_n5624_, new_n5625_, new_n5626_, new_n5627_, new_n5628_,
    new_n5629_, new_n5630_, new_n5631_, new_n5632_, new_n5633_, new_n5634_,
    new_n5636_, new_n5637_, new_n5638_, new_n5639_, new_n5640_, new_n5641_,
    new_n5642_, new_n5643_, new_n5644_, new_n5645_, new_n5646_, new_n5647_,
    new_n5648_, new_n5649_, new_n5650_, new_n5651_, new_n5652_, new_n5653_,
    new_n5654_, new_n5655_, new_n5656_, new_n5657_, new_n5658_, new_n5659_,
    new_n5660_, new_n5661_, new_n5662_, new_n5663_, new_n5664_, new_n5665_,
    new_n5666_, new_n5667_, new_n5668_, new_n5669_, new_n5670_, new_n5671_,
    new_n5672_, new_n5673_, new_n5674_, new_n5675_, new_n5676_, new_n5677_,
    new_n5678_, new_n5680_, new_n5681_, new_n5682_, new_n5683_, new_n5684_,
    new_n5685_, new_n5686_, new_n5687_, new_n5688_, new_n5689_, new_n5690_,
    new_n5691_, new_n5692_, new_n5693_, new_n5694_, new_n5695_, new_n5696_,
    new_n5697_, new_n5698_, new_n5699_, new_n5700_, new_n5701_, new_n5702_,
    new_n5703_, new_n5704_, new_n5705_, new_n5706_, new_n5707_, new_n5708_,
    new_n5709_, new_n5710_, new_n5711_, new_n5712_, new_n5713_, new_n5714_,
    new_n5715_, new_n5716_, new_n5717_, new_n5718_, new_n5719_, new_n5720_,
    new_n5721_, new_n5722_, new_n5724_, new_n5725_, new_n5726_, new_n5727_,
    new_n5728_, new_n5729_, new_n5730_, new_n5731_, new_n5732_, new_n5733_,
    new_n5734_, new_n5735_, new_n5736_, new_n5737_, new_n5738_, new_n5739_,
    new_n5740_, new_n5741_, new_n5742_, new_n5743_, new_n5744_, new_n5745_,
    new_n5746_, new_n5747_, new_n5748_, new_n5749_, new_n5750_, new_n5751_,
    new_n5752_, new_n5753_, new_n5754_, new_n5755_, new_n5756_, new_n5757_,
    new_n5758_, new_n5759_, new_n5760_, new_n5761_, new_n5762_, new_n5763_,
    new_n5764_, new_n5765_, new_n5766_, new_n5768_, new_n5769_, new_n5770_,
    new_n5771_, new_n5772_, new_n5773_, new_n5774_, new_n5775_, new_n5776_,
    new_n5777_, new_n5778_, new_n5779_, new_n5780_, new_n5781_, new_n5782_,
    new_n5783_, new_n5784_, new_n5785_, new_n5786_, new_n5787_, new_n5788_,
    new_n5789_, new_n5790_, new_n5791_, new_n5792_, new_n5793_, new_n5794_,
    new_n5795_, new_n5796_, new_n5797_, new_n5798_, new_n5799_, new_n5800_,
    new_n5801_, new_n5802_, new_n5803_, new_n5804_, new_n5805_, new_n5806_,
    new_n5807_, new_n5808_, new_n5809_, new_n5810_, new_n5812_, new_n5813_,
    new_n5814_, new_n5815_, new_n5816_, new_n5817_, new_n5818_, new_n5819_,
    new_n5820_, new_n5821_, new_n5822_, new_n5823_, new_n5824_, new_n5825_,
    new_n5826_, new_n5827_, new_n5828_, new_n5829_, new_n5830_, new_n5831_,
    new_n5832_, new_n5833_, new_n5834_, new_n5835_, new_n5836_, new_n5837_,
    new_n5838_, new_n5839_, new_n5840_, new_n5841_, new_n5842_, new_n5843_,
    new_n5844_, new_n5845_, new_n5846_, new_n5847_, new_n5848_, new_n5849_,
    new_n5850_, new_n5851_, new_n5852_, new_n5853_, new_n5854_, new_n5856_,
    new_n5857_, new_n5858_, new_n5859_, new_n5860_, new_n5861_, new_n5862_,
    new_n5863_, new_n5864_, new_n5865_, new_n5866_, new_n5867_, new_n5868_,
    new_n5869_, new_n5870_, new_n5871_, new_n5872_, new_n5873_, new_n5874_,
    new_n5875_, new_n5876_, new_n5877_, new_n5878_, new_n5879_, new_n5880_,
    new_n5881_, new_n5882_, new_n5883_, new_n5884_, new_n5885_, new_n5886_,
    new_n5887_, new_n5888_, new_n5889_, new_n5890_, new_n5891_, new_n5892_,
    new_n5893_, new_n5894_, new_n5895_, new_n5896_, new_n5897_, new_n5898_,
    new_n5900_, new_n5901_, new_n5902_, new_n5903_, new_n5904_, new_n5905_,
    new_n5906_, new_n5907_, new_n5908_, new_n5909_, new_n5910_, new_n5911_,
    new_n5912_, new_n5913_, new_n5914_, new_n5915_, new_n5916_, new_n5917_,
    new_n5918_, new_n5919_, new_n5920_, new_n5921_, new_n5922_, new_n5923_,
    new_n5924_, new_n5925_, new_n5926_, new_n5927_, new_n5928_, new_n5929_,
    new_n5930_, new_n5931_, new_n5932_, new_n5933_, new_n5934_, new_n5935_,
    new_n5936_, new_n5937_, new_n5938_, new_n5939_, new_n5940_, new_n5941_,
    new_n5942_, new_n5944_, new_n5945_, new_n5946_, new_n5947_, new_n5948_,
    new_n5949_, new_n5950_, new_n5951_, new_n5952_, new_n5953_, new_n5954_,
    new_n5955_, new_n5956_, new_n5957_, new_n5958_, new_n5959_, new_n5960_,
    new_n5961_, new_n5962_, new_n5963_, new_n5964_, new_n5965_, new_n5966_,
    new_n5967_, new_n5968_, new_n5969_, new_n5970_, new_n5971_, new_n5972_,
    new_n5973_, new_n5974_, new_n5975_, new_n5976_, new_n5977_, new_n5978_,
    new_n5979_, new_n5980_, new_n5981_, new_n5982_, new_n5983_, new_n5984_,
    new_n5985_, new_n5986_, new_n5988_, new_n5989_, new_n5990_, new_n5991_,
    new_n5992_, new_n5993_, new_n5994_, new_n5995_, new_n5996_, new_n5997_,
    new_n5998_, new_n5999_, new_n6000_, new_n6001_, new_n6002_, new_n6003_,
    new_n6004_, new_n6005_, new_n6006_, new_n6007_, new_n6008_, new_n6009_,
    new_n6010_, new_n6011_, new_n6012_, new_n6013_, new_n6014_, new_n6015_,
    new_n6016_, new_n6017_, new_n6018_, new_n6019_, new_n6020_, new_n6021_,
    new_n6022_, new_n6023_, new_n6024_, new_n6025_, new_n6026_, new_n6027_,
    new_n6028_, new_n6029_, new_n6030_, new_n6032_, new_n6033_, new_n6034_,
    new_n6035_, new_n6036_, new_n6037_, new_n6038_, new_n6039_, new_n6040_,
    new_n6041_, new_n6042_, new_n6043_, new_n6044_, new_n6045_, new_n6046_,
    new_n6047_, new_n6048_, new_n6049_, new_n6050_, new_n6051_, new_n6052_,
    new_n6053_, new_n6054_, new_n6055_, new_n6056_, new_n6057_, new_n6058_,
    new_n6059_, new_n6060_, new_n6061_, new_n6062_, new_n6063_, new_n6064_,
    new_n6065_, new_n6066_, new_n6067_, new_n6068_, new_n6069_, new_n6070_,
    new_n6071_, new_n6072_, new_n6073_, new_n6074_, new_n6076_, new_n6077_,
    new_n6078_, new_n6079_, new_n6080_, new_n6081_, new_n6082_, new_n6083_,
    new_n6084_, new_n6085_, new_n6086_, new_n6087_, new_n6088_, new_n6089_,
    new_n6090_, new_n6091_, new_n6092_, new_n6093_, new_n6094_, new_n6095_,
    new_n6096_, new_n6097_, new_n6098_, new_n6099_, new_n6100_, new_n6101_,
    new_n6102_, new_n6103_, new_n6104_, new_n6105_, new_n6106_, new_n6107_,
    new_n6108_, new_n6109_, new_n6110_, new_n6111_, new_n6112_, new_n6113_,
    new_n6114_, new_n6115_, new_n6116_, new_n6117_, new_n6118_, new_n6120_,
    new_n6121_, new_n6122_, new_n6123_, new_n6124_, new_n6125_, new_n6126_,
    new_n6127_, new_n6128_, new_n6129_, new_n6130_, new_n6131_, new_n6132_,
    new_n6133_, new_n6134_, new_n6135_, new_n6136_, new_n6137_, new_n6138_,
    new_n6139_, new_n6140_, new_n6141_, new_n6142_, new_n6143_, new_n6144_,
    new_n6145_, new_n6146_, new_n6147_, new_n6148_, new_n6149_, new_n6150_,
    new_n6151_, new_n6152_, new_n6153_, new_n6154_, new_n6155_, new_n6156_,
    new_n6157_, new_n6158_, new_n6159_, new_n6160_, new_n6161_, new_n6162_,
    new_n6164_, new_n6165_, new_n6166_, new_n6167_, new_n6168_, new_n6169_,
    new_n6170_, new_n6171_, new_n6172_, new_n6173_, new_n6174_, new_n6175_,
    new_n6176_, new_n6177_, new_n6178_, new_n6179_, new_n6180_, new_n6181_,
    new_n6182_, new_n6183_, new_n6184_, new_n6185_, new_n6186_, new_n6187_,
    new_n6188_, new_n6189_, new_n6190_, new_n6191_, new_n6192_, new_n6193_,
    new_n6194_, new_n6195_, new_n6196_, new_n6197_, new_n6198_, new_n6199_,
    new_n6200_, new_n6201_, new_n6202_, new_n6203_, new_n6204_, new_n6205_,
    new_n6206_, new_n6208_, new_n6209_, new_n6210_, new_n6211_, new_n6212_,
    new_n6213_, new_n6214_, new_n6215_, new_n6216_, new_n6217_, new_n6218_,
    new_n6219_, new_n6220_, new_n6221_, new_n6222_, new_n6223_, new_n6224_,
    new_n6225_, new_n6226_, new_n6227_, new_n6228_, new_n6229_, new_n6230_,
    new_n6231_, new_n6232_, new_n6233_, new_n6234_, new_n6235_, new_n6236_,
    new_n6237_, new_n6238_, new_n6239_, new_n6240_, new_n6241_, new_n6242_,
    new_n6243_, new_n6244_, new_n6245_, new_n6246_, new_n6247_, new_n6248_,
    new_n6249_, new_n6250_, new_n6252_, new_n6253_, new_n6254_, new_n6255_,
    new_n6256_, new_n6257_, new_n6258_, new_n6259_, new_n6260_, new_n6261_,
    new_n6262_, new_n6263_, new_n6264_, new_n6265_, new_n6266_, new_n6267_,
    new_n6268_, new_n6269_, new_n6270_, new_n6271_, new_n6272_, new_n6273_,
    new_n6274_, new_n6275_, new_n6276_, new_n6277_, new_n6278_, new_n6279_,
    new_n6280_, new_n6281_, new_n6282_, new_n6283_, new_n6284_, new_n6285_,
    new_n6286_, new_n6287_, new_n6288_, new_n6289_, new_n6290_, new_n6291_,
    new_n6292_, new_n6293_, new_n6294_, new_n6296_, new_n6297_, new_n6298_,
    new_n6299_, new_n6300_, new_n6301_, new_n6302_, new_n6303_, new_n6304_,
    new_n6305_, new_n6306_, new_n6307_, new_n6308_, new_n6309_, new_n6310_,
    new_n6311_, new_n6312_, new_n6313_, new_n6314_, new_n6315_, new_n6316_,
    new_n6317_, new_n6318_, new_n6319_, new_n6320_, new_n6321_, new_n6322_,
    new_n6323_, new_n6324_, new_n6325_, new_n6326_, new_n6327_, new_n6328_,
    new_n6329_, new_n6330_, new_n6331_, new_n6332_, new_n6333_, new_n6334_,
    new_n6335_, new_n6336_, new_n6337_, new_n6338_, new_n6340_, new_n6341_,
    new_n6342_, new_n6343_, new_n6344_, new_n6345_, new_n6346_, new_n6347_,
    new_n6348_, new_n6349_, new_n6350_, new_n6351_, new_n6352_, new_n6353_,
    new_n6354_, new_n6355_, new_n6356_, new_n6357_, new_n6358_, new_n6359_,
    new_n6360_, new_n6361_, new_n6362_, new_n6363_, new_n6364_, new_n6365_,
    new_n6366_, new_n6367_, new_n6368_, new_n6369_, new_n6370_, new_n6371_,
    new_n6372_, new_n6373_, new_n6374_, new_n6375_, new_n6376_, new_n6377_,
    new_n6378_, new_n6379_, new_n6380_, new_n6381_, new_n6382_, new_n6384_,
    new_n6385_, new_n6386_, new_n6387_, new_n6388_, new_n6389_, new_n6390_,
    new_n6391_, new_n6392_, new_n6393_, new_n6394_, new_n6395_, new_n6396_,
    new_n6397_, new_n6398_, new_n6399_, new_n6400_, new_n6401_, new_n6402_,
    new_n6403_, new_n6404_, new_n6405_, new_n6406_, new_n6407_, new_n6408_,
    new_n6409_, new_n6410_, new_n6411_, new_n6412_, new_n6413_, new_n6414_,
    new_n6415_, new_n6416_, new_n6417_, new_n6418_, new_n6419_, new_n6420_,
    new_n6421_, new_n6422_, new_n6423_, new_n6424_, new_n6425_, new_n6426_,
    new_n6428_, new_n6429_, new_n6430_, new_n6431_, new_n6432_, new_n6433_,
    new_n6434_, new_n6435_, new_n6436_, new_n6437_, new_n6438_, new_n6439_,
    new_n6440_, new_n6441_, new_n6442_, new_n6443_, new_n6444_, new_n6445_,
    new_n6446_, new_n6447_, new_n6448_, new_n6449_, new_n6450_, new_n6451_,
    new_n6452_, new_n6453_, new_n6454_, new_n6455_, new_n6456_, new_n6457_,
    new_n6458_, new_n6459_, new_n6460_, new_n6461_, new_n6462_, new_n6463_,
    new_n6464_, new_n6465_, new_n6466_, new_n6467_, new_n6468_, new_n6469_,
    new_n6470_, new_n6472_, new_n6473_, new_n6474_, new_n6475_, new_n6476_,
    new_n6477_, new_n6478_, new_n6479_, new_n6480_, new_n6481_, new_n6482_,
    new_n6483_, new_n6484_, new_n6485_, new_n6486_, new_n6487_, new_n6488_,
    new_n6489_, new_n6490_, new_n6491_, new_n6492_, new_n6493_, new_n6494_,
    new_n6495_, new_n6496_, new_n6497_, new_n6498_, new_n6499_, new_n6500_,
    new_n6501_, new_n6502_, new_n6503_, new_n6504_, new_n6505_, new_n6506_,
    new_n6507_, new_n6508_, new_n6509_, new_n6510_, new_n6511_, new_n6512_,
    new_n6513_, new_n6514_, new_n6516_, new_n6517_, new_n6518_, new_n6519_,
    new_n6520_, new_n6521_, new_n6522_, new_n6523_, new_n6524_, new_n6525_,
    new_n6526_, new_n6527_, new_n6528_, new_n6529_, new_n6530_, new_n6531_,
    new_n6532_, new_n6533_, new_n6534_, new_n6535_, new_n6536_, new_n6537_,
    new_n6538_, new_n6539_, new_n6540_, new_n6541_, new_n6542_, new_n6543_,
    new_n6544_, new_n6545_, new_n6546_, new_n6547_, new_n6548_, new_n6549_,
    new_n6550_, new_n6551_, new_n6552_, new_n6553_, new_n6554_, new_n6555_,
    new_n6556_, new_n6557_, new_n6558_, new_n6560_, new_n6561_, new_n6562_,
    new_n6563_, new_n6564_, new_n6565_, new_n6566_, new_n6567_, new_n6568_,
    new_n6569_, new_n6570_, new_n6571_, new_n6572_, new_n6573_, new_n6574_,
    new_n6575_, new_n6576_, new_n6577_, new_n6578_, new_n6579_, new_n6580_,
    new_n6581_, new_n6582_, new_n6583_, new_n6584_, new_n6585_, new_n6586_,
    new_n6587_, new_n6588_, new_n6589_, new_n6590_, new_n6591_, new_n6592_,
    new_n6593_, new_n6594_, new_n6595_, new_n6596_, new_n6597_, new_n6598_,
    new_n6599_, new_n6600_, new_n6601_, new_n6602_, new_n6604_, new_n6605_,
    new_n6606_, new_n6607_, new_n6608_, new_n6609_, new_n6610_, new_n6611_,
    new_n6612_, new_n6613_, new_n6614_, new_n6615_, new_n6616_, new_n6617_,
    new_n6618_, new_n6619_, new_n6620_, new_n6621_, new_n6622_, new_n6623_,
    new_n6624_, new_n6625_, new_n6626_, new_n6627_, new_n6628_, new_n6629_,
    new_n6630_, new_n6631_, new_n6632_, new_n6633_, new_n6634_, new_n6635_,
    new_n6636_, new_n6637_, new_n6638_, new_n6639_, new_n6640_, new_n6641_,
    new_n6642_, new_n6643_, new_n6644_, new_n6645_, new_n6646_, new_n6648_,
    new_n6649_, new_n6650_, new_n6651_, new_n6652_, new_n6653_, new_n6654_,
    new_n6655_, new_n6656_, new_n6657_, new_n6658_, new_n6659_, new_n6660_,
    new_n6661_, new_n6662_, new_n6663_, new_n6664_, new_n6665_, new_n6666_,
    new_n6667_, new_n6668_, new_n6669_, new_n6670_, new_n6671_, new_n6672_,
    new_n6673_, new_n6674_, new_n6675_, new_n6676_, new_n6677_, new_n6678_,
    new_n6679_, new_n6680_, new_n6681_, new_n6682_, new_n6683_, new_n6684_,
    new_n6685_, new_n6686_, new_n6687_, new_n6688_, new_n6689_, new_n6690_,
    new_n6692_, new_n6693_, new_n6694_, new_n6695_, new_n6696_, new_n6697_,
    new_n6698_, new_n6699_, new_n6700_, new_n6701_, new_n6702_, new_n6703_,
    new_n6704_, new_n6705_, new_n6706_, new_n6707_, new_n6708_, new_n6709_,
    new_n6710_, new_n6711_, new_n6712_, new_n6713_, new_n6714_, new_n6715_,
    new_n6716_, new_n6717_, new_n6718_, new_n6719_, new_n6720_, new_n6721_,
    new_n6722_, new_n6723_, new_n6724_, new_n6725_, new_n6726_, new_n6727_,
    new_n6728_, new_n6729_, new_n6730_, new_n6731_, new_n6732_, new_n6733_,
    new_n6734_, new_n6736_, new_n6737_, new_n6738_, new_n6739_, new_n6740_,
    new_n6741_, new_n6742_, new_n6743_, new_n6744_, new_n6745_, new_n6746_,
    new_n6747_, new_n6748_, new_n6749_, new_n6750_, new_n6751_, new_n6752_,
    new_n6753_, new_n6754_, new_n6755_, new_n6756_, new_n6757_, new_n6758_,
    new_n6759_, new_n6760_, new_n6761_, new_n6762_, new_n6763_, new_n6764_,
    new_n6765_, new_n6766_, new_n6767_, new_n6768_, new_n6769_, new_n6770_,
    new_n6771_, new_n6772_, new_n6773_, new_n6774_, new_n6775_, new_n6776_,
    new_n6777_, new_n6778_, new_n6780_, new_n6781_, new_n6782_, new_n6783_,
    new_n6784_, new_n6785_, new_n6786_, new_n6787_, new_n6788_, new_n6789_,
    new_n6790_, new_n6791_, new_n6792_, new_n6793_, new_n6794_, new_n6795_,
    new_n6796_, new_n6797_, new_n6798_, new_n6799_, new_n6800_, new_n6801_,
    new_n6802_, new_n6803_, new_n6804_, new_n6805_, new_n6806_, new_n6807_,
    new_n6808_, new_n6809_, new_n6810_, new_n6811_, new_n6812_, new_n6813_,
    new_n6814_, new_n6815_, new_n6816_, new_n6817_, new_n6818_, new_n6819_,
    new_n6820_, new_n6821_, new_n6822_, new_n6824_, new_n6825_, new_n6826_,
    new_n6827_, new_n6828_, new_n6829_, new_n6830_, new_n6831_, new_n6832_,
    new_n6833_, new_n6834_, new_n6835_, new_n6836_, new_n6837_, new_n6838_,
    new_n6839_, new_n6840_, new_n6841_, new_n6842_, new_n6843_, new_n6844_,
    new_n6845_, new_n6846_, new_n6847_, new_n6848_, new_n6849_, new_n6850_,
    new_n6851_, new_n6852_, new_n6853_, new_n6854_, new_n6855_, new_n6856_,
    new_n6857_, new_n6858_, new_n6859_, new_n6860_, new_n6861_, new_n6862_,
    new_n6863_, new_n6864_, new_n6865_, new_n6866_, new_n6868_, new_n6869_,
    new_n6870_, new_n6871_, new_n6872_, new_n6873_, new_n6874_, new_n6875_,
    new_n6876_, new_n6877_, new_n6878_, new_n6879_, new_n6880_, new_n6881_,
    new_n6882_, new_n6883_, new_n6884_, new_n6885_, new_n6886_, new_n6887_,
    new_n6888_, new_n6889_, new_n6890_, new_n6891_, new_n6892_, new_n6893_,
    new_n6894_, new_n6895_, new_n6896_, new_n6897_, new_n6898_, new_n6899_,
    new_n6900_, new_n6901_, new_n6902_, new_n6903_, new_n6904_, new_n6905_,
    new_n6906_, new_n6907_, new_n6908_, new_n6909_, new_n6910_, new_n6912_,
    new_n6913_, new_n6914_, new_n6915_, new_n6916_, new_n6917_, new_n6918_,
    new_n6919_, new_n6920_, new_n6921_, new_n6922_, new_n6923_, new_n6924_,
    new_n6925_, new_n6926_, new_n6927_, new_n6928_, new_n6929_, new_n6930_,
    new_n6931_, new_n6932_, new_n6933_, new_n6934_, new_n6935_, new_n6936_,
    new_n6937_, new_n6938_, new_n6939_, new_n6940_, new_n6941_, new_n6942_,
    new_n6943_, new_n6944_, new_n6945_, new_n6946_, new_n6947_, new_n6948_,
    new_n6949_, new_n6950_, new_n6951_, new_n6952_, new_n6953_, new_n6954_,
    new_n6956_, new_n6957_, new_n6958_, new_n6959_, new_n6960_, new_n6961_,
    new_n6962_, new_n6963_, new_n6964_, new_n6965_, new_n6966_, new_n6967_,
    new_n6968_, new_n6969_, new_n6970_, new_n6971_, new_n6972_, new_n6973_,
    new_n6974_, new_n6975_, new_n6976_, new_n6977_, new_n6978_, new_n6979_,
    new_n6980_, new_n6981_, new_n6982_, new_n6983_, new_n6984_, new_n6985_,
    new_n6986_, new_n6987_, new_n6988_, new_n6989_, new_n6990_, new_n6991_,
    new_n6992_, new_n6993_, new_n6994_, new_n6995_, new_n6996_, new_n6997_,
    new_n6998_, new_n7000_, new_n7001_, new_n7002_, new_n7003_, new_n7004_,
    new_n7005_, new_n7006_, new_n7007_, new_n7008_, new_n7009_, new_n7010_,
    new_n7011_, new_n7012_, new_n7013_, new_n7014_, new_n7015_, new_n7016_,
    new_n7017_, new_n7018_, new_n7019_, new_n7020_, new_n7021_, new_n7022_,
    new_n7023_, new_n7024_, new_n7025_, new_n7026_, new_n7027_, new_n7028_,
    new_n7029_, new_n7030_, new_n7031_, new_n7032_, new_n7033_, new_n7034_,
    new_n7035_, new_n7036_, new_n7037_, new_n7038_, new_n7039_, new_n7040_,
    new_n7041_, new_n7042_, new_n7044_, new_n7045_, new_n7046_, new_n7047_,
    new_n7048_, new_n7049_, new_n7050_, new_n7051_, new_n7052_, new_n7053_,
    new_n7054_, new_n7055_, new_n7056_, new_n7057_, new_n7058_, new_n7059_,
    new_n7060_, new_n7061_, new_n7062_, new_n7063_, new_n7064_, new_n7065_,
    new_n7066_, new_n7067_, new_n7068_, new_n7069_, new_n7070_, new_n7071_,
    new_n7072_, new_n7073_, new_n7074_, new_n7075_, new_n7076_, new_n7077_,
    new_n7078_, new_n7079_, new_n7080_, new_n7081_, new_n7082_, new_n7083_;
  INVX1    g0000(.A(\priority[1] ), .Y(new_n386_));
  INVX1    g0001(.A(\priority[2] ), .Y(new_n387_));
  OAI21X1  g0002(.A0(\req[1] ), .A1(new_n386_), .B0(new_n387_), .Y(new_n388_));
  NOR2X1   g0003(.A(\req[3] ), .B(\req[2] ), .Y(new_n389_));
  AND2X1   g0004(.A(new_n389_), .B(new_n388_), .Y(new_n390_));
  INVX1    g0005(.A(\priority[5] ), .Y(new_n391_));
  INVX1    g0006(.A(\req[3] ), .Y(new_n392_));
  AOI21X1  g0007(.A0(new_n392_), .A1(\priority[3] ), .B0(\priority[4] ), .Y(new_n393_));
  NAND2X1  g0008(.A(new_n393_), .B(new_n391_), .Y(new_n394_));
  OR2X1    g0009(.A(\req[6] ), .B(\req[5] ), .Y(new_n395_));
  AOI21X1  g0010(.A0(\req[4] ), .A1(new_n391_), .B0(new_n395_), .Y(new_n396_));
  OAI21X1  g0011(.A0(new_n394_), .A1(new_n390_), .B0(new_n396_), .Y(new_n397_));
  INVX1    g0012(.A(\priority[8] ), .Y(new_n398_));
  INVX1    g0013(.A(\req[6] ), .Y(new_n399_));
  AOI21X1  g0014(.A0(new_n399_), .A1(\priority[6] ), .B0(\priority[7] ), .Y(new_n400_));
  AND2X1   g0015(.A(new_n400_), .B(new_n398_), .Y(new_n401_));
  OR2X1    g0016(.A(\req[9] ), .B(\req[8] ), .Y(new_n402_));
  AOI21X1  g0017(.A0(\req[7] ), .A1(new_n398_), .B0(new_n402_), .Y(new_n403_));
  INVX1    g0018(.A(new_n403_), .Y(new_n404_));
  AOI21X1  g0019(.A0(new_n401_), .A1(new_n397_), .B0(new_n404_), .Y(new_n405_));
  INVX1    g0020(.A(\priority[11] ), .Y(new_n406_));
  INVX1    g0021(.A(\req[9] ), .Y(new_n407_));
  AOI21X1  g0022(.A0(new_n407_), .A1(\priority[9] ), .B0(\priority[10] ), .Y(new_n408_));
  NAND2X1  g0023(.A(new_n408_), .B(new_n406_), .Y(new_n409_));
  OR2X1    g0024(.A(\req[12] ), .B(\req[11] ), .Y(new_n410_));
  AOI21X1  g0025(.A0(\req[10] ), .A1(new_n406_), .B0(new_n410_), .Y(new_n411_));
  OAI21X1  g0026(.A0(new_n409_), .A1(new_n405_), .B0(new_n411_), .Y(new_n412_));
  INVX1    g0027(.A(\priority[14] ), .Y(new_n413_));
  INVX1    g0028(.A(\req[12] ), .Y(new_n414_));
  AOI21X1  g0029(.A0(new_n414_), .A1(\priority[12] ), .B0(\priority[13] ), .Y(new_n415_));
  AND2X1   g0030(.A(new_n415_), .B(new_n413_), .Y(new_n416_));
  OR2X1    g0031(.A(\req[15] ), .B(\req[14] ), .Y(new_n417_));
  AOI21X1  g0032(.A0(\req[13] ), .A1(new_n413_), .B0(new_n417_), .Y(new_n418_));
  INVX1    g0033(.A(new_n418_), .Y(new_n419_));
  AOI21X1  g0034(.A0(new_n416_), .A1(new_n412_), .B0(new_n419_), .Y(new_n420_));
  INVX1    g0035(.A(\priority[17] ), .Y(new_n421_));
  INVX1    g0036(.A(\req[15] ), .Y(new_n422_));
  AOI21X1  g0037(.A0(new_n422_), .A1(\priority[15] ), .B0(\priority[16] ), .Y(new_n423_));
  NAND2X1  g0038(.A(new_n423_), .B(new_n421_), .Y(new_n424_));
  OR2X1    g0039(.A(\req[18] ), .B(\req[17] ), .Y(new_n425_));
  AOI21X1  g0040(.A0(\req[16] ), .A1(new_n421_), .B0(new_n425_), .Y(new_n426_));
  OAI21X1  g0041(.A0(new_n424_), .A1(new_n420_), .B0(new_n426_), .Y(new_n427_));
  INVX1    g0042(.A(\priority[20] ), .Y(new_n428_));
  INVX1    g0043(.A(\req[18] ), .Y(new_n429_));
  AOI21X1  g0044(.A0(new_n429_), .A1(\priority[18] ), .B0(\priority[19] ), .Y(new_n430_));
  AND2X1   g0045(.A(new_n430_), .B(new_n428_), .Y(new_n431_));
  OR2X1    g0046(.A(\req[21] ), .B(\req[20] ), .Y(new_n432_));
  AOI21X1  g0047(.A0(\req[19] ), .A1(new_n428_), .B0(new_n432_), .Y(new_n433_));
  INVX1    g0048(.A(new_n433_), .Y(new_n434_));
  AOI21X1  g0049(.A0(new_n431_), .A1(new_n427_), .B0(new_n434_), .Y(new_n435_));
  INVX1    g0050(.A(\priority[23] ), .Y(new_n436_));
  INVX1    g0051(.A(\req[21] ), .Y(new_n437_));
  AOI21X1  g0052(.A0(new_n437_), .A1(\priority[21] ), .B0(\priority[22] ), .Y(new_n438_));
  NAND2X1  g0053(.A(new_n438_), .B(new_n436_), .Y(new_n439_));
  OR2X1    g0054(.A(\req[24] ), .B(\req[23] ), .Y(new_n440_));
  AOI21X1  g0055(.A0(\req[22] ), .A1(new_n436_), .B0(new_n440_), .Y(new_n441_));
  OAI21X1  g0056(.A0(new_n439_), .A1(new_n435_), .B0(new_n441_), .Y(new_n442_));
  INVX1    g0057(.A(\priority[26] ), .Y(new_n443_));
  INVX1    g0058(.A(\req[24] ), .Y(new_n444_));
  AOI21X1  g0059(.A0(new_n444_), .A1(\priority[24] ), .B0(\priority[25] ), .Y(new_n445_));
  AND2X1   g0060(.A(new_n445_), .B(new_n443_), .Y(new_n446_));
  OR2X1    g0061(.A(\req[27] ), .B(\req[26] ), .Y(new_n447_));
  AOI21X1  g0062(.A0(\req[25] ), .A1(new_n443_), .B0(new_n447_), .Y(new_n448_));
  INVX1    g0063(.A(new_n448_), .Y(new_n449_));
  AOI21X1  g0064(.A0(new_n446_), .A1(new_n442_), .B0(new_n449_), .Y(new_n450_));
  INVX1    g0065(.A(\priority[29] ), .Y(new_n451_));
  INVX1    g0066(.A(\req[27] ), .Y(new_n452_));
  AOI21X1  g0067(.A0(new_n452_), .A1(\priority[27] ), .B0(\priority[28] ), .Y(new_n453_));
  NAND2X1  g0068(.A(new_n453_), .B(new_n451_), .Y(new_n454_));
  OR2X1    g0069(.A(\req[30] ), .B(\req[29] ), .Y(new_n455_));
  AOI21X1  g0070(.A0(\req[28] ), .A1(new_n451_), .B0(new_n455_), .Y(new_n456_));
  OAI21X1  g0071(.A0(new_n454_), .A1(new_n450_), .B0(new_n456_), .Y(new_n457_));
  INVX1    g0072(.A(\priority[32] ), .Y(new_n458_));
  INVX1    g0073(.A(\req[30] ), .Y(new_n459_));
  AOI21X1  g0074(.A0(new_n459_), .A1(\priority[30] ), .B0(\priority[31] ), .Y(new_n460_));
  AND2X1   g0075(.A(new_n460_), .B(new_n458_), .Y(new_n461_));
  OR2X1    g0076(.A(\req[33] ), .B(\req[32] ), .Y(new_n462_));
  AOI21X1  g0077(.A0(\req[31] ), .A1(new_n458_), .B0(new_n462_), .Y(new_n463_));
  INVX1    g0078(.A(new_n463_), .Y(new_n464_));
  AOI21X1  g0079(.A0(new_n461_), .A1(new_n457_), .B0(new_n464_), .Y(new_n465_));
  INVX1    g0080(.A(\priority[35] ), .Y(new_n466_));
  INVX1    g0081(.A(\req[33] ), .Y(new_n467_));
  AOI21X1  g0082(.A0(new_n467_), .A1(\priority[33] ), .B0(\priority[34] ), .Y(new_n468_));
  NAND2X1  g0083(.A(new_n468_), .B(new_n466_), .Y(new_n469_));
  OR2X1    g0084(.A(\req[36] ), .B(\req[35] ), .Y(new_n470_));
  AOI21X1  g0085(.A0(\req[34] ), .A1(new_n466_), .B0(new_n470_), .Y(new_n471_));
  OAI21X1  g0086(.A0(new_n469_), .A1(new_n465_), .B0(new_n471_), .Y(new_n472_));
  INVX1    g0087(.A(\priority[38] ), .Y(new_n473_));
  INVX1    g0088(.A(\req[36] ), .Y(new_n474_));
  AOI21X1  g0089(.A0(new_n474_), .A1(\priority[36] ), .B0(\priority[37] ), .Y(new_n475_));
  AND2X1   g0090(.A(new_n475_), .B(new_n473_), .Y(new_n476_));
  OR2X1    g0091(.A(\req[39] ), .B(\req[38] ), .Y(new_n477_));
  AOI21X1  g0092(.A0(\req[37] ), .A1(new_n473_), .B0(new_n477_), .Y(new_n478_));
  INVX1    g0093(.A(new_n478_), .Y(new_n479_));
  AOI21X1  g0094(.A0(new_n476_), .A1(new_n472_), .B0(new_n479_), .Y(new_n480_));
  INVX1    g0095(.A(\priority[41] ), .Y(new_n481_));
  INVX1    g0096(.A(\req[39] ), .Y(new_n482_));
  AOI21X1  g0097(.A0(new_n482_), .A1(\priority[39] ), .B0(\priority[40] ), .Y(new_n483_));
  NAND2X1  g0098(.A(new_n483_), .B(new_n481_), .Y(new_n484_));
  OR2X1    g0099(.A(\req[42] ), .B(\req[41] ), .Y(new_n485_));
  AOI21X1  g0100(.A0(\req[40] ), .A1(new_n481_), .B0(new_n485_), .Y(new_n486_));
  OAI21X1  g0101(.A0(new_n484_), .A1(new_n480_), .B0(new_n486_), .Y(new_n487_));
  INVX1    g0102(.A(\priority[44] ), .Y(new_n488_));
  INVX1    g0103(.A(\req[42] ), .Y(new_n489_));
  AOI21X1  g0104(.A0(new_n489_), .A1(\priority[42] ), .B0(\priority[43] ), .Y(new_n490_));
  AND2X1   g0105(.A(new_n490_), .B(new_n488_), .Y(new_n491_));
  OR2X1    g0106(.A(\req[45] ), .B(\req[44] ), .Y(new_n492_));
  AOI21X1  g0107(.A0(\req[43] ), .A1(new_n488_), .B0(new_n492_), .Y(new_n493_));
  INVX1    g0108(.A(new_n493_), .Y(new_n494_));
  AOI21X1  g0109(.A0(new_n491_), .A1(new_n487_), .B0(new_n494_), .Y(new_n495_));
  INVX1    g0110(.A(\priority[47] ), .Y(new_n496_));
  INVX1    g0111(.A(\req[45] ), .Y(new_n497_));
  AOI21X1  g0112(.A0(new_n497_), .A1(\priority[45] ), .B0(\priority[46] ), .Y(new_n498_));
  NAND2X1  g0113(.A(new_n498_), .B(new_n496_), .Y(new_n499_));
  OR2X1    g0114(.A(\req[48] ), .B(\req[47] ), .Y(new_n500_));
  AOI21X1  g0115(.A0(\req[46] ), .A1(new_n496_), .B0(new_n500_), .Y(new_n501_));
  OAI21X1  g0116(.A0(new_n499_), .A1(new_n495_), .B0(new_n501_), .Y(new_n502_));
  INVX1    g0117(.A(\priority[50] ), .Y(new_n503_));
  INVX1    g0118(.A(\req[48] ), .Y(new_n504_));
  AOI21X1  g0119(.A0(new_n504_), .A1(\priority[48] ), .B0(\priority[49] ), .Y(new_n505_));
  AND2X1   g0120(.A(new_n505_), .B(new_n503_), .Y(new_n506_));
  OR2X1    g0121(.A(\req[51] ), .B(\req[50] ), .Y(new_n507_));
  AOI21X1  g0122(.A0(\req[49] ), .A1(new_n503_), .B0(new_n507_), .Y(new_n508_));
  INVX1    g0123(.A(new_n508_), .Y(new_n509_));
  AOI21X1  g0124(.A0(new_n506_), .A1(new_n502_), .B0(new_n509_), .Y(new_n510_));
  INVX1    g0125(.A(\priority[53] ), .Y(new_n511_));
  INVX1    g0126(.A(\req[51] ), .Y(new_n512_));
  AOI21X1  g0127(.A0(new_n512_), .A1(\priority[51] ), .B0(\priority[52] ), .Y(new_n513_));
  NAND2X1  g0128(.A(new_n513_), .B(new_n511_), .Y(new_n514_));
  OR2X1    g0129(.A(\req[54] ), .B(\req[53] ), .Y(new_n515_));
  AOI21X1  g0130(.A0(\req[52] ), .A1(new_n511_), .B0(new_n515_), .Y(new_n516_));
  OAI21X1  g0131(.A0(new_n514_), .A1(new_n510_), .B0(new_n516_), .Y(new_n517_));
  INVX1    g0132(.A(\priority[56] ), .Y(new_n518_));
  INVX1    g0133(.A(\req[54] ), .Y(new_n519_));
  AOI21X1  g0134(.A0(new_n519_), .A1(\priority[54] ), .B0(\priority[55] ), .Y(new_n520_));
  AND2X1   g0135(.A(new_n520_), .B(new_n518_), .Y(new_n521_));
  OR2X1    g0136(.A(\req[57] ), .B(\req[56] ), .Y(new_n522_));
  AOI21X1  g0137(.A0(\req[55] ), .A1(new_n518_), .B0(new_n522_), .Y(new_n523_));
  INVX1    g0138(.A(new_n523_), .Y(new_n524_));
  AOI21X1  g0139(.A0(new_n521_), .A1(new_n517_), .B0(new_n524_), .Y(new_n525_));
  INVX1    g0140(.A(\priority[59] ), .Y(new_n526_));
  INVX1    g0141(.A(\req[57] ), .Y(new_n527_));
  AOI21X1  g0142(.A0(new_n527_), .A1(\priority[57] ), .B0(\priority[58] ), .Y(new_n528_));
  NAND2X1  g0143(.A(new_n528_), .B(new_n526_), .Y(new_n529_));
  OR2X1    g0144(.A(\req[60] ), .B(\req[59] ), .Y(new_n530_));
  AOI21X1  g0145(.A0(\req[58] ), .A1(new_n526_), .B0(new_n530_), .Y(new_n531_));
  OAI21X1  g0146(.A0(new_n529_), .A1(new_n525_), .B0(new_n531_), .Y(new_n532_));
  INVX1    g0147(.A(\priority[62] ), .Y(new_n533_));
  INVX1    g0148(.A(\req[60] ), .Y(new_n534_));
  AOI21X1  g0149(.A0(new_n534_), .A1(\priority[60] ), .B0(\priority[61] ), .Y(new_n535_));
  AND2X1   g0150(.A(new_n535_), .B(new_n533_), .Y(new_n536_));
  OR2X1    g0151(.A(\req[63] ), .B(\req[62] ), .Y(new_n537_));
  AOI21X1  g0152(.A0(\req[61] ), .A1(new_n533_), .B0(new_n537_), .Y(new_n538_));
  INVX1    g0153(.A(new_n538_), .Y(new_n539_));
  AOI21X1  g0154(.A0(new_n536_), .A1(new_n532_), .B0(new_n539_), .Y(new_n540_));
  INVX1    g0155(.A(\priority[65] ), .Y(new_n541_));
  INVX1    g0156(.A(\req[63] ), .Y(new_n542_));
  AOI21X1  g0157(.A0(new_n542_), .A1(\priority[63] ), .B0(\priority[64] ), .Y(new_n543_));
  NAND2X1  g0158(.A(new_n543_), .B(new_n541_), .Y(new_n544_));
  OR2X1    g0159(.A(\req[66] ), .B(\req[65] ), .Y(new_n545_));
  AOI21X1  g0160(.A0(\req[64] ), .A1(new_n541_), .B0(new_n545_), .Y(new_n546_));
  OAI21X1  g0161(.A0(new_n544_), .A1(new_n540_), .B0(new_n546_), .Y(new_n547_));
  INVX1    g0162(.A(\priority[68] ), .Y(new_n548_));
  INVX1    g0163(.A(\req[66] ), .Y(new_n549_));
  AOI21X1  g0164(.A0(new_n549_), .A1(\priority[66] ), .B0(\priority[67] ), .Y(new_n550_));
  AND2X1   g0165(.A(new_n550_), .B(new_n548_), .Y(new_n551_));
  OR2X1    g0166(.A(\req[69] ), .B(\req[68] ), .Y(new_n552_));
  AOI21X1  g0167(.A0(\req[67] ), .A1(new_n548_), .B0(new_n552_), .Y(new_n553_));
  INVX1    g0168(.A(new_n553_), .Y(new_n554_));
  AOI21X1  g0169(.A0(new_n551_), .A1(new_n547_), .B0(new_n554_), .Y(new_n555_));
  INVX1    g0170(.A(\priority[71] ), .Y(new_n556_));
  INVX1    g0171(.A(\req[69] ), .Y(new_n557_));
  AOI21X1  g0172(.A0(new_n557_), .A1(\priority[69] ), .B0(\priority[70] ), .Y(new_n558_));
  NAND2X1  g0173(.A(new_n558_), .B(new_n556_), .Y(new_n559_));
  OR2X1    g0174(.A(\req[72] ), .B(\req[71] ), .Y(new_n560_));
  AOI21X1  g0175(.A0(\req[70] ), .A1(new_n556_), .B0(new_n560_), .Y(new_n561_));
  OAI21X1  g0176(.A0(new_n559_), .A1(new_n555_), .B0(new_n561_), .Y(new_n562_));
  INVX1    g0177(.A(\priority[74] ), .Y(new_n563_));
  INVX1    g0178(.A(\req[72] ), .Y(new_n564_));
  AOI21X1  g0179(.A0(new_n564_), .A1(\priority[72] ), .B0(\priority[73] ), .Y(new_n565_));
  AND2X1   g0180(.A(new_n565_), .B(new_n563_), .Y(new_n566_));
  OR2X1    g0181(.A(\req[75] ), .B(\req[74] ), .Y(new_n567_));
  AOI21X1  g0182(.A0(\req[73] ), .A1(new_n563_), .B0(new_n567_), .Y(new_n568_));
  INVX1    g0183(.A(new_n568_), .Y(new_n569_));
  AOI21X1  g0184(.A0(new_n566_), .A1(new_n562_), .B0(new_n569_), .Y(new_n570_));
  INVX1    g0185(.A(\priority[77] ), .Y(new_n571_));
  INVX1    g0186(.A(\req[75] ), .Y(new_n572_));
  AOI21X1  g0187(.A0(new_n572_), .A1(\priority[75] ), .B0(\priority[76] ), .Y(new_n573_));
  NAND2X1  g0188(.A(new_n573_), .B(new_n571_), .Y(new_n574_));
  OR2X1    g0189(.A(\req[78] ), .B(\req[77] ), .Y(new_n575_));
  AOI21X1  g0190(.A0(\req[76] ), .A1(new_n571_), .B0(new_n575_), .Y(new_n576_));
  OAI21X1  g0191(.A0(new_n574_), .A1(new_n570_), .B0(new_n576_), .Y(new_n577_));
  INVX1    g0192(.A(\priority[80] ), .Y(new_n578_));
  INVX1    g0193(.A(\req[78] ), .Y(new_n579_));
  AOI21X1  g0194(.A0(new_n579_), .A1(\priority[78] ), .B0(\priority[79] ), .Y(new_n580_));
  AND2X1   g0195(.A(new_n580_), .B(new_n578_), .Y(new_n581_));
  OR2X1    g0196(.A(\req[81] ), .B(\req[80] ), .Y(new_n582_));
  AOI21X1  g0197(.A0(\req[79] ), .A1(new_n578_), .B0(new_n582_), .Y(new_n583_));
  INVX1    g0198(.A(new_n583_), .Y(new_n584_));
  AOI21X1  g0199(.A0(new_n581_), .A1(new_n577_), .B0(new_n584_), .Y(new_n585_));
  INVX1    g0200(.A(\priority[83] ), .Y(new_n586_));
  INVX1    g0201(.A(\req[81] ), .Y(new_n587_));
  AOI21X1  g0202(.A0(new_n587_), .A1(\priority[81] ), .B0(\priority[82] ), .Y(new_n588_));
  NAND2X1  g0203(.A(new_n588_), .B(new_n586_), .Y(new_n589_));
  OR2X1    g0204(.A(\req[84] ), .B(\req[83] ), .Y(new_n590_));
  AOI21X1  g0205(.A0(\req[82] ), .A1(new_n586_), .B0(new_n590_), .Y(new_n591_));
  OAI21X1  g0206(.A0(new_n589_), .A1(new_n585_), .B0(new_n591_), .Y(new_n592_));
  INVX1    g0207(.A(\priority[86] ), .Y(new_n593_));
  INVX1    g0208(.A(\req[84] ), .Y(new_n594_));
  AOI21X1  g0209(.A0(new_n594_), .A1(\priority[84] ), .B0(\priority[85] ), .Y(new_n595_));
  AND2X1   g0210(.A(new_n595_), .B(new_n593_), .Y(new_n596_));
  OR2X1    g0211(.A(\req[87] ), .B(\req[86] ), .Y(new_n597_));
  AOI21X1  g0212(.A0(\req[85] ), .A1(new_n593_), .B0(new_n597_), .Y(new_n598_));
  INVX1    g0213(.A(new_n598_), .Y(new_n599_));
  AOI21X1  g0214(.A0(new_n596_), .A1(new_n592_), .B0(new_n599_), .Y(new_n600_));
  INVX1    g0215(.A(\priority[89] ), .Y(new_n601_));
  INVX1    g0216(.A(\req[87] ), .Y(new_n602_));
  AOI21X1  g0217(.A0(new_n602_), .A1(\priority[87] ), .B0(\priority[88] ), .Y(new_n603_));
  NAND2X1  g0218(.A(new_n603_), .B(new_n601_), .Y(new_n604_));
  OR2X1    g0219(.A(\req[90] ), .B(\req[89] ), .Y(new_n605_));
  AOI21X1  g0220(.A0(\req[88] ), .A1(new_n601_), .B0(new_n605_), .Y(new_n606_));
  OAI21X1  g0221(.A0(new_n604_), .A1(new_n600_), .B0(new_n606_), .Y(new_n607_));
  INVX1    g0222(.A(\priority[92] ), .Y(new_n608_));
  INVX1    g0223(.A(\req[90] ), .Y(new_n609_));
  AOI21X1  g0224(.A0(new_n609_), .A1(\priority[90] ), .B0(\priority[91] ), .Y(new_n610_));
  AND2X1   g0225(.A(new_n610_), .B(new_n608_), .Y(new_n611_));
  OR2X1    g0226(.A(\req[93] ), .B(\req[92] ), .Y(new_n612_));
  AOI21X1  g0227(.A0(\req[91] ), .A1(new_n608_), .B0(new_n612_), .Y(new_n613_));
  INVX1    g0228(.A(new_n613_), .Y(new_n614_));
  AOI21X1  g0229(.A0(new_n611_), .A1(new_n607_), .B0(new_n614_), .Y(new_n615_));
  INVX1    g0230(.A(\priority[95] ), .Y(new_n616_));
  INVX1    g0231(.A(\req[93] ), .Y(new_n617_));
  AOI21X1  g0232(.A0(new_n617_), .A1(\priority[93] ), .B0(\priority[94] ), .Y(new_n618_));
  NAND2X1  g0233(.A(new_n618_), .B(new_n616_), .Y(new_n619_));
  OR2X1    g0234(.A(\req[96] ), .B(\req[95] ), .Y(new_n620_));
  AOI21X1  g0235(.A0(\req[94] ), .A1(new_n616_), .B0(new_n620_), .Y(new_n621_));
  OAI21X1  g0236(.A0(new_n619_), .A1(new_n615_), .B0(new_n621_), .Y(new_n622_));
  INVX1    g0237(.A(\priority[98] ), .Y(new_n623_));
  INVX1    g0238(.A(\req[96] ), .Y(new_n624_));
  AOI21X1  g0239(.A0(new_n624_), .A1(\priority[96] ), .B0(\priority[97] ), .Y(new_n625_));
  AND2X1   g0240(.A(new_n625_), .B(new_n623_), .Y(new_n626_));
  OR2X1    g0241(.A(\req[99] ), .B(\req[98] ), .Y(new_n627_));
  AOI21X1  g0242(.A0(\req[97] ), .A1(new_n623_), .B0(new_n627_), .Y(new_n628_));
  INVX1    g0243(.A(new_n628_), .Y(new_n629_));
  AOI21X1  g0244(.A0(new_n626_), .A1(new_n622_), .B0(new_n629_), .Y(new_n630_));
  INVX1    g0245(.A(\priority[101] ), .Y(new_n631_));
  INVX1    g0246(.A(\req[99] ), .Y(new_n632_));
  AOI21X1  g0247(.A0(new_n632_), .A1(\priority[99] ), .B0(\priority[100] ), .Y(new_n633_));
  NAND2X1  g0248(.A(new_n633_), .B(new_n631_), .Y(new_n634_));
  OR2X1    g0249(.A(\req[102] ), .B(\req[101] ), .Y(new_n635_));
  AOI21X1  g0250(.A0(\req[100] ), .A1(new_n631_), .B0(new_n635_), .Y(new_n636_));
  OAI21X1  g0251(.A0(new_n634_), .A1(new_n630_), .B0(new_n636_), .Y(new_n637_));
  INVX1    g0252(.A(\priority[104] ), .Y(new_n638_));
  INVX1    g0253(.A(\req[102] ), .Y(new_n639_));
  AOI21X1  g0254(.A0(new_n639_), .A1(\priority[102] ), .B0(\priority[103] ), .Y(new_n640_));
  AND2X1   g0255(.A(new_n640_), .B(new_n638_), .Y(new_n641_));
  OR2X1    g0256(.A(\req[105] ), .B(\req[104] ), .Y(new_n642_));
  AOI21X1  g0257(.A0(\req[103] ), .A1(new_n638_), .B0(new_n642_), .Y(new_n643_));
  INVX1    g0258(.A(new_n643_), .Y(new_n644_));
  AOI21X1  g0259(.A0(new_n641_), .A1(new_n637_), .B0(new_n644_), .Y(new_n645_));
  INVX1    g0260(.A(\priority[107] ), .Y(new_n646_));
  INVX1    g0261(.A(\req[105] ), .Y(new_n647_));
  AOI21X1  g0262(.A0(new_n647_), .A1(\priority[105] ), .B0(\priority[106] ), .Y(new_n648_));
  NAND2X1  g0263(.A(new_n648_), .B(new_n646_), .Y(new_n649_));
  OR2X1    g0264(.A(\req[108] ), .B(\req[107] ), .Y(new_n650_));
  AOI21X1  g0265(.A0(\req[106] ), .A1(new_n646_), .B0(new_n650_), .Y(new_n651_));
  OAI21X1  g0266(.A0(new_n649_), .A1(new_n645_), .B0(new_n651_), .Y(new_n652_));
  INVX1    g0267(.A(\priority[110] ), .Y(new_n653_));
  INVX1    g0268(.A(\req[108] ), .Y(new_n654_));
  AOI21X1  g0269(.A0(new_n654_), .A1(\priority[108] ), .B0(\priority[109] ), .Y(new_n655_));
  AND2X1   g0270(.A(new_n655_), .B(new_n653_), .Y(new_n656_));
  OR2X1    g0271(.A(\req[111] ), .B(\req[110] ), .Y(new_n657_));
  AOI21X1  g0272(.A0(\req[109] ), .A1(new_n653_), .B0(new_n657_), .Y(new_n658_));
  INVX1    g0273(.A(new_n658_), .Y(new_n659_));
  AOI21X1  g0274(.A0(new_n656_), .A1(new_n652_), .B0(new_n659_), .Y(new_n660_));
  INVX1    g0275(.A(\priority[113] ), .Y(new_n661_));
  INVX1    g0276(.A(\req[111] ), .Y(new_n662_));
  AOI21X1  g0277(.A0(new_n662_), .A1(\priority[111] ), .B0(\priority[112] ), .Y(new_n663_));
  NAND2X1  g0278(.A(new_n663_), .B(new_n661_), .Y(new_n664_));
  OR2X1    g0279(.A(\req[114] ), .B(\req[113] ), .Y(new_n665_));
  AOI21X1  g0280(.A0(\req[112] ), .A1(new_n661_), .B0(new_n665_), .Y(new_n666_));
  OAI21X1  g0281(.A0(new_n664_), .A1(new_n660_), .B0(new_n666_), .Y(new_n667_));
  INVX1    g0282(.A(\priority[116] ), .Y(new_n668_));
  INVX1    g0283(.A(\req[114] ), .Y(new_n669_));
  AOI21X1  g0284(.A0(new_n669_), .A1(\priority[114] ), .B0(\priority[115] ), .Y(new_n670_));
  AND2X1   g0285(.A(new_n670_), .B(new_n668_), .Y(new_n671_));
  OR2X1    g0286(.A(\req[117] ), .B(\req[116] ), .Y(new_n672_));
  AOI21X1  g0287(.A0(\req[115] ), .A1(new_n668_), .B0(new_n672_), .Y(new_n673_));
  INVX1    g0288(.A(new_n673_), .Y(new_n674_));
  AOI21X1  g0289(.A0(new_n671_), .A1(new_n667_), .B0(new_n674_), .Y(new_n675_));
  INVX1    g0290(.A(\priority[119] ), .Y(new_n676_));
  INVX1    g0291(.A(\req[117] ), .Y(new_n677_));
  AOI21X1  g0292(.A0(new_n677_), .A1(\priority[117] ), .B0(\priority[118] ), .Y(new_n678_));
  NAND2X1  g0293(.A(new_n678_), .B(new_n676_), .Y(new_n679_));
  OR2X1    g0294(.A(\req[120] ), .B(\req[119] ), .Y(new_n680_));
  AOI21X1  g0295(.A0(\req[118] ), .A1(new_n676_), .B0(new_n680_), .Y(new_n681_));
  OAI21X1  g0296(.A0(new_n679_), .A1(new_n675_), .B0(new_n681_), .Y(new_n682_));
  INVX1    g0297(.A(\priority[122] ), .Y(new_n683_));
  INVX1    g0298(.A(\req[120] ), .Y(new_n684_));
  AOI21X1  g0299(.A0(new_n684_), .A1(\priority[120] ), .B0(\priority[121] ), .Y(new_n685_));
  AND2X1   g0300(.A(new_n685_), .B(new_n683_), .Y(new_n686_));
  OR2X1    g0301(.A(\req[123] ), .B(\req[122] ), .Y(new_n687_));
  AOI21X1  g0302(.A0(\req[121] ), .A1(new_n683_), .B0(new_n687_), .Y(new_n688_));
  INVX1    g0303(.A(new_n688_), .Y(new_n689_));
  AOI21X1  g0304(.A0(new_n686_), .A1(new_n682_), .B0(new_n689_), .Y(new_n690_));
  INVX1    g0305(.A(\priority[125] ), .Y(new_n691_));
  INVX1    g0306(.A(\req[123] ), .Y(new_n692_));
  AOI21X1  g0307(.A0(new_n692_), .A1(\priority[123] ), .B0(\priority[124] ), .Y(new_n693_));
  NAND2X1  g0308(.A(new_n693_), .B(new_n691_), .Y(new_n694_));
  OR2X1    g0309(.A(\req[126] ), .B(\req[125] ), .Y(new_n695_));
  AOI21X1  g0310(.A0(\req[124] ), .A1(new_n691_), .B0(new_n695_), .Y(new_n696_));
  OAI21X1  g0311(.A0(new_n694_), .A1(new_n690_), .B0(new_n696_), .Y(new_n697_));
  INVX1    g0312(.A(\priority[0] ), .Y(new_n698_));
  INVX1    g0313(.A(\req[126] ), .Y(new_n699_));
  AOI21X1  g0314(.A0(new_n699_), .A1(\priority[126] ), .B0(\priority[127] ), .Y(new_n700_));
  AND2X1   g0315(.A(new_n700_), .B(new_n698_), .Y(new_n701_));
  INVX1    g0316(.A(\req[127] ), .Y(new_n702_));
  OAI21X1  g0317(.A0(new_n702_), .A1(\priority[0] ), .B0(\req[0] ), .Y(new_n703_));
  AOI21X1  g0318(.A0(new_n701_), .A1(new_n697_), .B0(new_n703_), .Y(\grant[0] ));
  INVX1    g0319(.A(\priority[3] ), .Y(new_n705_));
  OAI21X1  g0320(.A0(\req[2] ), .A1(new_n387_), .B0(new_n705_), .Y(new_n706_));
  NOR2X1   g0321(.A(\req[4] ), .B(\req[3] ), .Y(new_n707_));
  AND2X1   g0322(.A(new_n707_), .B(new_n706_), .Y(new_n708_));
  INVX1    g0323(.A(\priority[6] ), .Y(new_n709_));
  INVX1    g0324(.A(\req[4] ), .Y(new_n710_));
  AOI21X1  g0325(.A0(new_n710_), .A1(\priority[4] ), .B0(\priority[5] ), .Y(new_n711_));
  NAND2X1  g0326(.A(new_n711_), .B(new_n709_), .Y(new_n712_));
  OR2X1    g0327(.A(\req[7] ), .B(\req[6] ), .Y(new_n713_));
  AOI21X1  g0328(.A0(\req[5] ), .A1(new_n709_), .B0(new_n713_), .Y(new_n714_));
  OAI21X1  g0329(.A0(new_n712_), .A1(new_n708_), .B0(new_n714_), .Y(new_n715_));
  INVX1    g0330(.A(\priority[9] ), .Y(new_n716_));
  INVX1    g0331(.A(\req[7] ), .Y(new_n717_));
  AOI21X1  g0332(.A0(new_n717_), .A1(\priority[7] ), .B0(\priority[8] ), .Y(new_n718_));
  AND2X1   g0333(.A(new_n718_), .B(new_n716_), .Y(new_n719_));
  OR2X1    g0334(.A(\req[10] ), .B(\req[9] ), .Y(new_n720_));
  AOI21X1  g0335(.A0(\req[8] ), .A1(new_n716_), .B0(new_n720_), .Y(new_n721_));
  INVX1    g0336(.A(new_n721_), .Y(new_n722_));
  AOI21X1  g0337(.A0(new_n719_), .A1(new_n715_), .B0(new_n722_), .Y(new_n723_));
  INVX1    g0338(.A(\priority[12] ), .Y(new_n724_));
  INVX1    g0339(.A(\req[10] ), .Y(new_n725_));
  AOI21X1  g0340(.A0(new_n725_), .A1(\priority[10] ), .B0(\priority[11] ), .Y(new_n726_));
  NAND2X1  g0341(.A(new_n726_), .B(new_n724_), .Y(new_n727_));
  OR2X1    g0342(.A(\req[13] ), .B(\req[12] ), .Y(new_n728_));
  AOI21X1  g0343(.A0(\req[11] ), .A1(new_n724_), .B0(new_n728_), .Y(new_n729_));
  OAI21X1  g0344(.A0(new_n727_), .A1(new_n723_), .B0(new_n729_), .Y(new_n730_));
  INVX1    g0345(.A(\priority[15] ), .Y(new_n731_));
  INVX1    g0346(.A(\req[13] ), .Y(new_n732_));
  AOI21X1  g0347(.A0(new_n732_), .A1(\priority[13] ), .B0(\priority[14] ), .Y(new_n733_));
  AND2X1   g0348(.A(new_n733_), .B(new_n731_), .Y(new_n734_));
  OR2X1    g0349(.A(\req[16] ), .B(\req[15] ), .Y(new_n735_));
  AOI21X1  g0350(.A0(\req[14] ), .A1(new_n731_), .B0(new_n735_), .Y(new_n736_));
  INVX1    g0351(.A(new_n736_), .Y(new_n737_));
  AOI21X1  g0352(.A0(new_n734_), .A1(new_n730_), .B0(new_n737_), .Y(new_n738_));
  INVX1    g0353(.A(\priority[18] ), .Y(new_n739_));
  INVX1    g0354(.A(\req[16] ), .Y(new_n740_));
  AOI21X1  g0355(.A0(new_n740_), .A1(\priority[16] ), .B0(\priority[17] ), .Y(new_n741_));
  NAND2X1  g0356(.A(new_n741_), .B(new_n739_), .Y(new_n742_));
  OR2X1    g0357(.A(\req[19] ), .B(\req[18] ), .Y(new_n743_));
  AOI21X1  g0358(.A0(\req[17] ), .A1(new_n739_), .B0(new_n743_), .Y(new_n744_));
  OAI21X1  g0359(.A0(new_n742_), .A1(new_n738_), .B0(new_n744_), .Y(new_n745_));
  INVX1    g0360(.A(\priority[21] ), .Y(new_n746_));
  INVX1    g0361(.A(\req[19] ), .Y(new_n747_));
  AOI21X1  g0362(.A0(new_n747_), .A1(\priority[19] ), .B0(\priority[20] ), .Y(new_n748_));
  AND2X1   g0363(.A(new_n748_), .B(new_n746_), .Y(new_n749_));
  OR2X1    g0364(.A(\req[22] ), .B(\req[21] ), .Y(new_n750_));
  AOI21X1  g0365(.A0(\req[20] ), .A1(new_n746_), .B0(new_n750_), .Y(new_n751_));
  INVX1    g0366(.A(new_n751_), .Y(new_n752_));
  AOI21X1  g0367(.A0(new_n749_), .A1(new_n745_), .B0(new_n752_), .Y(new_n753_));
  INVX1    g0368(.A(\priority[24] ), .Y(new_n754_));
  INVX1    g0369(.A(\req[22] ), .Y(new_n755_));
  AOI21X1  g0370(.A0(new_n755_), .A1(\priority[22] ), .B0(\priority[23] ), .Y(new_n756_));
  NAND2X1  g0371(.A(new_n756_), .B(new_n754_), .Y(new_n757_));
  OR2X1    g0372(.A(\req[25] ), .B(\req[24] ), .Y(new_n758_));
  AOI21X1  g0373(.A0(\req[23] ), .A1(new_n754_), .B0(new_n758_), .Y(new_n759_));
  OAI21X1  g0374(.A0(new_n757_), .A1(new_n753_), .B0(new_n759_), .Y(new_n760_));
  INVX1    g0375(.A(\priority[27] ), .Y(new_n761_));
  INVX1    g0376(.A(\req[25] ), .Y(new_n762_));
  AOI21X1  g0377(.A0(new_n762_), .A1(\priority[25] ), .B0(\priority[26] ), .Y(new_n763_));
  AND2X1   g0378(.A(new_n763_), .B(new_n761_), .Y(new_n764_));
  OR2X1    g0379(.A(\req[28] ), .B(\req[27] ), .Y(new_n765_));
  AOI21X1  g0380(.A0(\req[26] ), .A1(new_n761_), .B0(new_n765_), .Y(new_n766_));
  INVX1    g0381(.A(new_n766_), .Y(new_n767_));
  AOI21X1  g0382(.A0(new_n764_), .A1(new_n760_), .B0(new_n767_), .Y(new_n768_));
  INVX1    g0383(.A(\priority[30] ), .Y(new_n769_));
  INVX1    g0384(.A(\req[28] ), .Y(new_n770_));
  AOI21X1  g0385(.A0(new_n770_), .A1(\priority[28] ), .B0(\priority[29] ), .Y(new_n771_));
  NAND2X1  g0386(.A(new_n771_), .B(new_n769_), .Y(new_n772_));
  OR2X1    g0387(.A(\req[31] ), .B(\req[30] ), .Y(new_n773_));
  AOI21X1  g0388(.A0(\req[29] ), .A1(new_n769_), .B0(new_n773_), .Y(new_n774_));
  OAI21X1  g0389(.A0(new_n772_), .A1(new_n768_), .B0(new_n774_), .Y(new_n775_));
  INVX1    g0390(.A(\priority[33] ), .Y(new_n776_));
  INVX1    g0391(.A(\req[31] ), .Y(new_n777_));
  AOI21X1  g0392(.A0(new_n777_), .A1(\priority[31] ), .B0(\priority[32] ), .Y(new_n778_));
  AND2X1   g0393(.A(new_n778_), .B(new_n776_), .Y(new_n779_));
  OR2X1    g0394(.A(\req[34] ), .B(\req[33] ), .Y(new_n780_));
  AOI21X1  g0395(.A0(\req[32] ), .A1(new_n776_), .B0(new_n780_), .Y(new_n781_));
  INVX1    g0396(.A(new_n781_), .Y(new_n782_));
  AOI21X1  g0397(.A0(new_n779_), .A1(new_n775_), .B0(new_n782_), .Y(new_n783_));
  INVX1    g0398(.A(\priority[36] ), .Y(new_n784_));
  INVX1    g0399(.A(\req[34] ), .Y(new_n785_));
  AOI21X1  g0400(.A0(new_n785_), .A1(\priority[34] ), .B0(\priority[35] ), .Y(new_n786_));
  NAND2X1  g0401(.A(new_n786_), .B(new_n784_), .Y(new_n787_));
  OR2X1    g0402(.A(\req[37] ), .B(\req[36] ), .Y(new_n788_));
  AOI21X1  g0403(.A0(\req[35] ), .A1(new_n784_), .B0(new_n788_), .Y(new_n789_));
  OAI21X1  g0404(.A0(new_n787_), .A1(new_n783_), .B0(new_n789_), .Y(new_n790_));
  INVX1    g0405(.A(\priority[39] ), .Y(new_n791_));
  INVX1    g0406(.A(\req[37] ), .Y(new_n792_));
  AOI21X1  g0407(.A0(new_n792_), .A1(\priority[37] ), .B0(\priority[38] ), .Y(new_n793_));
  AND2X1   g0408(.A(new_n793_), .B(new_n791_), .Y(new_n794_));
  OR2X1    g0409(.A(\req[40] ), .B(\req[39] ), .Y(new_n795_));
  AOI21X1  g0410(.A0(\req[38] ), .A1(new_n791_), .B0(new_n795_), .Y(new_n796_));
  INVX1    g0411(.A(new_n796_), .Y(new_n797_));
  AOI21X1  g0412(.A0(new_n794_), .A1(new_n790_), .B0(new_n797_), .Y(new_n798_));
  INVX1    g0413(.A(\priority[42] ), .Y(new_n799_));
  INVX1    g0414(.A(\req[40] ), .Y(new_n800_));
  AOI21X1  g0415(.A0(new_n800_), .A1(\priority[40] ), .B0(\priority[41] ), .Y(new_n801_));
  NAND2X1  g0416(.A(new_n801_), .B(new_n799_), .Y(new_n802_));
  OR2X1    g0417(.A(\req[43] ), .B(\req[42] ), .Y(new_n803_));
  AOI21X1  g0418(.A0(\req[41] ), .A1(new_n799_), .B0(new_n803_), .Y(new_n804_));
  OAI21X1  g0419(.A0(new_n802_), .A1(new_n798_), .B0(new_n804_), .Y(new_n805_));
  INVX1    g0420(.A(\priority[45] ), .Y(new_n806_));
  INVX1    g0421(.A(\req[43] ), .Y(new_n807_));
  AOI21X1  g0422(.A0(new_n807_), .A1(\priority[43] ), .B0(\priority[44] ), .Y(new_n808_));
  AND2X1   g0423(.A(new_n808_), .B(new_n806_), .Y(new_n809_));
  OR2X1    g0424(.A(\req[46] ), .B(\req[45] ), .Y(new_n810_));
  AOI21X1  g0425(.A0(\req[44] ), .A1(new_n806_), .B0(new_n810_), .Y(new_n811_));
  INVX1    g0426(.A(new_n811_), .Y(new_n812_));
  AOI21X1  g0427(.A0(new_n809_), .A1(new_n805_), .B0(new_n812_), .Y(new_n813_));
  INVX1    g0428(.A(\priority[48] ), .Y(new_n814_));
  INVX1    g0429(.A(\req[46] ), .Y(new_n815_));
  AOI21X1  g0430(.A0(new_n815_), .A1(\priority[46] ), .B0(\priority[47] ), .Y(new_n816_));
  NAND2X1  g0431(.A(new_n816_), .B(new_n814_), .Y(new_n817_));
  OR2X1    g0432(.A(\req[49] ), .B(\req[48] ), .Y(new_n818_));
  AOI21X1  g0433(.A0(\req[47] ), .A1(new_n814_), .B0(new_n818_), .Y(new_n819_));
  OAI21X1  g0434(.A0(new_n817_), .A1(new_n813_), .B0(new_n819_), .Y(new_n820_));
  INVX1    g0435(.A(\priority[51] ), .Y(new_n821_));
  INVX1    g0436(.A(\req[49] ), .Y(new_n822_));
  AOI21X1  g0437(.A0(new_n822_), .A1(\priority[49] ), .B0(\priority[50] ), .Y(new_n823_));
  AND2X1   g0438(.A(new_n823_), .B(new_n821_), .Y(new_n824_));
  OR2X1    g0439(.A(\req[52] ), .B(\req[51] ), .Y(new_n825_));
  AOI21X1  g0440(.A0(\req[50] ), .A1(new_n821_), .B0(new_n825_), .Y(new_n826_));
  INVX1    g0441(.A(new_n826_), .Y(new_n827_));
  AOI21X1  g0442(.A0(new_n824_), .A1(new_n820_), .B0(new_n827_), .Y(new_n828_));
  INVX1    g0443(.A(\priority[54] ), .Y(new_n829_));
  INVX1    g0444(.A(\req[52] ), .Y(new_n830_));
  AOI21X1  g0445(.A0(new_n830_), .A1(\priority[52] ), .B0(\priority[53] ), .Y(new_n831_));
  NAND2X1  g0446(.A(new_n831_), .B(new_n829_), .Y(new_n832_));
  OR2X1    g0447(.A(\req[55] ), .B(\req[54] ), .Y(new_n833_));
  AOI21X1  g0448(.A0(\req[53] ), .A1(new_n829_), .B0(new_n833_), .Y(new_n834_));
  OAI21X1  g0449(.A0(new_n832_), .A1(new_n828_), .B0(new_n834_), .Y(new_n835_));
  INVX1    g0450(.A(\priority[57] ), .Y(new_n836_));
  INVX1    g0451(.A(\req[55] ), .Y(new_n837_));
  AOI21X1  g0452(.A0(new_n837_), .A1(\priority[55] ), .B0(\priority[56] ), .Y(new_n838_));
  AND2X1   g0453(.A(new_n838_), .B(new_n836_), .Y(new_n839_));
  OR2X1    g0454(.A(\req[58] ), .B(\req[57] ), .Y(new_n840_));
  AOI21X1  g0455(.A0(\req[56] ), .A1(new_n836_), .B0(new_n840_), .Y(new_n841_));
  INVX1    g0456(.A(new_n841_), .Y(new_n842_));
  AOI21X1  g0457(.A0(new_n839_), .A1(new_n835_), .B0(new_n842_), .Y(new_n843_));
  INVX1    g0458(.A(\priority[60] ), .Y(new_n844_));
  INVX1    g0459(.A(\req[58] ), .Y(new_n845_));
  AOI21X1  g0460(.A0(new_n845_), .A1(\priority[58] ), .B0(\priority[59] ), .Y(new_n846_));
  NAND2X1  g0461(.A(new_n846_), .B(new_n844_), .Y(new_n847_));
  OR2X1    g0462(.A(\req[61] ), .B(\req[60] ), .Y(new_n848_));
  AOI21X1  g0463(.A0(\req[59] ), .A1(new_n844_), .B0(new_n848_), .Y(new_n849_));
  OAI21X1  g0464(.A0(new_n847_), .A1(new_n843_), .B0(new_n849_), .Y(new_n850_));
  INVX1    g0465(.A(\priority[63] ), .Y(new_n851_));
  INVX1    g0466(.A(\req[61] ), .Y(new_n852_));
  AOI21X1  g0467(.A0(new_n852_), .A1(\priority[61] ), .B0(\priority[62] ), .Y(new_n853_));
  AND2X1   g0468(.A(new_n853_), .B(new_n851_), .Y(new_n854_));
  OR2X1    g0469(.A(\req[64] ), .B(\req[63] ), .Y(new_n855_));
  AOI21X1  g0470(.A0(\req[62] ), .A1(new_n851_), .B0(new_n855_), .Y(new_n856_));
  INVX1    g0471(.A(new_n856_), .Y(new_n857_));
  AOI21X1  g0472(.A0(new_n854_), .A1(new_n850_), .B0(new_n857_), .Y(new_n858_));
  INVX1    g0473(.A(\priority[66] ), .Y(new_n859_));
  INVX1    g0474(.A(\req[64] ), .Y(new_n860_));
  AOI21X1  g0475(.A0(new_n860_), .A1(\priority[64] ), .B0(\priority[65] ), .Y(new_n861_));
  NAND2X1  g0476(.A(new_n861_), .B(new_n859_), .Y(new_n862_));
  OR2X1    g0477(.A(\req[67] ), .B(\req[66] ), .Y(new_n863_));
  AOI21X1  g0478(.A0(\req[65] ), .A1(new_n859_), .B0(new_n863_), .Y(new_n864_));
  OAI21X1  g0479(.A0(new_n862_), .A1(new_n858_), .B0(new_n864_), .Y(new_n865_));
  INVX1    g0480(.A(\priority[69] ), .Y(new_n866_));
  INVX1    g0481(.A(\req[67] ), .Y(new_n867_));
  AOI21X1  g0482(.A0(new_n867_), .A1(\priority[67] ), .B0(\priority[68] ), .Y(new_n868_));
  AND2X1   g0483(.A(new_n868_), .B(new_n866_), .Y(new_n869_));
  OR2X1    g0484(.A(\req[70] ), .B(\req[69] ), .Y(new_n870_));
  AOI21X1  g0485(.A0(\req[68] ), .A1(new_n866_), .B0(new_n870_), .Y(new_n871_));
  INVX1    g0486(.A(new_n871_), .Y(new_n872_));
  AOI21X1  g0487(.A0(new_n869_), .A1(new_n865_), .B0(new_n872_), .Y(new_n873_));
  INVX1    g0488(.A(\priority[72] ), .Y(new_n874_));
  INVX1    g0489(.A(\req[70] ), .Y(new_n875_));
  AOI21X1  g0490(.A0(new_n875_), .A1(\priority[70] ), .B0(\priority[71] ), .Y(new_n876_));
  NAND2X1  g0491(.A(new_n876_), .B(new_n874_), .Y(new_n877_));
  OR2X1    g0492(.A(\req[73] ), .B(\req[72] ), .Y(new_n878_));
  AOI21X1  g0493(.A0(\req[71] ), .A1(new_n874_), .B0(new_n878_), .Y(new_n879_));
  OAI21X1  g0494(.A0(new_n877_), .A1(new_n873_), .B0(new_n879_), .Y(new_n880_));
  INVX1    g0495(.A(\priority[75] ), .Y(new_n881_));
  INVX1    g0496(.A(\req[73] ), .Y(new_n882_));
  AOI21X1  g0497(.A0(new_n882_), .A1(\priority[73] ), .B0(\priority[74] ), .Y(new_n883_));
  AND2X1   g0498(.A(new_n883_), .B(new_n881_), .Y(new_n884_));
  OR2X1    g0499(.A(\req[76] ), .B(\req[75] ), .Y(new_n885_));
  AOI21X1  g0500(.A0(\req[74] ), .A1(new_n881_), .B0(new_n885_), .Y(new_n886_));
  INVX1    g0501(.A(new_n886_), .Y(new_n887_));
  AOI21X1  g0502(.A0(new_n884_), .A1(new_n880_), .B0(new_n887_), .Y(new_n888_));
  INVX1    g0503(.A(\priority[78] ), .Y(new_n889_));
  INVX1    g0504(.A(\req[76] ), .Y(new_n890_));
  AOI21X1  g0505(.A0(new_n890_), .A1(\priority[76] ), .B0(\priority[77] ), .Y(new_n891_));
  NAND2X1  g0506(.A(new_n891_), .B(new_n889_), .Y(new_n892_));
  OR2X1    g0507(.A(\req[79] ), .B(\req[78] ), .Y(new_n893_));
  AOI21X1  g0508(.A0(\req[77] ), .A1(new_n889_), .B0(new_n893_), .Y(new_n894_));
  OAI21X1  g0509(.A0(new_n892_), .A1(new_n888_), .B0(new_n894_), .Y(new_n895_));
  INVX1    g0510(.A(\priority[81] ), .Y(new_n896_));
  INVX1    g0511(.A(\req[79] ), .Y(new_n897_));
  AOI21X1  g0512(.A0(new_n897_), .A1(\priority[79] ), .B0(\priority[80] ), .Y(new_n898_));
  AND2X1   g0513(.A(new_n898_), .B(new_n896_), .Y(new_n899_));
  OR2X1    g0514(.A(\req[82] ), .B(\req[81] ), .Y(new_n900_));
  AOI21X1  g0515(.A0(\req[80] ), .A1(new_n896_), .B0(new_n900_), .Y(new_n901_));
  INVX1    g0516(.A(new_n901_), .Y(new_n902_));
  AOI21X1  g0517(.A0(new_n899_), .A1(new_n895_), .B0(new_n902_), .Y(new_n903_));
  INVX1    g0518(.A(\priority[84] ), .Y(new_n904_));
  INVX1    g0519(.A(\req[82] ), .Y(new_n905_));
  AOI21X1  g0520(.A0(new_n905_), .A1(\priority[82] ), .B0(\priority[83] ), .Y(new_n906_));
  NAND2X1  g0521(.A(new_n906_), .B(new_n904_), .Y(new_n907_));
  OR2X1    g0522(.A(\req[85] ), .B(\req[84] ), .Y(new_n908_));
  AOI21X1  g0523(.A0(\req[83] ), .A1(new_n904_), .B0(new_n908_), .Y(new_n909_));
  OAI21X1  g0524(.A0(new_n907_), .A1(new_n903_), .B0(new_n909_), .Y(new_n910_));
  INVX1    g0525(.A(\priority[87] ), .Y(new_n911_));
  INVX1    g0526(.A(\req[85] ), .Y(new_n912_));
  AOI21X1  g0527(.A0(new_n912_), .A1(\priority[85] ), .B0(\priority[86] ), .Y(new_n913_));
  AND2X1   g0528(.A(new_n913_), .B(new_n911_), .Y(new_n914_));
  OR2X1    g0529(.A(\req[88] ), .B(\req[87] ), .Y(new_n915_));
  AOI21X1  g0530(.A0(\req[86] ), .A1(new_n911_), .B0(new_n915_), .Y(new_n916_));
  INVX1    g0531(.A(new_n916_), .Y(new_n917_));
  AOI21X1  g0532(.A0(new_n914_), .A1(new_n910_), .B0(new_n917_), .Y(new_n918_));
  INVX1    g0533(.A(\priority[90] ), .Y(new_n919_));
  INVX1    g0534(.A(\req[88] ), .Y(new_n920_));
  AOI21X1  g0535(.A0(new_n920_), .A1(\priority[88] ), .B0(\priority[89] ), .Y(new_n921_));
  NAND2X1  g0536(.A(new_n921_), .B(new_n919_), .Y(new_n922_));
  OR2X1    g0537(.A(\req[91] ), .B(\req[90] ), .Y(new_n923_));
  AOI21X1  g0538(.A0(\req[89] ), .A1(new_n919_), .B0(new_n923_), .Y(new_n924_));
  OAI21X1  g0539(.A0(new_n922_), .A1(new_n918_), .B0(new_n924_), .Y(new_n925_));
  INVX1    g0540(.A(\priority[93] ), .Y(new_n926_));
  INVX1    g0541(.A(\req[91] ), .Y(new_n927_));
  AOI21X1  g0542(.A0(new_n927_), .A1(\priority[91] ), .B0(\priority[92] ), .Y(new_n928_));
  AND2X1   g0543(.A(new_n928_), .B(new_n926_), .Y(new_n929_));
  OR2X1    g0544(.A(\req[94] ), .B(\req[93] ), .Y(new_n930_));
  AOI21X1  g0545(.A0(\req[92] ), .A1(new_n926_), .B0(new_n930_), .Y(new_n931_));
  INVX1    g0546(.A(new_n931_), .Y(new_n932_));
  AOI21X1  g0547(.A0(new_n929_), .A1(new_n925_), .B0(new_n932_), .Y(new_n933_));
  INVX1    g0548(.A(\priority[96] ), .Y(new_n934_));
  INVX1    g0549(.A(\req[94] ), .Y(new_n935_));
  AOI21X1  g0550(.A0(new_n935_), .A1(\priority[94] ), .B0(\priority[95] ), .Y(new_n936_));
  NAND2X1  g0551(.A(new_n936_), .B(new_n934_), .Y(new_n937_));
  OR2X1    g0552(.A(\req[97] ), .B(\req[96] ), .Y(new_n938_));
  AOI21X1  g0553(.A0(\req[95] ), .A1(new_n934_), .B0(new_n938_), .Y(new_n939_));
  OAI21X1  g0554(.A0(new_n937_), .A1(new_n933_), .B0(new_n939_), .Y(new_n940_));
  INVX1    g0555(.A(\priority[99] ), .Y(new_n941_));
  INVX1    g0556(.A(\req[97] ), .Y(new_n942_));
  AOI21X1  g0557(.A0(new_n942_), .A1(\priority[97] ), .B0(\priority[98] ), .Y(new_n943_));
  AND2X1   g0558(.A(new_n943_), .B(new_n941_), .Y(new_n944_));
  OR2X1    g0559(.A(\req[100] ), .B(\req[99] ), .Y(new_n945_));
  AOI21X1  g0560(.A0(\req[98] ), .A1(new_n941_), .B0(new_n945_), .Y(new_n946_));
  INVX1    g0561(.A(new_n946_), .Y(new_n947_));
  AOI21X1  g0562(.A0(new_n944_), .A1(new_n940_), .B0(new_n947_), .Y(new_n948_));
  INVX1    g0563(.A(\priority[102] ), .Y(new_n949_));
  INVX1    g0564(.A(\req[100] ), .Y(new_n950_));
  AOI21X1  g0565(.A0(new_n950_), .A1(\priority[100] ), .B0(\priority[101] ), .Y(new_n951_));
  NAND2X1  g0566(.A(new_n951_), .B(new_n949_), .Y(new_n952_));
  OR2X1    g0567(.A(\req[103] ), .B(\req[102] ), .Y(new_n953_));
  AOI21X1  g0568(.A0(\req[101] ), .A1(new_n949_), .B0(new_n953_), .Y(new_n954_));
  OAI21X1  g0569(.A0(new_n952_), .A1(new_n948_), .B0(new_n954_), .Y(new_n955_));
  INVX1    g0570(.A(\priority[105] ), .Y(new_n956_));
  INVX1    g0571(.A(\req[103] ), .Y(new_n957_));
  AOI21X1  g0572(.A0(new_n957_), .A1(\priority[103] ), .B0(\priority[104] ), .Y(new_n958_));
  AND2X1   g0573(.A(new_n958_), .B(new_n956_), .Y(new_n959_));
  OR2X1    g0574(.A(\req[106] ), .B(\req[105] ), .Y(new_n960_));
  AOI21X1  g0575(.A0(\req[104] ), .A1(new_n956_), .B0(new_n960_), .Y(new_n961_));
  INVX1    g0576(.A(new_n961_), .Y(new_n962_));
  AOI21X1  g0577(.A0(new_n959_), .A1(new_n955_), .B0(new_n962_), .Y(new_n963_));
  INVX1    g0578(.A(\priority[108] ), .Y(new_n964_));
  INVX1    g0579(.A(\req[106] ), .Y(new_n965_));
  AOI21X1  g0580(.A0(new_n965_), .A1(\priority[106] ), .B0(\priority[107] ), .Y(new_n966_));
  NAND2X1  g0581(.A(new_n966_), .B(new_n964_), .Y(new_n967_));
  OR2X1    g0582(.A(\req[109] ), .B(\req[108] ), .Y(new_n968_));
  AOI21X1  g0583(.A0(\req[107] ), .A1(new_n964_), .B0(new_n968_), .Y(new_n969_));
  OAI21X1  g0584(.A0(new_n967_), .A1(new_n963_), .B0(new_n969_), .Y(new_n970_));
  INVX1    g0585(.A(\priority[111] ), .Y(new_n971_));
  INVX1    g0586(.A(\req[109] ), .Y(new_n972_));
  AOI21X1  g0587(.A0(new_n972_), .A1(\priority[109] ), .B0(\priority[110] ), .Y(new_n973_));
  AND2X1   g0588(.A(new_n973_), .B(new_n971_), .Y(new_n974_));
  OR2X1    g0589(.A(\req[112] ), .B(\req[111] ), .Y(new_n975_));
  AOI21X1  g0590(.A0(\req[110] ), .A1(new_n971_), .B0(new_n975_), .Y(new_n976_));
  INVX1    g0591(.A(new_n976_), .Y(new_n977_));
  AOI21X1  g0592(.A0(new_n974_), .A1(new_n970_), .B0(new_n977_), .Y(new_n978_));
  INVX1    g0593(.A(\priority[114] ), .Y(new_n979_));
  INVX1    g0594(.A(\req[112] ), .Y(new_n980_));
  AOI21X1  g0595(.A0(new_n980_), .A1(\priority[112] ), .B0(\priority[113] ), .Y(new_n981_));
  NAND2X1  g0596(.A(new_n981_), .B(new_n979_), .Y(new_n982_));
  OR2X1    g0597(.A(\req[115] ), .B(\req[114] ), .Y(new_n983_));
  AOI21X1  g0598(.A0(\req[113] ), .A1(new_n979_), .B0(new_n983_), .Y(new_n984_));
  OAI21X1  g0599(.A0(new_n982_), .A1(new_n978_), .B0(new_n984_), .Y(new_n985_));
  INVX1    g0600(.A(\priority[117] ), .Y(new_n986_));
  INVX1    g0601(.A(\req[115] ), .Y(new_n987_));
  AOI21X1  g0602(.A0(new_n987_), .A1(\priority[115] ), .B0(\priority[116] ), .Y(new_n988_));
  AND2X1   g0603(.A(new_n988_), .B(new_n986_), .Y(new_n989_));
  OR2X1    g0604(.A(\req[118] ), .B(\req[117] ), .Y(new_n990_));
  AOI21X1  g0605(.A0(\req[116] ), .A1(new_n986_), .B0(new_n990_), .Y(new_n991_));
  INVX1    g0606(.A(new_n991_), .Y(new_n992_));
  AOI21X1  g0607(.A0(new_n989_), .A1(new_n985_), .B0(new_n992_), .Y(new_n993_));
  INVX1    g0608(.A(\priority[120] ), .Y(new_n994_));
  INVX1    g0609(.A(\req[118] ), .Y(new_n995_));
  AOI21X1  g0610(.A0(new_n995_), .A1(\priority[118] ), .B0(\priority[119] ), .Y(new_n996_));
  NAND2X1  g0611(.A(new_n996_), .B(new_n994_), .Y(new_n997_));
  OR2X1    g0612(.A(\req[121] ), .B(\req[120] ), .Y(new_n998_));
  AOI21X1  g0613(.A0(\req[119] ), .A1(new_n994_), .B0(new_n998_), .Y(new_n999_));
  OAI21X1  g0614(.A0(new_n997_), .A1(new_n993_), .B0(new_n999_), .Y(new_n1000_));
  INVX1    g0615(.A(\priority[123] ), .Y(new_n1001_));
  INVX1    g0616(.A(\req[121] ), .Y(new_n1002_));
  AOI21X1  g0617(.A0(new_n1002_), .A1(\priority[121] ), .B0(\priority[122] ), .Y(new_n1003_));
  AND2X1   g0618(.A(new_n1003_), .B(new_n1001_), .Y(new_n1004_));
  OR2X1    g0619(.A(\req[124] ), .B(\req[123] ), .Y(new_n1005_));
  AOI21X1  g0620(.A0(\req[122] ), .A1(new_n1001_), .B0(new_n1005_), .Y(new_n1006_));
  INVX1    g0621(.A(new_n1006_), .Y(new_n1007_));
  AOI21X1  g0622(.A0(new_n1004_), .A1(new_n1000_), .B0(new_n1007_), .Y(new_n1008_));
  INVX1    g0623(.A(\priority[126] ), .Y(new_n1009_));
  INVX1    g0624(.A(\req[124] ), .Y(new_n1010_));
  AOI21X1  g0625(.A0(new_n1010_), .A1(\priority[124] ), .B0(\priority[125] ), .Y(new_n1011_));
  NAND2X1  g0626(.A(new_n1011_), .B(new_n1009_), .Y(new_n1012_));
  OR2X1    g0627(.A(\req[127] ), .B(\req[126] ), .Y(new_n1013_));
  AOI21X1  g0628(.A0(\req[125] ), .A1(new_n1009_), .B0(new_n1013_), .Y(new_n1014_));
  OAI21X1  g0629(.A0(new_n1012_), .A1(new_n1008_), .B0(new_n1014_), .Y(new_n1015_));
  AOI21X1  g0630(.A0(new_n702_), .A1(\priority[127] ), .B0(\priority[0] ), .Y(new_n1016_));
  AND2X1   g0631(.A(new_n1016_), .B(new_n386_), .Y(new_n1017_));
  INVX1    g0632(.A(\req[0] ), .Y(new_n1018_));
  OAI21X1  g0633(.A0(new_n1018_), .A1(\priority[1] ), .B0(\req[1] ), .Y(new_n1019_));
  AOI21X1  g0634(.A0(new_n1017_), .A1(new_n1015_), .B0(new_n1019_), .Y(\grant[1] ));
  OR2X1    g0635(.A(\req[5] ), .B(\req[4] ), .Y(new_n1021_));
  NOR2X1   g0636(.A(new_n1021_), .B(new_n393_), .Y(new_n1022_));
  INVX1    g0637(.A(\priority[7] ), .Y(new_n1023_));
  INVX1    g0638(.A(\req[5] ), .Y(new_n1024_));
  AOI21X1  g0639(.A0(new_n1024_), .A1(\priority[5] ), .B0(\priority[6] ), .Y(new_n1025_));
  NAND2X1  g0640(.A(new_n1025_), .B(new_n1023_), .Y(new_n1026_));
  OR2X1    g0641(.A(\req[8] ), .B(\req[7] ), .Y(new_n1027_));
  AOI21X1  g0642(.A0(\req[6] ), .A1(new_n1023_), .B0(new_n1027_), .Y(new_n1028_));
  OAI21X1  g0643(.A0(new_n1026_), .A1(new_n1022_), .B0(new_n1028_), .Y(new_n1029_));
  INVX1    g0644(.A(\priority[10] ), .Y(new_n1030_));
  INVX1    g0645(.A(\req[8] ), .Y(new_n1031_));
  AOI21X1  g0646(.A0(new_n1031_), .A1(\priority[8] ), .B0(\priority[9] ), .Y(new_n1032_));
  AND2X1   g0647(.A(new_n1032_), .B(new_n1030_), .Y(new_n1033_));
  OR2X1    g0648(.A(\req[11] ), .B(\req[10] ), .Y(new_n1034_));
  AOI21X1  g0649(.A0(\req[9] ), .A1(new_n1030_), .B0(new_n1034_), .Y(new_n1035_));
  INVX1    g0650(.A(new_n1035_), .Y(new_n1036_));
  AOI21X1  g0651(.A0(new_n1033_), .A1(new_n1029_), .B0(new_n1036_), .Y(new_n1037_));
  INVX1    g0652(.A(\priority[13] ), .Y(new_n1038_));
  INVX1    g0653(.A(\req[11] ), .Y(new_n1039_));
  AOI21X1  g0654(.A0(new_n1039_), .A1(\priority[11] ), .B0(\priority[12] ), .Y(new_n1040_));
  NAND2X1  g0655(.A(new_n1040_), .B(new_n1038_), .Y(new_n1041_));
  OR2X1    g0656(.A(\req[14] ), .B(\req[13] ), .Y(new_n1042_));
  AOI21X1  g0657(.A0(\req[12] ), .A1(new_n1038_), .B0(new_n1042_), .Y(new_n1043_));
  OAI21X1  g0658(.A0(new_n1041_), .A1(new_n1037_), .B0(new_n1043_), .Y(new_n1044_));
  INVX1    g0659(.A(\priority[16] ), .Y(new_n1045_));
  INVX1    g0660(.A(\req[14] ), .Y(new_n1046_));
  AOI21X1  g0661(.A0(new_n1046_), .A1(\priority[14] ), .B0(\priority[15] ), .Y(new_n1047_));
  AND2X1   g0662(.A(new_n1047_), .B(new_n1045_), .Y(new_n1048_));
  OR2X1    g0663(.A(\req[17] ), .B(\req[16] ), .Y(new_n1049_));
  AOI21X1  g0664(.A0(\req[15] ), .A1(new_n1045_), .B0(new_n1049_), .Y(new_n1050_));
  INVX1    g0665(.A(new_n1050_), .Y(new_n1051_));
  AOI21X1  g0666(.A0(new_n1048_), .A1(new_n1044_), .B0(new_n1051_), .Y(new_n1052_));
  INVX1    g0667(.A(\priority[19] ), .Y(new_n1053_));
  INVX1    g0668(.A(\req[17] ), .Y(new_n1054_));
  AOI21X1  g0669(.A0(new_n1054_), .A1(\priority[17] ), .B0(\priority[18] ), .Y(new_n1055_));
  NAND2X1  g0670(.A(new_n1055_), .B(new_n1053_), .Y(new_n1056_));
  OR2X1    g0671(.A(\req[20] ), .B(\req[19] ), .Y(new_n1057_));
  AOI21X1  g0672(.A0(\req[18] ), .A1(new_n1053_), .B0(new_n1057_), .Y(new_n1058_));
  OAI21X1  g0673(.A0(new_n1056_), .A1(new_n1052_), .B0(new_n1058_), .Y(new_n1059_));
  INVX1    g0674(.A(\priority[22] ), .Y(new_n1060_));
  INVX1    g0675(.A(\req[20] ), .Y(new_n1061_));
  AOI21X1  g0676(.A0(new_n1061_), .A1(\priority[20] ), .B0(\priority[21] ), .Y(new_n1062_));
  AND2X1   g0677(.A(new_n1062_), .B(new_n1060_), .Y(new_n1063_));
  OR2X1    g0678(.A(\req[23] ), .B(\req[22] ), .Y(new_n1064_));
  AOI21X1  g0679(.A0(\req[21] ), .A1(new_n1060_), .B0(new_n1064_), .Y(new_n1065_));
  INVX1    g0680(.A(new_n1065_), .Y(new_n1066_));
  AOI21X1  g0681(.A0(new_n1063_), .A1(new_n1059_), .B0(new_n1066_), .Y(new_n1067_));
  INVX1    g0682(.A(\priority[25] ), .Y(new_n1068_));
  INVX1    g0683(.A(\req[23] ), .Y(new_n1069_));
  AOI21X1  g0684(.A0(new_n1069_), .A1(\priority[23] ), .B0(\priority[24] ), .Y(new_n1070_));
  NAND2X1  g0685(.A(new_n1070_), .B(new_n1068_), .Y(new_n1071_));
  OR2X1    g0686(.A(\req[26] ), .B(\req[25] ), .Y(new_n1072_));
  AOI21X1  g0687(.A0(\req[24] ), .A1(new_n1068_), .B0(new_n1072_), .Y(new_n1073_));
  OAI21X1  g0688(.A0(new_n1071_), .A1(new_n1067_), .B0(new_n1073_), .Y(new_n1074_));
  INVX1    g0689(.A(\priority[28] ), .Y(new_n1075_));
  INVX1    g0690(.A(\req[26] ), .Y(new_n1076_));
  AOI21X1  g0691(.A0(new_n1076_), .A1(\priority[26] ), .B0(\priority[27] ), .Y(new_n1077_));
  AND2X1   g0692(.A(new_n1077_), .B(new_n1075_), .Y(new_n1078_));
  OR2X1    g0693(.A(\req[29] ), .B(\req[28] ), .Y(new_n1079_));
  AOI21X1  g0694(.A0(\req[27] ), .A1(new_n1075_), .B0(new_n1079_), .Y(new_n1080_));
  INVX1    g0695(.A(new_n1080_), .Y(new_n1081_));
  AOI21X1  g0696(.A0(new_n1078_), .A1(new_n1074_), .B0(new_n1081_), .Y(new_n1082_));
  INVX1    g0697(.A(\priority[31] ), .Y(new_n1083_));
  INVX1    g0698(.A(\req[29] ), .Y(new_n1084_));
  AOI21X1  g0699(.A0(new_n1084_), .A1(\priority[29] ), .B0(\priority[30] ), .Y(new_n1085_));
  NAND2X1  g0700(.A(new_n1085_), .B(new_n1083_), .Y(new_n1086_));
  OR2X1    g0701(.A(\req[32] ), .B(\req[31] ), .Y(new_n1087_));
  AOI21X1  g0702(.A0(\req[30] ), .A1(new_n1083_), .B0(new_n1087_), .Y(new_n1088_));
  OAI21X1  g0703(.A0(new_n1086_), .A1(new_n1082_), .B0(new_n1088_), .Y(new_n1089_));
  INVX1    g0704(.A(\priority[34] ), .Y(new_n1090_));
  INVX1    g0705(.A(\req[32] ), .Y(new_n1091_));
  AOI21X1  g0706(.A0(new_n1091_), .A1(\priority[32] ), .B0(\priority[33] ), .Y(new_n1092_));
  AND2X1   g0707(.A(new_n1092_), .B(new_n1090_), .Y(new_n1093_));
  OR2X1    g0708(.A(\req[35] ), .B(\req[34] ), .Y(new_n1094_));
  AOI21X1  g0709(.A0(\req[33] ), .A1(new_n1090_), .B0(new_n1094_), .Y(new_n1095_));
  INVX1    g0710(.A(new_n1095_), .Y(new_n1096_));
  AOI21X1  g0711(.A0(new_n1093_), .A1(new_n1089_), .B0(new_n1096_), .Y(new_n1097_));
  INVX1    g0712(.A(\priority[37] ), .Y(new_n1098_));
  INVX1    g0713(.A(\req[35] ), .Y(new_n1099_));
  AOI21X1  g0714(.A0(new_n1099_), .A1(\priority[35] ), .B0(\priority[36] ), .Y(new_n1100_));
  NAND2X1  g0715(.A(new_n1100_), .B(new_n1098_), .Y(new_n1101_));
  OR2X1    g0716(.A(\req[38] ), .B(\req[37] ), .Y(new_n1102_));
  AOI21X1  g0717(.A0(\req[36] ), .A1(new_n1098_), .B0(new_n1102_), .Y(new_n1103_));
  OAI21X1  g0718(.A0(new_n1101_), .A1(new_n1097_), .B0(new_n1103_), .Y(new_n1104_));
  INVX1    g0719(.A(\priority[40] ), .Y(new_n1105_));
  INVX1    g0720(.A(\req[38] ), .Y(new_n1106_));
  AOI21X1  g0721(.A0(new_n1106_), .A1(\priority[38] ), .B0(\priority[39] ), .Y(new_n1107_));
  AND2X1   g0722(.A(new_n1107_), .B(new_n1105_), .Y(new_n1108_));
  OR2X1    g0723(.A(\req[41] ), .B(\req[40] ), .Y(new_n1109_));
  AOI21X1  g0724(.A0(\req[39] ), .A1(new_n1105_), .B0(new_n1109_), .Y(new_n1110_));
  INVX1    g0725(.A(new_n1110_), .Y(new_n1111_));
  AOI21X1  g0726(.A0(new_n1108_), .A1(new_n1104_), .B0(new_n1111_), .Y(new_n1112_));
  INVX1    g0727(.A(\priority[43] ), .Y(new_n1113_));
  INVX1    g0728(.A(\req[41] ), .Y(new_n1114_));
  AOI21X1  g0729(.A0(new_n1114_), .A1(\priority[41] ), .B0(\priority[42] ), .Y(new_n1115_));
  NAND2X1  g0730(.A(new_n1115_), .B(new_n1113_), .Y(new_n1116_));
  OR2X1    g0731(.A(\req[44] ), .B(\req[43] ), .Y(new_n1117_));
  AOI21X1  g0732(.A0(\req[42] ), .A1(new_n1113_), .B0(new_n1117_), .Y(new_n1118_));
  OAI21X1  g0733(.A0(new_n1116_), .A1(new_n1112_), .B0(new_n1118_), .Y(new_n1119_));
  INVX1    g0734(.A(\priority[46] ), .Y(new_n1120_));
  INVX1    g0735(.A(\req[44] ), .Y(new_n1121_));
  AOI21X1  g0736(.A0(new_n1121_), .A1(\priority[44] ), .B0(\priority[45] ), .Y(new_n1122_));
  AND2X1   g0737(.A(new_n1122_), .B(new_n1120_), .Y(new_n1123_));
  OR2X1    g0738(.A(\req[47] ), .B(\req[46] ), .Y(new_n1124_));
  AOI21X1  g0739(.A0(\req[45] ), .A1(new_n1120_), .B0(new_n1124_), .Y(new_n1125_));
  INVX1    g0740(.A(new_n1125_), .Y(new_n1126_));
  AOI21X1  g0741(.A0(new_n1123_), .A1(new_n1119_), .B0(new_n1126_), .Y(new_n1127_));
  INVX1    g0742(.A(\priority[49] ), .Y(new_n1128_));
  INVX1    g0743(.A(\req[47] ), .Y(new_n1129_));
  AOI21X1  g0744(.A0(new_n1129_), .A1(\priority[47] ), .B0(\priority[48] ), .Y(new_n1130_));
  NAND2X1  g0745(.A(new_n1130_), .B(new_n1128_), .Y(new_n1131_));
  OR2X1    g0746(.A(\req[50] ), .B(\req[49] ), .Y(new_n1132_));
  AOI21X1  g0747(.A0(\req[48] ), .A1(new_n1128_), .B0(new_n1132_), .Y(new_n1133_));
  OAI21X1  g0748(.A0(new_n1131_), .A1(new_n1127_), .B0(new_n1133_), .Y(new_n1134_));
  INVX1    g0749(.A(\priority[52] ), .Y(new_n1135_));
  INVX1    g0750(.A(\req[50] ), .Y(new_n1136_));
  AOI21X1  g0751(.A0(new_n1136_), .A1(\priority[50] ), .B0(\priority[51] ), .Y(new_n1137_));
  AND2X1   g0752(.A(new_n1137_), .B(new_n1135_), .Y(new_n1138_));
  OR2X1    g0753(.A(\req[53] ), .B(\req[52] ), .Y(new_n1139_));
  AOI21X1  g0754(.A0(\req[51] ), .A1(new_n1135_), .B0(new_n1139_), .Y(new_n1140_));
  INVX1    g0755(.A(new_n1140_), .Y(new_n1141_));
  AOI21X1  g0756(.A0(new_n1138_), .A1(new_n1134_), .B0(new_n1141_), .Y(new_n1142_));
  INVX1    g0757(.A(\priority[55] ), .Y(new_n1143_));
  INVX1    g0758(.A(\req[53] ), .Y(new_n1144_));
  AOI21X1  g0759(.A0(new_n1144_), .A1(\priority[53] ), .B0(\priority[54] ), .Y(new_n1145_));
  NAND2X1  g0760(.A(new_n1145_), .B(new_n1143_), .Y(new_n1146_));
  OR2X1    g0761(.A(\req[56] ), .B(\req[55] ), .Y(new_n1147_));
  AOI21X1  g0762(.A0(\req[54] ), .A1(new_n1143_), .B0(new_n1147_), .Y(new_n1148_));
  OAI21X1  g0763(.A0(new_n1146_), .A1(new_n1142_), .B0(new_n1148_), .Y(new_n1149_));
  INVX1    g0764(.A(\priority[58] ), .Y(new_n1150_));
  INVX1    g0765(.A(\req[56] ), .Y(new_n1151_));
  AOI21X1  g0766(.A0(new_n1151_), .A1(\priority[56] ), .B0(\priority[57] ), .Y(new_n1152_));
  AND2X1   g0767(.A(new_n1152_), .B(new_n1150_), .Y(new_n1153_));
  OR2X1    g0768(.A(\req[59] ), .B(\req[58] ), .Y(new_n1154_));
  AOI21X1  g0769(.A0(\req[57] ), .A1(new_n1150_), .B0(new_n1154_), .Y(new_n1155_));
  INVX1    g0770(.A(new_n1155_), .Y(new_n1156_));
  AOI21X1  g0771(.A0(new_n1153_), .A1(new_n1149_), .B0(new_n1156_), .Y(new_n1157_));
  INVX1    g0772(.A(\priority[61] ), .Y(new_n1158_));
  INVX1    g0773(.A(\req[59] ), .Y(new_n1159_));
  AOI21X1  g0774(.A0(new_n1159_), .A1(\priority[59] ), .B0(\priority[60] ), .Y(new_n1160_));
  NAND2X1  g0775(.A(new_n1160_), .B(new_n1158_), .Y(new_n1161_));
  OR2X1    g0776(.A(\req[62] ), .B(\req[61] ), .Y(new_n1162_));
  AOI21X1  g0777(.A0(\req[60] ), .A1(new_n1158_), .B0(new_n1162_), .Y(new_n1163_));
  OAI21X1  g0778(.A0(new_n1161_), .A1(new_n1157_), .B0(new_n1163_), .Y(new_n1164_));
  INVX1    g0779(.A(\priority[64] ), .Y(new_n1165_));
  INVX1    g0780(.A(\req[62] ), .Y(new_n1166_));
  AOI21X1  g0781(.A0(new_n1166_), .A1(\priority[62] ), .B0(\priority[63] ), .Y(new_n1167_));
  AND2X1   g0782(.A(new_n1167_), .B(new_n1165_), .Y(new_n1168_));
  OR2X1    g0783(.A(\req[65] ), .B(\req[64] ), .Y(new_n1169_));
  AOI21X1  g0784(.A0(\req[63] ), .A1(new_n1165_), .B0(new_n1169_), .Y(new_n1170_));
  INVX1    g0785(.A(new_n1170_), .Y(new_n1171_));
  AOI21X1  g0786(.A0(new_n1168_), .A1(new_n1164_), .B0(new_n1171_), .Y(new_n1172_));
  INVX1    g0787(.A(\priority[67] ), .Y(new_n1173_));
  INVX1    g0788(.A(\req[65] ), .Y(new_n1174_));
  AOI21X1  g0789(.A0(new_n1174_), .A1(\priority[65] ), .B0(\priority[66] ), .Y(new_n1175_));
  NAND2X1  g0790(.A(new_n1175_), .B(new_n1173_), .Y(new_n1176_));
  OR2X1    g0791(.A(\req[68] ), .B(\req[67] ), .Y(new_n1177_));
  AOI21X1  g0792(.A0(\req[66] ), .A1(new_n1173_), .B0(new_n1177_), .Y(new_n1178_));
  OAI21X1  g0793(.A0(new_n1176_), .A1(new_n1172_), .B0(new_n1178_), .Y(new_n1179_));
  INVX1    g0794(.A(\priority[70] ), .Y(new_n1180_));
  INVX1    g0795(.A(\req[68] ), .Y(new_n1181_));
  AOI21X1  g0796(.A0(new_n1181_), .A1(\priority[68] ), .B0(\priority[69] ), .Y(new_n1182_));
  AND2X1   g0797(.A(new_n1182_), .B(new_n1180_), .Y(new_n1183_));
  OR2X1    g0798(.A(\req[71] ), .B(\req[70] ), .Y(new_n1184_));
  AOI21X1  g0799(.A0(\req[69] ), .A1(new_n1180_), .B0(new_n1184_), .Y(new_n1185_));
  INVX1    g0800(.A(new_n1185_), .Y(new_n1186_));
  AOI21X1  g0801(.A0(new_n1183_), .A1(new_n1179_), .B0(new_n1186_), .Y(new_n1187_));
  INVX1    g0802(.A(\priority[73] ), .Y(new_n1188_));
  INVX1    g0803(.A(\req[71] ), .Y(new_n1189_));
  AOI21X1  g0804(.A0(new_n1189_), .A1(\priority[71] ), .B0(\priority[72] ), .Y(new_n1190_));
  NAND2X1  g0805(.A(new_n1190_), .B(new_n1188_), .Y(new_n1191_));
  OR2X1    g0806(.A(\req[74] ), .B(\req[73] ), .Y(new_n1192_));
  AOI21X1  g0807(.A0(\req[72] ), .A1(new_n1188_), .B0(new_n1192_), .Y(new_n1193_));
  OAI21X1  g0808(.A0(new_n1191_), .A1(new_n1187_), .B0(new_n1193_), .Y(new_n1194_));
  INVX1    g0809(.A(\priority[76] ), .Y(new_n1195_));
  INVX1    g0810(.A(\req[74] ), .Y(new_n1196_));
  AOI21X1  g0811(.A0(new_n1196_), .A1(\priority[74] ), .B0(\priority[75] ), .Y(new_n1197_));
  AND2X1   g0812(.A(new_n1197_), .B(new_n1195_), .Y(new_n1198_));
  OR2X1    g0813(.A(\req[77] ), .B(\req[76] ), .Y(new_n1199_));
  AOI21X1  g0814(.A0(\req[75] ), .A1(new_n1195_), .B0(new_n1199_), .Y(new_n1200_));
  INVX1    g0815(.A(new_n1200_), .Y(new_n1201_));
  AOI21X1  g0816(.A0(new_n1198_), .A1(new_n1194_), .B0(new_n1201_), .Y(new_n1202_));
  INVX1    g0817(.A(\priority[79] ), .Y(new_n1203_));
  INVX1    g0818(.A(\req[77] ), .Y(new_n1204_));
  AOI21X1  g0819(.A0(new_n1204_), .A1(\priority[77] ), .B0(\priority[78] ), .Y(new_n1205_));
  NAND2X1  g0820(.A(new_n1205_), .B(new_n1203_), .Y(new_n1206_));
  OR2X1    g0821(.A(\req[80] ), .B(\req[79] ), .Y(new_n1207_));
  AOI21X1  g0822(.A0(\req[78] ), .A1(new_n1203_), .B0(new_n1207_), .Y(new_n1208_));
  OAI21X1  g0823(.A0(new_n1206_), .A1(new_n1202_), .B0(new_n1208_), .Y(new_n1209_));
  INVX1    g0824(.A(\priority[82] ), .Y(new_n1210_));
  INVX1    g0825(.A(\req[80] ), .Y(new_n1211_));
  AOI21X1  g0826(.A0(new_n1211_), .A1(\priority[80] ), .B0(\priority[81] ), .Y(new_n1212_));
  AND2X1   g0827(.A(new_n1212_), .B(new_n1210_), .Y(new_n1213_));
  OR2X1    g0828(.A(\req[83] ), .B(\req[82] ), .Y(new_n1214_));
  AOI21X1  g0829(.A0(\req[81] ), .A1(new_n1210_), .B0(new_n1214_), .Y(new_n1215_));
  INVX1    g0830(.A(new_n1215_), .Y(new_n1216_));
  AOI21X1  g0831(.A0(new_n1213_), .A1(new_n1209_), .B0(new_n1216_), .Y(new_n1217_));
  INVX1    g0832(.A(\priority[85] ), .Y(new_n1218_));
  INVX1    g0833(.A(\req[83] ), .Y(new_n1219_));
  AOI21X1  g0834(.A0(new_n1219_), .A1(\priority[83] ), .B0(\priority[84] ), .Y(new_n1220_));
  NAND2X1  g0835(.A(new_n1220_), .B(new_n1218_), .Y(new_n1221_));
  OR2X1    g0836(.A(\req[86] ), .B(\req[85] ), .Y(new_n1222_));
  AOI21X1  g0837(.A0(\req[84] ), .A1(new_n1218_), .B0(new_n1222_), .Y(new_n1223_));
  OAI21X1  g0838(.A0(new_n1221_), .A1(new_n1217_), .B0(new_n1223_), .Y(new_n1224_));
  INVX1    g0839(.A(\priority[88] ), .Y(new_n1225_));
  INVX1    g0840(.A(\req[86] ), .Y(new_n1226_));
  AOI21X1  g0841(.A0(new_n1226_), .A1(\priority[86] ), .B0(\priority[87] ), .Y(new_n1227_));
  AND2X1   g0842(.A(new_n1227_), .B(new_n1225_), .Y(new_n1228_));
  OR2X1    g0843(.A(\req[89] ), .B(\req[88] ), .Y(new_n1229_));
  AOI21X1  g0844(.A0(\req[87] ), .A1(new_n1225_), .B0(new_n1229_), .Y(new_n1230_));
  INVX1    g0845(.A(new_n1230_), .Y(new_n1231_));
  AOI21X1  g0846(.A0(new_n1228_), .A1(new_n1224_), .B0(new_n1231_), .Y(new_n1232_));
  INVX1    g0847(.A(\priority[91] ), .Y(new_n1233_));
  INVX1    g0848(.A(\req[89] ), .Y(new_n1234_));
  AOI21X1  g0849(.A0(new_n1234_), .A1(\priority[89] ), .B0(\priority[90] ), .Y(new_n1235_));
  NAND2X1  g0850(.A(new_n1235_), .B(new_n1233_), .Y(new_n1236_));
  OR2X1    g0851(.A(\req[92] ), .B(\req[91] ), .Y(new_n1237_));
  AOI21X1  g0852(.A0(\req[90] ), .A1(new_n1233_), .B0(new_n1237_), .Y(new_n1238_));
  OAI21X1  g0853(.A0(new_n1236_), .A1(new_n1232_), .B0(new_n1238_), .Y(new_n1239_));
  INVX1    g0854(.A(\priority[94] ), .Y(new_n1240_));
  INVX1    g0855(.A(\req[92] ), .Y(new_n1241_));
  AOI21X1  g0856(.A0(new_n1241_), .A1(\priority[92] ), .B0(\priority[93] ), .Y(new_n1242_));
  AND2X1   g0857(.A(new_n1242_), .B(new_n1240_), .Y(new_n1243_));
  OR2X1    g0858(.A(\req[95] ), .B(\req[94] ), .Y(new_n1244_));
  AOI21X1  g0859(.A0(\req[93] ), .A1(new_n1240_), .B0(new_n1244_), .Y(new_n1245_));
  INVX1    g0860(.A(new_n1245_), .Y(new_n1246_));
  AOI21X1  g0861(.A0(new_n1243_), .A1(new_n1239_), .B0(new_n1246_), .Y(new_n1247_));
  INVX1    g0862(.A(\priority[97] ), .Y(new_n1248_));
  INVX1    g0863(.A(\req[95] ), .Y(new_n1249_));
  AOI21X1  g0864(.A0(new_n1249_), .A1(\priority[95] ), .B0(\priority[96] ), .Y(new_n1250_));
  NAND2X1  g0865(.A(new_n1250_), .B(new_n1248_), .Y(new_n1251_));
  OR2X1    g0866(.A(\req[98] ), .B(\req[97] ), .Y(new_n1252_));
  AOI21X1  g0867(.A0(\req[96] ), .A1(new_n1248_), .B0(new_n1252_), .Y(new_n1253_));
  OAI21X1  g0868(.A0(new_n1251_), .A1(new_n1247_), .B0(new_n1253_), .Y(new_n1254_));
  INVX1    g0869(.A(\priority[100] ), .Y(new_n1255_));
  INVX1    g0870(.A(\req[98] ), .Y(new_n1256_));
  AOI21X1  g0871(.A0(new_n1256_), .A1(\priority[98] ), .B0(\priority[99] ), .Y(new_n1257_));
  AND2X1   g0872(.A(new_n1257_), .B(new_n1255_), .Y(new_n1258_));
  OR2X1    g0873(.A(\req[101] ), .B(\req[100] ), .Y(new_n1259_));
  AOI21X1  g0874(.A0(\req[99] ), .A1(new_n1255_), .B0(new_n1259_), .Y(new_n1260_));
  INVX1    g0875(.A(new_n1260_), .Y(new_n1261_));
  AOI21X1  g0876(.A0(new_n1258_), .A1(new_n1254_), .B0(new_n1261_), .Y(new_n1262_));
  INVX1    g0877(.A(\priority[103] ), .Y(new_n1263_));
  INVX1    g0878(.A(\req[101] ), .Y(new_n1264_));
  AOI21X1  g0879(.A0(new_n1264_), .A1(\priority[101] ), .B0(\priority[102] ), .Y(new_n1265_));
  NAND2X1  g0880(.A(new_n1265_), .B(new_n1263_), .Y(new_n1266_));
  OR2X1    g0881(.A(\req[104] ), .B(\req[103] ), .Y(new_n1267_));
  AOI21X1  g0882(.A0(\req[102] ), .A1(new_n1263_), .B0(new_n1267_), .Y(new_n1268_));
  OAI21X1  g0883(.A0(new_n1266_), .A1(new_n1262_), .B0(new_n1268_), .Y(new_n1269_));
  INVX1    g0884(.A(\priority[106] ), .Y(new_n1270_));
  INVX1    g0885(.A(\req[104] ), .Y(new_n1271_));
  AOI21X1  g0886(.A0(new_n1271_), .A1(\priority[104] ), .B0(\priority[105] ), .Y(new_n1272_));
  AND2X1   g0887(.A(new_n1272_), .B(new_n1270_), .Y(new_n1273_));
  OR2X1    g0888(.A(\req[107] ), .B(\req[106] ), .Y(new_n1274_));
  AOI21X1  g0889(.A0(\req[105] ), .A1(new_n1270_), .B0(new_n1274_), .Y(new_n1275_));
  INVX1    g0890(.A(new_n1275_), .Y(new_n1276_));
  AOI21X1  g0891(.A0(new_n1273_), .A1(new_n1269_), .B0(new_n1276_), .Y(new_n1277_));
  INVX1    g0892(.A(\priority[109] ), .Y(new_n1278_));
  INVX1    g0893(.A(\req[107] ), .Y(new_n1279_));
  AOI21X1  g0894(.A0(new_n1279_), .A1(\priority[107] ), .B0(\priority[108] ), .Y(new_n1280_));
  NAND2X1  g0895(.A(new_n1280_), .B(new_n1278_), .Y(new_n1281_));
  OR2X1    g0896(.A(\req[110] ), .B(\req[109] ), .Y(new_n1282_));
  AOI21X1  g0897(.A0(\req[108] ), .A1(new_n1278_), .B0(new_n1282_), .Y(new_n1283_));
  OAI21X1  g0898(.A0(new_n1281_), .A1(new_n1277_), .B0(new_n1283_), .Y(new_n1284_));
  INVX1    g0899(.A(\priority[112] ), .Y(new_n1285_));
  INVX1    g0900(.A(\req[110] ), .Y(new_n1286_));
  AOI21X1  g0901(.A0(new_n1286_), .A1(\priority[110] ), .B0(\priority[111] ), .Y(new_n1287_));
  AND2X1   g0902(.A(new_n1287_), .B(new_n1285_), .Y(new_n1288_));
  OR2X1    g0903(.A(\req[113] ), .B(\req[112] ), .Y(new_n1289_));
  AOI21X1  g0904(.A0(\req[111] ), .A1(new_n1285_), .B0(new_n1289_), .Y(new_n1290_));
  INVX1    g0905(.A(new_n1290_), .Y(new_n1291_));
  AOI21X1  g0906(.A0(new_n1288_), .A1(new_n1284_), .B0(new_n1291_), .Y(new_n1292_));
  INVX1    g0907(.A(\priority[115] ), .Y(new_n1293_));
  INVX1    g0908(.A(\req[113] ), .Y(new_n1294_));
  AOI21X1  g0909(.A0(new_n1294_), .A1(\priority[113] ), .B0(\priority[114] ), .Y(new_n1295_));
  NAND2X1  g0910(.A(new_n1295_), .B(new_n1293_), .Y(new_n1296_));
  OR2X1    g0911(.A(\req[116] ), .B(\req[115] ), .Y(new_n1297_));
  AOI21X1  g0912(.A0(\req[114] ), .A1(new_n1293_), .B0(new_n1297_), .Y(new_n1298_));
  OAI21X1  g0913(.A0(new_n1296_), .A1(new_n1292_), .B0(new_n1298_), .Y(new_n1299_));
  INVX1    g0914(.A(\priority[118] ), .Y(new_n1300_));
  INVX1    g0915(.A(\req[116] ), .Y(new_n1301_));
  AOI21X1  g0916(.A0(new_n1301_), .A1(\priority[116] ), .B0(\priority[117] ), .Y(new_n1302_));
  AND2X1   g0917(.A(new_n1302_), .B(new_n1300_), .Y(new_n1303_));
  OR2X1    g0918(.A(\req[119] ), .B(\req[118] ), .Y(new_n1304_));
  AOI21X1  g0919(.A0(\req[117] ), .A1(new_n1300_), .B0(new_n1304_), .Y(new_n1305_));
  INVX1    g0920(.A(new_n1305_), .Y(new_n1306_));
  AOI21X1  g0921(.A0(new_n1303_), .A1(new_n1299_), .B0(new_n1306_), .Y(new_n1307_));
  INVX1    g0922(.A(\priority[121] ), .Y(new_n1308_));
  INVX1    g0923(.A(\req[119] ), .Y(new_n1309_));
  AOI21X1  g0924(.A0(new_n1309_), .A1(\priority[119] ), .B0(\priority[120] ), .Y(new_n1310_));
  NAND2X1  g0925(.A(new_n1310_), .B(new_n1308_), .Y(new_n1311_));
  OR2X1    g0926(.A(\req[122] ), .B(\req[121] ), .Y(new_n1312_));
  AOI21X1  g0927(.A0(\req[120] ), .A1(new_n1308_), .B0(new_n1312_), .Y(new_n1313_));
  OAI21X1  g0928(.A0(new_n1311_), .A1(new_n1307_), .B0(new_n1313_), .Y(new_n1314_));
  INVX1    g0929(.A(\priority[124] ), .Y(new_n1315_));
  INVX1    g0930(.A(\req[122] ), .Y(new_n1316_));
  AOI21X1  g0931(.A0(new_n1316_), .A1(\priority[122] ), .B0(\priority[123] ), .Y(new_n1317_));
  AND2X1   g0932(.A(new_n1317_), .B(new_n1315_), .Y(new_n1318_));
  OR2X1    g0933(.A(\req[125] ), .B(\req[124] ), .Y(new_n1319_));
  AOI21X1  g0934(.A0(\req[123] ), .A1(new_n1315_), .B0(new_n1319_), .Y(new_n1320_));
  INVX1    g0935(.A(new_n1320_), .Y(new_n1321_));
  AOI21X1  g0936(.A0(new_n1318_), .A1(new_n1314_), .B0(new_n1321_), .Y(new_n1322_));
  INVX1    g0937(.A(\priority[127] ), .Y(new_n1323_));
  INVX1    g0938(.A(\req[125] ), .Y(new_n1324_));
  AOI21X1  g0939(.A0(new_n1324_), .A1(\priority[125] ), .B0(\priority[126] ), .Y(new_n1325_));
  NAND2X1  g0940(.A(new_n1325_), .B(new_n1323_), .Y(new_n1326_));
  OR2X1    g0941(.A(\req[127] ), .B(\req[0] ), .Y(new_n1327_));
  AOI21X1  g0942(.A0(\req[126] ), .A1(new_n1323_), .B0(new_n1327_), .Y(new_n1328_));
  OAI21X1  g0943(.A0(new_n1326_), .A1(new_n1322_), .B0(new_n1328_), .Y(new_n1329_));
  AOI21X1  g0944(.A0(new_n1018_), .A1(\priority[0] ), .B0(\priority[1] ), .Y(new_n1330_));
  AND2X1   g0945(.A(new_n1330_), .B(new_n387_), .Y(new_n1331_));
  INVX1    g0946(.A(\req[1] ), .Y(new_n1332_));
  OAI21X1  g0947(.A0(new_n1332_), .A1(\priority[2] ), .B0(\req[2] ), .Y(new_n1333_));
  AOI21X1  g0948(.A0(new_n1331_), .A1(new_n1329_), .B0(new_n1333_), .Y(\grant[2] ));
  NAND2X1  g0949(.A(new_n700_), .B(new_n698_), .Y(new_n1335_));
  AND2X1   g0950(.A(new_n693_), .B(new_n691_), .Y(new_n1336_));
  INVX1    g0951(.A(new_n696_), .Y(new_n1337_));
  NAND2X1  g0952(.A(new_n685_), .B(new_n683_), .Y(new_n1338_));
  AND2X1   g0953(.A(new_n678_), .B(new_n676_), .Y(new_n1339_));
  INVX1    g0954(.A(new_n681_), .Y(new_n1340_));
  NAND2X1  g0955(.A(new_n670_), .B(new_n668_), .Y(new_n1341_));
  AND2X1   g0956(.A(new_n663_), .B(new_n661_), .Y(new_n1342_));
  INVX1    g0957(.A(new_n666_), .Y(new_n1343_));
  NAND2X1  g0958(.A(new_n655_), .B(new_n653_), .Y(new_n1344_));
  AND2X1   g0959(.A(new_n648_), .B(new_n646_), .Y(new_n1345_));
  INVX1    g0960(.A(new_n651_), .Y(new_n1346_));
  NAND2X1  g0961(.A(new_n640_), .B(new_n638_), .Y(new_n1347_));
  AND2X1   g0962(.A(new_n633_), .B(new_n631_), .Y(new_n1348_));
  INVX1    g0963(.A(new_n636_), .Y(new_n1349_));
  NAND2X1  g0964(.A(new_n625_), .B(new_n623_), .Y(new_n1350_));
  AND2X1   g0965(.A(new_n618_), .B(new_n616_), .Y(new_n1351_));
  INVX1    g0966(.A(new_n621_), .Y(new_n1352_));
  NAND2X1  g0967(.A(new_n610_), .B(new_n608_), .Y(new_n1353_));
  AND2X1   g0968(.A(new_n603_), .B(new_n601_), .Y(new_n1354_));
  INVX1    g0969(.A(new_n606_), .Y(new_n1355_));
  NAND2X1  g0970(.A(new_n595_), .B(new_n593_), .Y(new_n1356_));
  AND2X1   g0971(.A(new_n588_), .B(new_n586_), .Y(new_n1357_));
  INVX1    g0972(.A(new_n591_), .Y(new_n1358_));
  NAND2X1  g0973(.A(new_n580_), .B(new_n578_), .Y(new_n1359_));
  AND2X1   g0974(.A(new_n573_), .B(new_n571_), .Y(new_n1360_));
  INVX1    g0975(.A(new_n576_), .Y(new_n1361_));
  NAND2X1  g0976(.A(new_n565_), .B(new_n563_), .Y(new_n1362_));
  AND2X1   g0977(.A(new_n558_), .B(new_n556_), .Y(new_n1363_));
  INVX1    g0978(.A(new_n561_), .Y(new_n1364_));
  NAND2X1  g0979(.A(new_n550_), .B(new_n548_), .Y(new_n1365_));
  AND2X1   g0980(.A(new_n543_), .B(new_n541_), .Y(new_n1366_));
  INVX1    g0981(.A(new_n546_), .Y(new_n1367_));
  NAND2X1  g0982(.A(new_n535_), .B(new_n533_), .Y(new_n1368_));
  AND2X1   g0983(.A(new_n528_), .B(new_n526_), .Y(new_n1369_));
  INVX1    g0984(.A(new_n531_), .Y(new_n1370_));
  NAND2X1  g0985(.A(new_n520_), .B(new_n518_), .Y(new_n1371_));
  AND2X1   g0986(.A(new_n513_), .B(new_n511_), .Y(new_n1372_));
  INVX1    g0987(.A(new_n516_), .Y(new_n1373_));
  NAND2X1  g0988(.A(new_n505_), .B(new_n503_), .Y(new_n1374_));
  AND2X1   g0989(.A(new_n498_), .B(new_n496_), .Y(new_n1375_));
  INVX1    g0990(.A(new_n501_), .Y(new_n1376_));
  NAND2X1  g0991(.A(new_n490_), .B(new_n488_), .Y(new_n1377_));
  AND2X1   g0992(.A(new_n483_), .B(new_n481_), .Y(new_n1378_));
  INVX1    g0993(.A(new_n486_), .Y(new_n1379_));
  NAND2X1  g0994(.A(new_n475_), .B(new_n473_), .Y(new_n1380_));
  AND2X1   g0995(.A(new_n468_), .B(new_n466_), .Y(new_n1381_));
  INVX1    g0996(.A(new_n471_), .Y(new_n1382_));
  NAND2X1  g0997(.A(new_n460_), .B(new_n458_), .Y(new_n1383_));
  AND2X1   g0998(.A(new_n453_), .B(new_n451_), .Y(new_n1384_));
  INVX1    g0999(.A(new_n456_), .Y(new_n1385_));
  NAND2X1  g1000(.A(new_n445_), .B(new_n443_), .Y(new_n1386_));
  AND2X1   g1001(.A(new_n438_), .B(new_n436_), .Y(new_n1387_));
  INVX1    g1002(.A(new_n441_), .Y(new_n1388_));
  NAND2X1  g1003(.A(new_n430_), .B(new_n428_), .Y(new_n1389_));
  AND2X1   g1004(.A(new_n423_), .B(new_n421_), .Y(new_n1390_));
  INVX1    g1005(.A(new_n426_), .Y(new_n1391_));
  NAND2X1  g1006(.A(new_n415_), .B(new_n413_), .Y(new_n1392_));
  AND2X1   g1007(.A(new_n408_), .B(new_n406_), .Y(new_n1393_));
  INVX1    g1008(.A(new_n411_), .Y(new_n1394_));
  NAND2X1  g1009(.A(new_n400_), .B(new_n398_), .Y(new_n1395_));
  NOR2X1   g1010(.A(new_n711_), .B(new_n395_), .Y(new_n1396_));
  OAI21X1  g1011(.A0(new_n1396_), .A1(new_n1395_), .B0(new_n403_), .Y(new_n1397_));
  AOI21X1  g1012(.A0(new_n1397_), .A1(new_n1393_), .B0(new_n1394_), .Y(new_n1398_));
  OAI21X1  g1013(.A0(new_n1398_), .A1(new_n1392_), .B0(new_n418_), .Y(new_n1399_));
  AOI21X1  g1014(.A0(new_n1399_), .A1(new_n1390_), .B0(new_n1391_), .Y(new_n1400_));
  OAI21X1  g1015(.A0(new_n1400_), .A1(new_n1389_), .B0(new_n433_), .Y(new_n1401_));
  AOI21X1  g1016(.A0(new_n1401_), .A1(new_n1387_), .B0(new_n1388_), .Y(new_n1402_));
  OAI21X1  g1017(.A0(new_n1402_), .A1(new_n1386_), .B0(new_n448_), .Y(new_n1403_));
  AOI21X1  g1018(.A0(new_n1403_), .A1(new_n1384_), .B0(new_n1385_), .Y(new_n1404_));
  OAI21X1  g1019(.A0(new_n1404_), .A1(new_n1383_), .B0(new_n463_), .Y(new_n1405_));
  AOI21X1  g1020(.A0(new_n1405_), .A1(new_n1381_), .B0(new_n1382_), .Y(new_n1406_));
  OAI21X1  g1021(.A0(new_n1406_), .A1(new_n1380_), .B0(new_n478_), .Y(new_n1407_));
  AOI21X1  g1022(.A0(new_n1407_), .A1(new_n1378_), .B0(new_n1379_), .Y(new_n1408_));
  OAI21X1  g1023(.A0(new_n1408_), .A1(new_n1377_), .B0(new_n493_), .Y(new_n1409_));
  AOI21X1  g1024(.A0(new_n1409_), .A1(new_n1375_), .B0(new_n1376_), .Y(new_n1410_));
  OAI21X1  g1025(.A0(new_n1410_), .A1(new_n1374_), .B0(new_n508_), .Y(new_n1411_));
  AOI21X1  g1026(.A0(new_n1411_), .A1(new_n1372_), .B0(new_n1373_), .Y(new_n1412_));
  OAI21X1  g1027(.A0(new_n1412_), .A1(new_n1371_), .B0(new_n523_), .Y(new_n1413_));
  AOI21X1  g1028(.A0(new_n1413_), .A1(new_n1369_), .B0(new_n1370_), .Y(new_n1414_));
  OAI21X1  g1029(.A0(new_n1414_), .A1(new_n1368_), .B0(new_n538_), .Y(new_n1415_));
  AOI21X1  g1030(.A0(new_n1415_), .A1(new_n1366_), .B0(new_n1367_), .Y(new_n1416_));
  OAI21X1  g1031(.A0(new_n1416_), .A1(new_n1365_), .B0(new_n553_), .Y(new_n1417_));
  AOI21X1  g1032(.A0(new_n1417_), .A1(new_n1363_), .B0(new_n1364_), .Y(new_n1418_));
  OAI21X1  g1033(.A0(new_n1418_), .A1(new_n1362_), .B0(new_n568_), .Y(new_n1419_));
  AOI21X1  g1034(.A0(new_n1419_), .A1(new_n1360_), .B0(new_n1361_), .Y(new_n1420_));
  OAI21X1  g1035(.A0(new_n1420_), .A1(new_n1359_), .B0(new_n583_), .Y(new_n1421_));
  AOI21X1  g1036(.A0(new_n1421_), .A1(new_n1357_), .B0(new_n1358_), .Y(new_n1422_));
  OAI21X1  g1037(.A0(new_n1422_), .A1(new_n1356_), .B0(new_n598_), .Y(new_n1423_));
  AOI21X1  g1038(.A0(new_n1423_), .A1(new_n1354_), .B0(new_n1355_), .Y(new_n1424_));
  OAI21X1  g1039(.A0(new_n1424_), .A1(new_n1353_), .B0(new_n613_), .Y(new_n1425_));
  AOI21X1  g1040(.A0(new_n1425_), .A1(new_n1351_), .B0(new_n1352_), .Y(new_n1426_));
  OAI21X1  g1041(.A0(new_n1426_), .A1(new_n1350_), .B0(new_n628_), .Y(new_n1427_));
  AOI21X1  g1042(.A0(new_n1427_), .A1(new_n1348_), .B0(new_n1349_), .Y(new_n1428_));
  OAI21X1  g1043(.A0(new_n1428_), .A1(new_n1347_), .B0(new_n643_), .Y(new_n1429_));
  AOI21X1  g1044(.A0(new_n1429_), .A1(new_n1345_), .B0(new_n1346_), .Y(new_n1430_));
  OAI21X1  g1045(.A0(new_n1430_), .A1(new_n1344_), .B0(new_n658_), .Y(new_n1431_));
  AOI21X1  g1046(.A0(new_n1431_), .A1(new_n1342_), .B0(new_n1343_), .Y(new_n1432_));
  OAI21X1  g1047(.A0(new_n1432_), .A1(new_n1341_), .B0(new_n673_), .Y(new_n1433_));
  AOI21X1  g1048(.A0(new_n1433_), .A1(new_n1339_), .B0(new_n1340_), .Y(new_n1434_));
  OAI21X1  g1049(.A0(new_n1434_), .A1(new_n1338_), .B0(new_n688_), .Y(new_n1435_));
  AOI21X1  g1050(.A0(new_n1435_), .A1(new_n1336_), .B0(new_n1337_), .Y(new_n1436_));
  OR2X1    g1051(.A(\req[1] ), .B(\req[0] ), .Y(new_n1437_));
  AOI21X1  g1052(.A0(\req[127] ), .A1(new_n698_), .B0(new_n1437_), .Y(new_n1438_));
  OAI21X1  g1053(.A0(new_n1436_), .A1(new_n1335_), .B0(new_n1438_), .Y(new_n1439_));
  NOR2X1   g1054(.A(new_n388_), .B(\priority[3] ), .Y(new_n1440_));
  INVX1    g1055(.A(\req[2] ), .Y(new_n1441_));
  OAI21X1  g1056(.A0(new_n1441_), .A1(\priority[3] ), .B0(\req[3] ), .Y(new_n1442_));
  AOI21X1  g1057(.A0(new_n1440_), .A1(new_n1439_), .B0(new_n1442_), .Y(\grant[3] ));
  NAND2X1  g1058(.A(new_n1016_), .B(new_n386_), .Y(new_n1444_));
  AND2X1   g1059(.A(new_n1011_), .B(new_n1009_), .Y(new_n1445_));
  INVX1    g1060(.A(new_n1014_), .Y(new_n1446_));
  NAND2X1  g1061(.A(new_n1003_), .B(new_n1001_), .Y(new_n1447_));
  AND2X1   g1062(.A(new_n996_), .B(new_n994_), .Y(new_n1448_));
  INVX1    g1063(.A(new_n999_), .Y(new_n1449_));
  NAND2X1  g1064(.A(new_n988_), .B(new_n986_), .Y(new_n1450_));
  AND2X1   g1065(.A(new_n981_), .B(new_n979_), .Y(new_n1451_));
  INVX1    g1066(.A(new_n984_), .Y(new_n1452_));
  NAND2X1  g1067(.A(new_n973_), .B(new_n971_), .Y(new_n1453_));
  AND2X1   g1068(.A(new_n966_), .B(new_n964_), .Y(new_n1454_));
  INVX1    g1069(.A(new_n969_), .Y(new_n1455_));
  NAND2X1  g1070(.A(new_n958_), .B(new_n956_), .Y(new_n1456_));
  AND2X1   g1071(.A(new_n951_), .B(new_n949_), .Y(new_n1457_));
  INVX1    g1072(.A(new_n954_), .Y(new_n1458_));
  NAND2X1  g1073(.A(new_n943_), .B(new_n941_), .Y(new_n1459_));
  AND2X1   g1074(.A(new_n936_), .B(new_n934_), .Y(new_n1460_));
  INVX1    g1075(.A(new_n939_), .Y(new_n1461_));
  NAND2X1  g1076(.A(new_n928_), .B(new_n926_), .Y(new_n1462_));
  AND2X1   g1077(.A(new_n921_), .B(new_n919_), .Y(new_n1463_));
  INVX1    g1078(.A(new_n924_), .Y(new_n1464_));
  NAND2X1  g1079(.A(new_n913_), .B(new_n911_), .Y(new_n1465_));
  AND2X1   g1080(.A(new_n906_), .B(new_n904_), .Y(new_n1466_));
  INVX1    g1081(.A(new_n909_), .Y(new_n1467_));
  NAND2X1  g1082(.A(new_n898_), .B(new_n896_), .Y(new_n1468_));
  AND2X1   g1083(.A(new_n891_), .B(new_n889_), .Y(new_n1469_));
  INVX1    g1084(.A(new_n894_), .Y(new_n1470_));
  NAND2X1  g1085(.A(new_n883_), .B(new_n881_), .Y(new_n1471_));
  AND2X1   g1086(.A(new_n876_), .B(new_n874_), .Y(new_n1472_));
  INVX1    g1087(.A(new_n879_), .Y(new_n1473_));
  NAND2X1  g1088(.A(new_n868_), .B(new_n866_), .Y(new_n1474_));
  AND2X1   g1089(.A(new_n861_), .B(new_n859_), .Y(new_n1475_));
  INVX1    g1090(.A(new_n864_), .Y(new_n1476_));
  NAND2X1  g1091(.A(new_n853_), .B(new_n851_), .Y(new_n1477_));
  AND2X1   g1092(.A(new_n846_), .B(new_n844_), .Y(new_n1478_));
  INVX1    g1093(.A(new_n849_), .Y(new_n1479_));
  NAND2X1  g1094(.A(new_n838_), .B(new_n836_), .Y(new_n1480_));
  AND2X1   g1095(.A(new_n831_), .B(new_n829_), .Y(new_n1481_));
  INVX1    g1096(.A(new_n834_), .Y(new_n1482_));
  NAND2X1  g1097(.A(new_n823_), .B(new_n821_), .Y(new_n1483_));
  AND2X1   g1098(.A(new_n816_), .B(new_n814_), .Y(new_n1484_));
  INVX1    g1099(.A(new_n819_), .Y(new_n1485_));
  NAND2X1  g1100(.A(new_n808_), .B(new_n806_), .Y(new_n1486_));
  AND2X1   g1101(.A(new_n801_), .B(new_n799_), .Y(new_n1487_));
  INVX1    g1102(.A(new_n804_), .Y(new_n1488_));
  NAND2X1  g1103(.A(new_n793_), .B(new_n791_), .Y(new_n1489_));
  AND2X1   g1104(.A(new_n786_), .B(new_n784_), .Y(new_n1490_));
  INVX1    g1105(.A(new_n789_), .Y(new_n1491_));
  NAND2X1  g1106(.A(new_n778_), .B(new_n776_), .Y(new_n1492_));
  AND2X1   g1107(.A(new_n771_), .B(new_n769_), .Y(new_n1493_));
  INVX1    g1108(.A(new_n774_), .Y(new_n1494_));
  NAND2X1  g1109(.A(new_n763_), .B(new_n761_), .Y(new_n1495_));
  AND2X1   g1110(.A(new_n756_), .B(new_n754_), .Y(new_n1496_));
  INVX1    g1111(.A(new_n759_), .Y(new_n1497_));
  NAND2X1  g1112(.A(new_n748_), .B(new_n746_), .Y(new_n1498_));
  AND2X1   g1113(.A(new_n741_), .B(new_n739_), .Y(new_n1499_));
  INVX1    g1114(.A(new_n744_), .Y(new_n1500_));
  NAND2X1  g1115(.A(new_n733_), .B(new_n731_), .Y(new_n1501_));
  AND2X1   g1116(.A(new_n726_), .B(new_n724_), .Y(new_n1502_));
  INVX1    g1117(.A(new_n729_), .Y(new_n1503_));
  NAND2X1  g1118(.A(new_n718_), .B(new_n716_), .Y(new_n1504_));
  NOR2X1   g1119(.A(new_n1025_), .B(new_n713_), .Y(new_n1505_));
  OAI21X1  g1120(.A0(new_n1505_), .A1(new_n1504_), .B0(new_n721_), .Y(new_n1506_));
  AOI21X1  g1121(.A0(new_n1506_), .A1(new_n1502_), .B0(new_n1503_), .Y(new_n1507_));
  OAI21X1  g1122(.A0(new_n1507_), .A1(new_n1501_), .B0(new_n736_), .Y(new_n1508_));
  AOI21X1  g1123(.A0(new_n1508_), .A1(new_n1499_), .B0(new_n1500_), .Y(new_n1509_));
  OAI21X1  g1124(.A0(new_n1509_), .A1(new_n1498_), .B0(new_n751_), .Y(new_n1510_));
  AOI21X1  g1125(.A0(new_n1510_), .A1(new_n1496_), .B0(new_n1497_), .Y(new_n1511_));
  OAI21X1  g1126(.A0(new_n1511_), .A1(new_n1495_), .B0(new_n766_), .Y(new_n1512_));
  AOI21X1  g1127(.A0(new_n1512_), .A1(new_n1493_), .B0(new_n1494_), .Y(new_n1513_));
  OAI21X1  g1128(.A0(new_n1513_), .A1(new_n1492_), .B0(new_n781_), .Y(new_n1514_));
  AOI21X1  g1129(.A0(new_n1514_), .A1(new_n1490_), .B0(new_n1491_), .Y(new_n1515_));
  OAI21X1  g1130(.A0(new_n1515_), .A1(new_n1489_), .B0(new_n796_), .Y(new_n1516_));
  AOI21X1  g1131(.A0(new_n1516_), .A1(new_n1487_), .B0(new_n1488_), .Y(new_n1517_));
  OAI21X1  g1132(.A0(new_n1517_), .A1(new_n1486_), .B0(new_n811_), .Y(new_n1518_));
  AOI21X1  g1133(.A0(new_n1518_), .A1(new_n1484_), .B0(new_n1485_), .Y(new_n1519_));
  OAI21X1  g1134(.A0(new_n1519_), .A1(new_n1483_), .B0(new_n826_), .Y(new_n1520_));
  AOI21X1  g1135(.A0(new_n1520_), .A1(new_n1481_), .B0(new_n1482_), .Y(new_n1521_));
  OAI21X1  g1136(.A0(new_n1521_), .A1(new_n1480_), .B0(new_n841_), .Y(new_n1522_));
  AOI21X1  g1137(.A0(new_n1522_), .A1(new_n1478_), .B0(new_n1479_), .Y(new_n1523_));
  OAI21X1  g1138(.A0(new_n1523_), .A1(new_n1477_), .B0(new_n856_), .Y(new_n1524_));
  AOI21X1  g1139(.A0(new_n1524_), .A1(new_n1475_), .B0(new_n1476_), .Y(new_n1525_));
  OAI21X1  g1140(.A0(new_n1525_), .A1(new_n1474_), .B0(new_n871_), .Y(new_n1526_));
  AOI21X1  g1141(.A0(new_n1526_), .A1(new_n1472_), .B0(new_n1473_), .Y(new_n1527_));
  OAI21X1  g1142(.A0(new_n1527_), .A1(new_n1471_), .B0(new_n886_), .Y(new_n1528_));
  AOI21X1  g1143(.A0(new_n1528_), .A1(new_n1469_), .B0(new_n1470_), .Y(new_n1529_));
  OAI21X1  g1144(.A0(new_n1529_), .A1(new_n1468_), .B0(new_n901_), .Y(new_n1530_));
  AOI21X1  g1145(.A0(new_n1530_), .A1(new_n1466_), .B0(new_n1467_), .Y(new_n1531_));
  OAI21X1  g1146(.A0(new_n1531_), .A1(new_n1465_), .B0(new_n916_), .Y(new_n1532_));
  AOI21X1  g1147(.A0(new_n1532_), .A1(new_n1463_), .B0(new_n1464_), .Y(new_n1533_));
  OAI21X1  g1148(.A0(new_n1533_), .A1(new_n1462_), .B0(new_n931_), .Y(new_n1534_));
  AOI21X1  g1149(.A0(new_n1534_), .A1(new_n1460_), .B0(new_n1461_), .Y(new_n1535_));
  OAI21X1  g1150(.A0(new_n1535_), .A1(new_n1459_), .B0(new_n946_), .Y(new_n1536_));
  AOI21X1  g1151(.A0(new_n1536_), .A1(new_n1457_), .B0(new_n1458_), .Y(new_n1537_));
  OAI21X1  g1152(.A0(new_n1537_), .A1(new_n1456_), .B0(new_n961_), .Y(new_n1538_));
  AOI21X1  g1153(.A0(new_n1538_), .A1(new_n1454_), .B0(new_n1455_), .Y(new_n1539_));
  OAI21X1  g1154(.A0(new_n1539_), .A1(new_n1453_), .B0(new_n976_), .Y(new_n1540_));
  AOI21X1  g1155(.A0(new_n1540_), .A1(new_n1451_), .B0(new_n1452_), .Y(new_n1541_));
  OAI21X1  g1156(.A0(new_n1541_), .A1(new_n1450_), .B0(new_n991_), .Y(new_n1542_));
  AOI21X1  g1157(.A0(new_n1542_), .A1(new_n1448_), .B0(new_n1449_), .Y(new_n1543_));
  OAI21X1  g1158(.A0(new_n1543_), .A1(new_n1447_), .B0(new_n1006_), .Y(new_n1544_));
  AOI21X1  g1159(.A0(new_n1544_), .A1(new_n1445_), .B0(new_n1446_), .Y(new_n1545_));
  OR2X1    g1160(.A(\req[2] ), .B(\req[1] ), .Y(new_n1546_));
  AOI21X1  g1161(.A0(\req[0] ), .A1(new_n386_), .B0(new_n1546_), .Y(new_n1547_));
  OAI21X1  g1162(.A0(new_n1545_), .A1(new_n1444_), .B0(new_n1547_), .Y(new_n1548_));
  NOR2X1   g1163(.A(new_n706_), .B(\priority[4] ), .Y(new_n1549_));
  OAI21X1  g1164(.A0(new_n392_), .A1(\priority[4] ), .B0(\req[4] ), .Y(new_n1550_));
  AOI21X1  g1165(.A0(new_n1549_), .A1(new_n1548_), .B0(new_n1550_), .Y(\grant[4] ));
  AND2X1   g1166(.A(new_n393_), .B(new_n391_), .Y(new_n1552_));
  NAND2X1  g1167(.A(new_n1330_), .B(new_n387_), .Y(new_n1553_));
  AND2X1   g1168(.A(new_n1325_), .B(new_n1323_), .Y(new_n1554_));
  INVX1    g1169(.A(new_n1328_), .Y(new_n1555_));
  NAND2X1  g1170(.A(new_n1317_), .B(new_n1315_), .Y(new_n1556_));
  AND2X1   g1171(.A(new_n1310_), .B(new_n1308_), .Y(new_n1557_));
  INVX1    g1172(.A(new_n1313_), .Y(new_n1558_));
  NAND2X1  g1173(.A(new_n1302_), .B(new_n1300_), .Y(new_n1559_));
  AND2X1   g1174(.A(new_n1295_), .B(new_n1293_), .Y(new_n1560_));
  INVX1    g1175(.A(new_n1298_), .Y(new_n1561_));
  NAND2X1  g1176(.A(new_n1287_), .B(new_n1285_), .Y(new_n1562_));
  AND2X1   g1177(.A(new_n1280_), .B(new_n1278_), .Y(new_n1563_));
  INVX1    g1178(.A(new_n1283_), .Y(new_n1564_));
  NAND2X1  g1179(.A(new_n1272_), .B(new_n1270_), .Y(new_n1565_));
  AND2X1   g1180(.A(new_n1265_), .B(new_n1263_), .Y(new_n1566_));
  INVX1    g1181(.A(new_n1268_), .Y(new_n1567_));
  NAND2X1  g1182(.A(new_n1257_), .B(new_n1255_), .Y(new_n1568_));
  AND2X1   g1183(.A(new_n1250_), .B(new_n1248_), .Y(new_n1569_));
  INVX1    g1184(.A(new_n1253_), .Y(new_n1570_));
  NAND2X1  g1185(.A(new_n1242_), .B(new_n1240_), .Y(new_n1571_));
  AND2X1   g1186(.A(new_n1235_), .B(new_n1233_), .Y(new_n1572_));
  INVX1    g1187(.A(new_n1238_), .Y(new_n1573_));
  NAND2X1  g1188(.A(new_n1227_), .B(new_n1225_), .Y(new_n1574_));
  AND2X1   g1189(.A(new_n1220_), .B(new_n1218_), .Y(new_n1575_));
  INVX1    g1190(.A(new_n1223_), .Y(new_n1576_));
  NAND2X1  g1191(.A(new_n1212_), .B(new_n1210_), .Y(new_n1577_));
  AND2X1   g1192(.A(new_n1205_), .B(new_n1203_), .Y(new_n1578_));
  INVX1    g1193(.A(new_n1208_), .Y(new_n1579_));
  NAND2X1  g1194(.A(new_n1197_), .B(new_n1195_), .Y(new_n1580_));
  AND2X1   g1195(.A(new_n1190_), .B(new_n1188_), .Y(new_n1581_));
  INVX1    g1196(.A(new_n1193_), .Y(new_n1582_));
  NAND2X1  g1197(.A(new_n1182_), .B(new_n1180_), .Y(new_n1583_));
  AND2X1   g1198(.A(new_n1175_), .B(new_n1173_), .Y(new_n1584_));
  INVX1    g1199(.A(new_n1178_), .Y(new_n1585_));
  NAND2X1  g1200(.A(new_n1167_), .B(new_n1165_), .Y(new_n1586_));
  AND2X1   g1201(.A(new_n1160_), .B(new_n1158_), .Y(new_n1587_));
  INVX1    g1202(.A(new_n1163_), .Y(new_n1588_));
  NAND2X1  g1203(.A(new_n1152_), .B(new_n1150_), .Y(new_n1589_));
  AND2X1   g1204(.A(new_n1145_), .B(new_n1143_), .Y(new_n1590_));
  INVX1    g1205(.A(new_n1148_), .Y(new_n1591_));
  NAND2X1  g1206(.A(new_n1137_), .B(new_n1135_), .Y(new_n1592_));
  AND2X1   g1207(.A(new_n1130_), .B(new_n1128_), .Y(new_n1593_));
  INVX1    g1208(.A(new_n1133_), .Y(new_n1594_));
  NAND2X1  g1209(.A(new_n1122_), .B(new_n1120_), .Y(new_n1595_));
  AND2X1   g1210(.A(new_n1115_), .B(new_n1113_), .Y(new_n1596_));
  INVX1    g1211(.A(new_n1118_), .Y(new_n1597_));
  NAND2X1  g1212(.A(new_n1107_), .B(new_n1105_), .Y(new_n1598_));
  AND2X1   g1213(.A(new_n1100_), .B(new_n1098_), .Y(new_n1599_));
  INVX1    g1214(.A(new_n1103_), .Y(new_n1600_));
  NAND2X1  g1215(.A(new_n1092_), .B(new_n1090_), .Y(new_n1601_));
  AND2X1   g1216(.A(new_n1085_), .B(new_n1083_), .Y(new_n1602_));
  INVX1    g1217(.A(new_n1088_), .Y(new_n1603_));
  NAND2X1  g1218(.A(new_n1077_), .B(new_n1075_), .Y(new_n1604_));
  AND2X1   g1219(.A(new_n1070_), .B(new_n1068_), .Y(new_n1605_));
  INVX1    g1220(.A(new_n1073_), .Y(new_n1606_));
  NAND2X1  g1221(.A(new_n1062_), .B(new_n1060_), .Y(new_n1607_));
  AND2X1   g1222(.A(new_n1055_), .B(new_n1053_), .Y(new_n1608_));
  INVX1    g1223(.A(new_n1058_), .Y(new_n1609_));
  NAND2X1  g1224(.A(new_n1047_), .B(new_n1045_), .Y(new_n1610_));
  AND2X1   g1225(.A(new_n1040_), .B(new_n1038_), .Y(new_n1611_));
  INVX1    g1226(.A(new_n1043_), .Y(new_n1612_));
  NAND2X1  g1227(.A(new_n1032_), .B(new_n1030_), .Y(new_n1613_));
  NOR2X1   g1228(.A(new_n1027_), .B(new_n400_), .Y(new_n1614_));
  OAI21X1  g1229(.A0(new_n1614_), .A1(new_n1613_), .B0(new_n1035_), .Y(new_n1615_));
  AOI21X1  g1230(.A0(new_n1615_), .A1(new_n1611_), .B0(new_n1612_), .Y(new_n1616_));
  OAI21X1  g1231(.A0(new_n1616_), .A1(new_n1610_), .B0(new_n1050_), .Y(new_n1617_));
  AOI21X1  g1232(.A0(new_n1617_), .A1(new_n1608_), .B0(new_n1609_), .Y(new_n1618_));
  OAI21X1  g1233(.A0(new_n1618_), .A1(new_n1607_), .B0(new_n1065_), .Y(new_n1619_));
  AOI21X1  g1234(.A0(new_n1619_), .A1(new_n1605_), .B0(new_n1606_), .Y(new_n1620_));
  OAI21X1  g1235(.A0(new_n1620_), .A1(new_n1604_), .B0(new_n1080_), .Y(new_n1621_));
  AOI21X1  g1236(.A0(new_n1621_), .A1(new_n1602_), .B0(new_n1603_), .Y(new_n1622_));
  OAI21X1  g1237(.A0(new_n1622_), .A1(new_n1601_), .B0(new_n1095_), .Y(new_n1623_));
  AOI21X1  g1238(.A0(new_n1623_), .A1(new_n1599_), .B0(new_n1600_), .Y(new_n1624_));
  OAI21X1  g1239(.A0(new_n1624_), .A1(new_n1598_), .B0(new_n1110_), .Y(new_n1625_));
  AOI21X1  g1240(.A0(new_n1625_), .A1(new_n1596_), .B0(new_n1597_), .Y(new_n1626_));
  OAI21X1  g1241(.A0(new_n1626_), .A1(new_n1595_), .B0(new_n1125_), .Y(new_n1627_));
  AOI21X1  g1242(.A0(new_n1627_), .A1(new_n1593_), .B0(new_n1594_), .Y(new_n1628_));
  OAI21X1  g1243(.A0(new_n1628_), .A1(new_n1592_), .B0(new_n1140_), .Y(new_n1629_));
  AOI21X1  g1244(.A0(new_n1629_), .A1(new_n1590_), .B0(new_n1591_), .Y(new_n1630_));
  OAI21X1  g1245(.A0(new_n1630_), .A1(new_n1589_), .B0(new_n1155_), .Y(new_n1631_));
  AOI21X1  g1246(.A0(new_n1631_), .A1(new_n1587_), .B0(new_n1588_), .Y(new_n1632_));
  OAI21X1  g1247(.A0(new_n1632_), .A1(new_n1586_), .B0(new_n1170_), .Y(new_n1633_));
  AOI21X1  g1248(.A0(new_n1633_), .A1(new_n1584_), .B0(new_n1585_), .Y(new_n1634_));
  OAI21X1  g1249(.A0(new_n1634_), .A1(new_n1583_), .B0(new_n1185_), .Y(new_n1635_));
  AOI21X1  g1250(.A0(new_n1635_), .A1(new_n1581_), .B0(new_n1582_), .Y(new_n1636_));
  OAI21X1  g1251(.A0(new_n1636_), .A1(new_n1580_), .B0(new_n1200_), .Y(new_n1637_));
  AOI21X1  g1252(.A0(new_n1637_), .A1(new_n1578_), .B0(new_n1579_), .Y(new_n1638_));
  OAI21X1  g1253(.A0(new_n1638_), .A1(new_n1577_), .B0(new_n1215_), .Y(new_n1639_));
  AOI21X1  g1254(.A0(new_n1639_), .A1(new_n1575_), .B0(new_n1576_), .Y(new_n1640_));
  OAI21X1  g1255(.A0(new_n1640_), .A1(new_n1574_), .B0(new_n1230_), .Y(new_n1641_));
  AOI21X1  g1256(.A0(new_n1641_), .A1(new_n1572_), .B0(new_n1573_), .Y(new_n1642_));
  OAI21X1  g1257(.A0(new_n1642_), .A1(new_n1571_), .B0(new_n1245_), .Y(new_n1643_));
  AOI21X1  g1258(.A0(new_n1643_), .A1(new_n1569_), .B0(new_n1570_), .Y(new_n1644_));
  OAI21X1  g1259(.A0(new_n1644_), .A1(new_n1568_), .B0(new_n1260_), .Y(new_n1645_));
  AOI21X1  g1260(.A0(new_n1645_), .A1(new_n1566_), .B0(new_n1567_), .Y(new_n1646_));
  OAI21X1  g1261(.A0(new_n1646_), .A1(new_n1565_), .B0(new_n1275_), .Y(new_n1647_));
  AOI21X1  g1262(.A0(new_n1647_), .A1(new_n1563_), .B0(new_n1564_), .Y(new_n1648_));
  OAI21X1  g1263(.A0(new_n1648_), .A1(new_n1562_), .B0(new_n1290_), .Y(new_n1649_));
  AOI21X1  g1264(.A0(new_n1649_), .A1(new_n1560_), .B0(new_n1561_), .Y(new_n1650_));
  OAI21X1  g1265(.A0(new_n1650_), .A1(new_n1559_), .B0(new_n1305_), .Y(new_n1651_));
  AOI21X1  g1266(.A0(new_n1651_), .A1(new_n1557_), .B0(new_n1558_), .Y(new_n1652_));
  OAI21X1  g1267(.A0(new_n1652_), .A1(new_n1556_), .B0(new_n1320_), .Y(new_n1653_));
  AOI21X1  g1268(.A0(new_n1653_), .A1(new_n1554_), .B0(new_n1555_), .Y(new_n1654_));
  OR2X1    g1269(.A(\req[3] ), .B(\req[2] ), .Y(new_n1655_));
  AOI21X1  g1270(.A0(\req[1] ), .A1(new_n387_), .B0(new_n1655_), .Y(new_n1656_));
  OAI21X1  g1271(.A0(new_n1654_), .A1(new_n1553_), .B0(new_n1656_), .Y(new_n1657_));
  OAI21X1  g1272(.A0(new_n710_), .A1(\priority[5] ), .B0(\req[5] ), .Y(new_n1658_));
  AOI21X1  g1273(.A0(new_n1657_), .A1(new_n1552_), .B0(new_n1658_), .Y(\grant[5] ));
  AND2X1   g1274(.A(new_n711_), .B(new_n709_), .Y(new_n1660_));
  OR2X1    g1275(.A(new_n388_), .B(\priority[3] ), .Y(new_n1661_));
  INVX1    g1276(.A(new_n1438_), .Y(new_n1662_));
  NOR2X1   g1277(.A(new_n718_), .B(new_n402_), .Y(new_n1663_));
  OAI21X1  g1278(.A0(new_n1663_), .A1(new_n409_), .B0(new_n411_), .Y(new_n1664_));
  AOI21X1  g1279(.A0(new_n1664_), .A1(new_n416_), .B0(new_n419_), .Y(new_n1665_));
  OAI21X1  g1280(.A0(new_n1665_), .A1(new_n424_), .B0(new_n426_), .Y(new_n1666_));
  AOI21X1  g1281(.A0(new_n1666_), .A1(new_n431_), .B0(new_n434_), .Y(new_n1667_));
  OAI21X1  g1282(.A0(new_n1667_), .A1(new_n439_), .B0(new_n441_), .Y(new_n1668_));
  AOI21X1  g1283(.A0(new_n1668_), .A1(new_n446_), .B0(new_n449_), .Y(new_n1669_));
  OAI21X1  g1284(.A0(new_n1669_), .A1(new_n454_), .B0(new_n456_), .Y(new_n1670_));
  AOI21X1  g1285(.A0(new_n1670_), .A1(new_n461_), .B0(new_n464_), .Y(new_n1671_));
  OAI21X1  g1286(.A0(new_n1671_), .A1(new_n469_), .B0(new_n471_), .Y(new_n1672_));
  AOI21X1  g1287(.A0(new_n1672_), .A1(new_n476_), .B0(new_n479_), .Y(new_n1673_));
  OAI21X1  g1288(.A0(new_n1673_), .A1(new_n484_), .B0(new_n486_), .Y(new_n1674_));
  AOI21X1  g1289(.A0(new_n1674_), .A1(new_n491_), .B0(new_n494_), .Y(new_n1675_));
  OAI21X1  g1290(.A0(new_n1675_), .A1(new_n499_), .B0(new_n501_), .Y(new_n1676_));
  AOI21X1  g1291(.A0(new_n1676_), .A1(new_n506_), .B0(new_n509_), .Y(new_n1677_));
  OAI21X1  g1292(.A0(new_n1677_), .A1(new_n514_), .B0(new_n516_), .Y(new_n1678_));
  AOI21X1  g1293(.A0(new_n1678_), .A1(new_n521_), .B0(new_n524_), .Y(new_n1679_));
  OAI21X1  g1294(.A0(new_n1679_), .A1(new_n529_), .B0(new_n531_), .Y(new_n1680_));
  AOI21X1  g1295(.A0(new_n1680_), .A1(new_n536_), .B0(new_n539_), .Y(new_n1681_));
  OAI21X1  g1296(.A0(new_n1681_), .A1(new_n544_), .B0(new_n546_), .Y(new_n1682_));
  AOI21X1  g1297(.A0(new_n1682_), .A1(new_n551_), .B0(new_n554_), .Y(new_n1683_));
  OAI21X1  g1298(.A0(new_n1683_), .A1(new_n559_), .B0(new_n561_), .Y(new_n1684_));
  AOI21X1  g1299(.A0(new_n1684_), .A1(new_n566_), .B0(new_n569_), .Y(new_n1685_));
  OAI21X1  g1300(.A0(new_n1685_), .A1(new_n574_), .B0(new_n576_), .Y(new_n1686_));
  AOI21X1  g1301(.A0(new_n1686_), .A1(new_n581_), .B0(new_n584_), .Y(new_n1687_));
  OAI21X1  g1302(.A0(new_n1687_), .A1(new_n589_), .B0(new_n591_), .Y(new_n1688_));
  AOI21X1  g1303(.A0(new_n1688_), .A1(new_n596_), .B0(new_n599_), .Y(new_n1689_));
  OAI21X1  g1304(.A0(new_n1689_), .A1(new_n604_), .B0(new_n606_), .Y(new_n1690_));
  AOI21X1  g1305(.A0(new_n1690_), .A1(new_n611_), .B0(new_n614_), .Y(new_n1691_));
  OAI21X1  g1306(.A0(new_n1691_), .A1(new_n619_), .B0(new_n621_), .Y(new_n1692_));
  AOI21X1  g1307(.A0(new_n1692_), .A1(new_n626_), .B0(new_n629_), .Y(new_n1693_));
  OAI21X1  g1308(.A0(new_n1693_), .A1(new_n634_), .B0(new_n636_), .Y(new_n1694_));
  AOI21X1  g1309(.A0(new_n1694_), .A1(new_n641_), .B0(new_n644_), .Y(new_n1695_));
  OAI21X1  g1310(.A0(new_n1695_), .A1(new_n649_), .B0(new_n651_), .Y(new_n1696_));
  AOI21X1  g1311(.A0(new_n1696_), .A1(new_n656_), .B0(new_n659_), .Y(new_n1697_));
  OAI21X1  g1312(.A0(new_n1697_), .A1(new_n664_), .B0(new_n666_), .Y(new_n1698_));
  AOI21X1  g1313(.A0(new_n1698_), .A1(new_n671_), .B0(new_n674_), .Y(new_n1699_));
  OAI21X1  g1314(.A0(new_n1699_), .A1(new_n679_), .B0(new_n681_), .Y(new_n1700_));
  AOI21X1  g1315(.A0(new_n1700_), .A1(new_n686_), .B0(new_n689_), .Y(new_n1701_));
  OAI21X1  g1316(.A0(new_n1701_), .A1(new_n694_), .B0(new_n696_), .Y(new_n1702_));
  AOI21X1  g1317(.A0(new_n1702_), .A1(new_n701_), .B0(new_n1662_), .Y(new_n1703_));
  OR2X1    g1318(.A(\req[4] ), .B(\req[3] ), .Y(new_n1704_));
  AOI21X1  g1319(.A0(\req[2] ), .A1(new_n705_), .B0(new_n1704_), .Y(new_n1705_));
  OAI21X1  g1320(.A0(new_n1703_), .A1(new_n1661_), .B0(new_n1705_), .Y(new_n1706_));
  OAI21X1  g1321(.A0(new_n1024_), .A1(\priority[6] ), .B0(\req[6] ), .Y(new_n1707_));
  AOI21X1  g1322(.A0(new_n1706_), .A1(new_n1660_), .B0(new_n1707_), .Y(\grant[6] ));
  AND2X1   g1323(.A(new_n1025_), .B(new_n1023_), .Y(new_n1709_));
  OR2X1    g1324(.A(new_n706_), .B(\priority[4] ), .Y(new_n1710_));
  INVX1    g1325(.A(new_n1547_), .Y(new_n1711_));
  NOR2X1   g1326(.A(new_n1032_), .B(new_n720_), .Y(new_n1712_));
  OAI21X1  g1327(.A0(new_n1712_), .A1(new_n727_), .B0(new_n729_), .Y(new_n1713_));
  AOI21X1  g1328(.A0(new_n1713_), .A1(new_n734_), .B0(new_n737_), .Y(new_n1714_));
  OAI21X1  g1329(.A0(new_n1714_), .A1(new_n742_), .B0(new_n744_), .Y(new_n1715_));
  AOI21X1  g1330(.A0(new_n1715_), .A1(new_n749_), .B0(new_n752_), .Y(new_n1716_));
  OAI21X1  g1331(.A0(new_n1716_), .A1(new_n757_), .B0(new_n759_), .Y(new_n1717_));
  AOI21X1  g1332(.A0(new_n1717_), .A1(new_n764_), .B0(new_n767_), .Y(new_n1718_));
  OAI21X1  g1333(.A0(new_n1718_), .A1(new_n772_), .B0(new_n774_), .Y(new_n1719_));
  AOI21X1  g1334(.A0(new_n1719_), .A1(new_n779_), .B0(new_n782_), .Y(new_n1720_));
  OAI21X1  g1335(.A0(new_n1720_), .A1(new_n787_), .B0(new_n789_), .Y(new_n1721_));
  AOI21X1  g1336(.A0(new_n1721_), .A1(new_n794_), .B0(new_n797_), .Y(new_n1722_));
  OAI21X1  g1337(.A0(new_n1722_), .A1(new_n802_), .B0(new_n804_), .Y(new_n1723_));
  AOI21X1  g1338(.A0(new_n1723_), .A1(new_n809_), .B0(new_n812_), .Y(new_n1724_));
  OAI21X1  g1339(.A0(new_n1724_), .A1(new_n817_), .B0(new_n819_), .Y(new_n1725_));
  AOI21X1  g1340(.A0(new_n1725_), .A1(new_n824_), .B0(new_n827_), .Y(new_n1726_));
  OAI21X1  g1341(.A0(new_n1726_), .A1(new_n832_), .B0(new_n834_), .Y(new_n1727_));
  AOI21X1  g1342(.A0(new_n1727_), .A1(new_n839_), .B0(new_n842_), .Y(new_n1728_));
  OAI21X1  g1343(.A0(new_n1728_), .A1(new_n847_), .B0(new_n849_), .Y(new_n1729_));
  AOI21X1  g1344(.A0(new_n1729_), .A1(new_n854_), .B0(new_n857_), .Y(new_n1730_));
  OAI21X1  g1345(.A0(new_n1730_), .A1(new_n862_), .B0(new_n864_), .Y(new_n1731_));
  AOI21X1  g1346(.A0(new_n1731_), .A1(new_n869_), .B0(new_n872_), .Y(new_n1732_));
  OAI21X1  g1347(.A0(new_n1732_), .A1(new_n877_), .B0(new_n879_), .Y(new_n1733_));
  AOI21X1  g1348(.A0(new_n1733_), .A1(new_n884_), .B0(new_n887_), .Y(new_n1734_));
  OAI21X1  g1349(.A0(new_n1734_), .A1(new_n892_), .B0(new_n894_), .Y(new_n1735_));
  AOI21X1  g1350(.A0(new_n1735_), .A1(new_n899_), .B0(new_n902_), .Y(new_n1736_));
  OAI21X1  g1351(.A0(new_n1736_), .A1(new_n907_), .B0(new_n909_), .Y(new_n1737_));
  AOI21X1  g1352(.A0(new_n1737_), .A1(new_n914_), .B0(new_n917_), .Y(new_n1738_));
  OAI21X1  g1353(.A0(new_n1738_), .A1(new_n922_), .B0(new_n924_), .Y(new_n1739_));
  AOI21X1  g1354(.A0(new_n1739_), .A1(new_n929_), .B0(new_n932_), .Y(new_n1740_));
  OAI21X1  g1355(.A0(new_n1740_), .A1(new_n937_), .B0(new_n939_), .Y(new_n1741_));
  AOI21X1  g1356(.A0(new_n1741_), .A1(new_n944_), .B0(new_n947_), .Y(new_n1742_));
  OAI21X1  g1357(.A0(new_n1742_), .A1(new_n952_), .B0(new_n954_), .Y(new_n1743_));
  AOI21X1  g1358(.A0(new_n1743_), .A1(new_n959_), .B0(new_n962_), .Y(new_n1744_));
  OAI21X1  g1359(.A0(new_n1744_), .A1(new_n967_), .B0(new_n969_), .Y(new_n1745_));
  AOI21X1  g1360(.A0(new_n1745_), .A1(new_n974_), .B0(new_n977_), .Y(new_n1746_));
  OAI21X1  g1361(.A0(new_n1746_), .A1(new_n982_), .B0(new_n984_), .Y(new_n1747_));
  AOI21X1  g1362(.A0(new_n1747_), .A1(new_n989_), .B0(new_n992_), .Y(new_n1748_));
  OAI21X1  g1363(.A0(new_n1748_), .A1(new_n997_), .B0(new_n999_), .Y(new_n1749_));
  AOI21X1  g1364(.A0(new_n1749_), .A1(new_n1004_), .B0(new_n1007_), .Y(new_n1750_));
  OAI21X1  g1365(.A0(new_n1750_), .A1(new_n1012_), .B0(new_n1014_), .Y(new_n1751_));
  AOI21X1  g1366(.A0(new_n1751_), .A1(new_n1017_), .B0(new_n1711_), .Y(new_n1752_));
  INVX1    g1367(.A(\priority[4] ), .Y(new_n1753_));
  AOI21X1  g1368(.A0(\req[3] ), .A1(new_n1753_), .B0(new_n1021_), .Y(new_n1754_));
  OAI21X1  g1369(.A0(new_n1752_), .A1(new_n1710_), .B0(new_n1754_), .Y(new_n1755_));
  OAI21X1  g1370(.A0(new_n399_), .A1(\priority[7] ), .B0(\req[7] ), .Y(new_n1756_));
  AOI21X1  g1371(.A0(new_n1755_), .A1(new_n1709_), .B0(new_n1756_), .Y(\grant[7] ));
  INVX1    g1372(.A(new_n1656_), .Y(new_n1758_));
  NOR2X1   g1373(.A(new_n1034_), .B(new_n408_), .Y(new_n1759_));
  OAI21X1  g1374(.A0(new_n1759_), .A1(new_n1041_), .B0(new_n1043_), .Y(new_n1760_));
  AOI21X1  g1375(.A0(new_n1760_), .A1(new_n1048_), .B0(new_n1051_), .Y(new_n1761_));
  OAI21X1  g1376(.A0(new_n1761_), .A1(new_n1056_), .B0(new_n1058_), .Y(new_n1762_));
  AOI21X1  g1377(.A0(new_n1762_), .A1(new_n1063_), .B0(new_n1066_), .Y(new_n1763_));
  OAI21X1  g1378(.A0(new_n1763_), .A1(new_n1071_), .B0(new_n1073_), .Y(new_n1764_));
  AOI21X1  g1379(.A0(new_n1764_), .A1(new_n1078_), .B0(new_n1081_), .Y(new_n1765_));
  OAI21X1  g1380(.A0(new_n1765_), .A1(new_n1086_), .B0(new_n1088_), .Y(new_n1766_));
  AOI21X1  g1381(.A0(new_n1766_), .A1(new_n1093_), .B0(new_n1096_), .Y(new_n1767_));
  OAI21X1  g1382(.A0(new_n1767_), .A1(new_n1101_), .B0(new_n1103_), .Y(new_n1768_));
  AOI21X1  g1383(.A0(new_n1768_), .A1(new_n1108_), .B0(new_n1111_), .Y(new_n1769_));
  OAI21X1  g1384(.A0(new_n1769_), .A1(new_n1116_), .B0(new_n1118_), .Y(new_n1770_));
  AOI21X1  g1385(.A0(new_n1770_), .A1(new_n1123_), .B0(new_n1126_), .Y(new_n1771_));
  OAI21X1  g1386(.A0(new_n1771_), .A1(new_n1131_), .B0(new_n1133_), .Y(new_n1772_));
  AOI21X1  g1387(.A0(new_n1772_), .A1(new_n1138_), .B0(new_n1141_), .Y(new_n1773_));
  OAI21X1  g1388(.A0(new_n1773_), .A1(new_n1146_), .B0(new_n1148_), .Y(new_n1774_));
  AOI21X1  g1389(.A0(new_n1774_), .A1(new_n1153_), .B0(new_n1156_), .Y(new_n1775_));
  OAI21X1  g1390(.A0(new_n1775_), .A1(new_n1161_), .B0(new_n1163_), .Y(new_n1776_));
  AOI21X1  g1391(.A0(new_n1776_), .A1(new_n1168_), .B0(new_n1171_), .Y(new_n1777_));
  OAI21X1  g1392(.A0(new_n1777_), .A1(new_n1176_), .B0(new_n1178_), .Y(new_n1778_));
  AOI21X1  g1393(.A0(new_n1778_), .A1(new_n1183_), .B0(new_n1186_), .Y(new_n1779_));
  OAI21X1  g1394(.A0(new_n1779_), .A1(new_n1191_), .B0(new_n1193_), .Y(new_n1780_));
  AOI21X1  g1395(.A0(new_n1780_), .A1(new_n1198_), .B0(new_n1201_), .Y(new_n1781_));
  OAI21X1  g1396(.A0(new_n1781_), .A1(new_n1206_), .B0(new_n1208_), .Y(new_n1782_));
  AOI21X1  g1397(.A0(new_n1782_), .A1(new_n1213_), .B0(new_n1216_), .Y(new_n1783_));
  OAI21X1  g1398(.A0(new_n1783_), .A1(new_n1221_), .B0(new_n1223_), .Y(new_n1784_));
  AOI21X1  g1399(.A0(new_n1784_), .A1(new_n1228_), .B0(new_n1231_), .Y(new_n1785_));
  OAI21X1  g1400(.A0(new_n1785_), .A1(new_n1236_), .B0(new_n1238_), .Y(new_n1786_));
  AOI21X1  g1401(.A0(new_n1786_), .A1(new_n1243_), .B0(new_n1246_), .Y(new_n1787_));
  OAI21X1  g1402(.A0(new_n1787_), .A1(new_n1251_), .B0(new_n1253_), .Y(new_n1788_));
  AOI21X1  g1403(.A0(new_n1788_), .A1(new_n1258_), .B0(new_n1261_), .Y(new_n1789_));
  OAI21X1  g1404(.A0(new_n1789_), .A1(new_n1266_), .B0(new_n1268_), .Y(new_n1790_));
  AOI21X1  g1405(.A0(new_n1790_), .A1(new_n1273_), .B0(new_n1276_), .Y(new_n1791_));
  OAI21X1  g1406(.A0(new_n1791_), .A1(new_n1281_), .B0(new_n1283_), .Y(new_n1792_));
  AOI21X1  g1407(.A0(new_n1792_), .A1(new_n1288_), .B0(new_n1291_), .Y(new_n1793_));
  OAI21X1  g1408(.A0(new_n1793_), .A1(new_n1296_), .B0(new_n1298_), .Y(new_n1794_));
  AOI21X1  g1409(.A0(new_n1794_), .A1(new_n1303_), .B0(new_n1306_), .Y(new_n1795_));
  OAI21X1  g1410(.A0(new_n1795_), .A1(new_n1311_), .B0(new_n1313_), .Y(new_n1796_));
  AOI21X1  g1411(.A0(new_n1796_), .A1(new_n1318_), .B0(new_n1321_), .Y(new_n1797_));
  OAI21X1  g1412(.A0(new_n1797_), .A1(new_n1326_), .B0(new_n1328_), .Y(new_n1798_));
  AOI21X1  g1413(.A0(new_n1798_), .A1(new_n1331_), .B0(new_n1758_), .Y(new_n1799_));
  OAI21X1  g1414(.A0(new_n1799_), .A1(new_n394_), .B0(new_n396_), .Y(new_n1800_));
  OAI21X1  g1415(.A0(new_n717_), .A1(\priority[8] ), .B0(\req[8] ), .Y(new_n1801_));
  AOI21X1  g1416(.A0(new_n1800_), .A1(new_n401_), .B0(new_n1801_), .Y(\grant[8] ));
  INVX1    g1417(.A(new_n1705_), .Y(new_n1803_));
  NOR2X1   g1418(.A(new_n726_), .B(new_n410_), .Y(new_n1804_));
  OAI21X1  g1419(.A0(new_n1804_), .A1(new_n1392_), .B0(new_n418_), .Y(new_n1805_));
  AOI21X1  g1420(.A0(new_n1805_), .A1(new_n1390_), .B0(new_n1391_), .Y(new_n1806_));
  OAI21X1  g1421(.A0(new_n1806_), .A1(new_n1389_), .B0(new_n433_), .Y(new_n1807_));
  AOI21X1  g1422(.A0(new_n1807_), .A1(new_n1387_), .B0(new_n1388_), .Y(new_n1808_));
  OAI21X1  g1423(.A0(new_n1808_), .A1(new_n1386_), .B0(new_n448_), .Y(new_n1809_));
  AOI21X1  g1424(.A0(new_n1809_), .A1(new_n1384_), .B0(new_n1385_), .Y(new_n1810_));
  OAI21X1  g1425(.A0(new_n1810_), .A1(new_n1383_), .B0(new_n463_), .Y(new_n1811_));
  AOI21X1  g1426(.A0(new_n1811_), .A1(new_n1381_), .B0(new_n1382_), .Y(new_n1812_));
  OAI21X1  g1427(.A0(new_n1812_), .A1(new_n1380_), .B0(new_n478_), .Y(new_n1813_));
  AOI21X1  g1428(.A0(new_n1813_), .A1(new_n1378_), .B0(new_n1379_), .Y(new_n1814_));
  OAI21X1  g1429(.A0(new_n1814_), .A1(new_n1377_), .B0(new_n493_), .Y(new_n1815_));
  AOI21X1  g1430(.A0(new_n1815_), .A1(new_n1375_), .B0(new_n1376_), .Y(new_n1816_));
  OAI21X1  g1431(.A0(new_n1816_), .A1(new_n1374_), .B0(new_n508_), .Y(new_n1817_));
  AOI21X1  g1432(.A0(new_n1817_), .A1(new_n1372_), .B0(new_n1373_), .Y(new_n1818_));
  OAI21X1  g1433(.A0(new_n1818_), .A1(new_n1371_), .B0(new_n523_), .Y(new_n1819_));
  AOI21X1  g1434(.A0(new_n1819_), .A1(new_n1369_), .B0(new_n1370_), .Y(new_n1820_));
  OAI21X1  g1435(.A0(new_n1820_), .A1(new_n1368_), .B0(new_n538_), .Y(new_n1821_));
  AOI21X1  g1436(.A0(new_n1821_), .A1(new_n1366_), .B0(new_n1367_), .Y(new_n1822_));
  OAI21X1  g1437(.A0(new_n1822_), .A1(new_n1365_), .B0(new_n553_), .Y(new_n1823_));
  AOI21X1  g1438(.A0(new_n1823_), .A1(new_n1363_), .B0(new_n1364_), .Y(new_n1824_));
  OAI21X1  g1439(.A0(new_n1824_), .A1(new_n1362_), .B0(new_n568_), .Y(new_n1825_));
  AOI21X1  g1440(.A0(new_n1825_), .A1(new_n1360_), .B0(new_n1361_), .Y(new_n1826_));
  OAI21X1  g1441(.A0(new_n1826_), .A1(new_n1359_), .B0(new_n583_), .Y(new_n1827_));
  AOI21X1  g1442(.A0(new_n1827_), .A1(new_n1357_), .B0(new_n1358_), .Y(new_n1828_));
  OAI21X1  g1443(.A0(new_n1828_), .A1(new_n1356_), .B0(new_n598_), .Y(new_n1829_));
  AOI21X1  g1444(.A0(new_n1829_), .A1(new_n1354_), .B0(new_n1355_), .Y(new_n1830_));
  OAI21X1  g1445(.A0(new_n1830_), .A1(new_n1353_), .B0(new_n613_), .Y(new_n1831_));
  AOI21X1  g1446(.A0(new_n1831_), .A1(new_n1351_), .B0(new_n1352_), .Y(new_n1832_));
  OAI21X1  g1447(.A0(new_n1832_), .A1(new_n1350_), .B0(new_n628_), .Y(new_n1833_));
  AOI21X1  g1448(.A0(new_n1833_), .A1(new_n1348_), .B0(new_n1349_), .Y(new_n1834_));
  OAI21X1  g1449(.A0(new_n1834_), .A1(new_n1347_), .B0(new_n643_), .Y(new_n1835_));
  AOI21X1  g1450(.A0(new_n1835_), .A1(new_n1345_), .B0(new_n1346_), .Y(new_n1836_));
  OAI21X1  g1451(.A0(new_n1836_), .A1(new_n1344_), .B0(new_n658_), .Y(new_n1837_));
  AOI21X1  g1452(.A0(new_n1837_), .A1(new_n1342_), .B0(new_n1343_), .Y(new_n1838_));
  OAI21X1  g1453(.A0(new_n1838_), .A1(new_n1341_), .B0(new_n673_), .Y(new_n1839_));
  AOI21X1  g1454(.A0(new_n1839_), .A1(new_n1339_), .B0(new_n1340_), .Y(new_n1840_));
  OAI21X1  g1455(.A0(new_n1840_), .A1(new_n1338_), .B0(new_n688_), .Y(new_n1841_));
  AOI21X1  g1456(.A0(new_n1841_), .A1(new_n1336_), .B0(new_n1337_), .Y(new_n1842_));
  OAI21X1  g1457(.A0(new_n1842_), .A1(new_n1335_), .B0(new_n1438_), .Y(new_n1843_));
  AOI21X1  g1458(.A0(new_n1843_), .A1(new_n1440_), .B0(new_n1803_), .Y(new_n1844_));
  OAI21X1  g1459(.A0(new_n1844_), .A1(new_n712_), .B0(new_n714_), .Y(new_n1845_));
  OAI21X1  g1460(.A0(new_n1031_), .A1(\priority[9] ), .B0(\req[9] ), .Y(new_n1846_));
  AOI21X1  g1461(.A0(new_n1845_), .A1(new_n719_), .B0(new_n1846_), .Y(\grant[9] ));
  INVX1    g1462(.A(new_n1754_), .Y(new_n1848_));
  NOR2X1   g1463(.A(new_n1040_), .B(new_n728_), .Y(new_n1849_));
  OAI21X1  g1464(.A0(new_n1849_), .A1(new_n1501_), .B0(new_n736_), .Y(new_n1850_));
  AOI21X1  g1465(.A0(new_n1850_), .A1(new_n1499_), .B0(new_n1500_), .Y(new_n1851_));
  OAI21X1  g1466(.A0(new_n1851_), .A1(new_n1498_), .B0(new_n751_), .Y(new_n1852_));
  AOI21X1  g1467(.A0(new_n1852_), .A1(new_n1496_), .B0(new_n1497_), .Y(new_n1853_));
  OAI21X1  g1468(.A0(new_n1853_), .A1(new_n1495_), .B0(new_n766_), .Y(new_n1854_));
  AOI21X1  g1469(.A0(new_n1854_), .A1(new_n1493_), .B0(new_n1494_), .Y(new_n1855_));
  OAI21X1  g1470(.A0(new_n1855_), .A1(new_n1492_), .B0(new_n781_), .Y(new_n1856_));
  AOI21X1  g1471(.A0(new_n1856_), .A1(new_n1490_), .B0(new_n1491_), .Y(new_n1857_));
  OAI21X1  g1472(.A0(new_n1857_), .A1(new_n1489_), .B0(new_n796_), .Y(new_n1858_));
  AOI21X1  g1473(.A0(new_n1858_), .A1(new_n1487_), .B0(new_n1488_), .Y(new_n1859_));
  OAI21X1  g1474(.A0(new_n1859_), .A1(new_n1486_), .B0(new_n811_), .Y(new_n1860_));
  AOI21X1  g1475(.A0(new_n1860_), .A1(new_n1484_), .B0(new_n1485_), .Y(new_n1861_));
  OAI21X1  g1476(.A0(new_n1861_), .A1(new_n1483_), .B0(new_n826_), .Y(new_n1862_));
  AOI21X1  g1477(.A0(new_n1862_), .A1(new_n1481_), .B0(new_n1482_), .Y(new_n1863_));
  OAI21X1  g1478(.A0(new_n1863_), .A1(new_n1480_), .B0(new_n841_), .Y(new_n1864_));
  AOI21X1  g1479(.A0(new_n1864_), .A1(new_n1478_), .B0(new_n1479_), .Y(new_n1865_));
  OAI21X1  g1480(.A0(new_n1865_), .A1(new_n1477_), .B0(new_n856_), .Y(new_n1866_));
  AOI21X1  g1481(.A0(new_n1866_), .A1(new_n1475_), .B0(new_n1476_), .Y(new_n1867_));
  OAI21X1  g1482(.A0(new_n1867_), .A1(new_n1474_), .B0(new_n871_), .Y(new_n1868_));
  AOI21X1  g1483(.A0(new_n1868_), .A1(new_n1472_), .B0(new_n1473_), .Y(new_n1869_));
  OAI21X1  g1484(.A0(new_n1869_), .A1(new_n1471_), .B0(new_n886_), .Y(new_n1870_));
  AOI21X1  g1485(.A0(new_n1870_), .A1(new_n1469_), .B0(new_n1470_), .Y(new_n1871_));
  OAI21X1  g1486(.A0(new_n1871_), .A1(new_n1468_), .B0(new_n901_), .Y(new_n1872_));
  AOI21X1  g1487(.A0(new_n1872_), .A1(new_n1466_), .B0(new_n1467_), .Y(new_n1873_));
  OAI21X1  g1488(.A0(new_n1873_), .A1(new_n1465_), .B0(new_n916_), .Y(new_n1874_));
  AOI21X1  g1489(.A0(new_n1874_), .A1(new_n1463_), .B0(new_n1464_), .Y(new_n1875_));
  OAI21X1  g1490(.A0(new_n1875_), .A1(new_n1462_), .B0(new_n931_), .Y(new_n1876_));
  AOI21X1  g1491(.A0(new_n1876_), .A1(new_n1460_), .B0(new_n1461_), .Y(new_n1877_));
  OAI21X1  g1492(.A0(new_n1877_), .A1(new_n1459_), .B0(new_n946_), .Y(new_n1878_));
  AOI21X1  g1493(.A0(new_n1878_), .A1(new_n1457_), .B0(new_n1458_), .Y(new_n1879_));
  OAI21X1  g1494(.A0(new_n1879_), .A1(new_n1456_), .B0(new_n961_), .Y(new_n1880_));
  AOI21X1  g1495(.A0(new_n1880_), .A1(new_n1454_), .B0(new_n1455_), .Y(new_n1881_));
  OAI21X1  g1496(.A0(new_n1881_), .A1(new_n1453_), .B0(new_n976_), .Y(new_n1882_));
  AOI21X1  g1497(.A0(new_n1882_), .A1(new_n1451_), .B0(new_n1452_), .Y(new_n1883_));
  OAI21X1  g1498(.A0(new_n1883_), .A1(new_n1450_), .B0(new_n991_), .Y(new_n1884_));
  AOI21X1  g1499(.A0(new_n1884_), .A1(new_n1448_), .B0(new_n1449_), .Y(new_n1885_));
  OAI21X1  g1500(.A0(new_n1885_), .A1(new_n1447_), .B0(new_n1006_), .Y(new_n1886_));
  AOI21X1  g1501(.A0(new_n1886_), .A1(new_n1445_), .B0(new_n1446_), .Y(new_n1887_));
  OAI21X1  g1502(.A0(new_n1887_), .A1(new_n1444_), .B0(new_n1547_), .Y(new_n1888_));
  AOI21X1  g1503(.A0(new_n1888_), .A1(new_n1549_), .B0(new_n1848_), .Y(new_n1889_));
  OAI21X1  g1504(.A0(new_n1889_), .A1(new_n1026_), .B0(new_n1028_), .Y(new_n1890_));
  OAI21X1  g1505(.A0(new_n407_), .A1(\priority[10] ), .B0(\req[10] ), .Y(new_n1891_));
  AOI21X1  g1506(.A0(new_n1890_), .A1(new_n1033_), .B0(new_n1891_), .Y(\grant[10] ));
  INVX1    g1507(.A(new_n396_), .Y(new_n1893_));
  NOR2X1   g1508(.A(new_n1042_), .B(new_n415_), .Y(new_n1894_));
  OAI21X1  g1509(.A0(new_n1894_), .A1(new_n1610_), .B0(new_n1050_), .Y(new_n1895_));
  AOI21X1  g1510(.A0(new_n1895_), .A1(new_n1608_), .B0(new_n1609_), .Y(new_n1896_));
  OAI21X1  g1511(.A0(new_n1896_), .A1(new_n1607_), .B0(new_n1065_), .Y(new_n1897_));
  AOI21X1  g1512(.A0(new_n1897_), .A1(new_n1605_), .B0(new_n1606_), .Y(new_n1898_));
  OAI21X1  g1513(.A0(new_n1898_), .A1(new_n1604_), .B0(new_n1080_), .Y(new_n1899_));
  AOI21X1  g1514(.A0(new_n1899_), .A1(new_n1602_), .B0(new_n1603_), .Y(new_n1900_));
  OAI21X1  g1515(.A0(new_n1900_), .A1(new_n1601_), .B0(new_n1095_), .Y(new_n1901_));
  AOI21X1  g1516(.A0(new_n1901_), .A1(new_n1599_), .B0(new_n1600_), .Y(new_n1902_));
  OAI21X1  g1517(.A0(new_n1902_), .A1(new_n1598_), .B0(new_n1110_), .Y(new_n1903_));
  AOI21X1  g1518(.A0(new_n1903_), .A1(new_n1596_), .B0(new_n1597_), .Y(new_n1904_));
  OAI21X1  g1519(.A0(new_n1904_), .A1(new_n1595_), .B0(new_n1125_), .Y(new_n1905_));
  AOI21X1  g1520(.A0(new_n1905_), .A1(new_n1593_), .B0(new_n1594_), .Y(new_n1906_));
  OAI21X1  g1521(.A0(new_n1906_), .A1(new_n1592_), .B0(new_n1140_), .Y(new_n1907_));
  AOI21X1  g1522(.A0(new_n1907_), .A1(new_n1590_), .B0(new_n1591_), .Y(new_n1908_));
  OAI21X1  g1523(.A0(new_n1908_), .A1(new_n1589_), .B0(new_n1155_), .Y(new_n1909_));
  AOI21X1  g1524(.A0(new_n1909_), .A1(new_n1587_), .B0(new_n1588_), .Y(new_n1910_));
  OAI21X1  g1525(.A0(new_n1910_), .A1(new_n1586_), .B0(new_n1170_), .Y(new_n1911_));
  AOI21X1  g1526(.A0(new_n1911_), .A1(new_n1584_), .B0(new_n1585_), .Y(new_n1912_));
  OAI21X1  g1527(.A0(new_n1912_), .A1(new_n1583_), .B0(new_n1185_), .Y(new_n1913_));
  AOI21X1  g1528(.A0(new_n1913_), .A1(new_n1581_), .B0(new_n1582_), .Y(new_n1914_));
  OAI21X1  g1529(.A0(new_n1914_), .A1(new_n1580_), .B0(new_n1200_), .Y(new_n1915_));
  AOI21X1  g1530(.A0(new_n1915_), .A1(new_n1578_), .B0(new_n1579_), .Y(new_n1916_));
  OAI21X1  g1531(.A0(new_n1916_), .A1(new_n1577_), .B0(new_n1215_), .Y(new_n1917_));
  AOI21X1  g1532(.A0(new_n1917_), .A1(new_n1575_), .B0(new_n1576_), .Y(new_n1918_));
  OAI21X1  g1533(.A0(new_n1918_), .A1(new_n1574_), .B0(new_n1230_), .Y(new_n1919_));
  AOI21X1  g1534(.A0(new_n1919_), .A1(new_n1572_), .B0(new_n1573_), .Y(new_n1920_));
  OAI21X1  g1535(.A0(new_n1920_), .A1(new_n1571_), .B0(new_n1245_), .Y(new_n1921_));
  AOI21X1  g1536(.A0(new_n1921_), .A1(new_n1569_), .B0(new_n1570_), .Y(new_n1922_));
  OAI21X1  g1537(.A0(new_n1922_), .A1(new_n1568_), .B0(new_n1260_), .Y(new_n1923_));
  AOI21X1  g1538(.A0(new_n1923_), .A1(new_n1566_), .B0(new_n1567_), .Y(new_n1924_));
  OAI21X1  g1539(.A0(new_n1924_), .A1(new_n1565_), .B0(new_n1275_), .Y(new_n1925_));
  AOI21X1  g1540(.A0(new_n1925_), .A1(new_n1563_), .B0(new_n1564_), .Y(new_n1926_));
  OAI21X1  g1541(.A0(new_n1926_), .A1(new_n1562_), .B0(new_n1290_), .Y(new_n1927_));
  AOI21X1  g1542(.A0(new_n1927_), .A1(new_n1560_), .B0(new_n1561_), .Y(new_n1928_));
  OAI21X1  g1543(.A0(new_n1928_), .A1(new_n1559_), .B0(new_n1305_), .Y(new_n1929_));
  AOI21X1  g1544(.A0(new_n1929_), .A1(new_n1557_), .B0(new_n1558_), .Y(new_n1930_));
  OAI21X1  g1545(.A0(new_n1930_), .A1(new_n1556_), .B0(new_n1320_), .Y(new_n1931_));
  AOI21X1  g1546(.A0(new_n1931_), .A1(new_n1554_), .B0(new_n1555_), .Y(new_n1932_));
  OAI21X1  g1547(.A0(new_n1932_), .A1(new_n1553_), .B0(new_n1656_), .Y(new_n1933_));
  AOI21X1  g1548(.A0(new_n1933_), .A1(new_n1552_), .B0(new_n1893_), .Y(new_n1934_));
  OAI21X1  g1549(.A0(new_n1934_), .A1(new_n1395_), .B0(new_n403_), .Y(new_n1935_));
  OAI21X1  g1550(.A0(new_n725_), .A1(\priority[11] ), .B0(\req[11] ), .Y(new_n1936_));
  AOI21X1  g1551(.A0(new_n1935_), .A1(new_n1393_), .B0(new_n1936_), .Y(\grant[11] ));
  INVX1    g1552(.A(new_n714_), .Y(new_n1938_));
  NOR2X1   g1553(.A(new_n733_), .B(new_n417_), .Y(new_n1939_));
  OAI21X1  g1554(.A0(new_n1939_), .A1(new_n424_), .B0(new_n426_), .Y(new_n1940_));
  AOI21X1  g1555(.A0(new_n1940_), .A1(new_n431_), .B0(new_n434_), .Y(new_n1941_));
  OAI21X1  g1556(.A0(new_n1941_), .A1(new_n439_), .B0(new_n441_), .Y(new_n1942_));
  AOI21X1  g1557(.A0(new_n1942_), .A1(new_n446_), .B0(new_n449_), .Y(new_n1943_));
  OAI21X1  g1558(.A0(new_n1943_), .A1(new_n454_), .B0(new_n456_), .Y(new_n1944_));
  AOI21X1  g1559(.A0(new_n1944_), .A1(new_n461_), .B0(new_n464_), .Y(new_n1945_));
  OAI21X1  g1560(.A0(new_n1945_), .A1(new_n469_), .B0(new_n471_), .Y(new_n1946_));
  AOI21X1  g1561(.A0(new_n1946_), .A1(new_n476_), .B0(new_n479_), .Y(new_n1947_));
  OAI21X1  g1562(.A0(new_n1947_), .A1(new_n484_), .B0(new_n486_), .Y(new_n1948_));
  AOI21X1  g1563(.A0(new_n1948_), .A1(new_n491_), .B0(new_n494_), .Y(new_n1949_));
  OAI21X1  g1564(.A0(new_n1949_), .A1(new_n499_), .B0(new_n501_), .Y(new_n1950_));
  AOI21X1  g1565(.A0(new_n1950_), .A1(new_n506_), .B0(new_n509_), .Y(new_n1951_));
  OAI21X1  g1566(.A0(new_n1951_), .A1(new_n514_), .B0(new_n516_), .Y(new_n1952_));
  AOI21X1  g1567(.A0(new_n1952_), .A1(new_n521_), .B0(new_n524_), .Y(new_n1953_));
  OAI21X1  g1568(.A0(new_n1953_), .A1(new_n529_), .B0(new_n531_), .Y(new_n1954_));
  AOI21X1  g1569(.A0(new_n1954_), .A1(new_n536_), .B0(new_n539_), .Y(new_n1955_));
  OAI21X1  g1570(.A0(new_n1955_), .A1(new_n544_), .B0(new_n546_), .Y(new_n1956_));
  AOI21X1  g1571(.A0(new_n1956_), .A1(new_n551_), .B0(new_n554_), .Y(new_n1957_));
  OAI21X1  g1572(.A0(new_n1957_), .A1(new_n559_), .B0(new_n561_), .Y(new_n1958_));
  AOI21X1  g1573(.A0(new_n1958_), .A1(new_n566_), .B0(new_n569_), .Y(new_n1959_));
  OAI21X1  g1574(.A0(new_n1959_), .A1(new_n574_), .B0(new_n576_), .Y(new_n1960_));
  AOI21X1  g1575(.A0(new_n1960_), .A1(new_n581_), .B0(new_n584_), .Y(new_n1961_));
  OAI21X1  g1576(.A0(new_n1961_), .A1(new_n589_), .B0(new_n591_), .Y(new_n1962_));
  AOI21X1  g1577(.A0(new_n1962_), .A1(new_n596_), .B0(new_n599_), .Y(new_n1963_));
  OAI21X1  g1578(.A0(new_n1963_), .A1(new_n604_), .B0(new_n606_), .Y(new_n1964_));
  AOI21X1  g1579(.A0(new_n1964_), .A1(new_n611_), .B0(new_n614_), .Y(new_n1965_));
  OAI21X1  g1580(.A0(new_n1965_), .A1(new_n619_), .B0(new_n621_), .Y(new_n1966_));
  AOI21X1  g1581(.A0(new_n1966_), .A1(new_n626_), .B0(new_n629_), .Y(new_n1967_));
  OAI21X1  g1582(.A0(new_n1967_), .A1(new_n634_), .B0(new_n636_), .Y(new_n1968_));
  AOI21X1  g1583(.A0(new_n1968_), .A1(new_n641_), .B0(new_n644_), .Y(new_n1969_));
  OAI21X1  g1584(.A0(new_n1969_), .A1(new_n649_), .B0(new_n651_), .Y(new_n1970_));
  AOI21X1  g1585(.A0(new_n1970_), .A1(new_n656_), .B0(new_n659_), .Y(new_n1971_));
  OAI21X1  g1586(.A0(new_n1971_), .A1(new_n664_), .B0(new_n666_), .Y(new_n1972_));
  AOI21X1  g1587(.A0(new_n1972_), .A1(new_n671_), .B0(new_n674_), .Y(new_n1973_));
  OAI21X1  g1588(.A0(new_n1973_), .A1(new_n679_), .B0(new_n681_), .Y(new_n1974_));
  AOI21X1  g1589(.A0(new_n1974_), .A1(new_n686_), .B0(new_n689_), .Y(new_n1975_));
  OAI21X1  g1590(.A0(new_n1975_), .A1(new_n694_), .B0(new_n696_), .Y(new_n1976_));
  AOI21X1  g1591(.A0(new_n1976_), .A1(new_n701_), .B0(new_n1662_), .Y(new_n1977_));
  OAI21X1  g1592(.A0(new_n1977_), .A1(new_n1661_), .B0(new_n1705_), .Y(new_n1978_));
  AOI21X1  g1593(.A0(new_n1978_), .A1(new_n1660_), .B0(new_n1938_), .Y(new_n1979_));
  OAI21X1  g1594(.A0(new_n1979_), .A1(new_n1504_), .B0(new_n721_), .Y(new_n1980_));
  OAI21X1  g1595(.A0(new_n1039_), .A1(\priority[12] ), .B0(\req[12] ), .Y(new_n1981_));
  AOI21X1  g1596(.A0(new_n1980_), .A1(new_n1502_), .B0(new_n1981_), .Y(\grant[12] ));
  INVX1    g1597(.A(new_n1028_), .Y(new_n1983_));
  NOR2X1   g1598(.A(new_n1047_), .B(new_n735_), .Y(new_n1984_));
  OAI21X1  g1599(.A0(new_n1984_), .A1(new_n742_), .B0(new_n744_), .Y(new_n1985_));
  AOI21X1  g1600(.A0(new_n1985_), .A1(new_n749_), .B0(new_n752_), .Y(new_n1986_));
  OAI21X1  g1601(.A0(new_n1986_), .A1(new_n757_), .B0(new_n759_), .Y(new_n1987_));
  AOI21X1  g1602(.A0(new_n1987_), .A1(new_n764_), .B0(new_n767_), .Y(new_n1988_));
  OAI21X1  g1603(.A0(new_n1988_), .A1(new_n772_), .B0(new_n774_), .Y(new_n1989_));
  AOI21X1  g1604(.A0(new_n1989_), .A1(new_n779_), .B0(new_n782_), .Y(new_n1990_));
  OAI21X1  g1605(.A0(new_n1990_), .A1(new_n787_), .B0(new_n789_), .Y(new_n1991_));
  AOI21X1  g1606(.A0(new_n1991_), .A1(new_n794_), .B0(new_n797_), .Y(new_n1992_));
  OAI21X1  g1607(.A0(new_n1992_), .A1(new_n802_), .B0(new_n804_), .Y(new_n1993_));
  AOI21X1  g1608(.A0(new_n1993_), .A1(new_n809_), .B0(new_n812_), .Y(new_n1994_));
  OAI21X1  g1609(.A0(new_n1994_), .A1(new_n817_), .B0(new_n819_), .Y(new_n1995_));
  AOI21X1  g1610(.A0(new_n1995_), .A1(new_n824_), .B0(new_n827_), .Y(new_n1996_));
  OAI21X1  g1611(.A0(new_n1996_), .A1(new_n832_), .B0(new_n834_), .Y(new_n1997_));
  AOI21X1  g1612(.A0(new_n1997_), .A1(new_n839_), .B0(new_n842_), .Y(new_n1998_));
  OAI21X1  g1613(.A0(new_n1998_), .A1(new_n847_), .B0(new_n849_), .Y(new_n1999_));
  AOI21X1  g1614(.A0(new_n1999_), .A1(new_n854_), .B0(new_n857_), .Y(new_n2000_));
  OAI21X1  g1615(.A0(new_n2000_), .A1(new_n862_), .B0(new_n864_), .Y(new_n2001_));
  AOI21X1  g1616(.A0(new_n2001_), .A1(new_n869_), .B0(new_n872_), .Y(new_n2002_));
  OAI21X1  g1617(.A0(new_n2002_), .A1(new_n877_), .B0(new_n879_), .Y(new_n2003_));
  AOI21X1  g1618(.A0(new_n2003_), .A1(new_n884_), .B0(new_n887_), .Y(new_n2004_));
  OAI21X1  g1619(.A0(new_n2004_), .A1(new_n892_), .B0(new_n894_), .Y(new_n2005_));
  AOI21X1  g1620(.A0(new_n2005_), .A1(new_n899_), .B0(new_n902_), .Y(new_n2006_));
  OAI21X1  g1621(.A0(new_n2006_), .A1(new_n907_), .B0(new_n909_), .Y(new_n2007_));
  AOI21X1  g1622(.A0(new_n2007_), .A1(new_n914_), .B0(new_n917_), .Y(new_n2008_));
  OAI21X1  g1623(.A0(new_n2008_), .A1(new_n922_), .B0(new_n924_), .Y(new_n2009_));
  AOI21X1  g1624(.A0(new_n2009_), .A1(new_n929_), .B0(new_n932_), .Y(new_n2010_));
  OAI21X1  g1625(.A0(new_n2010_), .A1(new_n937_), .B0(new_n939_), .Y(new_n2011_));
  AOI21X1  g1626(.A0(new_n2011_), .A1(new_n944_), .B0(new_n947_), .Y(new_n2012_));
  OAI21X1  g1627(.A0(new_n2012_), .A1(new_n952_), .B0(new_n954_), .Y(new_n2013_));
  AOI21X1  g1628(.A0(new_n2013_), .A1(new_n959_), .B0(new_n962_), .Y(new_n2014_));
  OAI21X1  g1629(.A0(new_n2014_), .A1(new_n967_), .B0(new_n969_), .Y(new_n2015_));
  AOI21X1  g1630(.A0(new_n2015_), .A1(new_n974_), .B0(new_n977_), .Y(new_n2016_));
  OAI21X1  g1631(.A0(new_n2016_), .A1(new_n982_), .B0(new_n984_), .Y(new_n2017_));
  AOI21X1  g1632(.A0(new_n2017_), .A1(new_n989_), .B0(new_n992_), .Y(new_n2018_));
  OAI21X1  g1633(.A0(new_n2018_), .A1(new_n997_), .B0(new_n999_), .Y(new_n2019_));
  AOI21X1  g1634(.A0(new_n2019_), .A1(new_n1004_), .B0(new_n1007_), .Y(new_n2020_));
  OAI21X1  g1635(.A0(new_n2020_), .A1(new_n1012_), .B0(new_n1014_), .Y(new_n2021_));
  AOI21X1  g1636(.A0(new_n2021_), .A1(new_n1017_), .B0(new_n1711_), .Y(new_n2022_));
  OAI21X1  g1637(.A0(new_n2022_), .A1(new_n1710_), .B0(new_n1754_), .Y(new_n2023_));
  AOI21X1  g1638(.A0(new_n2023_), .A1(new_n1709_), .B0(new_n1983_), .Y(new_n2024_));
  OAI21X1  g1639(.A0(new_n2024_), .A1(new_n1613_), .B0(new_n1035_), .Y(new_n2025_));
  OAI21X1  g1640(.A0(new_n414_), .A1(\priority[13] ), .B0(\req[13] ), .Y(new_n2026_));
  AOI21X1  g1641(.A0(new_n2025_), .A1(new_n1611_), .B0(new_n2026_), .Y(\grant[13] ));
  NOR2X1   g1642(.A(new_n1049_), .B(new_n423_), .Y(new_n2028_));
  OAI21X1  g1643(.A0(new_n2028_), .A1(new_n1056_), .B0(new_n1058_), .Y(new_n2029_));
  AOI21X1  g1644(.A0(new_n2029_), .A1(new_n1063_), .B0(new_n1066_), .Y(new_n2030_));
  OAI21X1  g1645(.A0(new_n2030_), .A1(new_n1071_), .B0(new_n1073_), .Y(new_n2031_));
  AOI21X1  g1646(.A0(new_n2031_), .A1(new_n1078_), .B0(new_n1081_), .Y(new_n2032_));
  OAI21X1  g1647(.A0(new_n2032_), .A1(new_n1086_), .B0(new_n1088_), .Y(new_n2033_));
  AOI21X1  g1648(.A0(new_n2033_), .A1(new_n1093_), .B0(new_n1096_), .Y(new_n2034_));
  OAI21X1  g1649(.A0(new_n2034_), .A1(new_n1101_), .B0(new_n1103_), .Y(new_n2035_));
  AOI21X1  g1650(.A0(new_n2035_), .A1(new_n1108_), .B0(new_n1111_), .Y(new_n2036_));
  OAI21X1  g1651(.A0(new_n2036_), .A1(new_n1116_), .B0(new_n1118_), .Y(new_n2037_));
  AOI21X1  g1652(.A0(new_n2037_), .A1(new_n1123_), .B0(new_n1126_), .Y(new_n2038_));
  OAI21X1  g1653(.A0(new_n2038_), .A1(new_n1131_), .B0(new_n1133_), .Y(new_n2039_));
  AOI21X1  g1654(.A0(new_n2039_), .A1(new_n1138_), .B0(new_n1141_), .Y(new_n2040_));
  OAI21X1  g1655(.A0(new_n2040_), .A1(new_n1146_), .B0(new_n1148_), .Y(new_n2041_));
  AOI21X1  g1656(.A0(new_n2041_), .A1(new_n1153_), .B0(new_n1156_), .Y(new_n2042_));
  OAI21X1  g1657(.A0(new_n2042_), .A1(new_n1161_), .B0(new_n1163_), .Y(new_n2043_));
  AOI21X1  g1658(.A0(new_n2043_), .A1(new_n1168_), .B0(new_n1171_), .Y(new_n2044_));
  OAI21X1  g1659(.A0(new_n2044_), .A1(new_n1176_), .B0(new_n1178_), .Y(new_n2045_));
  AOI21X1  g1660(.A0(new_n2045_), .A1(new_n1183_), .B0(new_n1186_), .Y(new_n2046_));
  OAI21X1  g1661(.A0(new_n2046_), .A1(new_n1191_), .B0(new_n1193_), .Y(new_n2047_));
  AOI21X1  g1662(.A0(new_n2047_), .A1(new_n1198_), .B0(new_n1201_), .Y(new_n2048_));
  OAI21X1  g1663(.A0(new_n2048_), .A1(new_n1206_), .B0(new_n1208_), .Y(new_n2049_));
  AOI21X1  g1664(.A0(new_n2049_), .A1(new_n1213_), .B0(new_n1216_), .Y(new_n2050_));
  OAI21X1  g1665(.A0(new_n2050_), .A1(new_n1221_), .B0(new_n1223_), .Y(new_n2051_));
  AOI21X1  g1666(.A0(new_n2051_), .A1(new_n1228_), .B0(new_n1231_), .Y(new_n2052_));
  OAI21X1  g1667(.A0(new_n2052_), .A1(new_n1236_), .B0(new_n1238_), .Y(new_n2053_));
  AOI21X1  g1668(.A0(new_n2053_), .A1(new_n1243_), .B0(new_n1246_), .Y(new_n2054_));
  OAI21X1  g1669(.A0(new_n2054_), .A1(new_n1251_), .B0(new_n1253_), .Y(new_n2055_));
  AOI21X1  g1670(.A0(new_n2055_), .A1(new_n1258_), .B0(new_n1261_), .Y(new_n2056_));
  OAI21X1  g1671(.A0(new_n2056_), .A1(new_n1266_), .B0(new_n1268_), .Y(new_n2057_));
  AOI21X1  g1672(.A0(new_n2057_), .A1(new_n1273_), .B0(new_n1276_), .Y(new_n2058_));
  OAI21X1  g1673(.A0(new_n2058_), .A1(new_n1281_), .B0(new_n1283_), .Y(new_n2059_));
  AOI21X1  g1674(.A0(new_n2059_), .A1(new_n1288_), .B0(new_n1291_), .Y(new_n2060_));
  OAI21X1  g1675(.A0(new_n2060_), .A1(new_n1296_), .B0(new_n1298_), .Y(new_n2061_));
  AOI21X1  g1676(.A0(new_n2061_), .A1(new_n1303_), .B0(new_n1306_), .Y(new_n2062_));
  OAI21X1  g1677(.A0(new_n2062_), .A1(new_n1311_), .B0(new_n1313_), .Y(new_n2063_));
  AOI21X1  g1678(.A0(new_n2063_), .A1(new_n1318_), .B0(new_n1321_), .Y(new_n2064_));
  OAI21X1  g1679(.A0(new_n2064_), .A1(new_n1326_), .B0(new_n1328_), .Y(new_n2065_));
  AOI21X1  g1680(.A0(new_n2065_), .A1(new_n1331_), .B0(new_n1758_), .Y(new_n2066_));
  OAI21X1  g1681(.A0(new_n2066_), .A1(new_n394_), .B0(new_n396_), .Y(new_n2067_));
  AOI21X1  g1682(.A0(new_n2067_), .A1(new_n401_), .B0(new_n404_), .Y(new_n2068_));
  OAI21X1  g1683(.A0(new_n2068_), .A1(new_n409_), .B0(new_n411_), .Y(new_n2069_));
  OAI21X1  g1684(.A0(new_n732_), .A1(\priority[14] ), .B0(\req[14] ), .Y(new_n2070_));
  AOI21X1  g1685(.A0(new_n2069_), .A1(new_n416_), .B0(new_n2070_), .Y(\grant[14] ));
  NOR2X1   g1686(.A(new_n741_), .B(new_n425_), .Y(new_n2072_));
  OAI21X1  g1687(.A0(new_n2072_), .A1(new_n1389_), .B0(new_n433_), .Y(new_n2073_));
  AOI21X1  g1688(.A0(new_n2073_), .A1(new_n1387_), .B0(new_n1388_), .Y(new_n2074_));
  OAI21X1  g1689(.A0(new_n2074_), .A1(new_n1386_), .B0(new_n448_), .Y(new_n2075_));
  AOI21X1  g1690(.A0(new_n2075_), .A1(new_n1384_), .B0(new_n1385_), .Y(new_n2076_));
  OAI21X1  g1691(.A0(new_n2076_), .A1(new_n1383_), .B0(new_n463_), .Y(new_n2077_));
  AOI21X1  g1692(.A0(new_n2077_), .A1(new_n1381_), .B0(new_n1382_), .Y(new_n2078_));
  OAI21X1  g1693(.A0(new_n2078_), .A1(new_n1380_), .B0(new_n478_), .Y(new_n2079_));
  AOI21X1  g1694(.A0(new_n2079_), .A1(new_n1378_), .B0(new_n1379_), .Y(new_n2080_));
  OAI21X1  g1695(.A0(new_n2080_), .A1(new_n1377_), .B0(new_n493_), .Y(new_n2081_));
  AOI21X1  g1696(.A0(new_n2081_), .A1(new_n1375_), .B0(new_n1376_), .Y(new_n2082_));
  OAI21X1  g1697(.A0(new_n2082_), .A1(new_n1374_), .B0(new_n508_), .Y(new_n2083_));
  AOI21X1  g1698(.A0(new_n2083_), .A1(new_n1372_), .B0(new_n1373_), .Y(new_n2084_));
  OAI21X1  g1699(.A0(new_n2084_), .A1(new_n1371_), .B0(new_n523_), .Y(new_n2085_));
  AOI21X1  g1700(.A0(new_n2085_), .A1(new_n1369_), .B0(new_n1370_), .Y(new_n2086_));
  OAI21X1  g1701(.A0(new_n2086_), .A1(new_n1368_), .B0(new_n538_), .Y(new_n2087_));
  AOI21X1  g1702(.A0(new_n2087_), .A1(new_n1366_), .B0(new_n1367_), .Y(new_n2088_));
  OAI21X1  g1703(.A0(new_n2088_), .A1(new_n1365_), .B0(new_n553_), .Y(new_n2089_));
  AOI21X1  g1704(.A0(new_n2089_), .A1(new_n1363_), .B0(new_n1364_), .Y(new_n2090_));
  OAI21X1  g1705(.A0(new_n2090_), .A1(new_n1362_), .B0(new_n568_), .Y(new_n2091_));
  AOI21X1  g1706(.A0(new_n2091_), .A1(new_n1360_), .B0(new_n1361_), .Y(new_n2092_));
  OAI21X1  g1707(.A0(new_n2092_), .A1(new_n1359_), .B0(new_n583_), .Y(new_n2093_));
  AOI21X1  g1708(.A0(new_n2093_), .A1(new_n1357_), .B0(new_n1358_), .Y(new_n2094_));
  OAI21X1  g1709(.A0(new_n2094_), .A1(new_n1356_), .B0(new_n598_), .Y(new_n2095_));
  AOI21X1  g1710(.A0(new_n2095_), .A1(new_n1354_), .B0(new_n1355_), .Y(new_n2096_));
  OAI21X1  g1711(.A0(new_n2096_), .A1(new_n1353_), .B0(new_n613_), .Y(new_n2097_));
  AOI21X1  g1712(.A0(new_n2097_), .A1(new_n1351_), .B0(new_n1352_), .Y(new_n2098_));
  OAI21X1  g1713(.A0(new_n2098_), .A1(new_n1350_), .B0(new_n628_), .Y(new_n2099_));
  AOI21X1  g1714(.A0(new_n2099_), .A1(new_n1348_), .B0(new_n1349_), .Y(new_n2100_));
  OAI21X1  g1715(.A0(new_n2100_), .A1(new_n1347_), .B0(new_n643_), .Y(new_n2101_));
  AOI21X1  g1716(.A0(new_n2101_), .A1(new_n1345_), .B0(new_n1346_), .Y(new_n2102_));
  OAI21X1  g1717(.A0(new_n2102_), .A1(new_n1344_), .B0(new_n658_), .Y(new_n2103_));
  AOI21X1  g1718(.A0(new_n2103_), .A1(new_n1342_), .B0(new_n1343_), .Y(new_n2104_));
  OAI21X1  g1719(.A0(new_n2104_), .A1(new_n1341_), .B0(new_n673_), .Y(new_n2105_));
  AOI21X1  g1720(.A0(new_n2105_), .A1(new_n1339_), .B0(new_n1340_), .Y(new_n2106_));
  OAI21X1  g1721(.A0(new_n2106_), .A1(new_n1338_), .B0(new_n688_), .Y(new_n2107_));
  AOI21X1  g1722(.A0(new_n2107_), .A1(new_n1336_), .B0(new_n1337_), .Y(new_n2108_));
  OAI21X1  g1723(.A0(new_n2108_), .A1(new_n1335_), .B0(new_n1438_), .Y(new_n2109_));
  AOI21X1  g1724(.A0(new_n2109_), .A1(new_n1440_), .B0(new_n1803_), .Y(new_n2110_));
  OAI21X1  g1725(.A0(new_n2110_), .A1(new_n712_), .B0(new_n714_), .Y(new_n2111_));
  AOI21X1  g1726(.A0(new_n2111_), .A1(new_n719_), .B0(new_n722_), .Y(new_n2112_));
  OAI21X1  g1727(.A0(new_n2112_), .A1(new_n727_), .B0(new_n729_), .Y(new_n2113_));
  OAI21X1  g1728(.A0(new_n1046_), .A1(\priority[15] ), .B0(\req[15] ), .Y(new_n2114_));
  AOI21X1  g1729(.A0(new_n2113_), .A1(new_n734_), .B0(new_n2114_), .Y(\grant[15] ));
  NOR2X1   g1730(.A(new_n1055_), .B(new_n743_), .Y(new_n2116_));
  OAI21X1  g1731(.A0(new_n2116_), .A1(new_n1498_), .B0(new_n751_), .Y(new_n2117_));
  AOI21X1  g1732(.A0(new_n2117_), .A1(new_n1496_), .B0(new_n1497_), .Y(new_n2118_));
  OAI21X1  g1733(.A0(new_n2118_), .A1(new_n1495_), .B0(new_n766_), .Y(new_n2119_));
  AOI21X1  g1734(.A0(new_n2119_), .A1(new_n1493_), .B0(new_n1494_), .Y(new_n2120_));
  OAI21X1  g1735(.A0(new_n2120_), .A1(new_n1492_), .B0(new_n781_), .Y(new_n2121_));
  AOI21X1  g1736(.A0(new_n2121_), .A1(new_n1490_), .B0(new_n1491_), .Y(new_n2122_));
  OAI21X1  g1737(.A0(new_n2122_), .A1(new_n1489_), .B0(new_n796_), .Y(new_n2123_));
  AOI21X1  g1738(.A0(new_n2123_), .A1(new_n1487_), .B0(new_n1488_), .Y(new_n2124_));
  OAI21X1  g1739(.A0(new_n2124_), .A1(new_n1486_), .B0(new_n811_), .Y(new_n2125_));
  AOI21X1  g1740(.A0(new_n2125_), .A1(new_n1484_), .B0(new_n1485_), .Y(new_n2126_));
  OAI21X1  g1741(.A0(new_n2126_), .A1(new_n1483_), .B0(new_n826_), .Y(new_n2127_));
  AOI21X1  g1742(.A0(new_n2127_), .A1(new_n1481_), .B0(new_n1482_), .Y(new_n2128_));
  OAI21X1  g1743(.A0(new_n2128_), .A1(new_n1480_), .B0(new_n841_), .Y(new_n2129_));
  AOI21X1  g1744(.A0(new_n2129_), .A1(new_n1478_), .B0(new_n1479_), .Y(new_n2130_));
  OAI21X1  g1745(.A0(new_n2130_), .A1(new_n1477_), .B0(new_n856_), .Y(new_n2131_));
  AOI21X1  g1746(.A0(new_n2131_), .A1(new_n1475_), .B0(new_n1476_), .Y(new_n2132_));
  OAI21X1  g1747(.A0(new_n2132_), .A1(new_n1474_), .B0(new_n871_), .Y(new_n2133_));
  AOI21X1  g1748(.A0(new_n2133_), .A1(new_n1472_), .B0(new_n1473_), .Y(new_n2134_));
  OAI21X1  g1749(.A0(new_n2134_), .A1(new_n1471_), .B0(new_n886_), .Y(new_n2135_));
  AOI21X1  g1750(.A0(new_n2135_), .A1(new_n1469_), .B0(new_n1470_), .Y(new_n2136_));
  OAI21X1  g1751(.A0(new_n2136_), .A1(new_n1468_), .B0(new_n901_), .Y(new_n2137_));
  AOI21X1  g1752(.A0(new_n2137_), .A1(new_n1466_), .B0(new_n1467_), .Y(new_n2138_));
  OAI21X1  g1753(.A0(new_n2138_), .A1(new_n1465_), .B0(new_n916_), .Y(new_n2139_));
  AOI21X1  g1754(.A0(new_n2139_), .A1(new_n1463_), .B0(new_n1464_), .Y(new_n2140_));
  OAI21X1  g1755(.A0(new_n2140_), .A1(new_n1462_), .B0(new_n931_), .Y(new_n2141_));
  AOI21X1  g1756(.A0(new_n2141_), .A1(new_n1460_), .B0(new_n1461_), .Y(new_n2142_));
  OAI21X1  g1757(.A0(new_n2142_), .A1(new_n1459_), .B0(new_n946_), .Y(new_n2143_));
  AOI21X1  g1758(.A0(new_n2143_), .A1(new_n1457_), .B0(new_n1458_), .Y(new_n2144_));
  OAI21X1  g1759(.A0(new_n2144_), .A1(new_n1456_), .B0(new_n961_), .Y(new_n2145_));
  AOI21X1  g1760(.A0(new_n2145_), .A1(new_n1454_), .B0(new_n1455_), .Y(new_n2146_));
  OAI21X1  g1761(.A0(new_n2146_), .A1(new_n1453_), .B0(new_n976_), .Y(new_n2147_));
  AOI21X1  g1762(.A0(new_n2147_), .A1(new_n1451_), .B0(new_n1452_), .Y(new_n2148_));
  OAI21X1  g1763(.A0(new_n2148_), .A1(new_n1450_), .B0(new_n991_), .Y(new_n2149_));
  AOI21X1  g1764(.A0(new_n2149_), .A1(new_n1448_), .B0(new_n1449_), .Y(new_n2150_));
  OAI21X1  g1765(.A0(new_n2150_), .A1(new_n1447_), .B0(new_n1006_), .Y(new_n2151_));
  AOI21X1  g1766(.A0(new_n2151_), .A1(new_n1445_), .B0(new_n1446_), .Y(new_n2152_));
  OAI21X1  g1767(.A0(new_n2152_), .A1(new_n1444_), .B0(new_n1547_), .Y(new_n2153_));
  AOI21X1  g1768(.A0(new_n2153_), .A1(new_n1549_), .B0(new_n1848_), .Y(new_n2154_));
  OAI21X1  g1769(.A0(new_n2154_), .A1(new_n1026_), .B0(new_n1028_), .Y(new_n2155_));
  AOI21X1  g1770(.A0(new_n2155_), .A1(new_n1033_), .B0(new_n1036_), .Y(new_n2156_));
  OAI21X1  g1771(.A0(new_n2156_), .A1(new_n1041_), .B0(new_n1043_), .Y(new_n2157_));
  OAI21X1  g1772(.A0(new_n422_), .A1(\priority[16] ), .B0(\req[16] ), .Y(new_n2158_));
  AOI21X1  g1773(.A0(new_n2157_), .A1(new_n1048_), .B0(new_n2158_), .Y(\grant[16] ));
  NOR2X1   g1774(.A(new_n1057_), .B(new_n430_), .Y(new_n2160_));
  OAI21X1  g1775(.A0(new_n2160_), .A1(new_n1607_), .B0(new_n1065_), .Y(new_n2161_));
  AOI21X1  g1776(.A0(new_n2161_), .A1(new_n1605_), .B0(new_n1606_), .Y(new_n2162_));
  OAI21X1  g1777(.A0(new_n2162_), .A1(new_n1604_), .B0(new_n1080_), .Y(new_n2163_));
  AOI21X1  g1778(.A0(new_n2163_), .A1(new_n1602_), .B0(new_n1603_), .Y(new_n2164_));
  OAI21X1  g1779(.A0(new_n2164_), .A1(new_n1601_), .B0(new_n1095_), .Y(new_n2165_));
  AOI21X1  g1780(.A0(new_n2165_), .A1(new_n1599_), .B0(new_n1600_), .Y(new_n2166_));
  OAI21X1  g1781(.A0(new_n2166_), .A1(new_n1598_), .B0(new_n1110_), .Y(new_n2167_));
  AOI21X1  g1782(.A0(new_n2167_), .A1(new_n1596_), .B0(new_n1597_), .Y(new_n2168_));
  OAI21X1  g1783(.A0(new_n2168_), .A1(new_n1595_), .B0(new_n1125_), .Y(new_n2169_));
  AOI21X1  g1784(.A0(new_n2169_), .A1(new_n1593_), .B0(new_n1594_), .Y(new_n2170_));
  OAI21X1  g1785(.A0(new_n2170_), .A1(new_n1592_), .B0(new_n1140_), .Y(new_n2171_));
  AOI21X1  g1786(.A0(new_n2171_), .A1(new_n1590_), .B0(new_n1591_), .Y(new_n2172_));
  OAI21X1  g1787(.A0(new_n2172_), .A1(new_n1589_), .B0(new_n1155_), .Y(new_n2173_));
  AOI21X1  g1788(.A0(new_n2173_), .A1(new_n1587_), .B0(new_n1588_), .Y(new_n2174_));
  OAI21X1  g1789(.A0(new_n2174_), .A1(new_n1586_), .B0(new_n1170_), .Y(new_n2175_));
  AOI21X1  g1790(.A0(new_n2175_), .A1(new_n1584_), .B0(new_n1585_), .Y(new_n2176_));
  OAI21X1  g1791(.A0(new_n2176_), .A1(new_n1583_), .B0(new_n1185_), .Y(new_n2177_));
  AOI21X1  g1792(.A0(new_n2177_), .A1(new_n1581_), .B0(new_n1582_), .Y(new_n2178_));
  OAI21X1  g1793(.A0(new_n2178_), .A1(new_n1580_), .B0(new_n1200_), .Y(new_n2179_));
  AOI21X1  g1794(.A0(new_n2179_), .A1(new_n1578_), .B0(new_n1579_), .Y(new_n2180_));
  OAI21X1  g1795(.A0(new_n2180_), .A1(new_n1577_), .B0(new_n1215_), .Y(new_n2181_));
  AOI21X1  g1796(.A0(new_n2181_), .A1(new_n1575_), .B0(new_n1576_), .Y(new_n2182_));
  OAI21X1  g1797(.A0(new_n2182_), .A1(new_n1574_), .B0(new_n1230_), .Y(new_n2183_));
  AOI21X1  g1798(.A0(new_n2183_), .A1(new_n1572_), .B0(new_n1573_), .Y(new_n2184_));
  OAI21X1  g1799(.A0(new_n2184_), .A1(new_n1571_), .B0(new_n1245_), .Y(new_n2185_));
  AOI21X1  g1800(.A0(new_n2185_), .A1(new_n1569_), .B0(new_n1570_), .Y(new_n2186_));
  OAI21X1  g1801(.A0(new_n2186_), .A1(new_n1568_), .B0(new_n1260_), .Y(new_n2187_));
  AOI21X1  g1802(.A0(new_n2187_), .A1(new_n1566_), .B0(new_n1567_), .Y(new_n2188_));
  OAI21X1  g1803(.A0(new_n2188_), .A1(new_n1565_), .B0(new_n1275_), .Y(new_n2189_));
  AOI21X1  g1804(.A0(new_n2189_), .A1(new_n1563_), .B0(new_n1564_), .Y(new_n2190_));
  OAI21X1  g1805(.A0(new_n2190_), .A1(new_n1562_), .B0(new_n1290_), .Y(new_n2191_));
  AOI21X1  g1806(.A0(new_n2191_), .A1(new_n1560_), .B0(new_n1561_), .Y(new_n2192_));
  OAI21X1  g1807(.A0(new_n2192_), .A1(new_n1559_), .B0(new_n1305_), .Y(new_n2193_));
  AOI21X1  g1808(.A0(new_n2193_), .A1(new_n1557_), .B0(new_n1558_), .Y(new_n2194_));
  OAI21X1  g1809(.A0(new_n2194_), .A1(new_n1556_), .B0(new_n1320_), .Y(new_n2195_));
  AOI21X1  g1810(.A0(new_n2195_), .A1(new_n1554_), .B0(new_n1555_), .Y(new_n2196_));
  OAI21X1  g1811(.A0(new_n2196_), .A1(new_n1553_), .B0(new_n1656_), .Y(new_n2197_));
  AOI21X1  g1812(.A0(new_n2197_), .A1(new_n1552_), .B0(new_n1893_), .Y(new_n2198_));
  OAI21X1  g1813(.A0(new_n2198_), .A1(new_n1395_), .B0(new_n403_), .Y(new_n2199_));
  AOI21X1  g1814(.A0(new_n2199_), .A1(new_n1393_), .B0(new_n1394_), .Y(new_n2200_));
  OAI21X1  g1815(.A0(new_n2200_), .A1(new_n1392_), .B0(new_n418_), .Y(new_n2201_));
  OAI21X1  g1816(.A0(new_n740_), .A1(\priority[17] ), .B0(\req[17] ), .Y(new_n2202_));
  AOI21X1  g1817(.A0(new_n2201_), .A1(new_n1390_), .B0(new_n2202_), .Y(\grant[17] ));
  NOR2X1   g1818(.A(new_n748_), .B(new_n432_), .Y(new_n2204_));
  OAI21X1  g1819(.A0(new_n2204_), .A1(new_n439_), .B0(new_n441_), .Y(new_n2205_));
  AOI21X1  g1820(.A0(new_n2205_), .A1(new_n446_), .B0(new_n449_), .Y(new_n2206_));
  OAI21X1  g1821(.A0(new_n2206_), .A1(new_n454_), .B0(new_n456_), .Y(new_n2207_));
  AOI21X1  g1822(.A0(new_n2207_), .A1(new_n461_), .B0(new_n464_), .Y(new_n2208_));
  OAI21X1  g1823(.A0(new_n2208_), .A1(new_n469_), .B0(new_n471_), .Y(new_n2209_));
  AOI21X1  g1824(.A0(new_n2209_), .A1(new_n476_), .B0(new_n479_), .Y(new_n2210_));
  OAI21X1  g1825(.A0(new_n2210_), .A1(new_n484_), .B0(new_n486_), .Y(new_n2211_));
  AOI21X1  g1826(.A0(new_n2211_), .A1(new_n491_), .B0(new_n494_), .Y(new_n2212_));
  OAI21X1  g1827(.A0(new_n2212_), .A1(new_n499_), .B0(new_n501_), .Y(new_n2213_));
  AOI21X1  g1828(.A0(new_n2213_), .A1(new_n506_), .B0(new_n509_), .Y(new_n2214_));
  OAI21X1  g1829(.A0(new_n2214_), .A1(new_n514_), .B0(new_n516_), .Y(new_n2215_));
  AOI21X1  g1830(.A0(new_n2215_), .A1(new_n521_), .B0(new_n524_), .Y(new_n2216_));
  OAI21X1  g1831(.A0(new_n2216_), .A1(new_n529_), .B0(new_n531_), .Y(new_n2217_));
  AOI21X1  g1832(.A0(new_n2217_), .A1(new_n536_), .B0(new_n539_), .Y(new_n2218_));
  OAI21X1  g1833(.A0(new_n2218_), .A1(new_n544_), .B0(new_n546_), .Y(new_n2219_));
  AOI21X1  g1834(.A0(new_n2219_), .A1(new_n551_), .B0(new_n554_), .Y(new_n2220_));
  OAI21X1  g1835(.A0(new_n2220_), .A1(new_n559_), .B0(new_n561_), .Y(new_n2221_));
  AOI21X1  g1836(.A0(new_n2221_), .A1(new_n566_), .B0(new_n569_), .Y(new_n2222_));
  OAI21X1  g1837(.A0(new_n2222_), .A1(new_n574_), .B0(new_n576_), .Y(new_n2223_));
  AOI21X1  g1838(.A0(new_n2223_), .A1(new_n581_), .B0(new_n584_), .Y(new_n2224_));
  OAI21X1  g1839(.A0(new_n2224_), .A1(new_n589_), .B0(new_n591_), .Y(new_n2225_));
  AOI21X1  g1840(.A0(new_n2225_), .A1(new_n596_), .B0(new_n599_), .Y(new_n2226_));
  OAI21X1  g1841(.A0(new_n2226_), .A1(new_n604_), .B0(new_n606_), .Y(new_n2227_));
  AOI21X1  g1842(.A0(new_n2227_), .A1(new_n611_), .B0(new_n614_), .Y(new_n2228_));
  OAI21X1  g1843(.A0(new_n2228_), .A1(new_n619_), .B0(new_n621_), .Y(new_n2229_));
  AOI21X1  g1844(.A0(new_n2229_), .A1(new_n626_), .B0(new_n629_), .Y(new_n2230_));
  OAI21X1  g1845(.A0(new_n2230_), .A1(new_n634_), .B0(new_n636_), .Y(new_n2231_));
  AOI21X1  g1846(.A0(new_n2231_), .A1(new_n641_), .B0(new_n644_), .Y(new_n2232_));
  OAI21X1  g1847(.A0(new_n2232_), .A1(new_n649_), .B0(new_n651_), .Y(new_n2233_));
  AOI21X1  g1848(.A0(new_n2233_), .A1(new_n656_), .B0(new_n659_), .Y(new_n2234_));
  OAI21X1  g1849(.A0(new_n2234_), .A1(new_n664_), .B0(new_n666_), .Y(new_n2235_));
  AOI21X1  g1850(.A0(new_n2235_), .A1(new_n671_), .B0(new_n674_), .Y(new_n2236_));
  OAI21X1  g1851(.A0(new_n2236_), .A1(new_n679_), .B0(new_n681_), .Y(new_n2237_));
  AOI21X1  g1852(.A0(new_n2237_), .A1(new_n686_), .B0(new_n689_), .Y(new_n2238_));
  OAI21X1  g1853(.A0(new_n2238_), .A1(new_n694_), .B0(new_n696_), .Y(new_n2239_));
  AOI21X1  g1854(.A0(new_n2239_), .A1(new_n701_), .B0(new_n1662_), .Y(new_n2240_));
  OAI21X1  g1855(.A0(new_n2240_), .A1(new_n1661_), .B0(new_n1705_), .Y(new_n2241_));
  AOI21X1  g1856(.A0(new_n2241_), .A1(new_n1660_), .B0(new_n1938_), .Y(new_n2242_));
  OAI21X1  g1857(.A0(new_n2242_), .A1(new_n1504_), .B0(new_n721_), .Y(new_n2243_));
  AOI21X1  g1858(.A0(new_n2243_), .A1(new_n1502_), .B0(new_n1503_), .Y(new_n2244_));
  OAI21X1  g1859(.A0(new_n2244_), .A1(new_n1501_), .B0(new_n736_), .Y(new_n2245_));
  OAI21X1  g1860(.A0(new_n1054_), .A1(\priority[18] ), .B0(\req[18] ), .Y(new_n2246_));
  AOI21X1  g1861(.A0(new_n2245_), .A1(new_n1499_), .B0(new_n2246_), .Y(\grant[18] ));
  NOR2X1   g1862(.A(new_n1062_), .B(new_n750_), .Y(new_n2248_));
  OAI21X1  g1863(.A0(new_n2248_), .A1(new_n757_), .B0(new_n759_), .Y(new_n2249_));
  AOI21X1  g1864(.A0(new_n2249_), .A1(new_n764_), .B0(new_n767_), .Y(new_n2250_));
  OAI21X1  g1865(.A0(new_n2250_), .A1(new_n772_), .B0(new_n774_), .Y(new_n2251_));
  AOI21X1  g1866(.A0(new_n2251_), .A1(new_n779_), .B0(new_n782_), .Y(new_n2252_));
  OAI21X1  g1867(.A0(new_n2252_), .A1(new_n787_), .B0(new_n789_), .Y(new_n2253_));
  AOI21X1  g1868(.A0(new_n2253_), .A1(new_n794_), .B0(new_n797_), .Y(new_n2254_));
  OAI21X1  g1869(.A0(new_n2254_), .A1(new_n802_), .B0(new_n804_), .Y(new_n2255_));
  AOI21X1  g1870(.A0(new_n2255_), .A1(new_n809_), .B0(new_n812_), .Y(new_n2256_));
  OAI21X1  g1871(.A0(new_n2256_), .A1(new_n817_), .B0(new_n819_), .Y(new_n2257_));
  AOI21X1  g1872(.A0(new_n2257_), .A1(new_n824_), .B0(new_n827_), .Y(new_n2258_));
  OAI21X1  g1873(.A0(new_n2258_), .A1(new_n832_), .B0(new_n834_), .Y(new_n2259_));
  AOI21X1  g1874(.A0(new_n2259_), .A1(new_n839_), .B0(new_n842_), .Y(new_n2260_));
  OAI21X1  g1875(.A0(new_n2260_), .A1(new_n847_), .B0(new_n849_), .Y(new_n2261_));
  AOI21X1  g1876(.A0(new_n2261_), .A1(new_n854_), .B0(new_n857_), .Y(new_n2262_));
  OAI21X1  g1877(.A0(new_n2262_), .A1(new_n862_), .B0(new_n864_), .Y(new_n2263_));
  AOI21X1  g1878(.A0(new_n2263_), .A1(new_n869_), .B0(new_n872_), .Y(new_n2264_));
  OAI21X1  g1879(.A0(new_n2264_), .A1(new_n877_), .B0(new_n879_), .Y(new_n2265_));
  AOI21X1  g1880(.A0(new_n2265_), .A1(new_n884_), .B0(new_n887_), .Y(new_n2266_));
  OAI21X1  g1881(.A0(new_n2266_), .A1(new_n892_), .B0(new_n894_), .Y(new_n2267_));
  AOI21X1  g1882(.A0(new_n2267_), .A1(new_n899_), .B0(new_n902_), .Y(new_n2268_));
  OAI21X1  g1883(.A0(new_n2268_), .A1(new_n907_), .B0(new_n909_), .Y(new_n2269_));
  AOI21X1  g1884(.A0(new_n2269_), .A1(new_n914_), .B0(new_n917_), .Y(new_n2270_));
  OAI21X1  g1885(.A0(new_n2270_), .A1(new_n922_), .B0(new_n924_), .Y(new_n2271_));
  AOI21X1  g1886(.A0(new_n2271_), .A1(new_n929_), .B0(new_n932_), .Y(new_n2272_));
  OAI21X1  g1887(.A0(new_n2272_), .A1(new_n937_), .B0(new_n939_), .Y(new_n2273_));
  AOI21X1  g1888(.A0(new_n2273_), .A1(new_n944_), .B0(new_n947_), .Y(new_n2274_));
  OAI21X1  g1889(.A0(new_n2274_), .A1(new_n952_), .B0(new_n954_), .Y(new_n2275_));
  AOI21X1  g1890(.A0(new_n2275_), .A1(new_n959_), .B0(new_n962_), .Y(new_n2276_));
  OAI21X1  g1891(.A0(new_n2276_), .A1(new_n967_), .B0(new_n969_), .Y(new_n2277_));
  AOI21X1  g1892(.A0(new_n2277_), .A1(new_n974_), .B0(new_n977_), .Y(new_n2278_));
  OAI21X1  g1893(.A0(new_n2278_), .A1(new_n982_), .B0(new_n984_), .Y(new_n2279_));
  AOI21X1  g1894(.A0(new_n2279_), .A1(new_n989_), .B0(new_n992_), .Y(new_n2280_));
  OAI21X1  g1895(.A0(new_n2280_), .A1(new_n997_), .B0(new_n999_), .Y(new_n2281_));
  AOI21X1  g1896(.A0(new_n2281_), .A1(new_n1004_), .B0(new_n1007_), .Y(new_n2282_));
  OAI21X1  g1897(.A0(new_n2282_), .A1(new_n1012_), .B0(new_n1014_), .Y(new_n2283_));
  AOI21X1  g1898(.A0(new_n2283_), .A1(new_n1017_), .B0(new_n1711_), .Y(new_n2284_));
  OAI21X1  g1899(.A0(new_n2284_), .A1(new_n1710_), .B0(new_n1754_), .Y(new_n2285_));
  AOI21X1  g1900(.A0(new_n2285_), .A1(new_n1709_), .B0(new_n1983_), .Y(new_n2286_));
  OAI21X1  g1901(.A0(new_n2286_), .A1(new_n1613_), .B0(new_n1035_), .Y(new_n2287_));
  AOI21X1  g1902(.A0(new_n2287_), .A1(new_n1611_), .B0(new_n1612_), .Y(new_n2288_));
  OAI21X1  g1903(.A0(new_n2288_), .A1(new_n1610_), .B0(new_n1050_), .Y(new_n2289_));
  OAI21X1  g1904(.A0(new_n429_), .A1(\priority[19] ), .B0(\req[19] ), .Y(new_n2290_));
  AOI21X1  g1905(.A0(new_n2289_), .A1(new_n1608_), .B0(new_n2290_), .Y(\grant[19] ));
  NOR2X1   g1906(.A(new_n1064_), .B(new_n438_), .Y(new_n2292_));
  OAI21X1  g1907(.A0(new_n2292_), .A1(new_n1071_), .B0(new_n1073_), .Y(new_n2293_));
  AOI21X1  g1908(.A0(new_n2293_), .A1(new_n1078_), .B0(new_n1081_), .Y(new_n2294_));
  OAI21X1  g1909(.A0(new_n2294_), .A1(new_n1086_), .B0(new_n1088_), .Y(new_n2295_));
  AOI21X1  g1910(.A0(new_n2295_), .A1(new_n1093_), .B0(new_n1096_), .Y(new_n2296_));
  OAI21X1  g1911(.A0(new_n2296_), .A1(new_n1101_), .B0(new_n1103_), .Y(new_n2297_));
  AOI21X1  g1912(.A0(new_n2297_), .A1(new_n1108_), .B0(new_n1111_), .Y(new_n2298_));
  OAI21X1  g1913(.A0(new_n2298_), .A1(new_n1116_), .B0(new_n1118_), .Y(new_n2299_));
  AOI21X1  g1914(.A0(new_n2299_), .A1(new_n1123_), .B0(new_n1126_), .Y(new_n2300_));
  OAI21X1  g1915(.A0(new_n2300_), .A1(new_n1131_), .B0(new_n1133_), .Y(new_n2301_));
  AOI21X1  g1916(.A0(new_n2301_), .A1(new_n1138_), .B0(new_n1141_), .Y(new_n2302_));
  OAI21X1  g1917(.A0(new_n2302_), .A1(new_n1146_), .B0(new_n1148_), .Y(new_n2303_));
  AOI21X1  g1918(.A0(new_n2303_), .A1(new_n1153_), .B0(new_n1156_), .Y(new_n2304_));
  OAI21X1  g1919(.A0(new_n2304_), .A1(new_n1161_), .B0(new_n1163_), .Y(new_n2305_));
  AOI21X1  g1920(.A0(new_n2305_), .A1(new_n1168_), .B0(new_n1171_), .Y(new_n2306_));
  OAI21X1  g1921(.A0(new_n2306_), .A1(new_n1176_), .B0(new_n1178_), .Y(new_n2307_));
  AOI21X1  g1922(.A0(new_n2307_), .A1(new_n1183_), .B0(new_n1186_), .Y(new_n2308_));
  OAI21X1  g1923(.A0(new_n2308_), .A1(new_n1191_), .B0(new_n1193_), .Y(new_n2309_));
  AOI21X1  g1924(.A0(new_n2309_), .A1(new_n1198_), .B0(new_n1201_), .Y(new_n2310_));
  OAI21X1  g1925(.A0(new_n2310_), .A1(new_n1206_), .B0(new_n1208_), .Y(new_n2311_));
  AOI21X1  g1926(.A0(new_n2311_), .A1(new_n1213_), .B0(new_n1216_), .Y(new_n2312_));
  OAI21X1  g1927(.A0(new_n2312_), .A1(new_n1221_), .B0(new_n1223_), .Y(new_n2313_));
  AOI21X1  g1928(.A0(new_n2313_), .A1(new_n1228_), .B0(new_n1231_), .Y(new_n2314_));
  OAI21X1  g1929(.A0(new_n2314_), .A1(new_n1236_), .B0(new_n1238_), .Y(new_n2315_));
  AOI21X1  g1930(.A0(new_n2315_), .A1(new_n1243_), .B0(new_n1246_), .Y(new_n2316_));
  OAI21X1  g1931(.A0(new_n2316_), .A1(new_n1251_), .B0(new_n1253_), .Y(new_n2317_));
  AOI21X1  g1932(.A0(new_n2317_), .A1(new_n1258_), .B0(new_n1261_), .Y(new_n2318_));
  OAI21X1  g1933(.A0(new_n2318_), .A1(new_n1266_), .B0(new_n1268_), .Y(new_n2319_));
  AOI21X1  g1934(.A0(new_n2319_), .A1(new_n1273_), .B0(new_n1276_), .Y(new_n2320_));
  OAI21X1  g1935(.A0(new_n2320_), .A1(new_n1281_), .B0(new_n1283_), .Y(new_n2321_));
  AOI21X1  g1936(.A0(new_n2321_), .A1(new_n1288_), .B0(new_n1291_), .Y(new_n2322_));
  OAI21X1  g1937(.A0(new_n2322_), .A1(new_n1296_), .B0(new_n1298_), .Y(new_n2323_));
  AOI21X1  g1938(.A0(new_n2323_), .A1(new_n1303_), .B0(new_n1306_), .Y(new_n2324_));
  OAI21X1  g1939(.A0(new_n2324_), .A1(new_n1311_), .B0(new_n1313_), .Y(new_n2325_));
  AOI21X1  g1940(.A0(new_n2325_), .A1(new_n1318_), .B0(new_n1321_), .Y(new_n2326_));
  OAI21X1  g1941(.A0(new_n2326_), .A1(new_n1326_), .B0(new_n1328_), .Y(new_n2327_));
  AOI21X1  g1942(.A0(new_n2327_), .A1(new_n1331_), .B0(new_n1758_), .Y(new_n2328_));
  OAI21X1  g1943(.A0(new_n2328_), .A1(new_n394_), .B0(new_n396_), .Y(new_n2329_));
  AOI21X1  g1944(.A0(new_n2329_), .A1(new_n401_), .B0(new_n404_), .Y(new_n2330_));
  OAI21X1  g1945(.A0(new_n2330_), .A1(new_n409_), .B0(new_n411_), .Y(new_n2331_));
  AOI21X1  g1946(.A0(new_n2331_), .A1(new_n416_), .B0(new_n419_), .Y(new_n2332_));
  OAI21X1  g1947(.A0(new_n2332_), .A1(new_n424_), .B0(new_n426_), .Y(new_n2333_));
  OAI21X1  g1948(.A0(new_n747_), .A1(\priority[20] ), .B0(\req[20] ), .Y(new_n2334_));
  AOI21X1  g1949(.A0(new_n2333_), .A1(new_n431_), .B0(new_n2334_), .Y(\grant[20] ));
  NOR2X1   g1950(.A(new_n756_), .B(new_n440_), .Y(new_n2336_));
  OAI21X1  g1951(.A0(new_n2336_), .A1(new_n1386_), .B0(new_n448_), .Y(new_n2337_));
  AOI21X1  g1952(.A0(new_n2337_), .A1(new_n1384_), .B0(new_n1385_), .Y(new_n2338_));
  OAI21X1  g1953(.A0(new_n2338_), .A1(new_n1383_), .B0(new_n463_), .Y(new_n2339_));
  AOI21X1  g1954(.A0(new_n2339_), .A1(new_n1381_), .B0(new_n1382_), .Y(new_n2340_));
  OAI21X1  g1955(.A0(new_n2340_), .A1(new_n1380_), .B0(new_n478_), .Y(new_n2341_));
  AOI21X1  g1956(.A0(new_n2341_), .A1(new_n1378_), .B0(new_n1379_), .Y(new_n2342_));
  OAI21X1  g1957(.A0(new_n2342_), .A1(new_n1377_), .B0(new_n493_), .Y(new_n2343_));
  AOI21X1  g1958(.A0(new_n2343_), .A1(new_n1375_), .B0(new_n1376_), .Y(new_n2344_));
  OAI21X1  g1959(.A0(new_n2344_), .A1(new_n1374_), .B0(new_n508_), .Y(new_n2345_));
  AOI21X1  g1960(.A0(new_n2345_), .A1(new_n1372_), .B0(new_n1373_), .Y(new_n2346_));
  OAI21X1  g1961(.A0(new_n2346_), .A1(new_n1371_), .B0(new_n523_), .Y(new_n2347_));
  AOI21X1  g1962(.A0(new_n2347_), .A1(new_n1369_), .B0(new_n1370_), .Y(new_n2348_));
  OAI21X1  g1963(.A0(new_n2348_), .A1(new_n1368_), .B0(new_n538_), .Y(new_n2349_));
  AOI21X1  g1964(.A0(new_n2349_), .A1(new_n1366_), .B0(new_n1367_), .Y(new_n2350_));
  OAI21X1  g1965(.A0(new_n2350_), .A1(new_n1365_), .B0(new_n553_), .Y(new_n2351_));
  AOI21X1  g1966(.A0(new_n2351_), .A1(new_n1363_), .B0(new_n1364_), .Y(new_n2352_));
  OAI21X1  g1967(.A0(new_n2352_), .A1(new_n1362_), .B0(new_n568_), .Y(new_n2353_));
  AOI21X1  g1968(.A0(new_n2353_), .A1(new_n1360_), .B0(new_n1361_), .Y(new_n2354_));
  OAI21X1  g1969(.A0(new_n2354_), .A1(new_n1359_), .B0(new_n583_), .Y(new_n2355_));
  AOI21X1  g1970(.A0(new_n2355_), .A1(new_n1357_), .B0(new_n1358_), .Y(new_n2356_));
  OAI21X1  g1971(.A0(new_n2356_), .A1(new_n1356_), .B0(new_n598_), .Y(new_n2357_));
  AOI21X1  g1972(.A0(new_n2357_), .A1(new_n1354_), .B0(new_n1355_), .Y(new_n2358_));
  OAI21X1  g1973(.A0(new_n2358_), .A1(new_n1353_), .B0(new_n613_), .Y(new_n2359_));
  AOI21X1  g1974(.A0(new_n2359_), .A1(new_n1351_), .B0(new_n1352_), .Y(new_n2360_));
  OAI21X1  g1975(.A0(new_n2360_), .A1(new_n1350_), .B0(new_n628_), .Y(new_n2361_));
  AOI21X1  g1976(.A0(new_n2361_), .A1(new_n1348_), .B0(new_n1349_), .Y(new_n2362_));
  OAI21X1  g1977(.A0(new_n2362_), .A1(new_n1347_), .B0(new_n643_), .Y(new_n2363_));
  AOI21X1  g1978(.A0(new_n2363_), .A1(new_n1345_), .B0(new_n1346_), .Y(new_n2364_));
  OAI21X1  g1979(.A0(new_n2364_), .A1(new_n1344_), .B0(new_n658_), .Y(new_n2365_));
  AOI21X1  g1980(.A0(new_n2365_), .A1(new_n1342_), .B0(new_n1343_), .Y(new_n2366_));
  OAI21X1  g1981(.A0(new_n2366_), .A1(new_n1341_), .B0(new_n673_), .Y(new_n2367_));
  AOI21X1  g1982(.A0(new_n2367_), .A1(new_n1339_), .B0(new_n1340_), .Y(new_n2368_));
  OAI21X1  g1983(.A0(new_n2368_), .A1(new_n1338_), .B0(new_n688_), .Y(new_n2369_));
  AOI21X1  g1984(.A0(new_n2369_), .A1(new_n1336_), .B0(new_n1337_), .Y(new_n2370_));
  OAI21X1  g1985(.A0(new_n2370_), .A1(new_n1335_), .B0(new_n1438_), .Y(new_n2371_));
  AOI21X1  g1986(.A0(new_n2371_), .A1(new_n1440_), .B0(new_n1803_), .Y(new_n2372_));
  OAI21X1  g1987(.A0(new_n2372_), .A1(new_n712_), .B0(new_n714_), .Y(new_n2373_));
  AOI21X1  g1988(.A0(new_n2373_), .A1(new_n719_), .B0(new_n722_), .Y(new_n2374_));
  OAI21X1  g1989(.A0(new_n2374_), .A1(new_n727_), .B0(new_n729_), .Y(new_n2375_));
  AOI21X1  g1990(.A0(new_n2375_), .A1(new_n734_), .B0(new_n737_), .Y(new_n2376_));
  OAI21X1  g1991(.A0(new_n2376_), .A1(new_n742_), .B0(new_n744_), .Y(new_n2377_));
  OAI21X1  g1992(.A0(new_n1061_), .A1(\priority[21] ), .B0(\req[21] ), .Y(new_n2378_));
  AOI21X1  g1993(.A0(new_n2377_), .A1(new_n749_), .B0(new_n2378_), .Y(\grant[21] ));
  NOR2X1   g1994(.A(new_n1070_), .B(new_n758_), .Y(new_n2380_));
  OAI21X1  g1995(.A0(new_n2380_), .A1(new_n1495_), .B0(new_n766_), .Y(new_n2381_));
  AOI21X1  g1996(.A0(new_n2381_), .A1(new_n1493_), .B0(new_n1494_), .Y(new_n2382_));
  OAI21X1  g1997(.A0(new_n2382_), .A1(new_n1492_), .B0(new_n781_), .Y(new_n2383_));
  AOI21X1  g1998(.A0(new_n2383_), .A1(new_n1490_), .B0(new_n1491_), .Y(new_n2384_));
  OAI21X1  g1999(.A0(new_n2384_), .A1(new_n1489_), .B0(new_n796_), .Y(new_n2385_));
  AOI21X1  g2000(.A0(new_n2385_), .A1(new_n1487_), .B0(new_n1488_), .Y(new_n2386_));
  OAI21X1  g2001(.A0(new_n2386_), .A1(new_n1486_), .B0(new_n811_), .Y(new_n2387_));
  AOI21X1  g2002(.A0(new_n2387_), .A1(new_n1484_), .B0(new_n1485_), .Y(new_n2388_));
  OAI21X1  g2003(.A0(new_n2388_), .A1(new_n1483_), .B0(new_n826_), .Y(new_n2389_));
  AOI21X1  g2004(.A0(new_n2389_), .A1(new_n1481_), .B0(new_n1482_), .Y(new_n2390_));
  OAI21X1  g2005(.A0(new_n2390_), .A1(new_n1480_), .B0(new_n841_), .Y(new_n2391_));
  AOI21X1  g2006(.A0(new_n2391_), .A1(new_n1478_), .B0(new_n1479_), .Y(new_n2392_));
  OAI21X1  g2007(.A0(new_n2392_), .A1(new_n1477_), .B0(new_n856_), .Y(new_n2393_));
  AOI21X1  g2008(.A0(new_n2393_), .A1(new_n1475_), .B0(new_n1476_), .Y(new_n2394_));
  OAI21X1  g2009(.A0(new_n2394_), .A1(new_n1474_), .B0(new_n871_), .Y(new_n2395_));
  AOI21X1  g2010(.A0(new_n2395_), .A1(new_n1472_), .B0(new_n1473_), .Y(new_n2396_));
  OAI21X1  g2011(.A0(new_n2396_), .A1(new_n1471_), .B0(new_n886_), .Y(new_n2397_));
  AOI21X1  g2012(.A0(new_n2397_), .A1(new_n1469_), .B0(new_n1470_), .Y(new_n2398_));
  OAI21X1  g2013(.A0(new_n2398_), .A1(new_n1468_), .B0(new_n901_), .Y(new_n2399_));
  AOI21X1  g2014(.A0(new_n2399_), .A1(new_n1466_), .B0(new_n1467_), .Y(new_n2400_));
  OAI21X1  g2015(.A0(new_n2400_), .A1(new_n1465_), .B0(new_n916_), .Y(new_n2401_));
  AOI21X1  g2016(.A0(new_n2401_), .A1(new_n1463_), .B0(new_n1464_), .Y(new_n2402_));
  OAI21X1  g2017(.A0(new_n2402_), .A1(new_n1462_), .B0(new_n931_), .Y(new_n2403_));
  AOI21X1  g2018(.A0(new_n2403_), .A1(new_n1460_), .B0(new_n1461_), .Y(new_n2404_));
  OAI21X1  g2019(.A0(new_n2404_), .A1(new_n1459_), .B0(new_n946_), .Y(new_n2405_));
  AOI21X1  g2020(.A0(new_n2405_), .A1(new_n1457_), .B0(new_n1458_), .Y(new_n2406_));
  OAI21X1  g2021(.A0(new_n2406_), .A1(new_n1456_), .B0(new_n961_), .Y(new_n2407_));
  AOI21X1  g2022(.A0(new_n2407_), .A1(new_n1454_), .B0(new_n1455_), .Y(new_n2408_));
  OAI21X1  g2023(.A0(new_n2408_), .A1(new_n1453_), .B0(new_n976_), .Y(new_n2409_));
  AOI21X1  g2024(.A0(new_n2409_), .A1(new_n1451_), .B0(new_n1452_), .Y(new_n2410_));
  OAI21X1  g2025(.A0(new_n2410_), .A1(new_n1450_), .B0(new_n991_), .Y(new_n2411_));
  AOI21X1  g2026(.A0(new_n2411_), .A1(new_n1448_), .B0(new_n1449_), .Y(new_n2412_));
  OAI21X1  g2027(.A0(new_n2412_), .A1(new_n1447_), .B0(new_n1006_), .Y(new_n2413_));
  AOI21X1  g2028(.A0(new_n2413_), .A1(new_n1445_), .B0(new_n1446_), .Y(new_n2414_));
  OAI21X1  g2029(.A0(new_n2414_), .A1(new_n1444_), .B0(new_n1547_), .Y(new_n2415_));
  AOI21X1  g2030(.A0(new_n2415_), .A1(new_n1549_), .B0(new_n1848_), .Y(new_n2416_));
  OAI21X1  g2031(.A0(new_n2416_), .A1(new_n1026_), .B0(new_n1028_), .Y(new_n2417_));
  AOI21X1  g2032(.A0(new_n2417_), .A1(new_n1033_), .B0(new_n1036_), .Y(new_n2418_));
  OAI21X1  g2033(.A0(new_n2418_), .A1(new_n1041_), .B0(new_n1043_), .Y(new_n2419_));
  AOI21X1  g2034(.A0(new_n2419_), .A1(new_n1048_), .B0(new_n1051_), .Y(new_n2420_));
  OAI21X1  g2035(.A0(new_n2420_), .A1(new_n1056_), .B0(new_n1058_), .Y(new_n2421_));
  OAI21X1  g2036(.A0(new_n437_), .A1(\priority[22] ), .B0(\req[22] ), .Y(new_n2422_));
  AOI21X1  g2037(.A0(new_n2421_), .A1(new_n1063_), .B0(new_n2422_), .Y(\grant[22] ));
  NOR2X1   g2038(.A(new_n1072_), .B(new_n445_), .Y(new_n2424_));
  OAI21X1  g2039(.A0(new_n2424_), .A1(new_n1604_), .B0(new_n1080_), .Y(new_n2425_));
  AOI21X1  g2040(.A0(new_n2425_), .A1(new_n1602_), .B0(new_n1603_), .Y(new_n2426_));
  OAI21X1  g2041(.A0(new_n2426_), .A1(new_n1601_), .B0(new_n1095_), .Y(new_n2427_));
  AOI21X1  g2042(.A0(new_n2427_), .A1(new_n1599_), .B0(new_n1600_), .Y(new_n2428_));
  OAI21X1  g2043(.A0(new_n2428_), .A1(new_n1598_), .B0(new_n1110_), .Y(new_n2429_));
  AOI21X1  g2044(.A0(new_n2429_), .A1(new_n1596_), .B0(new_n1597_), .Y(new_n2430_));
  OAI21X1  g2045(.A0(new_n2430_), .A1(new_n1595_), .B0(new_n1125_), .Y(new_n2431_));
  AOI21X1  g2046(.A0(new_n2431_), .A1(new_n1593_), .B0(new_n1594_), .Y(new_n2432_));
  OAI21X1  g2047(.A0(new_n2432_), .A1(new_n1592_), .B0(new_n1140_), .Y(new_n2433_));
  AOI21X1  g2048(.A0(new_n2433_), .A1(new_n1590_), .B0(new_n1591_), .Y(new_n2434_));
  OAI21X1  g2049(.A0(new_n2434_), .A1(new_n1589_), .B0(new_n1155_), .Y(new_n2435_));
  AOI21X1  g2050(.A0(new_n2435_), .A1(new_n1587_), .B0(new_n1588_), .Y(new_n2436_));
  OAI21X1  g2051(.A0(new_n2436_), .A1(new_n1586_), .B0(new_n1170_), .Y(new_n2437_));
  AOI21X1  g2052(.A0(new_n2437_), .A1(new_n1584_), .B0(new_n1585_), .Y(new_n2438_));
  OAI21X1  g2053(.A0(new_n2438_), .A1(new_n1583_), .B0(new_n1185_), .Y(new_n2439_));
  AOI21X1  g2054(.A0(new_n2439_), .A1(new_n1581_), .B0(new_n1582_), .Y(new_n2440_));
  OAI21X1  g2055(.A0(new_n2440_), .A1(new_n1580_), .B0(new_n1200_), .Y(new_n2441_));
  AOI21X1  g2056(.A0(new_n2441_), .A1(new_n1578_), .B0(new_n1579_), .Y(new_n2442_));
  OAI21X1  g2057(.A0(new_n2442_), .A1(new_n1577_), .B0(new_n1215_), .Y(new_n2443_));
  AOI21X1  g2058(.A0(new_n2443_), .A1(new_n1575_), .B0(new_n1576_), .Y(new_n2444_));
  OAI21X1  g2059(.A0(new_n2444_), .A1(new_n1574_), .B0(new_n1230_), .Y(new_n2445_));
  AOI21X1  g2060(.A0(new_n2445_), .A1(new_n1572_), .B0(new_n1573_), .Y(new_n2446_));
  OAI21X1  g2061(.A0(new_n2446_), .A1(new_n1571_), .B0(new_n1245_), .Y(new_n2447_));
  AOI21X1  g2062(.A0(new_n2447_), .A1(new_n1569_), .B0(new_n1570_), .Y(new_n2448_));
  OAI21X1  g2063(.A0(new_n2448_), .A1(new_n1568_), .B0(new_n1260_), .Y(new_n2449_));
  AOI21X1  g2064(.A0(new_n2449_), .A1(new_n1566_), .B0(new_n1567_), .Y(new_n2450_));
  OAI21X1  g2065(.A0(new_n2450_), .A1(new_n1565_), .B0(new_n1275_), .Y(new_n2451_));
  AOI21X1  g2066(.A0(new_n2451_), .A1(new_n1563_), .B0(new_n1564_), .Y(new_n2452_));
  OAI21X1  g2067(.A0(new_n2452_), .A1(new_n1562_), .B0(new_n1290_), .Y(new_n2453_));
  AOI21X1  g2068(.A0(new_n2453_), .A1(new_n1560_), .B0(new_n1561_), .Y(new_n2454_));
  OAI21X1  g2069(.A0(new_n2454_), .A1(new_n1559_), .B0(new_n1305_), .Y(new_n2455_));
  AOI21X1  g2070(.A0(new_n2455_), .A1(new_n1557_), .B0(new_n1558_), .Y(new_n2456_));
  OAI21X1  g2071(.A0(new_n2456_), .A1(new_n1556_), .B0(new_n1320_), .Y(new_n2457_));
  AOI21X1  g2072(.A0(new_n2457_), .A1(new_n1554_), .B0(new_n1555_), .Y(new_n2458_));
  OAI21X1  g2073(.A0(new_n2458_), .A1(new_n1553_), .B0(new_n1656_), .Y(new_n2459_));
  AOI21X1  g2074(.A0(new_n2459_), .A1(new_n1552_), .B0(new_n1893_), .Y(new_n2460_));
  OAI21X1  g2075(.A0(new_n2460_), .A1(new_n1395_), .B0(new_n403_), .Y(new_n2461_));
  AOI21X1  g2076(.A0(new_n2461_), .A1(new_n1393_), .B0(new_n1394_), .Y(new_n2462_));
  OAI21X1  g2077(.A0(new_n2462_), .A1(new_n1392_), .B0(new_n418_), .Y(new_n2463_));
  AOI21X1  g2078(.A0(new_n2463_), .A1(new_n1390_), .B0(new_n1391_), .Y(new_n2464_));
  OAI21X1  g2079(.A0(new_n2464_), .A1(new_n1389_), .B0(new_n433_), .Y(new_n2465_));
  OAI21X1  g2080(.A0(new_n755_), .A1(\priority[23] ), .B0(\req[23] ), .Y(new_n2466_));
  AOI21X1  g2081(.A0(new_n2465_), .A1(new_n1387_), .B0(new_n2466_), .Y(\grant[23] ));
  NOR2X1   g2082(.A(new_n763_), .B(new_n447_), .Y(new_n2468_));
  OAI21X1  g2083(.A0(new_n2468_), .A1(new_n454_), .B0(new_n456_), .Y(new_n2469_));
  AOI21X1  g2084(.A0(new_n2469_), .A1(new_n461_), .B0(new_n464_), .Y(new_n2470_));
  OAI21X1  g2085(.A0(new_n2470_), .A1(new_n469_), .B0(new_n471_), .Y(new_n2471_));
  AOI21X1  g2086(.A0(new_n2471_), .A1(new_n476_), .B0(new_n479_), .Y(new_n2472_));
  OAI21X1  g2087(.A0(new_n2472_), .A1(new_n484_), .B0(new_n486_), .Y(new_n2473_));
  AOI21X1  g2088(.A0(new_n2473_), .A1(new_n491_), .B0(new_n494_), .Y(new_n2474_));
  OAI21X1  g2089(.A0(new_n2474_), .A1(new_n499_), .B0(new_n501_), .Y(new_n2475_));
  AOI21X1  g2090(.A0(new_n2475_), .A1(new_n506_), .B0(new_n509_), .Y(new_n2476_));
  OAI21X1  g2091(.A0(new_n2476_), .A1(new_n514_), .B0(new_n516_), .Y(new_n2477_));
  AOI21X1  g2092(.A0(new_n2477_), .A1(new_n521_), .B0(new_n524_), .Y(new_n2478_));
  OAI21X1  g2093(.A0(new_n2478_), .A1(new_n529_), .B0(new_n531_), .Y(new_n2479_));
  AOI21X1  g2094(.A0(new_n2479_), .A1(new_n536_), .B0(new_n539_), .Y(new_n2480_));
  OAI21X1  g2095(.A0(new_n2480_), .A1(new_n544_), .B0(new_n546_), .Y(new_n2481_));
  AOI21X1  g2096(.A0(new_n2481_), .A1(new_n551_), .B0(new_n554_), .Y(new_n2482_));
  OAI21X1  g2097(.A0(new_n2482_), .A1(new_n559_), .B0(new_n561_), .Y(new_n2483_));
  AOI21X1  g2098(.A0(new_n2483_), .A1(new_n566_), .B0(new_n569_), .Y(new_n2484_));
  OAI21X1  g2099(.A0(new_n2484_), .A1(new_n574_), .B0(new_n576_), .Y(new_n2485_));
  AOI21X1  g2100(.A0(new_n2485_), .A1(new_n581_), .B0(new_n584_), .Y(new_n2486_));
  OAI21X1  g2101(.A0(new_n2486_), .A1(new_n589_), .B0(new_n591_), .Y(new_n2487_));
  AOI21X1  g2102(.A0(new_n2487_), .A1(new_n596_), .B0(new_n599_), .Y(new_n2488_));
  OAI21X1  g2103(.A0(new_n2488_), .A1(new_n604_), .B0(new_n606_), .Y(new_n2489_));
  AOI21X1  g2104(.A0(new_n2489_), .A1(new_n611_), .B0(new_n614_), .Y(new_n2490_));
  OAI21X1  g2105(.A0(new_n2490_), .A1(new_n619_), .B0(new_n621_), .Y(new_n2491_));
  AOI21X1  g2106(.A0(new_n2491_), .A1(new_n626_), .B0(new_n629_), .Y(new_n2492_));
  OAI21X1  g2107(.A0(new_n2492_), .A1(new_n634_), .B0(new_n636_), .Y(new_n2493_));
  AOI21X1  g2108(.A0(new_n2493_), .A1(new_n641_), .B0(new_n644_), .Y(new_n2494_));
  OAI21X1  g2109(.A0(new_n2494_), .A1(new_n649_), .B0(new_n651_), .Y(new_n2495_));
  AOI21X1  g2110(.A0(new_n2495_), .A1(new_n656_), .B0(new_n659_), .Y(new_n2496_));
  OAI21X1  g2111(.A0(new_n2496_), .A1(new_n664_), .B0(new_n666_), .Y(new_n2497_));
  AOI21X1  g2112(.A0(new_n2497_), .A1(new_n671_), .B0(new_n674_), .Y(new_n2498_));
  OAI21X1  g2113(.A0(new_n2498_), .A1(new_n679_), .B0(new_n681_), .Y(new_n2499_));
  AOI21X1  g2114(.A0(new_n2499_), .A1(new_n686_), .B0(new_n689_), .Y(new_n2500_));
  OAI21X1  g2115(.A0(new_n2500_), .A1(new_n694_), .B0(new_n696_), .Y(new_n2501_));
  AOI21X1  g2116(.A0(new_n2501_), .A1(new_n701_), .B0(new_n1662_), .Y(new_n2502_));
  OAI21X1  g2117(.A0(new_n2502_), .A1(new_n1661_), .B0(new_n1705_), .Y(new_n2503_));
  AOI21X1  g2118(.A0(new_n2503_), .A1(new_n1660_), .B0(new_n1938_), .Y(new_n2504_));
  OAI21X1  g2119(.A0(new_n2504_), .A1(new_n1504_), .B0(new_n721_), .Y(new_n2505_));
  AOI21X1  g2120(.A0(new_n2505_), .A1(new_n1502_), .B0(new_n1503_), .Y(new_n2506_));
  OAI21X1  g2121(.A0(new_n2506_), .A1(new_n1501_), .B0(new_n736_), .Y(new_n2507_));
  AOI21X1  g2122(.A0(new_n2507_), .A1(new_n1499_), .B0(new_n1500_), .Y(new_n2508_));
  OAI21X1  g2123(.A0(new_n2508_), .A1(new_n1498_), .B0(new_n751_), .Y(new_n2509_));
  OAI21X1  g2124(.A0(new_n1069_), .A1(\priority[24] ), .B0(\req[24] ), .Y(new_n2510_));
  AOI21X1  g2125(.A0(new_n2509_), .A1(new_n1496_), .B0(new_n2510_), .Y(\grant[24] ));
  NOR2X1   g2126(.A(new_n1077_), .B(new_n765_), .Y(new_n2512_));
  OAI21X1  g2127(.A0(new_n2512_), .A1(new_n772_), .B0(new_n774_), .Y(new_n2513_));
  AOI21X1  g2128(.A0(new_n2513_), .A1(new_n779_), .B0(new_n782_), .Y(new_n2514_));
  OAI21X1  g2129(.A0(new_n2514_), .A1(new_n787_), .B0(new_n789_), .Y(new_n2515_));
  AOI21X1  g2130(.A0(new_n2515_), .A1(new_n794_), .B0(new_n797_), .Y(new_n2516_));
  OAI21X1  g2131(.A0(new_n2516_), .A1(new_n802_), .B0(new_n804_), .Y(new_n2517_));
  AOI21X1  g2132(.A0(new_n2517_), .A1(new_n809_), .B0(new_n812_), .Y(new_n2518_));
  OAI21X1  g2133(.A0(new_n2518_), .A1(new_n817_), .B0(new_n819_), .Y(new_n2519_));
  AOI21X1  g2134(.A0(new_n2519_), .A1(new_n824_), .B0(new_n827_), .Y(new_n2520_));
  OAI21X1  g2135(.A0(new_n2520_), .A1(new_n832_), .B0(new_n834_), .Y(new_n2521_));
  AOI21X1  g2136(.A0(new_n2521_), .A1(new_n839_), .B0(new_n842_), .Y(new_n2522_));
  OAI21X1  g2137(.A0(new_n2522_), .A1(new_n847_), .B0(new_n849_), .Y(new_n2523_));
  AOI21X1  g2138(.A0(new_n2523_), .A1(new_n854_), .B0(new_n857_), .Y(new_n2524_));
  OAI21X1  g2139(.A0(new_n2524_), .A1(new_n862_), .B0(new_n864_), .Y(new_n2525_));
  AOI21X1  g2140(.A0(new_n2525_), .A1(new_n869_), .B0(new_n872_), .Y(new_n2526_));
  OAI21X1  g2141(.A0(new_n2526_), .A1(new_n877_), .B0(new_n879_), .Y(new_n2527_));
  AOI21X1  g2142(.A0(new_n2527_), .A1(new_n884_), .B0(new_n887_), .Y(new_n2528_));
  OAI21X1  g2143(.A0(new_n2528_), .A1(new_n892_), .B0(new_n894_), .Y(new_n2529_));
  AOI21X1  g2144(.A0(new_n2529_), .A1(new_n899_), .B0(new_n902_), .Y(new_n2530_));
  OAI21X1  g2145(.A0(new_n2530_), .A1(new_n907_), .B0(new_n909_), .Y(new_n2531_));
  AOI21X1  g2146(.A0(new_n2531_), .A1(new_n914_), .B0(new_n917_), .Y(new_n2532_));
  OAI21X1  g2147(.A0(new_n2532_), .A1(new_n922_), .B0(new_n924_), .Y(new_n2533_));
  AOI21X1  g2148(.A0(new_n2533_), .A1(new_n929_), .B0(new_n932_), .Y(new_n2534_));
  OAI21X1  g2149(.A0(new_n2534_), .A1(new_n937_), .B0(new_n939_), .Y(new_n2535_));
  AOI21X1  g2150(.A0(new_n2535_), .A1(new_n944_), .B0(new_n947_), .Y(new_n2536_));
  OAI21X1  g2151(.A0(new_n2536_), .A1(new_n952_), .B0(new_n954_), .Y(new_n2537_));
  AOI21X1  g2152(.A0(new_n2537_), .A1(new_n959_), .B0(new_n962_), .Y(new_n2538_));
  OAI21X1  g2153(.A0(new_n2538_), .A1(new_n967_), .B0(new_n969_), .Y(new_n2539_));
  AOI21X1  g2154(.A0(new_n2539_), .A1(new_n974_), .B0(new_n977_), .Y(new_n2540_));
  OAI21X1  g2155(.A0(new_n2540_), .A1(new_n982_), .B0(new_n984_), .Y(new_n2541_));
  AOI21X1  g2156(.A0(new_n2541_), .A1(new_n989_), .B0(new_n992_), .Y(new_n2542_));
  OAI21X1  g2157(.A0(new_n2542_), .A1(new_n997_), .B0(new_n999_), .Y(new_n2543_));
  AOI21X1  g2158(.A0(new_n2543_), .A1(new_n1004_), .B0(new_n1007_), .Y(new_n2544_));
  OAI21X1  g2159(.A0(new_n2544_), .A1(new_n1012_), .B0(new_n1014_), .Y(new_n2545_));
  AOI21X1  g2160(.A0(new_n2545_), .A1(new_n1017_), .B0(new_n1711_), .Y(new_n2546_));
  OAI21X1  g2161(.A0(new_n2546_), .A1(new_n1710_), .B0(new_n1754_), .Y(new_n2547_));
  AOI21X1  g2162(.A0(new_n2547_), .A1(new_n1709_), .B0(new_n1983_), .Y(new_n2548_));
  OAI21X1  g2163(.A0(new_n2548_), .A1(new_n1613_), .B0(new_n1035_), .Y(new_n2549_));
  AOI21X1  g2164(.A0(new_n2549_), .A1(new_n1611_), .B0(new_n1612_), .Y(new_n2550_));
  OAI21X1  g2165(.A0(new_n2550_), .A1(new_n1610_), .B0(new_n1050_), .Y(new_n2551_));
  AOI21X1  g2166(.A0(new_n2551_), .A1(new_n1608_), .B0(new_n1609_), .Y(new_n2552_));
  OAI21X1  g2167(.A0(new_n2552_), .A1(new_n1607_), .B0(new_n1065_), .Y(new_n2553_));
  OAI21X1  g2168(.A0(new_n444_), .A1(\priority[25] ), .B0(\req[25] ), .Y(new_n2554_));
  AOI21X1  g2169(.A0(new_n2553_), .A1(new_n1605_), .B0(new_n2554_), .Y(\grant[25] ));
  NOR2X1   g2170(.A(new_n1079_), .B(new_n453_), .Y(new_n2556_));
  OAI21X1  g2171(.A0(new_n2556_), .A1(new_n1086_), .B0(new_n1088_), .Y(new_n2557_));
  AOI21X1  g2172(.A0(new_n2557_), .A1(new_n1093_), .B0(new_n1096_), .Y(new_n2558_));
  OAI21X1  g2173(.A0(new_n2558_), .A1(new_n1101_), .B0(new_n1103_), .Y(new_n2559_));
  AOI21X1  g2174(.A0(new_n2559_), .A1(new_n1108_), .B0(new_n1111_), .Y(new_n2560_));
  OAI21X1  g2175(.A0(new_n2560_), .A1(new_n1116_), .B0(new_n1118_), .Y(new_n2561_));
  AOI21X1  g2176(.A0(new_n2561_), .A1(new_n1123_), .B0(new_n1126_), .Y(new_n2562_));
  OAI21X1  g2177(.A0(new_n2562_), .A1(new_n1131_), .B0(new_n1133_), .Y(new_n2563_));
  AOI21X1  g2178(.A0(new_n2563_), .A1(new_n1138_), .B0(new_n1141_), .Y(new_n2564_));
  OAI21X1  g2179(.A0(new_n2564_), .A1(new_n1146_), .B0(new_n1148_), .Y(new_n2565_));
  AOI21X1  g2180(.A0(new_n2565_), .A1(new_n1153_), .B0(new_n1156_), .Y(new_n2566_));
  OAI21X1  g2181(.A0(new_n2566_), .A1(new_n1161_), .B0(new_n1163_), .Y(new_n2567_));
  AOI21X1  g2182(.A0(new_n2567_), .A1(new_n1168_), .B0(new_n1171_), .Y(new_n2568_));
  OAI21X1  g2183(.A0(new_n2568_), .A1(new_n1176_), .B0(new_n1178_), .Y(new_n2569_));
  AOI21X1  g2184(.A0(new_n2569_), .A1(new_n1183_), .B0(new_n1186_), .Y(new_n2570_));
  OAI21X1  g2185(.A0(new_n2570_), .A1(new_n1191_), .B0(new_n1193_), .Y(new_n2571_));
  AOI21X1  g2186(.A0(new_n2571_), .A1(new_n1198_), .B0(new_n1201_), .Y(new_n2572_));
  OAI21X1  g2187(.A0(new_n2572_), .A1(new_n1206_), .B0(new_n1208_), .Y(new_n2573_));
  AOI21X1  g2188(.A0(new_n2573_), .A1(new_n1213_), .B0(new_n1216_), .Y(new_n2574_));
  OAI21X1  g2189(.A0(new_n2574_), .A1(new_n1221_), .B0(new_n1223_), .Y(new_n2575_));
  AOI21X1  g2190(.A0(new_n2575_), .A1(new_n1228_), .B0(new_n1231_), .Y(new_n2576_));
  OAI21X1  g2191(.A0(new_n2576_), .A1(new_n1236_), .B0(new_n1238_), .Y(new_n2577_));
  AOI21X1  g2192(.A0(new_n2577_), .A1(new_n1243_), .B0(new_n1246_), .Y(new_n2578_));
  OAI21X1  g2193(.A0(new_n2578_), .A1(new_n1251_), .B0(new_n1253_), .Y(new_n2579_));
  AOI21X1  g2194(.A0(new_n2579_), .A1(new_n1258_), .B0(new_n1261_), .Y(new_n2580_));
  OAI21X1  g2195(.A0(new_n2580_), .A1(new_n1266_), .B0(new_n1268_), .Y(new_n2581_));
  AOI21X1  g2196(.A0(new_n2581_), .A1(new_n1273_), .B0(new_n1276_), .Y(new_n2582_));
  OAI21X1  g2197(.A0(new_n2582_), .A1(new_n1281_), .B0(new_n1283_), .Y(new_n2583_));
  AOI21X1  g2198(.A0(new_n2583_), .A1(new_n1288_), .B0(new_n1291_), .Y(new_n2584_));
  OAI21X1  g2199(.A0(new_n2584_), .A1(new_n1296_), .B0(new_n1298_), .Y(new_n2585_));
  AOI21X1  g2200(.A0(new_n2585_), .A1(new_n1303_), .B0(new_n1306_), .Y(new_n2586_));
  OAI21X1  g2201(.A0(new_n2586_), .A1(new_n1311_), .B0(new_n1313_), .Y(new_n2587_));
  AOI21X1  g2202(.A0(new_n2587_), .A1(new_n1318_), .B0(new_n1321_), .Y(new_n2588_));
  OAI21X1  g2203(.A0(new_n2588_), .A1(new_n1326_), .B0(new_n1328_), .Y(new_n2589_));
  AOI21X1  g2204(.A0(new_n2589_), .A1(new_n1331_), .B0(new_n1758_), .Y(new_n2590_));
  OAI21X1  g2205(.A0(new_n2590_), .A1(new_n394_), .B0(new_n396_), .Y(new_n2591_));
  AOI21X1  g2206(.A0(new_n2591_), .A1(new_n401_), .B0(new_n404_), .Y(new_n2592_));
  OAI21X1  g2207(.A0(new_n2592_), .A1(new_n409_), .B0(new_n411_), .Y(new_n2593_));
  AOI21X1  g2208(.A0(new_n2593_), .A1(new_n416_), .B0(new_n419_), .Y(new_n2594_));
  OAI21X1  g2209(.A0(new_n2594_), .A1(new_n424_), .B0(new_n426_), .Y(new_n2595_));
  AOI21X1  g2210(.A0(new_n2595_), .A1(new_n431_), .B0(new_n434_), .Y(new_n2596_));
  OAI21X1  g2211(.A0(new_n2596_), .A1(new_n439_), .B0(new_n441_), .Y(new_n2597_));
  OAI21X1  g2212(.A0(new_n762_), .A1(\priority[26] ), .B0(\req[26] ), .Y(new_n2598_));
  AOI21X1  g2213(.A0(new_n2597_), .A1(new_n446_), .B0(new_n2598_), .Y(\grant[26] ));
  NOR2X1   g2214(.A(new_n771_), .B(new_n455_), .Y(new_n2600_));
  OAI21X1  g2215(.A0(new_n2600_), .A1(new_n1383_), .B0(new_n463_), .Y(new_n2601_));
  AOI21X1  g2216(.A0(new_n2601_), .A1(new_n1381_), .B0(new_n1382_), .Y(new_n2602_));
  OAI21X1  g2217(.A0(new_n2602_), .A1(new_n1380_), .B0(new_n478_), .Y(new_n2603_));
  AOI21X1  g2218(.A0(new_n2603_), .A1(new_n1378_), .B0(new_n1379_), .Y(new_n2604_));
  OAI21X1  g2219(.A0(new_n2604_), .A1(new_n1377_), .B0(new_n493_), .Y(new_n2605_));
  AOI21X1  g2220(.A0(new_n2605_), .A1(new_n1375_), .B0(new_n1376_), .Y(new_n2606_));
  OAI21X1  g2221(.A0(new_n2606_), .A1(new_n1374_), .B0(new_n508_), .Y(new_n2607_));
  AOI21X1  g2222(.A0(new_n2607_), .A1(new_n1372_), .B0(new_n1373_), .Y(new_n2608_));
  OAI21X1  g2223(.A0(new_n2608_), .A1(new_n1371_), .B0(new_n523_), .Y(new_n2609_));
  AOI21X1  g2224(.A0(new_n2609_), .A1(new_n1369_), .B0(new_n1370_), .Y(new_n2610_));
  OAI21X1  g2225(.A0(new_n2610_), .A1(new_n1368_), .B0(new_n538_), .Y(new_n2611_));
  AOI21X1  g2226(.A0(new_n2611_), .A1(new_n1366_), .B0(new_n1367_), .Y(new_n2612_));
  OAI21X1  g2227(.A0(new_n2612_), .A1(new_n1365_), .B0(new_n553_), .Y(new_n2613_));
  AOI21X1  g2228(.A0(new_n2613_), .A1(new_n1363_), .B0(new_n1364_), .Y(new_n2614_));
  OAI21X1  g2229(.A0(new_n2614_), .A1(new_n1362_), .B0(new_n568_), .Y(new_n2615_));
  AOI21X1  g2230(.A0(new_n2615_), .A1(new_n1360_), .B0(new_n1361_), .Y(new_n2616_));
  OAI21X1  g2231(.A0(new_n2616_), .A1(new_n1359_), .B0(new_n583_), .Y(new_n2617_));
  AOI21X1  g2232(.A0(new_n2617_), .A1(new_n1357_), .B0(new_n1358_), .Y(new_n2618_));
  OAI21X1  g2233(.A0(new_n2618_), .A1(new_n1356_), .B0(new_n598_), .Y(new_n2619_));
  AOI21X1  g2234(.A0(new_n2619_), .A1(new_n1354_), .B0(new_n1355_), .Y(new_n2620_));
  OAI21X1  g2235(.A0(new_n2620_), .A1(new_n1353_), .B0(new_n613_), .Y(new_n2621_));
  AOI21X1  g2236(.A0(new_n2621_), .A1(new_n1351_), .B0(new_n1352_), .Y(new_n2622_));
  OAI21X1  g2237(.A0(new_n2622_), .A1(new_n1350_), .B0(new_n628_), .Y(new_n2623_));
  AOI21X1  g2238(.A0(new_n2623_), .A1(new_n1348_), .B0(new_n1349_), .Y(new_n2624_));
  OAI21X1  g2239(.A0(new_n2624_), .A1(new_n1347_), .B0(new_n643_), .Y(new_n2625_));
  AOI21X1  g2240(.A0(new_n2625_), .A1(new_n1345_), .B0(new_n1346_), .Y(new_n2626_));
  OAI21X1  g2241(.A0(new_n2626_), .A1(new_n1344_), .B0(new_n658_), .Y(new_n2627_));
  AOI21X1  g2242(.A0(new_n2627_), .A1(new_n1342_), .B0(new_n1343_), .Y(new_n2628_));
  OAI21X1  g2243(.A0(new_n2628_), .A1(new_n1341_), .B0(new_n673_), .Y(new_n2629_));
  AOI21X1  g2244(.A0(new_n2629_), .A1(new_n1339_), .B0(new_n1340_), .Y(new_n2630_));
  OAI21X1  g2245(.A0(new_n2630_), .A1(new_n1338_), .B0(new_n688_), .Y(new_n2631_));
  AOI21X1  g2246(.A0(new_n2631_), .A1(new_n1336_), .B0(new_n1337_), .Y(new_n2632_));
  OAI21X1  g2247(.A0(new_n2632_), .A1(new_n1335_), .B0(new_n1438_), .Y(new_n2633_));
  AOI21X1  g2248(.A0(new_n2633_), .A1(new_n1440_), .B0(new_n1803_), .Y(new_n2634_));
  OAI21X1  g2249(.A0(new_n2634_), .A1(new_n712_), .B0(new_n714_), .Y(new_n2635_));
  AOI21X1  g2250(.A0(new_n2635_), .A1(new_n719_), .B0(new_n722_), .Y(new_n2636_));
  OAI21X1  g2251(.A0(new_n2636_), .A1(new_n727_), .B0(new_n729_), .Y(new_n2637_));
  AOI21X1  g2252(.A0(new_n2637_), .A1(new_n734_), .B0(new_n737_), .Y(new_n2638_));
  OAI21X1  g2253(.A0(new_n2638_), .A1(new_n742_), .B0(new_n744_), .Y(new_n2639_));
  AOI21X1  g2254(.A0(new_n2639_), .A1(new_n749_), .B0(new_n752_), .Y(new_n2640_));
  OAI21X1  g2255(.A0(new_n2640_), .A1(new_n757_), .B0(new_n759_), .Y(new_n2641_));
  OAI21X1  g2256(.A0(new_n1076_), .A1(\priority[27] ), .B0(\req[27] ), .Y(new_n2642_));
  AOI21X1  g2257(.A0(new_n2641_), .A1(new_n764_), .B0(new_n2642_), .Y(\grant[27] ));
  NOR2X1   g2258(.A(new_n1085_), .B(new_n773_), .Y(new_n2644_));
  OAI21X1  g2259(.A0(new_n2644_), .A1(new_n1492_), .B0(new_n781_), .Y(new_n2645_));
  AOI21X1  g2260(.A0(new_n2645_), .A1(new_n1490_), .B0(new_n1491_), .Y(new_n2646_));
  OAI21X1  g2261(.A0(new_n2646_), .A1(new_n1489_), .B0(new_n796_), .Y(new_n2647_));
  AOI21X1  g2262(.A0(new_n2647_), .A1(new_n1487_), .B0(new_n1488_), .Y(new_n2648_));
  OAI21X1  g2263(.A0(new_n2648_), .A1(new_n1486_), .B0(new_n811_), .Y(new_n2649_));
  AOI21X1  g2264(.A0(new_n2649_), .A1(new_n1484_), .B0(new_n1485_), .Y(new_n2650_));
  OAI21X1  g2265(.A0(new_n2650_), .A1(new_n1483_), .B0(new_n826_), .Y(new_n2651_));
  AOI21X1  g2266(.A0(new_n2651_), .A1(new_n1481_), .B0(new_n1482_), .Y(new_n2652_));
  OAI21X1  g2267(.A0(new_n2652_), .A1(new_n1480_), .B0(new_n841_), .Y(new_n2653_));
  AOI21X1  g2268(.A0(new_n2653_), .A1(new_n1478_), .B0(new_n1479_), .Y(new_n2654_));
  OAI21X1  g2269(.A0(new_n2654_), .A1(new_n1477_), .B0(new_n856_), .Y(new_n2655_));
  AOI21X1  g2270(.A0(new_n2655_), .A1(new_n1475_), .B0(new_n1476_), .Y(new_n2656_));
  OAI21X1  g2271(.A0(new_n2656_), .A1(new_n1474_), .B0(new_n871_), .Y(new_n2657_));
  AOI21X1  g2272(.A0(new_n2657_), .A1(new_n1472_), .B0(new_n1473_), .Y(new_n2658_));
  OAI21X1  g2273(.A0(new_n2658_), .A1(new_n1471_), .B0(new_n886_), .Y(new_n2659_));
  AOI21X1  g2274(.A0(new_n2659_), .A1(new_n1469_), .B0(new_n1470_), .Y(new_n2660_));
  OAI21X1  g2275(.A0(new_n2660_), .A1(new_n1468_), .B0(new_n901_), .Y(new_n2661_));
  AOI21X1  g2276(.A0(new_n2661_), .A1(new_n1466_), .B0(new_n1467_), .Y(new_n2662_));
  OAI21X1  g2277(.A0(new_n2662_), .A1(new_n1465_), .B0(new_n916_), .Y(new_n2663_));
  AOI21X1  g2278(.A0(new_n2663_), .A1(new_n1463_), .B0(new_n1464_), .Y(new_n2664_));
  OAI21X1  g2279(.A0(new_n2664_), .A1(new_n1462_), .B0(new_n931_), .Y(new_n2665_));
  AOI21X1  g2280(.A0(new_n2665_), .A1(new_n1460_), .B0(new_n1461_), .Y(new_n2666_));
  OAI21X1  g2281(.A0(new_n2666_), .A1(new_n1459_), .B0(new_n946_), .Y(new_n2667_));
  AOI21X1  g2282(.A0(new_n2667_), .A1(new_n1457_), .B0(new_n1458_), .Y(new_n2668_));
  OAI21X1  g2283(.A0(new_n2668_), .A1(new_n1456_), .B0(new_n961_), .Y(new_n2669_));
  AOI21X1  g2284(.A0(new_n2669_), .A1(new_n1454_), .B0(new_n1455_), .Y(new_n2670_));
  OAI21X1  g2285(.A0(new_n2670_), .A1(new_n1453_), .B0(new_n976_), .Y(new_n2671_));
  AOI21X1  g2286(.A0(new_n2671_), .A1(new_n1451_), .B0(new_n1452_), .Y(new_n2672_));
  OAI21X1  g2287(.A0(new_n2672_), .A1(new_n1450_), .B0(new_n991_), .Y(new_n2673_));
  AOI21X1  g2288(.A0(new_n2673_), .A1(new_n1448_), .B0(new_n1449_), .Y(new_n2674_));
  OAI21X1  g2289(.A0(new_n2674_), .A1(new_n1447_), .B0(new_n1006_), .Y(new_n2675_));
  AOI21X1  g2290(.A0(new_n2675_), .A1(new_n1445_), .B0(new_n1446_), .Y(new_n2676_));
  OAI21X1  g2291(.A0(new_n2676_), .A1(new_n1444_), .B0(new_n1547_), .Y(new_n2677_));
  AOI21X1  g2292(.A0(new_n2677_), .A1(new_n1549_), .B0(new_n1848_), .Y(new_n2678_));
  OAI21X1  g2293(.A0(new_n2678_), .A1(new_n1026_), .B0(new_n1028_), .Y(new_n2679_));
  AOI21X1  g2294(.A0(new_n2679_), .A1(new_n1033_), .B0(new_n1036_), .Y(new_n2680_));
  OAI21X1  g2295(.A0(new_n2680_), .A1(new_n1041_), .B0(new_n1043_), .Y(new_n2681_));
  AOI21X1  g2296(.A0(new_n2681_), .A1(new_n1048_), .B0(new_n1051_), .Y(new_n2682_));
  OAI21X1  g2297(.A0(new_n2682_), .A1(new_n1056_), .B0(new_n1058_), .Y(new_n2683_));
  AOI21X1  g2298(.A0(new_n2683_), .A1(new_n1063_), .B0(new_n1066_), .Y(new_n2684_));
  OAI21X1  g2299(.A0(new_n2684_), .A1(new_n1071_), .B0(new_n1073_), .Y(new_n2685_));
  OAI21X1  g2300(.A0(new_n452_), .A1(\priority[28] ), .B0(\req[28] ), .Y(new_n2686_));
  AOI21X1  g2301(.A0(new_n2685_), .A1(new_n1078_), .B0(new_n2686_), .Y(\grant[28] ));
  NOR2X1   g2302(.A(new_n1087_), .B(new_n460_), .Y(new_n2688_));
  OAI21X1  g2303(.A0(new_n2688_), .A1(new_n1601_), .B0(new_n1095_), .Y(new_n2689_));
  AOI21X1  g2304(.A0(new_n2689_), .A1(new_n1599_), .B0(new_n1600_), .Y(new_n2690_));
  OAI21X1  g2305(.A0(new_n2690_), .A1(new_n1598_), .B0(new_n1110_), .Y(new_n2691_));
  AOI21X1  g2306(.A0(new_n2691_), .A1(new_n1596_), .B0(new_n1597_), .Y(new_n2692_));
  OAI21X1  g2307(.A0(new_n2692_), .A1(new_n1595_), .B0(new_n1125_), .Y(new_n2693_));
  AOI21X1  g2308(.A0(new_n2693_), .A1(new_n1593_), .B0(new_n1594_), .Y(new_n2694_));
  OAI21X1  g2309(.A0(new_n2694_), .A1(new_n1592_), .B0(new_n1140_), .Y(new_n2695_));
  AOI21X1  g2310(.A0(new_n2695_), .A1(new_n1590_), .B0(new_n1591_), .Y(new_n2696_));
  OAI21X1  g2311(.A0(new_n2696_), .A1(new_n1589_), .B0(new_n1155_), .Y(new_n2697_));
  AOI21X1  g2312(.A0(new_n2697_), .A1(new_n1587_), .B0(new_n1588_), .Y(new_n2698_));
  OAI21X1  g2313(.A0(new_n2698_), .A1(new_n1586_), .B0(new_n1170_), .Y(new_n2699_));
  AOI21X1  g2314(.A0(new_n2699_), .A1(new_n1584_), .B0(new_n1585_), .Y(new_n2700_));
  OAI21X1  g2315(.A0(new_n2700_), .A1(new_n1583_), .B0(new_n1185_), .Y(new_n2701_));
  AOI21X1  g2316(.A0(new_n2701_), .A1(new_n1581_), .B0(new_n1582_), .Y(new_n2702_));
  OAI21X1  g2317(.A0(new_n2702_), .A1(new_n1580_), .B0(new_n1200_), .Y(new_n2703_));
  AOI21X1  g2318(.A0(new_n2703_), .A1(new_n1578_), .B0(new_n1579_), .Y(new_n2704_));
  OAI21X1  g2319(.A0(new_n2704_), .A1(new_n1577_), .B0(new_n1215_), .Y(new_n2705_));
  AOI21X1  g2320(.A0(new_n2705_), .A1(new_n1575_), .B0(new_n1576_), .Y(new_n2706_));
  OAI21X1  g2321(.A0(new_n2706_), .A1(new_n1574_), .B0(new_n1230_), .Y(new_n2707_));
  AOI21X1  g2322(.A0(new_n2707_), .A1(new_n1572_), .B0(new_n1573_), .Y(new_n2708_));
  OAI21X1  g2323(.A0(new_n2708_), .A1(new_n1571_), .B0(new_n1245_), .Y(new_n2709_));
  AOI21X1  g2324(.A0(new_n2709_), .A1(new_n1569_), .B0(new_n1570_), .Y(new_n2710_));
  OAI21X1  g2325(.A0(new_n2710_), .A1(new_n1568_), .B0(new_n1260_), .Y(new_n2711_));
  AOI21X1  g2326(.A0(new_n2711_), .A1(new_n1566_), .B0(new_n1567_), .Y(new_n2712_));
  OAI21X1  g2327(.A0(new_n2712_), .A1(new_n1565_), .B0(new_n1275_), .Y(new_n2713_));
  AOI21X1  g2328(.A0(new_n2713_), .A1(new_n1563_), .B0(new_n1564_), .Y(new_n2714_));
  OAI21X1  g2329(.A0(new_n2714_), .A1(new_n1562_), .B0(new_n1290_), .Y(new_n2715_));
  AOI21X1  g2330(.A0(new_n2715_), .A1(new_n1560_), .B0(new_n1561_), .Y(new_n2716_));
  OAI21X1  g2331(.A0(new_n2716_), .A1(new_n1559_), .B0(new_n1305_), .Y(new_n2717_));
  AOI21X1  g2332(.A0(new_n2717_), .A1(new_n1557_), .B0(new_n1558_), .Y(new_n2718_));
  OAI21X1  g2333(.A0(new_n2718_), .A1(new_n1556_), .B0(new_n1320_), .Y(new_n2719_));
  AOI21X1  g2334(.A0(new_n2719_), .A1(new_n1554_), .B0(new_n1555_), .Y(new_n2720_));
  OAI21X1  g2335(.A0(new_n2720_), .A1(new_n1553_), .B0(new_n1656_), .Y(new_n2721_));
  AOI21X1  g2336(.A0(new_n2721_), .A1(new_n1552_), .B0(new_n1893_), .Y(new_n2722_));
  OAI21X1  g2337(.A0(new_n2722_), .A1(new_n1395_), .B0(new_n403_), .Y(new_n2723_));
  AOI21X1  g2338(.A0(new_n2723_), .A1(new_n1393_), .B0(new_n1394_), .Y(new_n2724_));
  OAI21X1  g2339(.A0(new_n2724_), .A1(new_n1392_), .B0(new_n418_), .Y(new_n2725_));
  AOI21X1  g2340(.A0(new_n2725_), .A1(new_n1390_), .B0(new_n1391_), .Y(new_n2726_));
  OAI21X1  g2341(.A0(new_n2726_), .A1(new_n1389_), .B0(new_n433_), .Y(new_n2727_));
  AOI21X1  g2342(.A0(new_n2727_), .A1(new_n1387_), .B0(new_n1388_), .Y(new_n2728_));
  OAI21X1  g2343(.A0(new_n2728_), .A1(new_n1386_), .B0(new_n448_), .Y(new_n2729_));
  OAI21X1  g2344(.A0(new_n770_), .A1(\priority[29] ), .B0(\req[29] ), .Y(new_n2730_));
  AOI21X1  g2345(.A0(new_n2729_), .A1(new_n1384_), .B0(new_n2730_), .Y(\grant[29] ));
  NOR2X1   g2346(.A(new_n778_), .B(new_n462_), .Y(new_n2732_));
  OAI21X1  g2347(.A0(new_n2732_), .A1(new_n469_), .B0(new_n471_), .Y(new_n2733_));
  AOI21X1  g2348(.A0(new_n2733_), .A1(new_n476_), .B0(new_n479_), .Y(new_n2734_));
  OAI21X1  g2349(.A0(new_n2734_), .A1(new_n484_), .B0(new_n486_), .Y(new_n2735_));
  AOI21X1  g2350(.A0(new_n2735_), .A1(new_n491_), .B0(new_n494_), .Y(new_n2736_));
  OAI21X1  g2351(.A0(new_n2736_), .A1(new_n499_), .B0(new_n501_), .Y(new_n2737_));
  AOI21X1  g2352(.A0(new_n2737_), .A1(new_n506_), .B0(new_n509_), .Y(new_n2738_));
  OAI21X1  g2353(.A0(new_n2738_), .A1(new_n514_), .B0(new_n516_), .Y(new_n2739_));
  AOI21X1  g2354(.A0(new_n2739_), .A1(new_n521_), .B0(new_n524_), .Y(new_n2740_));
  OAI21X1  g2355(.A0(new_n2740_), .A1(new_n529_), .B0(new_n531_), .Y(new_n2741_));
  AOI21X1  g2356(.A0(new_n2741_), .A1(new_n536_), .B0(new_n539_), .Y(new_n2742_));
  OAI21X1  g2357(.A0(new_n2742_), .A1(new_n544_), .B0(new_n546_), .Y(new_n2743_));
  AOI21X1  g2358(.A0(new_n2743_), .A1(new_n551_), .B0(new_n554_), .Y(new_n2744_));
  OAI21X1  g2359(.A0(new_n2744_), .A1(new_n559_), .B0(new_n561_), .Y(new_n2745_));
  AOI21X1  g2360(.A0(new_n2745_), .A1(new_n566_), .B0(new_n569_), .Y(new_n2746_));
  OAI21X1  g2361(.A0(new_n2746_), .A1(new_n574_), .B0(new_n576_), .Y(new_n2747_));
  AOI21X1  g2362(.A0(new_n2747_), .A1(new_n581_), .B0(new_n584_), .Y(new_n2748_));
  OAI21X1  g2363(.A0(new_n2748_), .A1(new_n589_), .B0(new_n591_), .Y(new_n2749_));
  AOI21X1  g2364(.A0(new_n2749_), .A1(new_n596_), .B0(new_n599_), .Y(new_n2750_));
  OAI21X1  g2365(.A0(new_n2750_), .A1(new_n604_), .B0(new_n606_), .Y(new_n2751_));
  AOI21X1  g2366(.A0(new_n2751_), .A1(new_n611_), .B0(new_n614_), .Y(new_n2752_));
  OAI21X1  g2367(.A0(new_n2752_), .A1(new_n619_), .B0(new_n621_), .Y(new_n2753_));
  AOI21X1  g2368(.A0(new_n2753_), .A1(new_n626_), .B0(new_n629_), .Y(new_n2754_));
  OAI21X1  g2369(.A0(new_n2754_), .A1(new_n634_), .B0(new_n636_), .Y(new_n2755_));
  AOI21X1  g2370(.A0(new_n2755_), .A1(new_n641_), .B0(new_n644_), .Y(new_n2756_));
  OAI21X1  g2371(.A0(new_n2756_), .A1(new_n649_), .B0(new_n651_), .Y(new_n2757_));
  AOI21X1  g2372(.A0(new_n2757_), .A1(new_n656_), .B0(new_n659_), .Y(new_n2758_));
  OAI21X1  g2373(.A0(new_n2758_), .A1(new_n664_), .B0(new_n666_), .Y(new_n2759_));
  AOI21X1  g2374(.A0(new_n2759_), .A1(new_n671_), .B0(new_n674_), .Y(new_n2760_));
  OAI21X1  g2375(.A0(new_n2760_), .A1(new_n679_), .B0(new_n681_), .Y(new_n2761_));
  AOI21X1  g2376(.A0(new_n2761_), .A1(new_n686_), .B0(new_n689_), .Y(new_n2762_));
  OAI21X1  g2377(.A0(new_n2762_), .A1(new_n694_), .B0(new_n696_), .Y(new_n2763_));
  AOI21X1  g2378(.A0(new_n2763_), .A1(new_n701_), .B0(new_n1662_), .Y(new_n2764_));
  OAI21X1  g2379(.A0(new_n2764_), .A1(new_n1661_), .B0(new_n1705_), .Y(new_n2765_));
  AOI21X1  g2380(.A0(new_n2765_), .A1(new_n1660_), .B0(new_n1938_), .Y(new_n2766_));
  OAI21X1  g2381(.A0(new_n2766_), .A1(new_n1504_), .B0(new_n721_), .Y(new_n2767_));
  AOI21X1  g2382(.A0(new_n2767_), .A1(new_n1502_), .B0(new_n1503_), .Y(new_n2768_));
  OAI21X1  g2383(.A0(new_n2768_), .A1(new_n1501_), .B0(new_n736_), .Y(new_n2769_));
  AOI21X1  g2384(.A0(new_n2769_), .A1(new_n1499_), .B0(new_n1500_), .Y(new_n2770_));
  OAI21X1  g2385(.A0(new_n2770_), .A1(new_n1498_), .B0(new_n751_), .Y(new_n2771_));
  AOI21X1  g2386(.A0(new_n2771_), .A1(new_n1496_), .B0(new_n1497_), .Y(new_n2772_));
  OAI21X1  g2387(.A0(new_n2772_), .A1(new_n1495_), .B0(new_n766_), .Y(new_n2773_));
  OAI21X1  g2388(.A0(new_n1084_), .A1(\priority[30] ), .B0(\req[30] ), .Y(new_n2774_));
  AOI21X1  g2389(.A0(new_n2773_), .A1(new_n1493_), .B0(new_n2774_), .Y(\grant[30] ));
  NOR2X1   g2390(.A(new_n1092_), .B(new_n780_), .Y(new_n2776_));
  OAI21X1  g2391(.A0(new_n2776_), .A1(new_n787_), .B0(new_n789_), .Y(new_n2777_));
  AOI21X1  g2392(.A0(new_n2777_), .A1(new_n794_), .B0(new_n797_), .Y(new_n2778_));
  OAI21X1  g2393(.A0(new_n2778_), .A1(new_n802_), .B0(new_n804_), .Y(new_n2779_));
  AOI21X1  g2394(.A0(new_n2779_), .A1(new_n809_), .B0(new_n812_), .Y(new_n2780_));
  OAI21X1  g2395(.A0(new_n2780_), .A1(new_n817_), .B0(new_n819_), .Y(new_n2781_));
  AOI21X1  g2396(.A0(new_n2781_), .A1(new_n824_), .B0(new_n827_), .Y(new_n2782_));
  OAI21X1  g2397(.A0(new_n2782_), .A1(new_n832_), .B0(new_n834_), .Y(new_n2783_));
  AOI21X1  g2398(.A0(new_n2783_), .A1(new_n839_), .B0(new_n842_), .Y(new_n2784_));
  OAI21X1  g2399(.A0(new_n2784_), .A1(new_n847_), .B0(new_n849_), .Y(new_n2785_));
  AOI21X1  g2400(.A0(new_n2785_), .A1(new_n854_), .B0(new_n857_), .Y(new_n2786_));
  OAI21X1  g2401(.A0(new_n2786_), .A1(new_n862_), .B0(new_n864_), .Y(new_n2787_));
  AOI21X1  g2402(.A0(new_n2787_), .A1(new_n869_), .B0(new_n872_), .Y(new_n2788_));
  OAI21X1  g2403(.A0(new_n2788_), .A1(new_n877_), .B0(new_n879_), .Y(new_n2789_));
  AOI21X1  g2404(.A0(new_n2789_), .A1(new_n884_), .B0(new_n887_), .Y(new_n2790_));
  OAI21X1  g2405(.A0(new_n2790_), .A1(new_n892_), .B0(new_n894_), .Y(new_n2791_));
  AOI21X1  g2406(.A0(new_n2791_), .A1(new_n899_), .B0(new_n902_), .Y(new_n2792_));
  OAI21X1  g2407(.A0(new_n2792_), .A1(new_n907_), .B0(new_n909_), .Y(new_n2793_));
  AOI21X1  g2408(.A0(new_n2793_), .A1(new_n914_), .B0(new_n917_), .Y(new_n2794_));
  OAI21X1  g2409(.A0(new_n2794_), .A1(new_n922_), .B0(new_n924_), .Y(new_n2795_));
  AOI21X1  g2410(.A0(new_n2795_), .A1(new_n929_), .B0(new_n932_), .Y(new_n2796_));
  OAI21X1  g2411(.A0(new_n2796_), .A1(new_n937_), .B0(new_n939_), .Y(new_n2797_));
  AOI21X1  g2412(.A0(new_n2797_), .A1(new_n944_), .B0(new_n947_), .Y(new_n2798_));
  OAI21X1  g2413(.A0(new_n2798_), .A1(new_n952_), .B0(new_n954_), .Y(new_n2799_));
  AOI21X1  g2414(.A0(new_n2799_), .A1(new_n959_), .B0(new_n962_), .Y(new_n2800_));
  OAI21X1  g2415(.A0(new_n2800_), .A1(new_n967_), .B0(new_n969_), .Y(new_n2801_));
  AOI21X1  g2416(.A0(new_n2801_), .A1(new_n974_), .B0(new_n977_), .Y(new_n2802_));
  OAI21X1  g2417(.A0(new_n2802_), .A1(new_n982_), .B0(new_n984_), .Y(new_n2803_));
  AOI21X1  g2418(.A0(new_n2803_), .A1(new_n989_), .B0(new_n992_), .Y(new_n2804_));
  OAI21X1  g2419(.A0(new_n2804_), .A1(new_n997_), .B0(new_n999_), .Y(new_n2805_));
  AOI21X1  g2420(.A0(new_n2805_), .A1(new_n1004_), .B0(new_n1007_), .Y(new_n2806_));
  OAI21X1  g2421(.A0(new_n2806_), .A1(new_n1012_), .B0(new_n1014_), .Y(new_n2807_));
  AOI21X1  g2422(.A0(new_n2807_), .A1(new_n1017_), .B0(new_n1711_), .Y(new_n2808_));
  OAI21X1  g2423(.A0(new_n2808_), .A1(new_n1710_), .B0(new_n1754_), .Y(new_n2809_));
  AOI21X1  g2424(.A0(new_n2809_), .A1(new_n1709_), .B0(new_n1983_), .Y(new_n2810_));
  OAI21X1  g2425(.A0(new_n2810_), .A1(new_n1613_), .B0(new_n1035_), .Y(new_n2811_));
  AOI21X1  g2426(.A0(new_n2811_), .A1(new_n1611_), .B0(new_n1612_), .Y(new_n2812_));
  OAI21X1  g2427(.A0(new_n2812_), .A1(new_n1610_), .B0(new_n1050_), .Y(new_n2813_));
  AOI21X1  g2428(.A0(new_n2813_), .A1(new_n1608_), .B0(new_n1609_), .Y(new_n2814_));
  OAI21X1  g2429(.A0(new_n2814_), .A1(new_n1607_), .B0(new_n1065_), .Y(new_n2815_));
  AOI21X1  g2430(.A0(new_n2815_), .A1(new_n1605_), .B0(new_n1606_), .Y(new_n2816_));
  OAI21X1  g2431(.A0(new_n2816_), .A1(new_n1604_), .B0(new_n1080_), .Y(new_n2817_));
  OAI21X1  g2432(.A0(new_n459_), .A1(\priority[31] ), .B0(\req[31] ), .Y(new_n2818_));
  AOI21X1  g2433(.A0(new_n2817_), .A1(new_n1602_), .B0(new_n2818_), .Y(\grant[31] ));
  NOR2X1   g2434(.A(new_n1094_), .B(new_n468_), .Y(new_n2820_));
  OAI21X1  g2435(.A0(new_n2820_), .A1(new_n1101_), .B0(new_n1103_), .Y(new_n2821_));
  AOI21X1  g2436(.A0(new_n2821_), .A1(new_n1108_), .B0(new_n1111_), .Y(new_n2822_));
  OAI21X1  g2437(.A0(new_n2822_), .A1(new_n1116_), .B0(new_n1118_), .Y(new_n2823_));
  AOI21X1  g2438(.A0(new_n2823_), .A1(new_n1123_), .B0(new_n1126_), .Y(new_n2824_));
  OAI21X1  g2439(.A0(new_n2824_), .A1(new_n1131_), .B0(new_n1133_), .Y(new_n2825_));
  AOI21X1  g2440(.A0(new_n2825_), .A1(new_n1138_), .B0(new_n1141_), .Y(new_n2826_));
  OAI21X1  g2441(.A0(new_n2826_), .A1(new_n1146_), .B0(new_n1148_), .Y(new_n2827_));
  AOI21X1  g2442(.A0(new_n2827_), .A1(new_n1153_), .B0(new_n1156_), .Y(new_n2828_));
  OAI21X1  g2443(.A0(new_n2828_), .A1(new_n1161_), .B0(new_n1163_), .Y(new_n2829_));
  AOI21X1  g2444(.A0(new_n2829_), .A1(new_n1168_), .B0(new_n1171_), .Y(new_n2830_));
  OAI21X1  g2445(.A0(new_n2830_), .A1(new_n1176_), .B0(new_n1178_), .Y(new_n2831_));
  AOI21X1  g2446(.A0(new_n2831_), .A1(new_n1183_), .B0(new_n1186_), .Y(new_n2832_));
  OAI21X1  g2447(.A0(new_n2832_), .A1(new_n1191_), .B0(new_n1193_), .Y(new_n2833_));
  AOI21X1  g2448(.A0(new_n2833_), .A1(new_n1198_), .B0(new_n1201_), .Y(new_n2834_));
  OAI21X1  g2449(.A0(new_n2834_), .A1(new_n1206_), .B0(new_n1208_), .Y(new_n2835_));
  AOI21X1  g2450(.A0(new_n2835_), .A1(new_n1213_), .B0(new_n1216_), .Y(new_n2836_));
  OAI21X1  g2451(.A0(new_n2836_), .A1(new_n1221_), .B0(new_n1223_), .Y(new_n2837_));
  AOI21X1  g2452(.A0(new_n2837_), .A1(new_n1228_), .B0(new_n1231_), .Y(new_n2838_));
  OAI21X1  g2453(.A0(new_n2838_), .A1(new_n1236_), .B0(new_n1238_), .Y(new_n2839_));
  AOI21X1  g2454(.A0(new_n2839_), .A1(new_n1243_), .B0(new_n1246_), .Y(new_n2840_));
  OAI21X1  g2455(.A0(new_n2840_), .A1(new_n1251_), .B0(new_n1253_), .Y(new_n2841_));
  AOI21X1  g2456(.A0(new_n2841_), .A1(new_n1258_), .B0(new_n1261_), .Y(new_n2842_));
  OAI21X1  g2457(.A0(new_n2842_), .A1(new_n1266_), .B0(new_n1268_), .Y(new_n2843_));
  AOI21X1  g2458(.A0(new_n2843_), .A1(new_n1273_), .B0(new_n1276_), .Y(new_n2844_));
  OAI21X1  g2459(.A0(new_n2844_), .A1(new_n1281_), .B0(new_n1283_), .Y(new_n2845_));
  AOI21X1  g2460(.A0(new_n2845_), .A1(new_n1288_), .B0(new_n1291_), .Y(new_n2846_));
  OAI21X1  g2461(.A0(new_n2846_), .A1(new_n1296_), .B0(new_n1298_), .Y(new_n2847_));
  AOI21X1  g2462(.A0(new_n2847_), .A1(new_n1303_), .B0(new_n1306_), .Y(new_n2848_));
  OAI21X1  g2463(.A0(new_n2848_), .A1(new_n1311_), .B0(new_n1313_), .Y(new_n2849_));
  AOI21X1  g2464(.A0(new_n2849_), .A1(new_n1318_), .B0(new_n1321_), .Y(new_n2850_));
  OAI21X1  g2465(.A0(new_n2850_), .A1(new_n1326_), .B0(new_n1328_), .Y(new_n2851_));
  AOI21X1  g2466(.A0(new_n2851_), .A1(new_n1331_), .B0(new_n1758_), .Y(new_n2852_));
  OAI21X1  g2467(.A0(new_n2852_), .A1(new_n394_), .B0(new_n396_), .Y(new_n2853_));
  AOI21X1  g2468(.A0(new_n2853_), .A1(new_n401_), .B0(new_n404_), .Y(new_n2854_));
  OAI21X1  g2469(.A0(new_n2854_), .A1(new_n409_), .B0(new_n411_), .Y(new_n2855_));
  AOI21X1  g2470(.A0(new_n2855_), .A1(new_n416_), .B0(new_n419_), .Y(new_n2856_));
  OAI21X1  g2471(.A0(new_n2856_), .A1(new_n424_), .B0(new_n426_), .Y(new_n2857_));
  AOI21X1  g2472(.A0(new_n2857_), .A1(new_n431_), .B0(new_n434_), .Y(new_n2858_));
  OAI21X1  g2473(.A0(new_n2858_), .A1(new_n439_), .B0(new_n441_), .Y(new_n2859_));
  AOI21X1  g2474(.A0(new_n2859_), .A1(new_n446_), .B0(new_n449_), .Y(new_n2860_));
  OAI21X1  g2475(.A0(new_n2860_), .A1(new_n454_), .B0(new_n456_), .Y(new_n2861_));
  OAI21X1  g2476(.A0(new_n777_), .A1(\priority[32] ), .B0(\req[32] ), .Y(new_n2862_));
  AOI21X1  g2477(.A0(new_n2861_), .A1(new_n461_), .B0(new_n2862_), .Y(\grant[32] ));
  NOR2X1   g2478(.A(new_n786_), .B(new_n470_), .Y(new_n2864_));
  OAI21X1  g2479(.A0(new_n2864_), .A1(new_n1380_), .B0(new_n478_), .Y(new_n2865_));
  AOI21X1  g2480(.A0(new_n2865_), .A1(new_n1378_), .B0(new_n1379_), .Y(new_n2866_));
  OAI21X1  g2481(.A0(new_n2866_), .A1(new_n1377_), .B0(new_n493_), .Y(new_n2867_));
  AOI21X1  g2482(.A0(new_n2867_), .A1(new_n1375_), .B0(new_n1376_), .Y(new_n2868_));
  OAI21X1  g2483(.A0(new_n2868_), .A1(new_n1374_), .B0(new_n508_), .Y(new_n2869_));
  AOI21X1  g2484(.A0(new_n2869_), .A1(new_n1372_), .B0(new_n1373_), .Y(new_n2870_));
  OAI21X1  g2485(.A0(new_n2870_), .A1(new_n1371_), .B0(new_n523_), .Y(new_n2871_));
  AOI21X1  g2486(.A0(new_n2871_), .A1(new_n1369_), .B0(new_n1370_), .Y(new_n2872_));
  OAI21X1  g2487(.A0(new_n2872_), .A1(new_n1368_), .B0(new_n538_), .Y(new_n2873_));
  AOI21X1  g2488(.A0(new_n2873_), .A1(new_n1366_), .B0(new_n1367_), .Y(new_n2874_));
  OAI21X1  g2489(.A0(new_n2874_), .A1(new_n1365_), .B0(new_n553_), .Y(new_n2875_));
  AOI21X1  g2490(.A0(new_n2875_), .A1(new_n1363_), .B0(new_n1364_), .Y(new_n2876_));
  OAI21X1  g2491(.A0(new_n2876_), .A1(new_n1362_), .B0(new_n568_), .Y(new_n2877_));
  AOI21X1  g2492(.A0(new_n2877_), .A1(new_n1360_), .B0(new_n1361_), .Y(new_n2878_));
  OAI21X1  g2493(.A0(new_n2878_), .A1(new_n1359_), .B0(new_n583_), .Y(new_n2879_));
  AOI21X1  g2494(.A0(new_n2879_), .A1(new_n1357_), .B0(new_n1358_), .Y(new_n2880_));
  OAI21X1  g2495(.A0(new_n2880_), .A1(new_n1356_), .B0(new_n598_), .Y(new_n2881_));
  AOI21X1  g2496(.A0(new_n2881_), .A1(new_n1354_), .B0(new_n1355_), .Y(new_n2882_));
  OAI21X1  g2497(.A0(new_n2882_), .A1(new_n1353_), .B0(new_n613_), .Y(new_n2883_));
  AOI21X1  g2498(.A0(new_n2883_), .A1(new_n1351_), .B0(new_n1352_), .Y(new_n2884_));
  OAI21X1  g2499(.A0(new_n2884_), .A1(new_n1350_), .B0(new_n628_), .Y(new_n2885_));
  AOI21X1  g2500(.A0(new_n2885_), .A1(new_n1348_), .B0(new_n1349_), .Y(new_n2886_));
  OAI21X1  g2501(.A0(new_n2886_), .A1(new_n1347_), .B0(new_n643_), .Y(new_n2887_));
  AOI21X1  g2502(.A0(new_n2887_), .A1(new_n1345_), .B0(new_n1346_), .Y(new_n2888_));
  OAI21X1  g2503(.A0(new_n2888_), .A1(new_n1344_), .B0(new_n658_), .Y(new_n2889_));
  AOI21X1  g2504(.A0(new_n2889_), .A1(new_n1342_), .B0(new_n1343_), .Y(new_n2890_));
  OAI21X1  g2505(.A0(new_n2890_), .A1(new_n1341_), .B0(new_n673_), .Y(new_n2891_));
  AOI21X1  g2506(.A0(new_n2891_), .A1(new_n1339_), .B0(new_n1340_), .Y(new_n2892_));
  OAI21X1  g2507(.A0(new_n2892_), .A1(new_n1338_), .B0(new_n688_), .Y(new_n2893_));
  AOI21X1  g2508(.A0(new_n2893_), .A1(new_n1336_), .B0(new_n1337_), .Y(new_n2894_));
  OAI21X1  g2509(.A0(new_n2894_), .A1(new_n1335_), .B0(new_n1438_), .Y(new_n2895_));
  AOI21X1  g2510(.A0(new_n2895_), .A1(new_n1440_), .B0(new_n1803_), .Y(new_n2896_));
  OAI21X1  g2511(.A0(new_n2896_), .A1(new_n712_), .B0(new_n714_), .Y(new_n2897_));
  AOI21X1  g2512(.A0(new_n2897_), .A1(new_n719_), .B0(new_n722_), .Y(new_n2898_));
  OAI21X1  g2513(.A0(new_n2898_), .A1(new_n727_), .B0(new_n729_), .Y(new_n2899_));
  AOI21X1  g2514(.A0(new_n2899_), .A1(new_n734_), .B0(new_n737_), .Y(new_n2900_));
  OAI21X1  g2515(.A0(new_n2900_), .A1(new_n742_), .B0(new_n744_), .Y(new_n2901_));
  AOI21X1  g2516(.A0(new_n2901_), .A1(new_n749_), .B0(new_n752_), .Y(new_n2902_));
  OAI21X1  g2517(.A0(new_n2902_), .A1(new_n757_), .B0(new_n759_), .Y(new_n2903_));
  AOI21X1  g2518(.A0(new_n2903_), .A1(new_n764_), .B0(new_n767_), .Y(new_n2904_));
  OAI21X1  g2519(.A0(new_n2904_), .A1(new_n772_), .B0(new_n774_), .Y(new_n2905_));
  OAI21X1  g2520(.A0(new_n1091_), .A1(\priority[33] ), .B0(\req[33] ), .Y(new_n2906_));
  AOI21X1  g2521(.A0(new_n2905_), .A1(new_n779_), .B0(new_n2906_), .Y(\grant[33] ));
  NOR2X1   g2522(.A(new_n1100_), .B(new_n788_), .Y(new_n2908_));
  OAI21X1  g2523(.A0(new_n2908_), .A1(new_n1489_), .B0(new_n796_), .Y(new_n2909_));
  AOI21X1  g2524(.A0(new_n2909_), .A1(new_n1487_), .B0(new_n1488_), .Y(new_n2910_));
  OAI21X1  g2525(.A0(new_n2910_), .A1(new_n1486_), .B0(new_n811_), .Y(new_n2911_));
  AOI21X1  g2526(.A0(new_n2911_), .A1(new_n1484_), .B0(new_n1485_), .Y(new_n2912_));
  OAI21X1  g2527(.A0(new_n2912_), .A1(new_n1483_), .B0(new_n826_), .Y(new_n2913_));
  AOI21X1  g2528(.A0(new_n2913_), .A1(new_n1481_), .B0(new_n1482_), .Y(new_n2914_));
  OAI21X1  g2529(.A0(new_n2914_), .A1(new_n1480_), .B0(new_n841_), .Y(new_n2915_));
  AOI21X1  g2530(.A0(new_n2915_), .A1(new_n1478_), .B0(new_n1479_), .Y(new_n2916_));
  OAI21X1  g2531(.A0(new_n2916_), .A1(new_n1477_), .B0(new_n856_), .Y(new_n2917_));
  AOI21X1  g2532(.A0(new_n2917_), .A1(new_n1475_), .B0(new_n1476_), .Y(new_n2918_));
  OAI21X1  g2533(.A0(new_n2918_), .A1(new_n1474_), .B0(new_n871_), .Y(new_n2919_));
  AOI21X1  g2534(.A0(new_n2919_), .A1(new_n1472_), .B0(new_n1473_), .Y(new_n2920_));
  OAI21X1  g2535(.A0(new_n2920_), .A1(new_n1471_), .B0(new_n886_), .Y(new_n2921_));
  AOI21X1  g2536(.A0(new_n2921_), .A1(new_n1469_), .B0(new_n1470_), .Y(new_n2922_));
  OAI21X1  g2537(.A0(new_n2922_), .A1(new_n1468_), .B0(new_n901_), .Y(new_n2923_));
  AOI21X1  g2538(.A0(new_n2923_), .A1(new_n1466_), .B0(new_n1467_), .Y(new_n2924_));
  OAI21X1  g2539(.A0(new_n2924_), .A1(new_n1465_), .B0(new_n916_), .Y(new_n2925_));
  AOI21X1  g2540(.A0(new_n2925_), .A1(new_n1463_), .B0(new_n1464_), .Y(new_n2926_));
  OAI21X1  g2541(.A0(new_n2926_), .A1(new_n1462_), .B0(new_n931_), .Y(new_n2927_));
  AOI21X1  g2542(.A0(new_n2927_), .A1(new_n1460_), .B0(new_n1461_), .Y(new_n2928_));
  OAI21X1  g2543(.A0(new_n2928_), .A1(new_n1459_), .B0(new_n946_), .Y(new_n2929_));
  AOI21X1  g2544(.A0(new_n2929_), .A1(new_n1457_), .B0(new_n1458_), .Y(new_n2930_));
  OAI21X1  g2545(.A0(new_n2930_), .A1(new_n1456_), .B0(new_n961_), .Y(new_n2931_));
  AOI21X1  g2546(.A0(new_n2931_), .A1(new_n1454_), .B0(new_n1455_), .Y(new_n2932_));
  OAI21X1  g2547(.A0(new_n2932_), .A1(new_n1453_), .B0(new_n976_), .Y(new_n2933_));
  AOI21X1  g2548(.A0(new_n2933_), .A1(new_n1451_), .B0(new_n1452_), .Y(new_n2934_));
  OAI21X1  g2549(.A0(new_n2934_), .A1(new_n1450_), .B0(new_n991_), .Y(new_n2935_));
  AOI21X1  g2550(.A0(new_n2935_), .A1(new_n1448_), .B0(new_n1449_), .Y(new_n2936_));
  OAI21X1  g2551(.A0(new_n2936_), .A1(new_n1447_), .B0(new_n1006_), .Y(new_n2937_));
  AOI21X1  g2552(.A0(new_n2937_), .A1(new_n1445_), .B0(new_n1446_), .Y(new_n2938_));
  OAI21X1  g2553(.A0(new_n2938_), .A1(new_n1444_), .B0(new_n1547_), .Y(new_n2939_));
  AOI21X1  g2554(.A0(new_n2939_), .A1(new_n1549_), .B0(new_n1848_), .Y(new_n2940_));
  OAI21X1  g2555(.A0(new_n2940_), .A1(new_n1026_), .B0(new_n1028_), .Y(new_n2941_));
  AOI21X1  g2556(.A0(new_n2941_), .A1(new_n1033_), .B0(new_n1036_), .Y(new_n2942_));
  OAI21X1  g2557(.A0(new_n2942_), .A1(new_n1041_), .B0(new_n1043_), .Y(new_n2943_));
  AOI21X1  g2558(.A0(new_n2943_), .A1(new_n1048_), .B0(new_n1051_), .Y(new_n2944_));
  OAI21X1  g2559(.A0(new_n2944_), .A1(new_n1056_), .B0(new_n1058_), .Y(new_n2945_));
  AOI21X1  g2560(.A0(new_n2945_), .A1(new_n1063_), .B0(new_n1066_), .Y(new_n2946_));
  OAI21X1  g2561(.A0(new_n2946_), .A1(new_n1071_), .B0(new_n1073_), .Y(new_n2947_));
  AOI21X1  g2562(.A0(new_n2947_), .A1(new_n1078_), .B0(new_n1081_), .Y(new_n2948_));
  OAI21X1  g2563(.A0(new_n2948_), .A1(new_n1086_), .B0(new_n1088_), .Y(new_n2949_));
  OAI21X1  g2564(.A0(new_n467_), .A1(\priority[34] ), .B0(\req[34] ), .Y(new_n2950_));
  AOI21X1  g2565(.A0(new_n2949_), .A1(new_n1093_), .B0(new_n2950_), .Y(\grant[34] ));
  NOR2X1   g2566(.A(new_n1102_), .B(new_n475_), .Y(new_n2952_));
  OAI21X1  g2567(.A0(new_n2952_), .A1(new_n1598_), .B0(new_n1110_), .Y(new_n2953_));
  AOI21X1  g2568(.A0(new_n2953_), .A1(new_n1596_), .B0(new_n1597_), .Y(new_n2954_));
  OAI21X1  g2569(.A0(new_n2954_), .A1(new_n1595_), .B0(new_n1125_), .Y(new_n2955_));
  AOI21X1  g2570(.A0(new_n2955_), .A1(new_n1593_), .B0(new_n1594_), .Y(new_n2956_));
  OAI21X1  g2571(.A0(new_n2956_), .A1(new_n1592_), .B0(new_n1140_), .Y(new_n2957_));
  AOI21X1  g2572(.A0(new_n2957_), .A1(new_n1590_), .B0(new_n1591_), .Y(new_n2958_));
  OAI21X1  g2573(.A0(new_n2958_), .A1(new_n1589_), .B0(new_n1155_), .Y(new_n2959_));
  AOI21X1  g2574(.A0(new_n2959_), .A1(new_n1587_), .B0(new_n1588_), .Y(new_n2960_));
  OAI21X1  g2575(.A0(new_n2960_), .A1(new_n1586_), .B0(new_n1170_), .Y(new_n2961_));
  AOI21X1  g2576(.A0(new_n2961_), .A1(new_n1584_), .B0(new_n1585_), .Y(new_n2962_));
  OAI21X1  g2577(.A0(new_n2962_), .A1(new_n1583_), .B0(new_n1185_), .Y(new_n2963_));
  AOI21X1  g2578(.A0(new_n2963_), .A1(new_n1581_), .B0(new_n1582_), .Y(new_n2964_));
  OAI21X1  g2579(.A0(new_n2964_), .A1(new_n1580_), .B0(new_n1200_), .Y(new_n2965_));
  AOI21X1  g2580(.A0(new_n2965_), .A1(new_n1578_), .B0(new_n1579_), .Y(new_n2966_));
  OAI21X1  g2581(.A0(new_n2966_), .A1(new_n1577_), .B0(new_n1215_), .Y(new_n2967_));
  AOI21X1  g2582(.A0(new_n2967_), .A1(new_n1575_), .B0(new_n1576_), .Y(new_n2968_));
  OAI21X1  g2583(.A0(new_n2968_), .A1(new_n1574_), .B0(new_n1230_), .Y(new_n2969_));
  AOI21X1  g2584(.A0(new_n2969_), .A1(new_n1572_), .B0(new_n1573_), .Y(new_n2970_));
  OAI21X1  g2585(.A0(new_n2970_), .A1(new_n1571_), .B0(new_n1245_), .Y(new_n2971_));
  AOI21X1  g2586(.A0(new_n2971_), .A1(new_n1569_), .B0(new_n1570_), .Y(new_n2972_));
  OAI21X1  g2587(.A0(new_n2972_), .A1(new_n1568_), .B0(new_n1260_), .Y(new_n2973_));
  AOI21X1  g2588(.A0(new_n2973_), .A1(new_n1566_), .B0(new_n1567_), .Y(new_n2974_));
  OAI21X1  g2589(.A0(new_n2974_), .A1(new_n1565_), .B0(new_n1275_), .Y(new_n2975_));
  AOI21X1  g2590(.A0(new_n2975_), .A1(new_n1563_), .B0(new_n1564_), .Y(new_n2976_));
  OAI21X1  g2591(.A0(new_n2976_), .A1(new_n1562_), .B0(new_n1290_), .Y(new_n2977_));
  AOI21X1  g2592(.A0(new_n2977_), .A1(new_n1560_), .B0(new_n1561_), .Y(new_n2978_));
  OAI21X1  g2593(.A0(new_n2978_), .A1(new_n1559_), .B0(new_n1305_), .Y(new_n2979_));
  AOI21X1  g2594(.A0(new_n2979_), .A1(new_n1557_), .B0(new_n1558_), .Y(new_n2980_));
  OAI21X1  g2595(.A0(new_n2980_), .A1(new_n1556_), .B0(new_n1320_), .Y(new_n2981_));
  AOI21X1  g2596(.A0(new_n2981_), .A1(new_n1554_), .B0(new_n1555_), .Y(new_n2982_));
  OAI21X1  g2597(.A0(new_n2982_), .A1(new_n1553_), .B0(new_n1656_), .Y(new_n2983_));
  AOI21X1  g2598(.A0(new_n2983_), .A1(new_n1552_), .B0(new_n1893_), .Y(new_n2984_));
  OAI21X1  g2599(.A0(new_n2984_), .A1(new_n1395_), .B0(new_n403_), .Y(new_n2985_));
  AOI21X1  g2600(.A0(new_n2985_), .A1(new_n1393_), .B0(new_n1394_), .Y(new_n2986_));
  OAI21X1  g2601(.A0(new_n2986_), .A1(new_n1392_), .B0(new_n418_), .Y(new_n2987_));
  AOI21X1  g2602(.A0(new_n2987_), .A1(new_n1390_), .B0(new_n1391_), .Y(new_n2988_));
  OAI21X1  g2603(.A0(new_n2988_), .A1(new_n1389_), .B0(new_n433_), .Y(new_n2989_));
  AOI21X1  g2604(.A0(new_n2989_), .A1(new_n1387_), .B0(new_n1388_), .Y(new_n2990_));
  OAI21X1  g2605(.A0(new_n2990_), .A1(new_n1386_), .B0(new_n448_), .Y(new_n2991_));
  AOI21X1  g2606(.A0(new_n2991_), .A1(new_n1384_), .B0(new_n1385_), .Y(new_n2992_));
  OAI21X1  g2607(.A0(new_n2992_), .A1(new_n1383_), .B0(new_n463_), .Y(new_n2993_));
  OAI21X1  g2608(.A0(new_n785_), .A1(\priority[35] ), .B0(\req[35] ), .Y(new_n2994_));
  AOI21X1  g2609(.A0(new_n2993_), .A1(new_n1381_), .B0(new_n2994_), .Y(\grant[35] ));
  NOR2X1   g2610(.A(new_n793_), .B(new_n477_), .Y(new_n2996_));
  OAI21X1  g2611(.A0(new_n2996_), .A1(new_n484_), .B0(new_n486_), .Y(new_n2997_));
  AOI21X1  g2612(.A0(new_n2997_), .A1(new_n491_), .B0(new_n494_), .Y(new_n2998_));
  OAI21X1  g2613(.A0(new_n2998_), .A1(new_n499_), .B0(new_n501_), .Y(new_n2999_));
  AOI21X1  g2614(.A0(new_n2999_), .A1(new_n506_), .B0(new_n509_), .Y(new_n3000_));
  OAI21X1  g2615(.A0(new_n3000_), .A1(new_n514_), .B0(new_n516_), .Y(new_n3001_));
  AOI21X1  g2616(.A0(new_n3001_), .A1(new_n521_), .B0(new_n524_), .Y(new_n3002_));
  OAI21X1  g2617(.A0(new_n3002_), .A1(new_n529_), .B0(new_n531_), .Y(new_n3003_));
  AOI21X1  g2618(.A0(new_n3003_), .A1(new_n536_), .B0(new_n539_), .Y(new_n3004_));
  OAI21X1  g2619(.A0(new_n3004_), .A1(new_n544_), .B0(new_n546_), .Y(new_n3005_));
  AOI21X1  g2620(.A0(new_n3005_), .A1(new_n551_), .B0(new_n554_), .Y(new_n3006_));
  OAI21X1  g2621(.A0(new_n3006_), .A1(new_n559_), .B0(new_n561_), .Y(new_n3007_));
  AOI21X1  g2622(.A0(new_n3007_), .A1(new_n566_), .B0(new_n569_), .Y(new_n3008_));
  OAI21X1  g2623(.A0(new_n3008_), .A1(new_n574_), .B0(new_n576_), .Y(new_n3009_));
  AOI21X1  g2624(.A0(new_n3009_), .A1(new_n581_), .B0(new_n584_), .Y(new_n3010_));
  OAI21X1  g2625(.A0(new_n3010_), .A1(new_n589_), .B0(new_n591_), .Y(new_n3011_));
  AOI21X1  g2626(.A0(new_n3011_), .A1(new_n596_), .B0(new_n599_), .Y(new_n3012_));
  OAI21X1  g2627(.A0(new_n3012_), .A1(new_n604_), .B0(new_n606_), .Y(new_n3013_));
  AOI21X1  g2628(.A0(new_n3013_), .A1(new_n611_), .B0(new_n614_), .Y(new_n3014_));
  OAI21X1  g2629(.A0(new_n3014_), .A1(new_n619_), .B0(new_n621_), .Y(new_n3015_));
  AOI21X1  g2630(.A0(new_n3015_), .A1(new_n626_), .B0(new_n629_), .Y(new_n3016_));
  OAI21X1  g2631(.A0(new_n3016_), .A1(new_n634_), .B0(new_n636_), .Y(new_n3017_));
  AOI21X1  g2632(.A0(new_n3017_), .A1(new_n641_), .B0(new_n644_), .Y(new_n3018_));
  OAI21X1  g2633(.A0(new_n3018_), .A1(new_n649_), .B0(new_n651_), .Y(new_n3019_));
  AOI21X1  g2634(.A0(new_n3019_), .A1(new_n656_), .B0(new_n659_), .Y(new_n3020_));
  OAI21X1  g2635(.A0(new_n3020_), .A1(new_n664_), .B0(new_n666_), .Y(new_n3021_));
  AOI21X1  g2636(.A0(new_n3021_), .A1(new_n671_), .B0(new_n674_), .Y(new_n3022_));
  OAI21X1  g2637(.A0(new_n3022_), .A1(new_n679_), .B0(new_n681_), .Y(new_n3023_));
  AOI21X1  g2638(.A0(new_n3023_), .A1(new_n686_), .B0(new_n689_), .Y(new_n3024_));
  OAI21X1  g2639(.A0(new_n3024_), .A1(new_n694_), .B0(new_n696_), .Y(new_n3025_));
  AOI21X1  g2640(.A0(new_n3025_), .A1(new_n701_), .B0(new_n1662_), .Y(new_n3026_));
  OAI21X1  g2641(.A0(new_n3026_), .A1(new_n1661_), .B0(new_n1705_), .Y(new_n3027_));
  AOI21X1  g2642(.A0(new_n3027_), .A1(new_n1660_), .B0(new_n1938_), .Y(new_n3028_));
  OAI21X1  g2643(.A0(new_n3028_), .A1(new_n1504_), .B0(new_n721_), .Y(new_n3029_));
  AOI21X1  g2644(.A0(new_n3029_), .A1(new_n1502_), .B0(new_n1503_), .Y(new_n3030_));
  OAI21X1  g2645(.A0(new_n3030_), .A1(new_n1501_), .B0(new_n736_), .Y(new_n3031_));
  AOI21X1  g2646(.A0(new_n3031_), .A1(new_n1499_), .B0(new_n1500_), .Y(new_n3032_));
  OAI21X1  g2647(.A0(new_n3032_), .A1(new_n1498_), .B0(new_n751_), .Y(new_n3033_));
  AOI21X1  g2648(.A0(new_n3033_), .A1(new_n1496_), .B0(new_n1497_), .Y(new_n3034_));
  OAI21X1  g2649(.A0(new_n3034_), .A1(new_n1495_), .B0(new_n766_), .Y(new_n3035_));
  AOI21X1  g2650(.A0(new_n3035_), .A1(new_n1493_), .B0(new_n1494_), .Y(new_n3036_));
  OAI21X1  g2651(.A0(new_n3036_), .A1(new_n1492_), .B0(new_n781_), .Y(new_n3037_));
  OAI21X1  g2652(.A0(new_n1099_), .A1(\priority[36] ), .B0(\req[36] ), .Y(new_n3038_));
  AOI21X1  g2653(.A0(new_n3037_), .A1(new_n1490_), .B0(new_n3038_), .Y(\grant[36] ));
  NOR2X1   g2654(.A(new_n1107_), .B(new_n795_), .Y(new_n3040_));
  OAI21X1  g2655(.A0(new_n3040_), .A1(new_n802_), .B0(new_n804_), .Y(new_n3041_));
  AOI21X1  g2656(.A0(new_n3041_), .A1(new_n809_), .B0(new_n812_), .Y(new_n3042_));
  OAI21X1  g2657(.A0(new_n3042_), .A1(new_n817_), .B0(new_n819_), .Y(new_n3043_));
  AOI21X1  g2658(.A0(new_n3043_), .A1(new_n824_), .B0(new_n827_), .Y(new_n3044_));
  OAI21X1  g2659(.A0(new_n3044_), .A1(new_n832_), .B0(new_n834_), .Y(new_n3045_));
  AOI21X1  g2660(.A0(new_n3045_), .A1(new_n839_), .B0(new_n842_), .Y(new_n3046_));
  OAI21X1  g2661(.A0(new_n3046_), .A1(new_n847_), .B0(new_n849_), .Y(new_n3047_));
  AOI21X1  g2662(.A0(new_n3047_), .A1(new_n854_), .B0(new_n857_), .Y(new_n3048_));
  OAI21X1  g2663(.A0(new_n3048_), .A1(new_n862_), .B0(new_n864_), .Y(new_n3049_));
  AOI21X1  g2664(.A0(new_n3049_), .A1(new_n869_), .B0(new_n872_), .Y(new_n3050_));
  OAI21X1  g2665(.A0(new_n3050_), .A1(new_n877_), .B0(new_n879_), .Y(new_n3051_));
  AOI21X1  g2666(.A0(new_n3051_), .A1(new_n884_), .B0(new_n887_), .Y(new_n3052_));
  OAI21X1  g2667(.A0(new_n3052_), .A1(new_n892_), .B0(new_n894_), .Y(new_n3053_));
  AOI21X1  g2668(.A0(new_n3053_), .A1(new_n899_), .B0(new_n902_), .Y(new_n3054_));
  OAI21X1  g2669(.A0(new_n3054_), .A1(new_n907_), .B0(new_n909_), .Y(new_n3055_));
  AOI21X1  g2670(.A0(new_n3055_), .A1(new_n914_), .B0(new_n917_), .Y(new_n3056_));
  OAI21X1  g2671(.A0(new_n3056_), .A1(new_n922_), .B0(new_n924_), .Y(new_n3057_));
  AOI21X1  g2672(.A0(new_n3057_), .A1(new_n929_), .B0(new_n932_), .Y(new_n3058_));
  OAI21X1  g2673(.A0(new_n3058_), .A1(new_n937_), .B0(new_n939_), .Y(new_n3059_));
  AOI21X1  g2674(.A0(new_n3059_), .A1(new_n944_), .B0(new_n947_), .Y(new_n3060_));
  OAI21X1  g2675(.A0(new_n3060_), .A1(new_n952_), .B0(new_n954_), .Y(new_n3061_));
  AOI21X1  g2676(.A0(new_n3061_), .A1(new_n959_), .B0(new_n962_), .Y(new_n3062_));
  OAI21X1  g2677(.A0(new_n3062_), .A1(new_n967_), .B0(new_n969_), .Y(new_n3063_));
  AOI21X1  g2678(.A0(new_n3063_), .A1(new_n974_), .B0(new_n977_), .Y(new_n3064_));
  OAI21X1  g2679(.A0(new_n3064_), .A1(new_n982_), .B0(new_n984_), .Y(new_n3065_));
  AOI21X1  g2680(.A0(new_n3065_), .A1(new_n989_), .B0(new_n992_), .Y(new_n3066_));
  OAI21X1  g2681(.A0(new_n3066_), .A1(new_n997_), .B0(new_n999_), .Y(new_n3067_));
  AOI21X1  g2682(.A0(new_n3067_), .A1(new_n1004_), .B0(new_n1007_), .Y(new_n3068_));
  OAI21X1  g2683(.A0(new_n3068_), .A1(new_n1012_), .B0(new_n1014_), .Y(new_n3069_));
  AOI21X1  g2684(.A0(new_n3069_), .A1(new_n1017_), .B0(new_n1711_), .Y(new_n3070_));
  OAI21X1  g2685(.A0(new_n3070_), .A1(new_n1710_), .B0(new_n1754_), .Y(new_n3071_));
  AOI21X1  g2686(.A0(new_n3071_), .A1(new_n1709_), .B0(new_n1983_), .Y(new_n3072_));
  OAI21X1  g2687(.A0(new_n3072_), .A1(new_n1613_), .B0(new_n1035_), .Y(new_n3073_));
  AOI21X1  g2688(.A0(new_n3073_), .A1(new_n1611_), .B0(new_n1612_), .Y(new_n3074_));
  OAI21X1  g2689(.A0(new_n3074_), .A1(new_n1610_), .B0(new_n1050_), .Y(new_n3075_));
  AOI21X1  g2690(.A0(new_n3075_), .A1(new_n1608_), .B0(new_n1609_), .Y(new_n3076_));
  OAI21X1  g2691(.A0(new_n3076_), .A1(new_n1607_), .B0(new_n1065_), .Y(new_n3077_));
  AOI21X1  g2692(.A0(new_n3077_), .A1(new_n1605_), .B0(new_n1606_), .Y(new_n3078_));
  OAI21X1  g2693(.A0(new_n3078_), .A1(new_n1604_), .B0(new_n1080_), .Y(new_n3079_));
  AOI21X1  g2694(.A0(new_n3079_), .A1(new_n1602_), .B0(new_n1603_), .Y(new_n3080_));
  OAI21X1  g2695(.A0(new_n3080_), .A1(new_n1601_), .B0(new_n1095_), .Y(new_n3081_));
  OAI21X1  g2696(.A0(new_n474_), .A1(\priority[37] ), .B0(\req[37] ), .Y(new_n3082_));
  AOI21X1  g2697(.A0(new_n3081_), .A1(new_n1599_), .B0(new_n3082_), .Y(\grant[37] ));
  NOR2X1   g2698(.A(new_n1109_), .B(new_n483_), .Y(new_n3084_));
  OAI21X1  g2699(.A0(new_n3084_), .A1(new_n1116_), .B0(new_n1118_), .Y(new_n3085_));
  AOI21X1  g2700(.A0(new_n3085_), .A1(new_n1123_), .B0(new_n1126_), .Y(new_n3086_));
  OAI21X1  g2701(.A0(new_n3086_), .A1(new_n1131_), .B0(new_n1133_), .Y(new_n3087_));
  AOI21X1  g2702(.A0(new_n3087_), .A1(new_n1138_), .B0(new_n1141_), .Y(new_n3088_));
  OAI21X1  g2703(.A0(new_n3088_), .A1(new_n1146_), .B0(new_n1148_), .Y(new_n3089_));
  AOI21X1  g2704(.A0(new_n3089_), .A1(new_n1153_), .B0(new_n1156_), .Y(new_n3090_));
  OAI21X1  g2705(.A0(new_n3090_), .A1(new_n1161_), .B0(new_n1163_), .Y(new_n3091_));
  AOI21X1  g2706(.A0(new_n3091_), .A1(new_n1168_), .B0(new_n1171_), .Y(new_n3092_));
  OAI21X1  g2707(.A0(new_n3092_), .A1(new_n1176_), .B0(new_n1178_), .Y(new_n3093_));
  AOI21X1  g2708(.A0(new_n3093_), .A1(new_n1183_), .B0(new_n1186_), .Y(new_n3094_));
  OAI21X1  g2709(.A0(new_n3094_), .A1(new_n1191_), .B0(new_n1193_), .Y(new_n3095_));
  AOI21X1  g2710(.A0(new_n3095_), .A1(new_n1198_), .B0(new_n1201_), .Y(new_n3096_));
  OAI21X1  g2711(.A0(new_n3096_), .A1(new_n1206_), .B0(new_n1208_), .Y(new_n3097_));
  AOI21X1  g2712(.A0(new_n3097_), .A1(new_n1213_), .B0(new_n1216_), .Y(new_n3098_));
  OAI21X1  g2713(.A0(new_n3098_), .A1(new_n1221_), .B0(new_n1223_), .Y(new_n3099_));
  AOI21X1  g2714(.A0(new_n3099_), .A1(new_n1228_), .B0(new_n1231_), .Y(new_n3100_));
  OAI21X1  g2715(.A0(new_n3100_), .A1(new_n1236_), .B0(new_n1238_), .Y(new_n3101_));
  AOI21X1  g2716(.A0(new_n3101_), .A1(new_n1243_), .B0(new_n1246_), .Y(new_n3102_));
  OAI21X1  g2717(.A0(new_n3102_), .A1(new_n1251_), .B0(new_n1253_), .Y(new_n3103_));
  AOI21X1  g2718(.A0(new_n3103_), .A1(new_n1258_), .B0(new_n1261_), .Y(new_n3104_));
  OAI21X1  g2719(.A0(new_n3104_), .A1(new_n1266_), .B0(new_n1268_), .Y(new_n3105_));
  AOI21X1  g2720(.A0(new_n3105_), .A1(new_n1273_), .B0(new_n1276_), .Y(new_n3106_));
  OAI21X1  g2721(.A0(new_n3106_), .A1(new_n1281_), .B0(new_n1283_), .Y(new_n3107_));
  AOI21X1  g2722(.A0(new_n3107_), .A1(new_n1288_), .B0(new_n1291_), .Y(new_n3108_));
  OAI21X1  g2723(.A0(new_n3108_), .A1(new_n1296_), .B0(new_n1298_), .Y(new_n3109_));
  AOI21X1  g2724(.A0(new_n3109_), .A1(new_n1303_), .B0(new_n1306_), .Y(new_n3110_));
  OAI21X1  g2725(.A0(new_n3110_), .A1(new_n1311_), .B0(new_n1313_), .Y(new_n3111_));
  AOI21X1  g2726(.A0(new_n3111_), .A1(new_n1318_), .B0(new_n1321_), .Y(new_n3112_));
  OAI21X1  g2727(.A0(new_n3112_), .A1(new_n1326_), .B0(new_n1328_), .Y(new_n3113_));
  AOI21X1  g2728(.A0(new_n3113_), .A1(new_n1331_), .B0(new_n1758_), .Y(new_n3114_));
  OAI21X1  g2729(.A0(new_n3114_), .A1(new_n394_), .B0(new_n396_), .Y(new_n3115_));
  AOI21X1  g2730(.A0(new_n3115_), .A1(new_n401_), .B0(new_n404_), .Y(new_n3116_));
  OAI21X1  g2731(.A0(new_n3116_), .A1(new_n409_), .B0(new_n411_), .Y(new_n3117_));
  AOI21X1  g2732(.A0(new_n3117_), .A1(new_n416_), .B0(new_n419_), .Y(new_n3118_));
  OAI21X1  g2733(.A0(new_n3118_), .A1(new_n424_), .B0(new_n426_), .Y(new_n3119_));
  AOI21X1  g2734(.A0(new_n3119_), .A1(new_n431_), .B0(new_n434_), .Y(new_n3120_));
  OAI21X1  g2735(.A0(new_n3120_), .A1(new_n439_), .B0(new_n441_), .Y(new_n3121_));
  AOI21X1  g2736(.A0(new_n3121_), .A1(new_n446_), .B0(new_n449_), .Y(new_n3122_));
  OAI21X1  g2737(.A0(new_n3122_), .A1(new_n454_), .B0(new_n456_), .Y(new_n3123_));
  AOI21X1  g2738(.A0(new_n3123_), .A1(new_n461_), .B0(new_n464_), .Y(new_n3124_));
  OAI21X1  g2739(.A0(new_n3124_), .A1(new_n469_), .B0(new_n471_), .Y(new_n3125_));
  OAI21X1  g2740(.A0(new_n792_), .A1(\priority[38] ), .B0(\req[38] ), .Y(new_n3126_));
  AOI21X1  g2741(.A0(new_n3125_), .A1(new_n476_), .B0(new_n3126_), .Y(\grant[38] ));
  NOR2X1   g2742(.A(new_n801_), .B(new_n485_), .Y(new_n3128_));
  OAI21X1  g2743(.A0(new_n3128_), .A1(new_n1377_), .B0(new_n493_), .Y(new_n3129_));
  AOI21X1  g2744(.A0(new_n3129_), .A1(new_n1375_), .B0(new_n1376_), .Y(new_n3130_));
  OAI21X1  g2745(.A0(new_n3130_), .A1(new_n1374_), .B0(new_n508_), .Y(new_n3131_));
  AOI21X1  g2746(.A0(new_n3131_), .A1(new_n1372_), .B0(new_n1373_), .Y(new_n3132_));
  OAI21X1  g2747(.A0(new_n3132_), .A1(new_n1371_), .B0(new_n523_), .Y(new_n3133_));
  AOI21X1  g2748(.A0(new_n3133_), .A1(new_n1369_), .B0(new_n1370_), .Y(new_n3134_));
  OAI21X1  g2749(.A0(new_n3134_), .A1(new_n1368_), .B0(new_n538_), .Y(new_n3135_));
  AOI21X1  g2750(.A0(new_n3135_), .A1(new_n1366_), .B0(new_n1367_), .Y(new_n3136_));
  OAI21X1  g2751(.A0(new_n3136_), .A1(new_n1365_), .B0(new_n553_), .Y(new_n3137_));
  AOI21X1  g2752(.A0(new_n3137_), .A1(new_n1363_), .B0(new_n1364_), .Y(new_n3138_));
  OAI21X1  g2753(.A0(new_n3138_), .A1(new_n1362_), .B0(new_n568_), .Y(new_n3139_));
  AOI21X1  g2754(.A0(new_n3139_), .A1(new_n1360_), .B0(new_n1361_), .Y(new_n3140_));
  OAI21X1  g2755(.A0(new_n3140_), .A1(new_n1359_), .B0(new_n583_), .Y(new_n3141_));
  AOI21X1  g2756(.A0(new_n3141_), .A1(new_n1357_), .B0(new_n1358_), .Y(new_n3142_));
  OAI21X1  g2757(.A0(new_n3142_), .A1(new_n1356_), .B0(new_n598_), .Y(new_n3143_));
  AOI21X1  g2758(.A0(new_n3143_), .A1(new_n1354_), .B0(new_n1355_), .Y(new_n3144_));
  OAI21X1  g2759(.A0(new_n3144_), .A1(new_n1353_), .B0(new_n613_), .Y(new_n3145_));
  AOI21X1  g2760(.A0(new_n3145_), .A1(new_n1351_), .B0(new_n1352_), .Y(new_n3146_));
  OAI21X1  g2761(.A0(new_n3146_), .A1(new_n1350_), .B0(new_n628_), .Y(new_n3147_));
  AOI21X1  g2762(.A0(new_n3147_), .A1(new_n1348_), .B0(new_n1349_), .Y(new_n3148_));
  OAI21X1  g2763(.A0(new_n3148_), .A1(new_n1347_), .B0(new_n643_), .Y(new_n3149_));
  AOI21X1  g2764(.A0(new_n3149_), .A1(new_n1345_), .B0(new_n1346_), .Y(new_n3150_));
  OAI21X1  g2765(.A0(new_n3150_), .A1(new_n1344_), .B0(new_n658_), .Y(new_n3151_));
  AOI21X1  g2766(.A0(new_n3151_), .A1(new_n1342_), .B0(new_n1343_), .Y(new_n3152_));
  OAI21X1  g2767(.A0(new_n3152_), .A1(new_n1341_), .B0(new_n673_), .Y(new_n3153_));
  AOI21X1  g2768(.A0(new_n3153_), .A1(new_n1339_), .B0(new_n1340_), .Y(new_n3154_));
  OAI21X1  g2769(.A0(new_n3154_), .A1(new_n1338_), .B0(new_n688_), .Y(new_n3155_));
  AOI21X1  g2770(.A0(new_n3155_), .A1(new_n1336_), .B0(new_n1337_), .Y(new_n3156_));
  OAI21X1  g2771(.A0(new_n3156_), .A1(new_n1335_), .B0(new_n1438_), .Y(new_n3157_));
  AOI21X1  g2772(.A0(new_n3157_), .A1(new_n1440_), .B0(new_n1803_), .Y(new_n3158_));
  OAI21X1  g2773(.A0(new_n3158_), .A1(new_n712_), .B0(new_n714_), .Y(new_n3159_));
  AOI21X1  g2774(.A0(new_n3159_), .A1(new_n719_), .B0(new_n722_), .Y(new_n3160_));
  OAI21X1  g2775(.A0(new_n3160_), .A1(new_n727_), .B0(new_n729_), .Y(new_n3161_));
  AOI21X1  g2776(.A0(new_n3161_), .A1(new_n734_), .B0(new_n737_), .Y(new_n3162_));
  OAI21X1  g2777(.A0(new_n3162_), .A1(new_n742_), .B0(new_n744_), .Y(new_n3163_));
  AOI21X1  g2778(.A0(new_n3163_), .A1(new_n749_), .B0(new_n752_), .Y(new_n3164_));
  OAI21X1  g2779(.A0(new_n3164_), .A1(new_n757_), .B0(new_n759_), .Y(new_n3165_));
  AOI21X1  g2780(.A0(new_n3165_), .A1(new_n764_), .B0(new_n767_), .Y(new_n3166_));
  OAI21X1  g2781(.A0(new_n3166_), .A1(new_n772_), .B0(new_n774_), .Y(new_n3167_));
  AOI21X1  g2782(.A0(new_n3167_), .A1(new_n779_), .B0(new_n782_), .Y(new_n3168_));
  OAI21X1  g2783(.A0(new_n3168_), .A1(new_n787_), .B0(new_n789_), .Y(new_n3169_));
  OAI21X1  g2784(.A0(new_n1106_), .A1(\priority[39] ), .B0(\req[39] ), .Y(new_n3170_));
  AOI21X1  g2785(.A0(new_n3169_), .A1(new_n794_), .B0(new_n3170_), .Y(\grant[39] ));
  NOR2X1   g2786(.A(new_n1115_), .B(new_n803_), .Y(new_n3172_));
  OAI21X1  g2787(.A0(new_n3172_), .A1(new_n1486_), .B0(new_n811_), .Y(new_n3173_));
  AOI21X1  g2788(.A0(new_n3173_), .A1(new_n1484_), .B0(new_n1485_), .Y(new_n3174_));
  OAI21X1  g2789(.A0(new_n3174_), .A1(new_n1483_), .B0(new_n826_), .Y(new_n3175_));
  AOI21X1  g2790(.A0(new_n3175_), .A1(new_n1481_), .B0(new_n1482_), .Y(new_n3176_));
  OAI21X1  g2791(.A0(new_n3176_), .A1(new_n1480_), .B0(new_n841_), .Y(new_n3177_));
  AOI21X1  g2792(.A0(new_n3177_), .A1(new_n1478_), .B0(new_n1479_), .Y(new_n3178_));
  OAI21X1  g2793(.A0(new_n3178_), .A1(new_n1477_), .B0(new_n856_), .Y(new_n3179_));
  AOI21X1  g2794(.A0(new_n3179_), .A1(new_n1475_), .B0(new_n1476_), .Y(new_n3180_));
  OAI21X1  g2795(.A0(new_n3180_), .A1(new_n1474_), .B0(new_n871_), .Y(new_n3181_));
  AOI21X1  g2796(.A0(new_n3181_), .A1(new_n1472_), .B0(new_n1473_), .Y(new_n3182_));
  OAI21X1  g2797(.A0(new_n3182_), .A1(new_n1471_), .B0(new_n886_), .Y(new_n3183_));
  AOI21X1  g2798(.A0(new_n3183_), .A1(new_n1469_), .B0(new_n1470_), .Y(new_n3184_));
  OAI21X1  g2799(.A0(new_n3184_), .A1(new_n1468_), .B0(new_n901_), .Y(new_n3185_));
  AOI21X1  g2800(.A0(new_n3185_), .A1(new_n1466_), .B0(new_n1467_), .Y(new_n3186_));
  OAI21X1  g2801(.A0(new_n3186_), .A1(new_n1465_), .B0(new_n916_), .Y(new_n3187_));
  AOI21X1  g2802(.A0(new_n3187_), .A1(new_n1463_), .B0(new_n1464_), .Y(new_n3188_));
  OAI21X1  g2803(.A0(new_n3188_), .A1(new_n1462_), .B0(new_n931_), .Y(new_n3189_));
  AOI21X1  g2804(.A0(new_n3189_), .A1(new_n1460_), .B0(new_n1461_), .Y(new_n3190_));
  OAI21X1  g2805(.A0(new_n3190_), .A1(new_n1459_), .B0(new_n946_), .Y(new_n3191_));
  AOI21X1  g2806(.A0(new_n3191_), .A1(new_n1457_), .B0(new_n1458_), .Y(new_n3192_));
  OAI21X1  g2807(.A0(new_n3192_), .A1(new_n1456_), .B0(new_n961_), .Y(new_n3193_));
  AOI21X1  g2808(.A0(new_n3193_), .A1(new_n1454_), .B0(new_n1455_), .Y(new_n3194_));
  OAI21X1  g2809(.A0(new_n3194_), .A1(new_n1453_), .B0(new_n976_), .Y(new_n3195_));
  AOI21X1  g2810(.A0(new_n3195_), .A1(new_n1451_), .B0(new_n1452_), .Y(new_n3196_));
  OAI21X1  g2811(.A0(new_n3196_), .A1(new_n1450_), .B0(new_n991_), .Y(new_n3197_));
  AOI21X1  g2812(.A0(new_n3197_), .A1(new_n1448_), .B0(new_n1449_), .Y(new_n3198_));
  OAI21X1  g2813(.A0(new_n3198_), .A1(new_n1447_), .B0(new_n1006_), .Y(new_n3199_));
  AOI21X1  g2814(.A0(new_n3199_), .A1(new_n1445_), .B0(new_n1446_), .Y(new_n3200_));
  OAI21X1  g2815(.A0(new_n3200_), .A1(new_n1444_), .B0(new_n1547_), .Y(new_n3201_));
  AOI21X1  g2816(.A0(new_n3201_), .A1(new_n1549_), .B0(new_n1848_), .Y(new_n3202_));
  OAI21X1  g2817(.A0(new_n3202_), .A1(new_n1026_), .B0(new_n1028_), .Y(new_n3203_));
  AOI21X1  g2818(.A0(new_n3203_), .A1(new_n1033_), .B0(new_n1036_), .Y(new_n3204_));
  OAI21X1  g2819(.A0(new_n3204_), .A1(new_n1041_), .B0(new_n1043_), .Y(new_n3205_));
  AOI21X1  g2820(.A0(new_n3205_), .A1(new_n1048_), .B0(new_n1051_), .Y(new_n3206_));
  OAI21X1  g2821(.A0(new_n3206_), .A1(new_n1056_), .B0(new_n1058_), .Y(new_n3207_));
  AOI21X1  g2822(.A0(new_n3207_), .A1(new_n1063_), .B0(new_n1066_), .Y(new_n3208_));
  OAI21X1  g2823(.A0(new_n3208_), .A1(new_n1071_), .B0(new_n1073_), .Y(new_n3209_));
  AOI21X1  g2824(.A0(new_n3209_), .A1(new_n1078_), .B0(new_n1081_), .Y(new_n3210_));
  OAI21X1  g2825(.A0(new_n3210_), .A1(new_n1086_), .B0(new_n1088_), .Y(new_n3211_));
  AOI21X1  g2826(.A0(new_n3211_), .A1(new_n1093_), .B0(new_n1096_), .Y(new_n3212_));
  OAI21X1  g2827(.A0(new_n3212_), .A1(new_n1101_), .B0(new_n1103_), .Y(new_n3213_));
  OAI21X1  g2828(.A0(new_n482_), .A1(\priority[40] ), .B0(\req[40] ), .Y(new_n3214_));
  AOI21X1  g2829(.A0(new_n3213_), .A1(new_n1108_), .B0(new_n3214_), .Y(\grant[40] ));
  NOR2X1   g2830(.A(new_n1117_), .B(new_n490_), .Y(new_n3216_));
  OAI21X1  g2831(.A0(new_n3216_), .A1(new_n1595_), .B0(new_n1125_), .Y(new_n3217_));
  AOI21X1  g2832(.A0(new_n3217_), .A1(new_n1593_), .B0(new_n1594_), .Y(new_n3218_));
  OAI21X1  g2833(.A0(new_n3218_), .A1(new_n1592_), .B0(new_n1140_), .Y(new_n3219_));
  AOI21X1  g2834(.A0(new_n3219_), .A1(new_n1590_), .B0(new_n1591_), .Y(new_n3220_));
  OAI21X1  g2835(.A0(new_n3220_), .A1(new_n1589_), .B0(new_n1155_), .Y(new_n3221_));
  AOI21X1  g2836(.A0(new_n3221_), .A1(new_n1587_), .B0(new_n1588_), .Y(new_n3222_));
  OAI21X1  g2837(.A0(new_n3222_), .A1(new_n1586_), .B0(new_n1170_), .Y(new_n3223_));
  AOI21X1  g2838(.A0(new_n3223_), .A1(new_n1584_), .B0(new_n1585_), .Y(new_n3224_));
  OAI21X1  g2839(.A0(new_n3224_), .A1(new_n1583_), .B0(new_n1185_), .Y(new_n3225_));
  AOI21X1  g2840(.A0(new_n3225_), .A1(new_n1581_), .B0(new_n1582_), .Y(new_n3226_));
  OAI21X1  g2841(.A0(new_n3226_), .A1(new_n1580_), .B0(new_n1200_), .Y(new_n3227_));
  AOI21X1  g2842(.A0(new_n3227_), .A1(new_n1578_), .B0(new_n1579_), .Y(new_n3228_));
  OAI21X1  g2843(.A0(new_n3228_), .A1(new_n1577_), .B0(new_n1215_), .Y(new_n3229_));
  AOI21X1  g2844(.A0(new_n3229_), .A1(new_n1575_), .B0(new_n1576_), .Y(new_n3230_));
  OAI21X1  g2845(.A0(new_n3230_), .A1(new_n1574_), .B0(new_n1230_), .Y(new_n3231_));
  AOI21X1  g2846(.A0(new_n3231_), .A1(new_n1572_), .B0(new_n1573_), .Y(new_n3232_));
  OAI21X1  g2847(.A0(new_n3232_), .A1(new_n1571_), .B0(new_n1245_), .Y(new_n3233_));
  AOI21X1  g2848(.A0(new_n3233_), .A1(new_n1569_), .B0(new_n1570_), .Y(new_n3234_));
  OAI21X1  g2849(.A0(new_n3234_), .A1(new_n1568_), .B0(new_n1260_), .Y(new_n3235_));
  AOI21X1  g2850(.A0(new_n3235_), .A1(new_n1566_), .B0(new_n1567_), .Y(new_n3236_));
  OAI21X1  g2851(.A0(new_n3236_), .A1(new_n1565_), .B0(new_n1275_), .Y(new_n3237_));
  AOI21X1  g2852(.A0(new_n3237_), .A1(new_n1563_), .B0(new_n1564_), .Y(new_n3238_));
  OAI21X1  g2853(.A0(new_n3238_), .A1(new_n1562_), .B0(new_n1290_), .Y(new_n3239_));
  AOI21X1  g2854(.A0(new_n3239_), .A1(new_n1560_), .B0(new_n1561_), .Y(new_n3240_));
  OAI21X1  g2855(.A0(new_n3240_), .A1(new_n1559_), .B0(new_n1305_), .Y(new_n3241_));
  AOI21X1  g2856(.A0(new_n3241_), .A1(new_n1557_), .B0(new_n1558_), .Y(new_n3242_));
  OAI21X1  g2857(.A0(new_n3242_), .A1(new_n1556_), .B0(new_n1320_), .Y(new_n3243_));
  AOI21X1  g2858(.A0(new_n3243_), .A1(new_n1554_), .B0(new_n1555_), .Y(new_n3244_));
  OAI21X1  g2859(.A0(new_n3244_), .A1(new_n1553_), .B0(new_n1656_), .Y(new_n3245_));
  AOI21X1  g2860(.A0(new_n3245_), .A1(new_n1552_), .B0(new_n1893_), .Y(new_n3246_));
  OAI21X1  g2861(.A0(new_n3246_), .A1(new_n1395_), .B0(new_n403_), .Y(new_n3247_));
  AOI21X1  g2862(.A0(new_n3247_), .A1(new_n1393_), .B0(new_n1394_), .Y(new_n3248_));
  OAI21X1  g2863(.A0(new_n3248_), .A1(new_n1392_), .B0(new_n418_), .Y(new_n3249_));
  AOI21X1  g2864(.A0(new_n3249_), .A1(new_n1390_), .B0(new_n1391_), .Y(new_n3250_));
  OAI21X1  g2865(.A0(new_n3250_), .A1(new_n1389_), .B0(new_n433_), .Y(new_n3251_));
  AOI21X1  g2866(.A0(new_n3251_), .A1(new_n1387_), .B0(new_n1388_), .Y(new_n3252_));
  OAI21X1  g2867(.A0(new_n3252_), .A1(new_n1386_), .B0(new_n448_), .Y(new_n3253_));
  AOI21X1  g2868(.A0(new_n3253_), .A1(new_n1384_), .B0(new_n1385_), .Y(new_n3254_));
  OAI21X1  g2869(.A0(new_n3254_), .A1(new_n1383_), .B0(new_n463_), .Y(new_n3255_));
  AOI21X1  g2870(.A0(new_n3255_), .A1(new_n1381_), .B0(new_n1382_), .Y(new_n3256_));
  OAI21X1  g2871(.A0(new_n3256_), .A1(new_n1380_), .B0(new_n478_), .Y(new_n3257_));
  OAI21X1  g2872(.A0(new_n800_), .A1(\priority[41] ), .B0(\req[41] ), .Y(new_n3258_));
  AOI21X1  g2873(.A0(new_n3257_), .A1(new_n1378_), .B0(new_n3258_), .Y(\grant[41] ));
  NOR2X1   g2874(.A(new_n808_), .B(new_n492_), .Y(new_n3260_));
  OAI21X1  g2875(.A0(new_n3260_), .A1(new_n499_), .B0(new_n501_), .Y(new_n3261_));
  AOI21X1  g2876(.A0(new_n3261_), .A1(new_n506_), .B0(new_n509_), .Y(new_n3262_));
  OAI21X1  g2877(.A0(new_n3262_), .A1(new_n514_), .B0(new_n516_), .Y(new_n3263_));
  AOI21X1  g2878(.A0(new_n3263_), .A1(new_n521_), .B0(new_n524_), .Y(new_n3264_));
  OAI21X1  g2879(.A0(new_n3264_), .A1(new_n529_), .B0(new_n531_), .Y(new_n3265_));
  AOI21X1  g2880(.A0(new_n3265_), .A1(new_n536_), .B0(new_n539_), .Y(new_n3266_));
  OAI21X1  g2881(.A0(new_n3266_), .A1(new_n544_), .B0(new_n546_), .Y(new_n3267_));
  AOI21X1  g2882(.A0(new_n3267_), .A1(new_n551_), .B0(new_n554_), .Y(new_n3268_));
  OAI21X1  g2883(.A0(new_n3268_), .A1(new_n559_), .B0(new_n561_), .Y(new_n3269_));
  AOI21X1  g2884(.A0(new_n3269_), .A1(new_n566_), .B0(new_n569_), .Y(new_n3270_));
  OAI21X1  g2885(.A0(new_n3270_), .A1(new_n574_), .B0(new_n576_), .Y(new_n3271_));
  AOI21X1  g2886(.A0(new_n3271_), .A1(new_n581_), .B0(new_n584_), .Y(new_n3272_));
  OAI21X1  g2887(.A0(new_n3272_), .A1(new_n589_), .B0(new_n591_), .Y(new_n3273_));
  AOI21X1  g2888(.A0(new_n3273_), .A1(new_n596_), .B0(new_n599_), .Y(new_n3274_));
  OAI21X1  g2889(.A0(new_n3274_), .A1(new_n604_), .B0(new_n606_), .Y(new_n3275_));
  AOI21X1  g2890(.A0(new_n3275_), .A1(new_n611_), .B0(new_n614_), .Y(new_n3276_));
  OAI21X1  g2891(.A0(new_n3276_), .A1(new_n619_), .B0(new_n621_), .Y(new_n3277_));
  AOI21X1  g2892(.A0(new_n3277_), .A1(new_n626_), .B0(new_n629_), .Y(new_n3278_));
  OAI21X1  g2893(.A0(new_n3278_), .A1(new_n634_), .B0(new_n636_), .Y(new_n3279_));
  AOI21X1  g2894(.A0(new_n3279_), .A1(new_n641_), .B0(new_n644_), .Y(new_n3280_));
  OAI21X1  g2895(.A0(new_n3280_), .A1(new_n649_), .B0(new_n651_), .Y(new_n3281_));
  AOI21X1  g2896(.A0(new_n3281_), .A1(new_n656_), .B0(new_n659_), .Y(new_n3282_));
  OAI21X1  g2897(.A0(new_n3282_), .A1(new_n664_), .B0(new_n666_), .Y(new_n3283_));
  AOI21X1  g2898(.A0(new_n3283_), .A1(new_n671_), .B0(new_n674_), .Y(new_n3284_));
  OAI21X1  g2899(.A0(new_n3284_), .A1(new_n679_), .B0(new_n681_), .Y(new_n3285_));
  AOI21X1  g2900(.A0(new_n3285_), .A1(new_n686_), .B0(new_n689_), .Y(new_n3286_));
  OAI21X1  g2901(.A0(new_n3286_), .A1(new_n694_), .B0(new_n696_), .Y(new_n3287_));
  AOI21X1  g2902(.A0(new_n3287_), .A1(new_n701_), .B0(new_n1662_), .Y(new_n3288_));
  OAI21X1  g2903(.A0(new_n3288_), .A1(new_n1661_), .B0(new_n1705_), .Y(new_n3289_));
  AOI21X1  g2904(.A0(new_n3289_), .A1(new_n1660_), .B0(new_n1938_), .Y(new_n3290_));
  OAI21X1  g2905(.A0(new_n3290_), .A1(new_n1504_), .B0(new_n721_), .Y(new_n3291_));
  AOI21X1  g2906(.A0(new_n3291_), .A1(new_n1502_), .B0(new_n1503_), .Y(new_n3292_));
  OAI21X1  g2907(.A0(new_n3292_), .A1(new_n1501_), .B0(new_n736_), .Y(new_n3293_));
  AOI21X1  g2908(.A0(new_n3293_), .A1(new_n1499_), .B0(new_n1500_), .Y(new_n3294_));
  OAI21X1  g2909(.A0(new_n3294_), .A1(new_n1498_), .B0(new_n751_), .Y(new_n3295_));
  AOI21X1  g2910(.A0(new_n3295_), .A1(new_n1496_), .B0(new_n1497_), .Y(new_n3296_));
  OAI21X1  g2911(.A0(new_n3296_), .A1(new_n1495_), .B0(new_n766_), .Y(new_n3297_));
  AOI21X1  g2912(.A0(new_n3297_), .A1(new_n1493_), .B0(new_n1494_), .Y(new_n3298_));
  OAI21X1  g2913(.A0(new_n3298_), .A1(new_n1492_), .B0(new_n781_), .Y(new_n3299_));
  AOI21X1  g2914(.A0(new_n3299_), .A1(new_n1490_), .B0(new_n1491_), .Y(new_n3300_));
  OAI21X1  g2915(.A0(new_n3300_), .A1(new_n1489_), .B0(new_n796_), .Y(new_n3301_));
  OAI21X1  g2916(.A0(new_n1114_), .A1(\priority[42] ), .B0(\req[42] ), .Y(new_n3302_));
  AOI21X1  g2917(.A0(new_n3301_), .A1(new_n1487_), .B0(new_n3302_), .Y(\grant[42] ));
  NOR2X1   g2918(.A(new_n1122_), .B(new_n810_), .Y(new_n3304_));
  OAI21X1  g2919(.A0(new_n3304_), .A1(new_n817_), .B0(new_n819_), .Y(new_n3305_));
  AOI21X1  g2920(.A0(new_n3305_), .A1(new_n824_), .B0(new_n827_), .Y(new_n3306_));
  OAI21X1  g2921(.A0(new_n3306_), .A1(new_n832_), .B0(new_n834_), .Y(new_n3307_));
  AOI21X1  g2922(.A0(new_n3307_), .A1(new_n839_), .B0(new_n842_), .Y(new_n3308_));
  OAI21X1  g2923(.A0(new_n3308_), .A1(new_n847_), .B0(new_n849_), .Y(new_n3309_));
  AOI21X1  g2924(.A0(new_n3309_), .A1(new_n854_), .B0(new_n857_), .Y(new_n3310_));
  OAI21X1  g2925(.A0(new_n3310_), .A1(new_n862_), .B0(new_n864_), .Y(new_n3311_));
  AOI21X1  g2926(.A0(new_n3311_), .A1(new_n869_), .B0(new_n872_), .Y(new_n3312_));
  OAI21X1  g2927(.A0(new_n3312_), .A1(new_n877_), .B0(new_n879_), .Y(new_n3313_));
  AOI21X1  g2928(.A0(new_n3313_), .A1(new_n884_), .B0(new_n887_), .Y(new_n3314_));
  OAI21X1  g2929(.A0(new_n3314_), .A1(new_n892_), .B0(new_n894_), .Y(new_n3315_));
  AOI21X1  g2930(.A0(new_n3315_), .A1(new_n899_), .B0(new_n902_), .Y(new_n3316_));
  OAI21X1  g2931(.A0(new_n3316_), .A1(new_n907_), .B0(new_n909_), .Y(new_n3317_));
  AOI21X1  g2932(.A0(new_n3317_), .A1(new_n914_), .B0(new_n917_), .Y(new_n3318_));
  OAI21X1  g2933(.A0(new_n3318_), .A1(new_n922_), .B0(new_n924_), .Y(new_n3319_));
  AOI21X1  g2934(.A0(new_n3319_), .A1(new_n929_), .B0(new_n932_), .Y(new_n3320_));
  OAI21X1  g2935(.A0(new_n3320_), .A1(new_n937_), .B0(new_n939_), .Y(new_n3321_));
  AOI21X1  g2936(.A0(new_n3321_), .A1(new_n944_), .B0(new_n947_), .Y(new_n3322_));
  OAI21X1  g2937(.A0(new_n3322_), .A1(new_n952_), .B0(new_n954_), .Y(new_n3323_));
  AOI21X1  g2938(.A0(new_n3323_), .A1(new_n959_), .B0(new_n962_), .Y(new_n3324_));
  OAI21X1  g2939(.A0(new_n3324_), .A1(new_n967_), .B0(new_n969_), .Y(new_n3325_));
  AOI21X1  g2940(.A0(new_n3325_), .A1(new_n974_), .B0(new_n977_), .Y(new_n3326_));
  OAI21X1  g2941(.A0(new_n3326_), .A1(new_n982_), .B0(new_n984_), .Y(new_n3327_));
  AOI21X1  g2942(.A0(new_n3327_), .A1(new_n989_), .B0(new_n992_), .Y(new_n3328_));
  OAI21X1  g2943(.A0(new_n3328_), .A1(new_n997_), .B0(new_n999_), .Y(new_n3329_));
  AOI21X1  g2944(.A0(new_n3329_), .A1(new_n1004_), .B0(new_n1007_), .Y(new_n3330_));
  OAI21X1  g2945(.A0(new_n3330_), .A1(new_n1012_), .B0(new_n1014_), .Y(new_n3331_));
  AOI21X1  g2946(.A0(new_n3331_), .A1(new_n1017_), .B0(new_n1711_), .Y(new_n3332_));
  OAI21X1  g2947(.A0(new_n3332_), .A1(new_n1710_), .B0(new_n1754_), .Y(new_n3333_));
  AOI21X1  g2948(.A0(new_n3333_), .A1(new_n1709_), .B0(new_n1983_), .Y(new_n3334_));
  OAI21X1  g2949(.A0(new_n3334_), .A1(new_n1613_), .B0(new_n1035_), .Y(new_n3335_));
  AOI21X1  g2950(.A0(new_n3335_), .A1(new_n1611_), .B0(new_n1612_), .Y(new_n3336_));
  OAI21X1  g2951(.A0(new_n3336_), .A1(new_n1610_), .B0(new_n1050_), .Y(new_n3337_));
  AOI21X1  g2952(.A0(new_n3337_), .A1(new_n1608_), .B0(new_n1609_), .Y(new_n3338_));
  OAI21X1  g2953(.A0(new_n3338_), .A1(new_n1607_), .B0(new_n1065_), .Y(new_n3339_));
  AOI21X1  g2954(.A0(new_n3339_), .A1(new_n1605_), .B0(new_n1606_), .Y(new_n3340_));
  OAI21X1  g2955(.A0(new_n3340_), .A1(new_n1604_), .B0(new_n1080_), .Y(new_n3341_));
  AOI21X1  g2956(.A0(new_n3341_), .A1(new_n1602_), .B0(new_n1603_), .Y(new_n3342_));
  OAI21X1  g2957(.A0(new_n3342_), .A1(new_n1601_), .B0(new_n1095_), .Y(new_n3343_));
  AOI21X1  g2958(.A0(new_n3343_), .A1(new_n1599_), .B0(new_n1600_), .Y(new_n3344_));
  OAI21X1  g2959(.A0(new_n3344_), .A1(new_n1598_), .B0(new_n1110_), .Y(new_n3345_));
  OAI21X1  g2960(.A0(new_n489_), .A1(\priority[43] ), .B0(\req[43] ), .Y(new_n3346_));
  AOI21X1  g2961(.A0(new_n3345_), .A1(new_n1596_), .B0(new_n3346_), .Y(\grant[43] ));
  NOR2X1   g2962(.A(new_n1124_), .B(new_n498_), .Y(new_n3348_));
  OAI21X1  g2963(.A0(new_n3348_), .A1(new_n1131_), .B0(new_n1133_), .Y(new_n3349_));
  AOI21X1  g2964(.A0(new_n3349_), .A1(new_n1138_), .B0(new_n1141_), .Y(new_n3350_));
  OAI21X1  g2965(.A0(new_n3350_), .A1(new_n1146_), .B0(new_n1148_), .Y(new_n3351_));
  AOI21X1  g2966(.A0(new_n3351_), .A1(new_n1153_), .B0(new_n1156_), .Y(new_n3352_));
  OAI21X1  g2967(.A0(new_n3352_), .A1(new_n1161_), .B0(new_n1163_), .Y(new_n3353_));
  AOI21X1  g2968(.A0(new_n3353_), .A1(new_n1168_), .B0(new_n1171_), .Y(new_n3354_));
  OAI21X1  g2969(.A0(new_n3354_), .A1(new_n1176_), .B0(new_n1178_), .Y(new_n3355_));
  AOI21X1  g2970(.A0(new_n3355_), .A1(new_n1183_), .B0(new_n1186_), .Y(new_n3356_));
  OAI21X1  g2971(.A0(new_n3356_), .A1(new_n1191_), .B0(new_n1193_), .Y(new_n3357_));
  AOI21X1  g2972(.A0(new_n3357_), .A1(new_n1198_), .B0(new_n1201_), .Y(new_n3358_));
  OAI21X1  g2973(.A0(new_n3358_), .A1(new_n1206_), .B0(new_n1208_), .Y(new_n3359_));
  AOI21X1  g2974(.A0(new_n3359_), .A1(new_n1213_), .B0(new_n1216_), .Y(new_n3360_));
  OAI21X1  g2975(.A0(new_n3360_), .A1(new_n1221_), .B0(new_n1223_), .Y(new_n3361_));
  AOI21X1  g2976(.A0(new_n3361_), .A1(new_n1228_), .B0(new_n1231_), .Y(new_n3362_));
  OAI21X1  g2977(.A0(new_n3362_), .A1(new_n1236_), .B0(new_n1238_), .Y(new_n3363_));
  AOI21X1  g2978(.A0(new_n3363_), .A1(new_n1243_), .B0(new_n1246_), .Y(new_n3364_));
  OAI21X1  g2979(.A0(new_n3364_), .A1(new_n1251_), .B0(new_n1253_), .Y(new_n3365_));
  AOI21X1  g2980(.A0(new_n3365_), .A1(new_n1258_), .B0(new_n1261_), .Y(new_n3366_));
  OAI21X1  g2981(.A0(new_n3366_), .A1(new_n1266_), .B0(new_n1268_), .Y(new_n3367_));
  AOI21X1  g2982(.A0(new_n3367_), .A1(new_n1273_), .B0(new_n1276_), .Y(new_n3368_));
  OAI21X1  g2983(.A0(new_n3368_), .A1(new_n1281_), .B0(new_n1283_), .Y(new_n3369_));
  AOI21X1  g2984(.A0(new_n3369_), .A1(new_n1288_), .B0(new_n1291_), .Y(new_n3370_));
  OAI21X1  g2985(.A0(new_n3370_), .A1(new_n1296_), .B0(new_n1298_), .Y(new_n3371_));
  AOI21X1  g2986(.A0(new_n3371_), .A1(new_n1303_), .B0(new_n1306_), .Y(new_n3372_));
  OAI21X1  g2987(.A0(new_n3372_), .A1(new_n1311_), .B0(new_n1313_), .Y(new_n3373_));
  AOI21X1  g2988(.A0(new_n3373_), .A1(new_n1318_), .B0(new_n1321_), .Y(new_n3374_));
  OAI21X1  g2989(.A0(new_n3374_), .A1(new_n1326_), .B0(new_n1328_), .Y(new_n3375_));
  AOI21X1  g2990(.A0(new_n3375_), .A1(new_n1331_), .B0(new_n1758_), .Y(new_n3376_));
  OAI21X1  g2991(.A0(new_n3376_), .A1(new_n394_), .B0(new_n396_), .Y(new_n3377_));
  AOI21X1  g2992(.A0(new_n3377_), .A1(new_n401_), .B0(new_n404_), .Y(new_n3378_));
  OAI21X1  g2993(.A0(new_n3378_), .A1(new_n409_), .B0(new_n411_), .Y(new_n3379_));
  AOI21X1  g2994(.A0(new_n3379_), .A1(new_n416_), .B0(new_n419_), .Y(new_n3380_));
  OAI21X1  g2995(.A0(new_n3380_), .A1(new_n424_), .B0(new_n426_), .Y(new_n3381_));
  AOI21X1  g2996(.A0(new_n3381_), .A1(new_n431_), .B0(new_n434_), .Y(new_n3382_));
  OAI21X1  g2997(.A0(new_n3382_), .A1(new_n439_), .B0(new_n441_), .Y(new_n3383_));
  AOI21X1  g2998(.A0(new_n3383_), .A1(new_n446_), .B0(new_n449_), .Y(new_n3384_));
  OAI21X1  g2999(.A0(new_n3384_), .A1(new_n454_), .B0(new_n456_), .Y(new_n3385_));
  AOI21X1  g3000(.A0(new_n3385_), .A1(new_n461_), .B0(new_n464_), .Y(new_n3386_));
  OAI21X1  g3001(.A0(new_n3386_), .A1(new_n469_), .B0(new_n471_), .Y(new_n3387_));
  AOI21X1  g3002(.A0(new_n3387_), .A1(new_n476_), .B0(new_n479_), .Y(new_n3388_));
  OAI21X1  g3003(.A0(new_n3388_), .A1(new_n484_), .B0(new_n486_), .Y(new_n3389_));
  OAI21X1  g3004(.A0(new_n807_), .A1(\priority[44] ), .B0(\req[44] ), .Y(new_n3390_));
  AOI21X1  g3005(.A0(new_n3389_), .A1(new_n491_), .B0(new_n3390_), .Y(\grant[44] ));
  NOR2X1   g3006(.A(new_n816_), .B(new_n500_), .Y(new_n3392_));
  OAI21X1  g3007(.A0(new_n3392_), .A1(new_n1374_), .B0(new_n508_), .Y(new_n3393_));
  AOI21X1  g3008(.A0(new_n3393_), .A1(new_n1372_), .B0(new_n1373_), .Y(new_n3394_));
  OAI21X1  g3009(.A0(new_n3394_), .A1(new_n1371_), .B0(new_n523_), .Y(new_n3395_));
  AOI21X1  g3010(.A0(new_n3395_), .A1(new_n1369_), .B0(new_n1370_), .Y(new_n3396_));
  OAI21X1  g3011(.A0(new_n3396_), .A1(new_n1368_), .B0(new_n538_), .Y(new_n3397_));
  AOI21X1  g3012(.A0(new_n3397_), .A1(new_n1366_), .B0(new_n1367_), .Y(new_n3398_));
  OAI21X1  g3013(.A0(new_n3398_), .A1(new_n1365_), .B0(new_n553_), .Y(new_n3399_));
  AOI21X1  g3014(.A0(new_n3399_), .A1(new_n1363_), .B0(new_n1364_), .Y(new_n3400_));
  OAI21X1  g3015(.A0(new_n3400_), .A1(new_n1362_), .B0(new_n568_), .Y(new_n3401_));
  AOI21X1  g3016(.A0(new_n3401_), .A1(new_n1360_), .B0(new_n1361_), .Y(new_n3402_));
  OAI21X1  g3017(.A0(new_n3402_), .A1(new_n1359_), .B0(new_n583_), .Y(new_n3403_));
  AOI21X1  g3018(.A0(new_n3403_), .A1(new_n1357_), .B0(new_n1358_), .Y(new_n3404_));
  OAI21X1  g3019(.A0(new_n3404_), .A1(new_n1356_), .B0(new_n598_), .Y(new_n3405_));
  AOI21X1  g3020(.A0(new_n3405_), .A1(new_n1354_), .B0(new_n1355_), .Y(new_n3406_));
  OAI21X1  g3021(.A0(new_n3406_), .A1(new_n1353_), .B0(new_n613_), .Y(new_n3407_));
  AOI21X1  g3022(.A0(new_n3407_), .A1(new_n1351_), .B0(new_n1352_), .Y(new_n3408_));
  OAI21X1  g3023(.A0(new_n3408_), .A1(new_n1350_), .B0(new_n628_), .Y(new_n3409_));
  AOI21X1  g3024(.A0(new_n3409_), .A1(new_n1348_), .B0(new_n1349_), .Y(new_n3410_));
  OAI21X1  g3025(.A0(new_n3410_), .A1(new_n1347_), .B0(new_n643_), .Y(new_n3411_));
  AOI21X1  g3026(.A0(new_n3411_), .A1(new_n1345_), .B0(new_n1346_), .Y(new_n3412_));
  OAI21X1  g3027(.A0(new_n3412_), .A1(new_n1344_), .B0(new_n658_), .Y(new_n3413_));
  AOI21X1  g3028(.A0(new_n3413_), .A1(new_n1342_), .B0(new_n1343_), .Y(new_n3414_));
  OAI21X1  g3029(.A0(new_n3414_), .A1(new_n1341_), .B0(new_n673_), .Y(new_n3415_));
  AOI21X1  g3030(.A0(new_n3415_), .A1(new_n1339_), .B0(new_n1340_), .Y(new_n3416_));
  OAI21X1  g3031(.A0(new_n3416_), .A1(new_n1338_), .B0(new_n688_), .Y(new_n3417_));
  AOI21X1  g3032(.A0(new_n3417_), .A1(new_n1336_), .B0(new_n1337_), .Y(new_n3418_));
  OAI21X1  g3033(.A0(new_n3418_), .A1(new_n1335_), .B0(new_n1438_), .Y(new_n3419_));
  AOI21X1  g3034(.A0(new_n3419_), .A1(new_n1440_), .B0(new_n1803_), .Y(new_n3420_));
  OAI21X1  g3035(.A0(new_n3420_), .A1(new_n712_), .B0(new_n714_), .Y(new_n3421_));
  AOI21X1  g3036(.A0(new_n3421_), .A1(new_n719_), .B0(new_n722_), .Y(new_n3422_));
  OAI21X1  g3037(.A0(new_n3422_), .A1(new_n727_), .B0(new_n729_), .Y(new_n3423_));
  AOI21X1  g3038(.A0(new_n3423_), .A1(new_n734_), .B0(new_n737_), .Y(new_n3424_));
  OAI21X1  g3039(.A0(new_n3424_), .A1(new_n742_), .B0(new_n744_), .Y(new_n3425_));
  AOI21X1  g3040(.A0(new_n3425_), .A1(new_n749_), .B0(new_n752_), .Y(new_n3426_));
  OAI21X1  g3041(.A0(new_n3426_), .A1(new_n757_), .B0(new_n759_), .Y(new_n3427_));
  AOI21X1  g3042(.A0(new_n3427_), .A1(new_n764_), .B0(new_n767_), .Y(new_n3428_));
  OAI21X1  g3043(.A0(new_n3428_), .A1(new_n772_), .B0(new_n774_), .Y(new_n3429_));
  AOI21X1  g3044(.A0(new_n3429_), .A1(new_n779_), .B0(new_n782_), .Y(new_n3430_));
  OAI21X1  g3045(.A0(new_n3430_), .A1(new_n787_), .B0(new_n789_), .Y(new_n3431_));
  AOI21X1  g3046(.A0(new_n3431_), .A1(new_n794_), .B0(new_n797_), .Y(new_n3432_));
  OAI21X1  g3047(.A0(new_n3432_), .A1(new_n802_), .B0(new_n804_), .Y(new_n3433_));
  OAI21X1  g3048(.A0(new_n1121_), .A1(\priority[45] ), .B0(\req[45] ), .Y(new_n3434_));
  AOI21X1  g3049(.A0(new_n3433_), .A1(new_n809_), .B0(new_n3434_), .Y(\grant[45] ));
  NOR2X1   g3050(.A(new_n1130_), .B(new_n818_), .Y(new_n3436_));
  OAI21X1  g3051(.A0(new_n3436_), .A1(new_n1483_), .B0(new_n826_), .Y(new_n3437_));
  AOI21X1  g3052(.A0(new_n3437_), .A1(new_n1481_), .B0(new_n1482_), .Y(new_n3438_));
  OAI21X1  g3053(.A0(new_n3438_), .A1(new_n1480_), .B0(new_n841_), .Y(new_n3439_));
  AOI21X1  g3054(.A0(new_n3439_), .A1(new_n1478_), .B0(new_n1479_), .Y(new_n3440_));
  OAI21X1  g3055(.A0(new_n3440_), .A1(new_n1477_), .B0(new_n856_), .Y(new_n3441_));
  AOI21X1  g3056(.A0(new_n3441_), .A1(new_n1475_), .B0(new_n1476_), .Y(new_n3442_));
  OAI21X1  g3057(.A0(new_n3442_), .A1(new_n1474_), .B0(new_n871_), .Y(new_n3443_));
  AOI21X1  g3058(.A0(new_n3443_), .A1(new_n1472_), .B0(new_n1473_), .Y(new_n3444_));
  OAI21X1  g3059(.A0(new_n3444_), .A1(new_n1471_), .B0(new_n886_), .Y(new_n3445_));
  AOI21X1  g3060(.A0(new_n3445_), .A1(new_n1469_), .B0(new_n1470_), .Y(new_n3446_));
  OAI21X1  g3061(.A0(new_n3446_), .A1(new_n1468_), .B0(new_n901_), .Y(new_n3447_));
  AOI21X1  g3062(.A0(new_n3447_), .A1(new_n1466_), .B0(new_n1467_), .Y(new_n3448_));
  OAI21X1  g3063(.A0(new_n3448_), .A1(new_n1465_), .B0(new_n916_), .Y(new_n3449_));
  AOI21X1  g3064(.A0(new_n3449_), .A1(new_n1463_), .B0(new_n1464_), .Y(new_n3450_));
  OAI21X1  g3065(.A0(new_n3450_), .A1(new_n1462_), .B0(new_n931_), .Y(new_n3451_));
  AOI21X1  g3066(.A0(new_n3451_), .A1(new_n1460_), .B0(new_n1461_), .Y(new_n3452_));
  OAI21X1  g3067(.A0(new_n3452_), .A1(new_n1459_), .B0(new_n946_), .Y(new_n3453_));
  AOI21X1  g3068(.A0(new_n3453_), .A1(new_n1457_), .B0(new_n1458_), .Y(new_n3454_));
  OAI21X1  g3069(.A0(new_n3454_), .A1(new_n1456_), .B0(new_n961_), .Y(new_n3455_));
  AOI21X1  g3070(.A0(new_n3455_), .A1(new_n1454_), .B0(new_n1455_), .Y(new_n3456_));
  OAI21X1  g3071(.A0(new_n3456_), .A1(new_n1453_), .B0(new_n976_), .Y(new_n3457_));
  AOI21X1  g3072(.A0(new_n3457_), .A1(new_n1451_), .B0(new_n1452_), .Y(new_n3458_));
  OAI21X1  g3073(.A0(new_n3458_), .A1(new_n1450_), .B0(new_n991_), .Y(new_n3459_));
  AOI21X1  g3074(.A0(new_n3459_), .A1(new_n1448_), .B0(new_n1449_), .Y(new_n3460_));
  OAI21X1  g3075(.A0(new_n3460_), .A1(new_n1447_), .B0(new_n1006_), .Y(new_n3461_));
  AOI21X1  g3076(.A0(new_n3461_), .A1(new_n1445_), .B0(new_n1446_), .Y(new_n3462_));
  OAI21X1  g3077(.A0(new_n3462_), .A1(new_n1444_), .B0(new_n1547_), .Y(new_n3463_));
  AOI21X1  g3078(.A0(new_n3463_), .A1(new_n1549_), .B0(new_n1848_), .Y(new_n3464_));
  OAI21X1  g3079(.A0(new_n3464_), .A1(new_n1026_), .B0(new_n1028_), .Y(new_n3465_));
  AOI21X1  g3080(.A0(new_n3465_), .A1(new_n1033_), .B0(new_n1036_), .Y(new_n3466_));
  OAI21X1  g3081(.A0(new_n3466_), .A1(new_n1041_), .B0(new_n1043_), .Y(new_n3467_));
  AOI21X1  g3082(.A0(new_n3467_), .A1(new_n1048_), .B0(new_n1051_), .Y(new_n3468_));
  OAI21X1  g3083(.A0(new_n3468_), .A1(new_n1056_), .B0(new_n1058_), .Y(new_n3469_));
  AOI21X1  g3084(.A0(new_n3469_), .A1(new_n1063_), .B0(new_n1066_), .Y(new_n3470_));
  OAI21X1  g3085(.A0(new_n3470_), .A1(new_n1071_), .B0(new_n1073_), .Y(new_n3471_));
  AOI21X1  g3086(.A0(new_n3471_), .A1(new_n1078_), .B0(new_n1081_), .Y(new_n3472_));
  OAI21X1  g3087(.A0(new_n3472_), .A1(new_n1086_), .B0(new_n1088_), .Y(new_n3473_));
  AOI21X1  g3088(.A0(new_n3473_), .A1(new_n1093_), .B0(new_n1096_), .Y(new_n3474_));
  OAI21X1  g3089(.A0(new_n3474_), .A1(new_n1101_), .B0(new_n1103_), .Y(new_n3475_));
  AOI21X1  g3090(.A0(new_n3475_), .A1(new_n1108_), .B0(new_n1111_), .Y(new_n3476_));
  OAI21X1  g3091(.A0(new_n3476_), .A1(new_n1116_), .B0(new_n1118_), .Y(new_n3477_));
  OAI21X1  g3092(.A0(new_n497_), .A1(\priority[46] ), .B0(\req[46] ), .Y(new_n3478_));
  AOI21X1  g3093(.A0(new_n3477_), .A1(new_n1123_), .B0(new_n3478_), .Y(\grant[46] ));
  NOR2X1   g3094(.A(new_n1132_), .B(new_n505_), .Y(new_n3480_));
  OAI21X1  g3095(.A0(new_n3480_), .A1(new_n1592_), .B0(new_n1140_), .Y(new_n3481_));
  AOI21X1  g3096(.A0(new_n3481_), .A1(new_n1590_), .B0(new_n1591_), .Y(new_n3482_));
  OAI21X1  g3097(.A0(new_n3482_), .A1(new_n1589_), .B0(new_n1155_), .Y(new_n3483_));
  AOI21X1  g3098(.A0(new_n3483_), .A1(new_n1587_), .B0(new_n1588_), .Y(new_n3484_));
  OAI21X1  g3099(.A0(new_n3484_), .A1(new_n1586_), .B0(new_n1170_), .Y(new_n3485_));
  AOI21X1  g3100(.A0(new_n3485_), .A1(new_n1584_), .B0(new_n1585_), .Y(new_n3486_));
  OAI21X1  g3101(.A0(new_n3486_), .A1(new_n1583_), .B0(new_n1185_), .Y(new_n3487_));
  AOI21X1  g3102(.A0(new_n3487_), .A1(new_n1581_), .B0(new_n1582_), .Y(new_n3488_));
  OAI21X1  g3103(.A0(new_n3488_), .A1(new_n1580_), .B0(new_n1200_), .Y(new_n3489_));
  AOI21X1  g3104(.A0(new_n3489_), .A1(new_n1578_), .B0(new_n1579_), .Y(new_n3490_));
  OAI21X1  g3105(.A0(new_n3490_), .A1(new_n1577_), .B0(new_n1215_), .Y(new_n3491_));
  AOI21X1  g3106(.A0(new_n3491_), .A1(new_n1575_), .B0(new_n1576_), .Y(new_n3492_));
  OAI21X1  g3107(.A0(new_n3492_), .A1(new_n1574_), .B0(new_n1230_), .Y(new_n3493_));
  AOI21X1  g3108(.A0(new_n3493_), .A1(new_n1572_), .B0(new_n1573_), .Y(new_n3494_));
  OAI21X1  g3109(.A0(new_n3494_), .A1(new_n1571_), .B0(new_n1245_), .Y(new_n3495_));
  AOI21X1  g3110(.A0(new_n3495_), .A1(new_n1569_), .B0(new_n1570_), .Y(new_n3496_));
  OAI21X1  g3111(.A0(new_n3496_), .A1(new_n1568_), .B0(new_n1260_), .Y(new_n3497_));
  AOI21X1  g3112(.A0(new_n3497_), .A1(new_n1566_), .B0(new_n1567_), .Y(new_n3498_));
  OAI21X1  g3113(.A0(new_n3498_), .A1(new_n1565_), .B0(new_n1275_), .Y(new_n3499_));
  AOI21X1  g3114(.A0(new_n3499_), .A1(new_n1563_), .B0(new_n1564_), .Y(new_n3500_));
  OAI21X1  g3115(.A0(new_n3500_), .A1(new_n1562_), .B0(new_n1290_), .Y(new_n3501_));
  AOI21X1  g3116(.A0(new_n3501_), .A1(new_n1560_), .B0(new_n1561_), .Y(new_n3502_));
  OAI21X1  g3117(.A0(new_n3502_), .A1(new_n1559_), .B0(new_n1305_), .Y(new_n3503_));
  AOI21X1  g3118(.A0(new_n3503_), .A1(new_n1557_), .B0(new_n1558_), .Y(new_n3504_));
  OAI21X1  g3119(.A0(new_n3504_), .A1(new_n1556_), .B0(new_n1320_), .Y(new_n3505_));
  AOI21X1  g3120(.A0(new_n3505_), .A1(new_n1554_), .B0(new_n1555_), .Y(new_n3506_));
  OAI21X1  g3121(.A0(new_n3506_), .A1(new_n1553_), .B0(new_n1656_), .Y(new_n3507_));
  AOI21X1  g3122(.A0(new_n3507_), .A1(new_n1552_), .B0(new_n1893_), .Y(new_n3508_));
  OAI21X1  g3123(.A0(new_n3508_), .A1(new_n1395_), .B0(new_n403_), .Y(new_n3509_));
  AOI21X1  g3124(.A0(new_n3509_), .A1(new_n1393_), .B0(new_n1394_), .Y(new_n3510_));
  OAI21X1  g3125(.A0(new_n3510_), .A1(new_n1392_), .B0(new_n418_), .Y(new_n3511_));
  AOI21X1  g3126(.A0(new_n3511_), .A1(new_n1390_), .B0(new_n1391_), .Y(new_n3512_));
  OAI21X1  g3127(.A0(new_n3512_), .A1(new_n1389_), .B0(new_n433_), .Y(new_n3513_));
  AOI21X1  g3128(.A0(new_n3513_), .A1(new_n1387_), .B0(new_n1388_), .Y(new_n3514_));
  OAI21X1  g3129(.A0(new_n3514_), .A1(new_n1386_), .B0(new_n448_), .Y(new_n3515_));
  AOI21X1  g3130(.A0(new_n3515_), .A1(new_n1384_), .B0(new_n1385_), .Y(new_n3516_));
  OAI21X1  g3131(.A0(new_n3516_), .A1(new_n1383_), .B0(new_n463_), .Y(new_n3517_));
  AOI21X1  g3132(.A0(new_n3517_), .A1(new_n1381_), .B0(new_n1382_), .Y(new_n3518_));
  OAI21X1  g3133(.A0(new_n3518_), .A1(new_n1380_), .B0(new_n478_), .Y(new_n3519_));
  AOI21X1  g3134(.A0(new_n3519_), .A1(new_n1378_), .B0(new_n1379_), .Y(new_n3520_));
  OAI21X1  g3135(.A0(new_n3520_), .A1(new_n1377_), .B0(new_n493_), .Y(new_n3521_));
  OAI21X1  g3136(.A0(new_n815_), .A1(\priority[47] ), .B0(\req[47] ), .Y(new_n3522_));
  AOI21X1  g3137(.A0(new_n3521_), .A1(new_n1375_), .B0(new_n3522_), .Y(\grant[47] ));
  NOR2X1   g3138(.A(new_n823_), .B(new_n507_), .Y(new_n3524_));
  OAI21X1  g3139(.A0(new_n3524_), .A1(new_n514_), .B0(new_n516_), .Y(new_n3525_));
  AOI21X1  g3140(.A0(new_n3525_), .A1(new_n521_), .B0(new_n524_), .Y(new_n3526_));
  OAI21X1  g3141(.A0(new_n3526_), .A1(new_n529_), .B0(new_n531_), .Y(new_n3527_));
  AOI21X1  g3142(.A0(new_n3527_), .A1(new_n536_), .B0(new_n539_), .Y(new_n3528_));
  OAI21X1  g3143(.A0(new_n3528_), .A1(new_n544_), .B0(new_n546_), .Y(new_n3529_));
  AOI21X1  g3144(.A0(new_n3529_), .A1(new_n551_), .B0(new_n554_), .Y(new_n3530_));
  OAI21X1  g3145(.A0(new_n3530_), .A1(new_n559_), .B0(new_n561_), .Y(new_n3531_));
  AOI21X1  g3146(.A0(new_n3531_), .A1(new_n566_), .B0(new_n569_), .Y(new_n3532_));
  OAI21X1  g3147(.A0(new_n3532_), .A1(new_n574_), .B0(new_n576_), .Y(new_n3533_));
  AOI21X1  g3148(.A0(new_n3533_), .A1(new_n581_), .B0(new_n584_), .Y(new_n3534_));
  OAI21X1  g3149(.A0(new_n3534_), .A1(new_n589_), .B0(new_n591_), .Y(new_n3535_));
  AOI21X1  g3150(.A0(new_n3535_), .A1(new_n596_), .B0(new_n599_), .Y(new_n3536_));
  OAI21X1  g3151(.A0(new_n3536_), .A1(new_n604_), .B0(new_n606_), .Y(new_n3537_));
  AOI21X1  g3152(.A0(new_n3537_), .A1(new_n611_), .B0(new_n614_), .Y(new_n3538_));
  OAI21X1  g3153(.A0(new_n3538_), .A1(new_n619_), .B0(new_n621_), .Y(new_n3539_));
  AOI21X1  g3154(.A0(new_n3539_), .A1(new_n626_), .B0(new_n629_), .Y(new_n3540_));
  OAI21X1  g3155(.A0(new_n3540_), .A1(new_n634_), .B0(new_n636_), .Y(new_n3541_));
  AOI21X1  g3156(.A0(new_n3541_), .A1(new_n641_), .B0(new_n644_), .Y(new_n3542_));
  OAI21X1  g3157(.A0(new_n3542_), .A1(new_n649_), .B0(new_n651_), .Y(new_n3543_));
  AOI21X1  g3158(.A0(new_n3543_), .A1(new_n656_), .B0(new_n659_), .Y(new_n3544_));
  OAI21X1  g3159(.A0(new_n3544_), .A1(new_n664_), .B0(new_n666_), .Y(new_n3545_));
  AOI21X1  g3160(.A0(new_n3545_), .A1(new_n671_), .B0(new_n674_), .Y(new_n3546_));
  OAI21X1  g3161(.A0(new_n3546_), .A1(new_n679_), .B0(new_n681_), .Y(new_n3547_));
  AOI21X1  g3162(.A0(new_n3547_), .A1(new_n686_), .B0(new_n689_), .Y(new_n3548_));
  OAI21X1  g3163(.A0(new_n3548_), .A1(new_n694_), .B0(new_n696_), .Y(new_n3549_));
  AOI21X1  g3164(.A0(new_n3549_), .A1(new_n701_), .B0(new_n1662_), .Y(new_n3550_));
  OAI21X1  g3165(.A0(new_n3550_), .A1(new_n1661_), .B0(new_n1705_), .Y(new_n3551_));
  AOI21X1  g3166(.A0(new_n3551_), .A1(new_n1660_), .B0(new_n1938_), .Y(new_n3552_));
  OAI21X1  g3167(.A0(new_n3552_), .A1(new_n1504_), .B0(new_n721_), .Y(new_n3553_));
  AOI21X1  g3168(.A0(new_n3553_), .A1(new_n1502_), .B0(new_n1503_), .Y(new_n3554_));
  OAI21X1  g3169(.A0(new_n3554_), .A1(new_n1501_), .B0(new_n736_), .Y(new_n3555_));
  AOI21X1  g3170(.A0(new_n3555_), .A1(new_n1499_), .B0(new_n1500_), .Y(new_n3556_));
  OAI21X1  g3171(.A0(new_n3556_), .A1(new_n1498_), .B0(new_n751_), .Y(new_n3557_));
  AOI21X1  g3172(.A0(new_n3557_), .A1(new_n1496_), .B0(new_n1497_), .Y(new_n3558_));
  OAI21X1  g3173(.A0(new_n3558_), .A1(new_n1495_), .B0(new_n766_), .Y(new_n3559_));
  AOI21X1  g3174(.A0(new_n3559_), .A1(new_n1493_), .B0(new_n1494_), .Y(new_n3560_));
  OAI21X1  g3175(.A0(new_n3560_), .A1(new_n1492_), .B0(new_n781_), .Y(new_n3561_));
  AOI21X1  g3176(.A0(new_n3561_), .A1(new_n1490_), .B0(new_n1491_), .Y(new_n3562_));
  OAI21X1  g3177(.A0(new_n3562_), .A1(new_n1489_), .B0(new_n796_), .Y(new_n3563_));
  AOI21X1  g3178(.A0(new_n3563_), .A1(new_n1487_), .B0(new_n1488_), .Y(new_n3564_));
  OAI21X1  g3179(.A0(new_n3564_), .A1(new_n1486_), .B0(new_n811_), .Y(new_n3565_));
  OAI21X1  g3180(.A0(new_n1129_), .A1(\priority[48] ), .B0(\req[48] ), .Y(new_n3566_));
  AOI21X1  g3181(.A0(new_n3565_), .A1(new_n1484_), .B0(new_n3566_), .Y(\grant[48] ));
  NOR2X1   g3182(.A(new_n1137_), .B(new_n825_), .Y(new_n3568_));
  OAI21X1  g3183(.A0(new_n3568_), .A1(new_n832_), .B0(new_n834_), .Y(new_n3569_));
  AOI21X1  g3184(.A0(new_n3569_), .A1(new_n839_), .B0(new_n842_), .Y(new_n3570_));
  OAI21X1  g3185(.A0(new_n3570_), .A1(new_n847_), .B0(new_n849_), .Y(new_n3571_));
  AOI21X1  g3186(.A0(new_n3571_), .A1(new_n854_), .B0(new_n857_), .Y(new_n3572_));
  OAI21X1  g3187(.A0(new_n3572_), .A1(new_n862_), .B0(new_n864_), .Y(new_n3573_));
  AOI21X1  g3188(.A0(new_n3573_), .A1(new_n869_), .B0(new_n872_), .Y(new_n3574_));
  OAI21X1  g3189(.A0(new_n3574_), .A1(new_n877_), .B0(new_n879_), .Y(new_n3575_));
  AOI21X1  g3190(.A0(new_n3575_), .A1(new_n884_), .B0(new_n887_), .Y(new_n3576_));
  OAI21X1  g3191(.A0(new_n3576_), .A1(new_n892_), .B0(new_n894_), .Y(new_n3577_));
  AOI21X1  g3192(.A0(new_n3577_), .A1(new_n899_), .B0(new_n902_), .Y(new_n3578_));
  OAI21X1  g3193(.A0(new_n3578_), .A1(new_n907_), .B0(new_n909_), .Y(new_n3579_));
  AOI21X1  g3194(.A0(new_n3579_), .A1(new_n914_), .B0(new_n917_), .Y(new_n3580_));
  OAI21X1  g3195(.A0(new_n3580_), .A1(new_n922_), .B0(new_n924_), .Y(new_n3581_));
  AOI21X1  g3196(.A0(new_n3581_), .A1(new_n929_), .B0(new_n932_), .Y(new_n3582_));
  OAI21X1  g3197(.A0(new_n3582_), .A1(new_n937_), .B0(new_n939_), .Y(new_n3583_));
  AOI21X1  g3198(.A0(new_n3583_), .A1(new_n944_), .B0(new_n947_), .Y(new_n3584_));
  OAI21X1  g3199(.A0(new_n3584_), .A1(new_n952_), .B0(new_n954_), .Y(new_n3585_));
  AOI21X1  g3200(.A0(new_n3585_), .A1(new_n959_), .B0(new_n962_), .Y(new_n3586_));
  OAI21X1  g3201(.A0(new_n3586_), .A1(new_n967_), .B0(new_n969_), .Y(new_n3587_));
  AOI21X1  g3202(.A0(new_n3587_), .A1(new_n974_), .B0(new_n977_), .Y(new_n3588_));
  OAI21X1  g3203(.A0(new_n3588_), .A1(new_n982_), .B0(new_n984_), .Y(new_n3589_));
  AOI21X1  g3204(.A0(new_n3589_), .A1(new_n989_), .B0(new_n992_), .Y(new_n3590_));
  OAI21X1  g3205(.A0(new_n3590_), .A1(new_n997_), .B0(new_n999_), .Y(new_n3591_));
  AOI21X1  g3206(.A0(new_n3591_), .A1(new_n1004_), .B0(new_n1007_), .Y(new_n3592_));
  OAI21X1  g3207(.A0(new_n3592_), .A1(new_n1012_), .B0(new_n1014_), .Y(new_n3593_));
  AOI21X1  g3208(.A0(new_n3593_), .A1(new_n1017_), .B0(new_n1711_), .Y(new_n3594_));
  OAI21X1  g3209(.A0(new_n3594_), .A1(new_n1710_), .B0(new_n1754_), .Y(new_n3595_));
  AOI21X1  g3210(.A0(new_n3595_), .A1(new_n1709_), .B0(new_n1983_), .Y(new_n3596_));
  OAI21X1  g3211(.A0(new_n3596_), .A1(new_n1613_), .B0(new_n1035_), .Y(new_n3597_));
  AOI21X1  g3212(.A0(new_n3597_), .A1(new_n1611_), .B0(new_n1612_), .Y(new_n3598_));
  OAI21X1  g3213(.A0(new_n3598_), .A1(new_n1610_), .B0(new_n1050_), .Y(new_n3599_));
  AOI21X1  g3214(.A0(new_n3599_), .A1(new_n1608_), .B0(new_n1609_), .Y(new_n3600_));
  OAI21X1  g3215(.A0(new_n3600_), .A1(new_n1607_), .B0(new_n1065_), .Y(new_n3601_));
  AOI21X1  g3216(.A0(new_n3601_), .A1(new_n1605_), .B0(new_n1606_), .Y(new_n3602_));
  OAI21X1  g3217(.A0(new_n3602_), .A1(new_n1604_), .B0(new_n1080_), .Y(new_n3603_));
  AOI21X1  g3218(.A0(new_n3603_), .A1(new_n1602_), .B0(new_n1603_), .Y(new_n3604_));
  OAI21X1  g3219(.A0(new_n3604_), .A1(new_n1601_), .B0(new_n1095_), .Y(new_n3605_));
  AOI21X1  g3220(.A0(new_n3605_), .A1(new_n1599_), .B0(new_n1600_), .Y(new_n3606_));
  OAI21X1  g3221(.A0(new_n3606_), .A1(new_n1598_), .B0(new_n1110_), .Y(new_n3607_));
  AOI21X1  g3222(.A0(new_n3607_), .A1(new_n1596_), .B0(new_n1597_), .Y(new_n3608_));
  OAI21X1  g3223(.A0(new_n3608_), .A1(new_n1595_), .B0(new_n1125_), .Y(new_n3609_));
  OAI21X1  g3224(.A0(new_n504_), .A1(\priority[49] ), .B0(\req[49] ), .Y(new_n3610_));
  AOI21X1  g3225(.A0(new_n3609_), .A1(new_n1593_), .B0(new_n3610_), .Y(\grant[49] ));
  NOR2X1   g3226(.A(new_n1139_), .B(new_n513_), .Y(new_n3612_));
  OAI21X1  g3227(.A0(new_n3612_), .A1(new_n1146_), .B0(new_n1148_), .Y(new_n3613_));
  AOI21X1  g3228(.A0(new_n3613_), .A1(new_n1153_), .B0(new_n1156_), .Y(new_n3614_));
  OAI21X1  g3229(.A0(new_n3614_), .A1(new_n1161_), .B0(new_n1163_), .Y(new_n3615_));
  AOI21X1  g3230(.A0(new_n3615_), .A1(new_n1168_), .B0(new_n1171_), .Y(new_n3616_));
  OAI21X1  g3231(.A0(new_n3616_), .A1(new_n1176_), .B0(new_n1178_), .Y(new_n3617_));
  AOI21X1  g3232(.A0(new_n3617_), .A1(new_n1183_), .B0(new_n1186_), .Y(new_n3618_));
  OAI21X1  g3233(.A0(new_n3618_), .A1(new_n1191_), .B0(new_n1193_), .Y(new_n3619_));
  AOI21X1  g3234(.A0(new_n3619_), .A1(new_n1198_), .B0(new_n1201_), .Y(new_n3620_));
  OAI21X1  g3235(.A0(new_n3620_), .A1(new_n1206_), .B0(new_n1208_), .Y(new_n3621_));
  AOI21X1  g3236(.A0(new_n3621_), .A1(new_n1213_), .B0(new_n1216_), .Y(new_n3622_));
  OAI21X1  g3237(.A0(new_n3622_), .A1(new_n1221_), .B0(new_n1223_), .Y(new_n3623_));
  AOI21X1  g3238(.A0(new_n3623_), .A1(new_n1228_), .B0(new_n1231_), .Y(new_n3624_));
  OAI21X1  g3239(.A0(new_n3624_), .A1(new_n1236_), .B0(new_n1238_), .Y(new_n3625_));
  AOI21X1  g3240(.A0(new_n3625_), .A1(new_n1243_), .B0(new_n1246_), .Y(new_n3626_));
  OAI21X1  g3241(.A0(new_n3626_), .A1(new_n1251_), .B0(new_n1253_), .Y(new_n3627_));
  AOI21X1  g3242(.A0(new_n3627_), .A1(new_n1258_), .B0(new_n1261_), .Y(new_n3628_));
  OAI21X1  g3243(.A0(new_n3628_), .A1(new_n1266_), .B0(new_n1268_), .Y(new_n3629_));
  AOI21X1  g3244(.A0(new_n3629_), .A1(new_n1273_), .B0(new_n1276_), .Y(new_n3630_));
  OAI21X1  g3245(.A0(new_n3630_), .A1(new_n1281_), .B0(new_n1283_), .Y(new_n3631_));
  AOI21X1  g3246(.A0(new_n3631_), .A1(new_n1288_), .B0(new_n1291_), .Y(new_n3632_));
  OAI21X1  g3247(.A0(new_n3632_), .A1(new_n1296_), .B0(new_n1298_), .Y(new_n3633_));
  AOI21X1  g3248(.A0(new_n3633_), .A1(new_n1303_), .B0(new_n1306_), .Y(new_n3634_));
  OAI21X1  g3249(.A0(new_n3634_), .A1(new_n1311_), .B0(new_n1313_), .Y(new_n3635_));
  AOI21X1  g3250(.A0(new_n3635_), .A1(new_n1318_), .B0(new_n1321_), .Y(new_n3636_));
  OAI21X1  g3251(.A0(new_n3636_), .A1(new_n1326_), .B0(new_n1328_), .Y(new_n3637_));
  AOI21X1  g3252(.A0(new_n3637_), .A1(new_n1331_), .B0(new_n1758_), .Y(new_n3638_));
  OAI21X1  g3253(.A0(new_n3638_), .A1(new_n394_), .B0(new_n396_), .Y(new_n3639_));
  AOI21X1  g3254(.A0(new_n3639_), .A1(new_n401_), .B0(new_n404_), .Y(new_n3640_));
  OAI21X1  g3255(.A0(new_n3640_), .A1(new_n409_), .B0(new_n411_), .Y(new_n3641_));
  AOI21X1  g3256(.A0(new_n3641_), .A1(new_n416_), .B0(new_n419_), .Y(new_n3642_));
  OAI21X1  g3257(.A0(new_n3642_), .A1(new_n424_), .B0(new_n426_), .Y(new_n3643_));
  AOI21X1  g3258(.A0(new_n3643_), .A1(new_n431_), .B0(new_n434_), .Y(new_n3644_));
  OAI21X1  g3259(.A0(new_n3644_), .A1(new_n439_), .B0(new_n441_), .Y(new_n3645_));
  AOI21X1  g3260(.A0(new_n3645_), .A1(new_n446_), .B0(new_n449_), .Y(new_n3646_));
  OAI21X1  g3261(.A0(new_n3646_), .A1(new_n454_), .B0(new_n456_), .Y(new_n3647_));
  AOI21X1  g3262(.A0(new_n3647_), .A1(new_n461_), .B0(new_n464_), .Y(new_n3648_));
  OAI21X1  g3263(.A0(new_n3648_), .A1(new_n469_), .B0(new_n471_), .Y(new_n3649_));
  AOI21X1  g3264(.A0(new_n3649_), .A1(new_n476_), .B0(new_n479_), .Y(new_n3650_));
  OAI21X1  g3265(.A0(new_n3650_), .A1(new_n484_), .B0(new_n486_), .Y(new_n3651_));
  AOI21X1  g3266(.A0(new_n3651_), .A1(new_n491_), .B0(new_n494_), .Y(new_n3652_));
  OAI21X1  g3267(.A0(new_n3652_), .A1(new_n499_), .B0(new_n501_), .Y(new_n3653_));
  OAI21X1  g3268(.A0(new_n822_), .A1(\priority[50] ), .B0(\req[50] ), .Y(new_n3654_));
  AOI21X1  g3269(.A0(new_n3653_), .A1(new_n506_), .B0(new_n3654_), .Y(\grant[50] ));
  NOR2X1   g3270(.A(new_n831_), .B(new_n515_), .Y(new_n3656_));
  OAI21X1  g3271(.A0(new_n3656_), .A1(new_n1371_), .B0(new_n523_), .Y(new_n3657_));
  AOI21X1  g3272(.A0(new_n3657_), .A1(new_n1369_), .B0(new_n1370_), .Y(new_n3658_));
  OAI21X1  g3273(.A0(new_n3658_), .A1(new_n1368_), .B0(new_n538_), .Y(new_n3659_));
  AOI21X1  g3274(.A0(new_n3659_), .A1(new_n1366_), .B0(new_n1367_), .Y(new_n3660_));
  OAI21X1  g3275(.A0(new_n3660_), .A1(new_n1365_), .B0(new_n553_), .Y(new_n3661_));
  AOI21X1  g3276(.A0(new_n3661_), .A1(new_n1363_), .B0(new_n1364_), .Y(new_n3662_));
  OAI21X1  g3277(.A0(new_n3662_), .A1(new_n1362_), .B0(new_n568_), .Y(new_n3663_));
  AOI21X1  g3278(.A0(new_n3663_), .A1(new_n1360_), .B0(new_n1361_), .Y(new_n3664_));
  OAI21X1  g3279(.A0(new_n3664_), .A1(new_n1359_), .B0(new_n583_), .Y(new_n3665_));
  AOI21X1  g3280(.A0(new_n3665_), .A1(new_n1357_), .B0(new_n1358_), .Y(new_n3666_));
  OAI21X1  g3281(.A0(new_n3666_), .A1(new_n1356_), .B0(new_n598_), .Y(new_n3667_));
  AOI21X1  g3282(.A0(new_n3667_), .A1(new_n1354_), .B0(new_n1355_), .Y(new_n3668_));
  OAI21X1  g3283(.A0(new_n3668_), .A1(new_n1353_), .B0(new_n613_), .Y(new_n3669_));
  AOI21X1  g3284(.A0(new_n3669_), .A1(new_n1351_), .B0(new_n1352_), .Y(new_n3670_));
  OAI21X1  g3285(.A0(new_n3670_), .A1(new_n1350_), .B0(new_n628_), .Y(new_n3671_));
  AOI21X1  g3286(.A0(new_n3671_), .A1(new_n1348_), .B0(new_n1349_), .Y(new_n3672_));
  OAI21X1  g3287(.A0(new_n3672_), .A1(new_n1347_), .B0(new_n643_), .Y(new_n3673_));
  AOI21X1  g3288(.A0(new_n3673_), .A1(new_n1345_), .B0(new_n1346_), .Y(new_n3674_));
  OAI21X1  g3289(.A0(new_n3674_), .A1(new_n1344_), .B0(new_n658_), .Y(new_n3675_));
  AOI21X1  g3290(.A0(new_n3675_), .A1(new_n1342_), .B0(new_n1343_), .Y(new_n3676_));
  OAI21X1  g3291(.A0(new_n3676_), .A1(new_n1341_), .B0(new_n673_), .Y(new_n3677_));
  AOI21X1  g3292(.A0(new_n3677_), .A1(new_n1339_), .B0(new_n1340_), .Y(new_n3678_));
  OAI21X1  g3293(.A0(new_n3678_), .A1(new_n1338_), .B0(new_n688_), .Y(new_n3679_));
  AOI21X1  g3294(.A0(new_n3679_), .A1(new_n1336_), .B0(new_n1337_), .Y(new_n3680_));
  OAI21X1  g3295(.A0(new_n3680_), .A1(new_n1335_), .B0(new_n1438_), .Y(new_n3681_));
  AOI21X1  g3296(.A0(new_n3681_), .A1(new_n1440_), .B0(new_n1803_), .Y(new_n3682_));
  OAI21X1  g3297(.A0(new_n3682_), .A1(new_n712_), .B0(new_n714_), .Y(new_n3683_));
  AOI21X1  g3298(.A0(new_n3683_), .A1(new_n719_), .B0(new_n722_), .Y(new_n3684_));
  OAI21X1  g3299(.A0(new_n3684_), .A1(new_n727_), .B0(new_n729_), .Y(new_n3685_));
  AOI21X1  g3300(.A0(new_n3685_), .A1(new_n734_), .B0(new_n737_), .Y(new_n3686_));
  OAI21X1  g3301(.A0(new_n3686_), .A1(new_n742_), .B0(new_n744_), .Y(new_n3687_));
  AOI21X1  g3302(.A0(new_n3687_), .A1(new_n749_), .B0(new_n752_), .Y(new_n3688_));
  OAI21X1  g3303(.A0(new_n3688_), .A1(new_n757_), .B0(new_n759_), .Y(new_n3689_));
  AOI21X1  g3304(.A0(new_n3689_), .A1(new_n764_), .B0(new_n767_), .Y(new_n3690_));
  OAI21X1  g3305(.A0(new_n3690_), .A1(new_n772_), .B0(new_n774_), .Y(new_n3691_));
  AOI21X1  g3306(.A0(new_n3691_), .A1(new_n779_), .B0(new_n782_), .Y(new_n3692_));
  OAI21X1  g3307(.A0(new_n3692_), .A1(new_n787_), .B0(new_n789_), .Y(new_n3693_));
  AOI21X1  g3308(.A0(new_n3693_), .A1(new_n794_), .B0(new_n797_), .Y(new_n3694_));
  OAI21X1  g3309(.A0(new_n3694_), .A1(new_n802_), .B0(new_n804_), .Y(new_n3695_));
  AOI21X1  g3310(.A0(new_n3695_), .A1(new_n809_), .B0(new_n812_), .Y(new_n3696_));
  OAI21X1  g3311(.A0(new_n3696_), .A1(new_n817_), .B0(new_n819_), .Y(new_n3697_));
  OAI21X1  g3312(.A0(new_n1136_), .A1(\priority[51] ), .B0(\req[51] ), .Y(new_n3698_));
  AOI21X1  g3313(.A0(new_n3697_), .A1(new_n824_), .B0(new_n3698_), .Y(\grant[51] ));
  NOR2X1   g3314(.A(new_n1145_), .B(new_n833_), .Y(new_n3700_));
  OAI21X1  g3315(.A0(new_n3700_), .A1(new_n1480_), .B0(new_n841_), .Y(new_n3701_));
  AOI21X1  g3316(.A0(new_n3701_), .A1(new_n1478_), .B0(new_n1479_), .Y(new_n3702_));
  OAI21X1  g3317(.A0(new_n3702_), .A1(new_n1477_), .B0(new_n856_), .Y(new_n3703_));
  AOI21X1  g3318(.A0(new_n3703_), .A1(new_n1475_), .B0(new_n1476_), .Y(new_n3704_));
  OAI21X1  g3319(.A0(new_n3704_), .A1(new_n1474_), .B0(new_n871_), .Y(new_n3705_));
  AOI21X1  g3320(.A0(new_n3705_), .A1(new_n1472_), .B0(new_n1473_), .Y(new_n3706_));
  OAI21X1  g3321(.A0(new_n3706_), .A1(new_n1471_), .B0(new_n886_), .Y(new_n3707_));
  AOI21X1  g3322(.A0(new_n3707_), .A1(new_n1469_), .B0(new_n1470_), .Y(new_n3708_));
  OAI21X1  g3323(.A0(new_n3708_), .A1(new_n1468_), .B0(new_n901_), .Y(new_n3709_));
  AOI21X1  g3324(.A0(new_n3709_), .A1(new_n1466_), .B0(new_n1467_), .Y(new_n3710_));
  OAI21X1  g3325(.A0(new_n3710_), .A1(new_n1465_), .B0(new_n916_), .Y(new_n3711_));
  AOI21X1  g3326(.A0(new_n3711_), .A1(new_n1463_), .B0(new_n1464_), .Y(new_n3712_));
  OAI21X1  g3327(.A0(new_n3712_), .A1(new_n1462_), .B0(new_n931_), .Y(new_n3713_));
  AOI21X1  g3328(.A0(new_n3713_), .A1(new_n1460_), .B0(new_n1461_), .Y(new_n3714_));
  OAI21X1  g3329(.A0(new_n3714_), .A1(new_n1459_), .B0(new_n946_), .Y(new_n3715_));
  AOI21X1  g3330(.A0(new_n3715_), .A1(new_n1457_), .B0(new_n1458_), .Y(new_n3716_));
  OAI21X1  g3331(.A0(new_n3716_), .A1(new_n1456_), .B0(new_n961_), .Y(new_n3717_));
  AOI21X1  g3332(.A0(new_n3717_), .A1(new_n1454_), .B0(new_n1455_), .Y(new_n3718_));
  OAI21X1  g3333(.A0(new_n3718_), .A1(new_n1453_), .B0(new_n976_), .Y(new_n3719_));
  AOI21X1  g3334(.A0(new_n3719_), .A1(new_n1451_), .B0(new_n1452_), .Y(new_n3720_));
  OAI21X1  g3335(.A0(new_n3720_), .A1(new_n1450_), .B0(new_n991_), .Y(new_n3721_));
  AOI21X1  g3336(.A0(new_n3721_), .A1(new_n1448_), .B0(new_n1449_), .Y(new_n3722_));
  OAI21X1  g3337(.A0(new_n3722_), .A1(new_n1447_), .B0(new_n1006_), .Y(new_n3723_));
  AOI21X1  g3338(.A0(new_n3723_), .A1(new_n1445_), .B0(new_n1446_), .Y(new_n3724_));
  OAI21X1  g3339(.A0(new_n3724_), .A1(new_n1444_), .B0(new_n1547_), .Y(new_n3725_));
  AOI21X1  g3340(.A0(new_n3725_), .A1(new_n1549_), .B0(new_n1848_), .Y(new_n3726_));
  OAI21X1  g3341(.A0(new_n3726_), .A1(new_n1026_), .B0(new_n1028_), .Y(new_n3727_));
  AOI21X1  g3342(.A0(new_n3727_), .A1(new_n1033_), .B0(new_n1036_), .Y(new_n3728_));
  OAI21X1  g3343(.A0(new_n3728_), .A1(new_n1041_), .B0(new_n1043_), .Y(new_n3729_));
  AOI21X1  g3344(.A0(new_n3729_), .A1(new_n1048_), .B0(new_n1051_), .Y(new_n3730_));
  OAI21X1  g3345(.A0(new_n3730_), .A1(new_n1056_), .B0(new_n1058_), .Y(new_n3731_));
  AOI21X1  g3346(.A0(new_n3731_), .A1(new_n1063_), .B0(new_n1066_), .Y(new_n3732_));
  OAI21X1  g3347(.A0(new_n3732_), .A1(new_n1071_), .B0(new_n1073_), .Y(new_n3733_));
  AOI21X1  g3348(.A0(new_n3733_), .A1(new_n1078_), .B0(new_n1081_), .Y(new_n3734_));
  OAI21X1  g3349(.A0(new_n3734_), .A1(new_n1086_), .B0(new_n1088_), .Y(new_n3735_));
  AOI21X1  g3350(.A0(new_n3735_), .A1(new_n1093_), .B0(new_n1096_), .Y(new_n3736_));
  OAI21X1  g3351(.A0(new_n3736_), .A1(new_n1101_), .B0(new_n1103_), .Y(new_n3737_));
  AOI21X1  g3352(.A0(new_n3737_), .A1(new_n1108_), .B0(new_n1111_), .Y(new_n3738_));
  OAI21X1  g3353(.A0(new_n3738_), .A1(new_n1116_), .B0(new_n1118_), .Y(new_n3739_));
  AOI21X1  g3354(.A0(new_n3739_), .A1(new_n1123_), .B0(new_n1126_), .Y(new_n3740_));
  OAI21X1  g3355(.A0(new_n3740_), .A1(new_n1131_), .B0(new_n1133_), .Y(new_n3741_));
  OAI21X1  g3356(.A0(new_n512_), .A1(\priority[52] ), .B0(\req[52] ), .Y(new_n3742_));
  AOI21X1  g3357(.A0(new_n3741_), .A1(new_n1138_), .B0(new_n3742_), .Y(\grant[52] ));
  NOR2X1   g3358(.A(new_n1147_), .B(new_n520_), .Y(new_n3744_));
  OAI21X1  g3359(.A0(new_n3744_), .A1(new_n1589_), .B0(new_n1155_), .Y(new_n3745_));
  AOI21X1  g3360(.A0(new_n3745_), .A1(new_n1587_), .B0(new_n1588_), .Y(new_n3746_));
  OAI21X1  g3361(.A0(new_n3746_), .A1(new_n1586_), .B0(new_n1170_), .Y(new_n3747_));
  AOI21X1  g3362(.A0(new_n3747_), .A1(new_n1584_), .B0(new_n1585_), .Y(new_n3748_));
  OAI21X1  g3363(.A0(new_n3748_), .A1(new_n1583_), .B0(new_n1185_), .Y(new_n3749_));
  AOI21X1  g3364(.A0(new_n3749_), .A1(new_n1581_), .B0(new_n1582_), .Y(new_n3750_));
  OAI21X1  g3365(.A0(new_n3750_), .A1(new_n1580_), .B0(new_n1200_), .Y(new_n3751_));
  AOI21X1  g3366(.A0(new_n3751_), .A1(new_n1578_), .B0(new_n1579_), .Y(new_n3752_));
  OAI21X1  g3367(.A0(new_n3752_), .A1(new_n1577_), .B0(new_n1215_), .Y(new_n3753_));
  AOI21X1  g3368(.A0(new_n3753_), .A1(new_n1575_), .B0(new_n1576_), .Y(new_n3754_));
  OAI21X1  g3369(.A0(new_n3754_), .A1(new_n1574_), .B0(new_n1230_), .Y(new_n3755_));
  AOI21X1  g3370(.A0(new_n3755_), .A1(new_n1572_), .B0(new_n1573_), .Y(new_n3756_));
  OAI21X1  g3371(.A0(new_n3756_), .A1(new_n1571_), .B0(new_n1245_), .Y(new_n3757_));
  AOI21X1  g3372(.A0(new_n3757_), .A1(new_n1569_), .B0(new_n1570_), .Y(new_n3758_));
  OAI21X1  g3373(.A0(new_n3758_), .A1(new_n1568_), .B0(new_n1260_), .Y(new_n3759_));
  AOI21X1  g3374(.A0(new_n3759_), .A1(new_n1566_), .B0(new_n1567_), .Y(new_n3760_));
  OAI21X1  g3375(.A0(new_n3760_), .A1(new_n1565_), .B0(new_n1275_), .Y(new_n3761_));
  AOI21X1  g3376(.A0(new_n3761_), .A1(new_n1563_), .B0(new_n1564_), .Y(new_n3762_));
  OAI21X1  g3377(.A0(new_n3762_), .A1(new_n1562_), .B0(new_n1290_), .Y(new_n3763_));
  AOI21X1  g3378(.A0(new_n3763_), .A1(new_n1560_), .B0(new_n1561_), .Y(new_n3764_));
  OAI21X1  g3379(.A0(new_n3764_), .A1(new_n1559_), .B0(new_n1305_), .Y(new_n3765_));
  AOI21X1  g3380(.A0(new_n3765_), .A1(new_n1557_), .B0(new_n1558_), .Y(new_n3766_));
  OAI21X1  g3381(.A0(new_n3766_), .A1(new_n1556_), .B0(new_n1320_), .Y(new_n3767_));
  AOI21X1  g3382(.A0(new_n3767_), .A1(new_n1554_), .B0(new_n1555_), .Y(new_n3768_));
  OAI21X1  g3383(.A0(new_n3768_), .A1(new_n1553_), .B0(new_n1656_), .Y(new_n3769_));
  AOI21X1  g3384(.A0(new_n3769_), .A1(new_n1552_), .B0(new_n1893_), .Y(new_n3770_));
  OAI21X1  g3385(.A0(new_n3770_), .A1(new_n1395_), .B0(new_n403_), .Y(new_n3771_));
  AOI21X1  g3386(.A0(new_n3771_), .A1(new_n1393_), .B0(new_n1394_), .Y(new_n3772_));
  OAI21X1  g3387(.A0(new_n3772_), .A1(new_n1392_), .B0(new_n418_), .Y(new_n3773_));
  AOI21X1  g3388(.A0(new_n3773_), .A1(new_n1390_), .B0(new_n1391_), .Y(new_n3774_));
  OAI21X1  g3389(.A0(new_n3774_), .A1(new_n1389_), .B0(new_n433_), .Y(new_n3775_));
  AOI21X1  g3390(.A0(new_n3775_), .A1(new_n1387_), .B0(new_n1388_), .Y(new_n3776_));
  OAI21X1  g3391(.A0(new_n3776_), .A1(new_n1386_), .B0(new_n448_), .Y(new_n3777_));
  AOI21X1  g3392(.A0(new_n3777_), .A1(new_n1384_), .B0(new_n1385_), .Y(new_n3778_));
  OAI21X1  g3393(.A0(new_n3778_), .A1(new_n1383_), .B0(new_n463_), .Y(new_n3779_));
  AOI21X1  g3394(.A0(new_n3779_), .A1(new_n1381_), .B0(new_n1382_), .Y(new_n3780_));
  OAI21X1  g3395(.A0(new_n3780_), .A1(new_n1380_), .B0(new_n478_), .Y(new_n3781_));
  AOI21X1  g3396(.A0(new_n3781_), .A1(new_n1378_), .B0(new_n1379_), .Y(new_n3782_));
  OAI21X1  g3397(.A0(new_n3782_), .A1(new_n1377_), .B0(new_n493_), .Y(new_n3783_));
  AOI21X1  g3398(.A0(new_n3783_), .A1(new_n1375_), .B0(new_n1376_), .Y(new_n3784_));
  OAI21X1  g3399(.A0(new_n3784_), .A1(new_n1374_), .B0(new_n508_), .Y(new_n3785_));
  OAI21X1  g3400(.A0(new_n830_), .A1(\priority[53] ), .B0(\req[53] ), .Y(new_n3786_));
  AOI21X1  g3401(.A0(new_n3785_), .A1(new_n1372_), .B0(new_n3786_), .Y(\grant[53] ));
  NOR2X1   g3402(.A(new_n838_), .B(new_n522_), .Y(new_n3788_));
  OAI21X1  g3403(.A0(new_n3788_), .A1(new_n529_), .B0(new_n531_), .Y(new_n3789_));
  AOI21X1  g3404(.A0(new_n3789_), .A1(new_n536_), .B0(new_n539_), .Y(new_n3790_));
  OAI21X1  g3405(.A0(new_n3790_), .A1(new_n544_), .B0(new_n546_), .Y(new_n3791_));
  AOI21X1  g3406(.A0(new_n3791_), .A1(new_n551_), .B0(new_n554_), .Y(new_n3792_));
  OAI21X1  g3407(.A0(new_n3792_), .A1(new_n559_), .B0(new_n561_), .Y(new_n3793_));
  AOI21X1  g3408(.A0(new_n3793_), .A1(new_n566_), .B0(new_n569_), .Y(new_n3794_));
  OAI21X1  g3409(.A0(new_n3794_), .A1(new_n574_), .B0(new_n576_), .Y(new_n3795_));
  AOI21X1  g3410(.A0(new_n3795_), .A1(new_n581_), .B0(new_n584_), .Y(new_n3796_));
  OAI21X1  g3411(.A0(new_n3796_), .A1(new_n589_), .B0(new_n591_), .Y(new_n3797_));
  AOI21X1  g3412(.A0(new_n3797_), .A1(new_n596_), .B0(new_n599_), .Y(new_n3798_));
  OAI21X1  g3413(.A0(new_n3798_), .A1(new_n604_), .B0(new_n606_), .Y(new_n3799_));
  AOI21X1  g3414(.A0(new_n3799_), .A1(new_n611_), .B0(new_n614_), .Y(new_n3800_));
  OAI21X1  g3415(.A0(new_n3800_), .A1(new_n619_), .B0(new_n621_), .Y(new_n3801_));
  AOI21X1  g3416(.A0(new_n3801_), .A1(new_n626_), .B0(new_n629_), .Y(new_n3802_));
  OAI21X1  g3417(.A0(new_n3802_), .A1(new_n634_), .B0(new_n636_), .Y(new_n3803_));
  AOI21X1  g3418(.A0(new_n3803_), .A1(new_n641_), .B0(new_n644_), .Y(new_n3804_));
  OAI21X1  g3419(.A0(new_n3804_), .A1(new_n649_), .B0(new_n651_), .Y(new_n3805_));
  AOI21X1  g3420(.A0(new_n3805_), .A1(new_n656_), .B0(new_n659_), .Y(new_n3806_));
  OAI21X1  g3421(.A0(new_n3806_), .A1(new_n664_), .B0(new_n666_), .Y(new_n3807_));
  AOI21X1  g3422(.A0(new_n3807_), .A1(new_n671_), .B0(new_n674_), .Y(new_n3808_));
  OAI21X1  g3423(.A0(new_n3808_), .A1(new_n679_), .B0(new_n681_), .Y(new_n3809_));
  AOI21X1  g3424(.A0(new_n3809_), .A1(new_n686_), .B0(new_n689_), .Y(new_n3810_));
  OAI21X1  g3425(.A0(new_n3810_), .A1(new_n694_), .B0(new_n696_), .Y(new_n3811_));
  AOI21X1  g3426(.A0(new_n3811_), .A1(new_n701_), .B0(new_n1662_), .Y(new_n3812_));
  OAI21X1  g3427(.A0(new_n3812_), .A1(new_n1661_), .B0(new_n1705_), .Y(new_n3813_));
  AOI21X1  g3428(.A0(new_n3813_), .A1(new_n1660_), .B0(new_n1938_), .Y(new_n3814_));
  OAI21X1  g3429(.A0(new_n3814_), .A1(new_n1504_), .B0(new_n721_), .Y(new_n3815_));
  AOI21X1  g3430(.A0(new_n3815_), .A1(new_n1502_), .B0(new_n1503_), .Y(new_n3816_));
  OAI21X1  g3431(.A0(new_n3816_), .A1(new_n1501_), .B0(new_n736_), .Y(new_n3817_));
  AOI21X1  g3432(.A0(new_n3817_), .A1(new_n1499_), .B0(new_n1500_), .Y(new_n3818_));
  OAI21X1  g3433(.A0(new_n3818_), .A1(new_n1498_), .B0(new_n751_), .Y(new_n3819_));
  AOI21X1  g3434(.A0(new_n3819_), .A1(new_n1496_), .B0(new_n1497_), .Y(new_n3820_));
  OAI21X1  g3435(.A0(new_n3820_), .A1(new_n1495_), .B0(new_n766_), .Y(new_n3821_));
  AOI21X1  g3436(.A0(new_n3821_), .A1(new_n1493_), .B0(new_n1494_), .Y(new_n3822_));
  OAI21X1  g3437(.A0(new_n3822_), .A1(new_n1492_), .B0(new_n781_), .Y(new_n3823_));
  AOI21X1  g3438(.A0(new_n3823_), .A1(new_n1490_), .B0(new_n1491_), .Y(new_n3824_));
  OAI21X1  g3439(.A0(new_n3824_), .A1(new_n1489_), .B0(new_n796_), .Y(new_n3825_));
  AOI21X1  g3440(.A0(new_n3825_), .A1(new_n1487_), .B0(new_n1488_), .Y(new_n3826_));
  OAI21X1  g3441(.A0(new_n3826_), .A1(new_n1486_), .B0(new_n811_), .Y(new_n3827_));
  AOI21X1  g3442(.A0(new_n3827_), .A1(new_n1484_), .B0(new_n1485_), .Y(new_n3828_));
  OAI21X1  g3443(.A0(new_n3828_), .A1(new_n1483_), .B0(new_n826_), .Y(new_n3829_));
  OAI21X1  g3444(.A0(new_n1144_), .A1(\priority[54] ), .B0(\req[54] ), .Y(new_n3830_));
  AOI21X1  g3445(.A0(new_n3829_), .A1(new_n1481_), .B0(new_n3830_), .Y(\grant[54] ));
  NOR2X1   g3446(.A(new_n1152_), .B(new_n840_), .Y(new_n3832_));
  OAI21X1  g3447(.A0(new_n3832_), .A1(new_n847_), .B0(new_n849_), .Y(new_n3833_));
  AOI21X1  g3448(.A0(new_n3833_), .A1(new_n854_), .B0(new_n857_), .Y(new_n3834_));
  OAI21X1  g3449(.A0(new_n3834_), .A1(new_n862_), .B0(new_n864_), .Y(new_n3835_));
  AOI21X1  g3450(.A0(new_n3835_), .A1(new_n869_), .B0(new_n872_), .Y(new_n3836_));
  OAI21X1  g3451(.A0(new_n3836_), .A1(new_n877_), .B0(new_n879_), .Y(new_n3837_));
  AOI21X1  g3452(.A0(new_n3837_), .A1(new_n884_), .B0(new_n887_), .Y(new_n3838_));
  OAI21X1  g3453(.A0(new_n3838_), .A1(new_n892_), .B0(new_n894_), .Y(new_n3839_));
  AOI21X1  g3454(.A0(new_n3839_), .A1(new_n899_), .B0(new_n902_), .Y(new_n3840_));
  OAI21X1  g3455(.A0(new_n3840_), .A1(new_n907_), .B0(new_n909_), .Y(new_n3841_));
  AOI21X1  g3456(.A0(new_n3841_), .A1(new_n914_), .B0(new_n917_), .Y(new_n3842_));
  OAI21X1  g3457(.A0(new_n3842_), .A1(new_n922_), .B0(new_n924_), .Y(new_n3843_));
  AOI21X1  g3458(.A0(new_n3843_), .A1(new_n929_), .B0(new_n932_), .Y(new_n3844_));
  OAI21X1  g3459(.A0(new_n3844_), .A1(new_n937_), .B0(new_n939_), .Y(new_n3845_));
  AOI21X1  g3460(.A0(new_n3845_), .A1(new_n944_), .B0(new_n947_), .Y(new_n3846_));
  OAI21X1  g3461(.A0(new_n3846_), .A1(new_n952_), .B0(new_n954_), .Y(new_n3847_));
  AOI21X1  g3462(.A0(new_n3847_), .A1(new_n959_), .B0(new_n962_), .Y(new_n3848_));
  OAI21X1  g3463(.A0(new_n3848_), .A1(new_n967_), .B0(new_n969_), .Y(new_n3849_));
  AOI21X1  g3464(.A0(new_n3849_), .A1(new_n974_), .B0(new_n977_), .Y(new_n3850_));
  OAI21X1  g3465(.A0(new_n3850_), .A1(new_n982_), .B0(new_n984_), .Y(new_n3851_));
  AOI21X1  g3466(.A0(new_n3851_), .A1(new_n989_), .B0(new_n992_), .Y(new_n3852_));
  OAI21X1  g3467(.A0(new_n3852_), .A1(new_n997_), .B0(new_n999_), .Y(new_n3853_));
  AOI21X1  g3468(.A0(new_n3853_), .A1(new_n1004_), .B0(new_n1007_), .Y(new_n3854_));
  OAI21X1  g3469(.A0(new_n3854_), .A1(new_n1012_), .B0(new_n1014_), .Y(new_n3855_));
  AOI21X1  g3470(.A0(new_n3855_), .A1(new_n1017_), .B0(new_n1711_), .Y(new_n3856_));
  OAI21X1  g3471(.A0(new_n3856_), .A1(new_n1710_), .B0(new_n1754_), .Y(new_n3857_));
  AOI21X1  g3472(.A0(new_n3857_), .A1(new_n1709_), .B0(new_n1983_), .Y(new_n3858_));
  OAI21X1  g3473(.A0(new_n3858_), .A1(new_n1613_), .B0(new_n1035_), .Y(new_n3859_));
  AOI21X1  g3474(.A0(new_n3859_), .A1(new_n1611_), .B0(new_n1612_), .Y(new_n3860_));
  OAI21X1  g3475(.A0(new_n3860_), .A1(new_n1610_), .B0(new_n1050_), .Y(new_n3861_));
  AOI21X1  g3476(.A0(new_n3861_), .A1(new_n1608_), .B0(new_n1609_), .Y(new_n3862_));
  OAI21X1  g3477(.A0(new_n3862_), .A1(new_n1607_), .B0(new_n1065_), .Y(new_n3863_));
  AOI21X1  g3478(.A0(new_n3863_), .A1(new_n1605_), .B0(new_n1606_), .Y(new_n3864_));
  OAI21X1  g3479(.A0(new_n3864_), .A1(new_n1604_), .B0(new_n1080_), .Y(new_n3865_));
  AOI21X1  g3480(.A0(new_n3865_), .A1(new_n1602_), .B0(new_n1603_), .Y(new_n3866_));
  OAI21X1  g3481(.A0(new_n3866_), .A1(new_n1601_), .B0(new_n1095_), .Y(new_n3867_));
  AOI21X1  g3482(.A0(new_n3867_), .A1(new_n1599_), .B0(new_n1600_), .Y(new_n3868_));
  OAI21X1  g3483(.A0(new_n3868_), .A1(new_n1598_), .B0(new_n1110_), .Y(new_n3869_));
  AOI21X1  g3484(.A0(new_n3869_), .A1(new_n1596_), .B0(new_n1597_), .Y(new_n3870_));
  OAI21X1  g3485(.A0(new_n3870_), .A1(new_n1595_), .B0(new_n1125_), .Y(new_n3871_));
  AOI21X1  g3486(.A0(new_n3871_), .A1(new_n1593_), .B0(new_n1594_), .Y(new_n3872_));
  OAI21X1  g3487(.A0(new_n3872_), .A1(new_n1592_), .B0(new_n1140_), .Y(new_n3873_));
  OAI21X1  g3488(.A0(new_n519_), .A1(\priority[55] ), .B0(\req[55] ), .Y(new_n3874_));
  AOI21X1  g3489(.A0(new_n3873_), .A1(new_n1590_), .B0(new_n3874_), .Y(\grant[55] ));
  NOR2X1   g3490(.A(new_n1154_), .B(new_n528_), .Y(new_n3876_));
  OAI21X1  g3491(.A0(new_n3876_), .A1(new_n1161_), .B0(new_n1163_), .Y(new_n3877_));
  AOI21X1  g3492(.A0(new_n3877_), .A1(new_n1168_), .B0(new_n1171_), .Y(new_n3878_));
  OAI21X1  g3493(.A0(new_n3878_), .A1(new_n1176_), .B0(new_n1178_), .Y(new_n3879_));
  AOI21X1  g3494(.A0(new_n3879_), .A1(new_n1183_), .B0(new_n1186_), .Y(new_n3880_));
  OAI21X1  g3495(.A0(new_n3880_), .A1(new_n1191_), .B0(new_n1193_), .Y(new_n3881_));
  AOI21X1  g3496(.A0(new_n3881_), .A1(new_n1198_), .B0(new_n1201_), .Y(new_n3882_));
  OAI21X1  g3497(.A0(new_n3882_), .A1(new_n1206_), .B0(new_n1208_), .Y(new_n3883_));
  AOI21X1  g3498(.A0(new_n3883_), .A1(new_n1213_), .B0(new_n1216_), .Y(new_n3884_));
  OAI21X1  g3499(.A0(new_n3884_), .A1(new_n1221_), .B0(new_n1223_), .Y(new_n3885_));
  AOI21X1  g3500(.A0(new_n3885_), .A1(new_n1228_), .B0(new_n1231_), .Y(new_n3886_));
  OAI21X1  g3501(.A0(new_n3886_), .A1(new_n1236_), .B0(new_n1238_), .Y(new_n3887_));
  AOI21X1  g3502(.A0(new_n3887_), .A1(new_n1243_), .B0(new_n1246_), .Y(new_n3888_));
  OAI21X1  g3503(.A0(new_n3888_), .A1(new_n1251_), .B0(new_n1253_), .Y(new_n3889_));
  AOI21X1  g3504(.A0(new_n3889_), .A1(new_n1258_), .B0(new_n1261_), .Y(new_n3890_));
  OAI21X1  g3505(.A0(new_n3890_), .A1(new_n1266_), .B0(new_n1268_), .Y(new_n3891_));
  AOI21X1  g3506(.A0(new_n3891_), .A1(new_n1273_), .B0(new_n1276_), .Y(new_n3892_));
  OAI21X1  g3507(.A0(new_n3892_), .A1(new_n1281_), .B0(new_n1283_), .Y(new_n3893_));
  AOI21X1  g3508(.A0(new_n3893_), .A1(new_n1288_), .B0(new_n1291_), .Y(new_n3894_));
  OAI21X1  g3509(.A0(new_n3894_), .A1(new_n1296_), .B0(new_n1298_), .Y(new_n3895_));
  AOI21X1  g3510(.A0(new_n3895_), .A1(new_n1303_), .B0(new_n1306_), .Y(new_n3896_));
  OAI21X1  g3511(.A0(new_n3896_), .A1(new_n1311_), .B0(new_n1313_), .Y(new_n3897_));
  AOI21X1  g3512(.A0(new_n3897_), .A1(new_n1318_), .B0(new_n1321_), .Y(new_n3898_));
  OAI21X1  g3513(.A0(new_n3898_), .A1(new_n1326_), .B0(new_n1328_), .Y(new_n3899_));
  AOI21X1  g3514(.A0(new_n3899_), .A1(new_n1331_), .B0(new_n1758_), .Y(new_n3900_));
  OAI21X1  g3515(.A0(new_n3900_), .A1(new_n394_), .B0(new_n396_), .Y(new_n3901_));
  AOI21X1  g3516(.A0(new_n3901_), .A1(new_n401_), .B0(new_n404_), .Y(new_n3902_));
  OAI21X1  g3517(.A0(new_n3902_), .A1(new_n409_), .B0(new_n411_), .Y(new_n3903_));
  AOI21X1  g3518(.A0(new_n3903_), .A1(new_n416_), .B0(new_n419_), .Y(new_n3904_));
  OAI21X1  g3519(.A0(new_n3904_), .A1(new_n424_), .B0(new_n426_), .Y(new_n3905_));
  AOI21X1  g3520(.A0(new_n3905_), .A1(new_n431_), .B0(new_n434_), .Y(new_n3906_));
  OAI21X1  g3521(.A0(new_n3906_), .A1(new_n439_), .B0(new_n441_), .Y(new_n3907_));
  AOI21X1  g3522(.A0(new_n3907_), .A1(new_n446_), .B0(new_n449_), .Y(new_n3908_));
  OAI21X1  g3523(.A0(new_n3908_), .A1(new_n454_), .B0(new_n456_), .Y(new_n3909_));
  AOI21X1  g3524(.A0(new_n3909_), .A1(new_n461_), .B0(new_n464_), .Y(new_n3910_));
  OAI21X1  g3525(.A0(new_n3910_), .A1(new_n469_), .B0(new_n471_), .Y(new_n3911_));
  AOI21X1  g3526(.A0(new_n3911_), .A1(new_n476_), .B0(new_n479_), .Y(new_n3912_));
  OAI21X1  g3527(.A0(new_n3912_), .A1(new_n484_), .B0(new_n486_), .Y(new_n3913_));
  AOI21X1  g3528(.A0(new_n3913_), .A1(new_n491_), .B0(new_n494_), .Y(new_n3914_));
  OAI21X1  g3529(.A0(new_n3914_), .A1(new_n499_), .B0(new_n501_), .Y(new_n3915_));
  AOI21X1  g3530(.A0(new_n3915_), .A1(new_n506_), .B0(new_n509_), .Y(new_n3916_));
  OAI21X1  g3531(.A0(new_n3916_), .A1(new_n514_), .B0(new_n516_), .Y(new_n3917_));
  OAI21X1  g3532(.A0(new_n837_), .A1(\priority[56] ), .B0(\req[56] ), .Y(new_n3918_));
  AOI21X1  g3533(.A0(new_n3917_), .A1(new_n521_), .B0(new_n3918_), .Y(\grant[56] ));
  NOR2X1   g3534(.A(new_n846_), .B(new_n530_), .Y(new_n3920_));
  OAI21X1  g3535(.A0(new_n3920_), .A1(new_n1368_), .B0(new_n538_), .Y(new_n3921_));
  AOI21X1  g3536(.A0(new_n3921_), .A1(new_n1366_), .B0(new_n1367_), .Y(new_n3922_));
  OAI21X1  g3537(.A0(new_n3922_), .A1(new_n1365_), .B0(new_n553_), .Y(new_n3923_));
  AOI21X1  g3538(.A0(new_n3923_), .A1(new_n1363_), .B0(new_n1364_), .Y(new_n3924_));
  OAI21X1  g3539(.A0(new_n3924_), .A1(new_n1362_), .B0(new_n568_), .Y(new_n3925_));
  AOI21X1  g3540(.A0(new_n3925_), .A1(new_n1360_), .B0(new_n1361_), .Y(new_n3926_));
  OAI21X1  g3541(.A0(new_n3926_), .A1(new_n1359_), .B0(new_n583_), .Y(new_n3927_));
  AOI21X1  g3542(.A0(new_n3927_), .A1(new_n1357_), .B0(new_n1358_), .Y(new_n3928_));
  OAI21X1  g3543(.A0(new_n3928_), .A1(new_n1356_), .B0(new_n598_), .Y(new_n3929_));
  AOI21X1  g3544(.A0(new_n3929_), .A1(new_n1354_), .B0(new_n1355_), .Y(new_n3930_));
  OAI21X1  g3545(.A0(new_n3930_), .A1(new_n1353_), .B0(new_n613_), .Y(new_n3931_));
  AOI21X1  g3546(.A0(new_n3931_), .A1(new_n1351_), .B0(new_n1352_), .Y(new_n3932_));
  OAI21X1  g3547(.A0(new_n3932_), .A1(new_n1350_), .B0(new_n628_), .Y(new_n3933_));
  AOI21X1  g3548(.A0(new_n3933_), .A1(new_n1348_), .B0(new_n1349_), .Y(new_n3934_));
  OAI21X1  g3549(.A0(new_n3934_), .A1(new_n1347_), .B0(new_n643_), .Y(new_n3935_));
  AOI21X1  g3550(.A0(new_n3935_), .A1(new_n1345_), .B0(new_n1346_), .Y(new_n3936_));
  OAI21X1  g3551(.A0(new_n3936_), .A1(new_n1344_), .B0(new_n658_), .Y(new_n3937_));
  AOI21X1  g3552(.A0(new_n3937_), .A1(new_n1342_), .B0(new_n1343_), .Y(new_n3938_));
  OAI21X1  g3553(.A0(new_n3938_), .A1(new_n1341_), .B0(new_n673_), .Y(new_n3939_));
  AOI21X1  g3554(.A0(new_n3939_), .A1(new_n1339_), .B0(new_n1340_), .Y(new_n3940_));
  OAI21X1  g3555(.A0(new_n3940_), .A1(new_n1338_), .B0(new_n688_), .Y(new_n3941_));
  AOI21X1  g3556(.A0(new_n3941_), .A1(new_n1336_), .B0(new_n1337_), .Y(new_n3942_));
  OAI21X1  g3557(.A0(new_n3942_), .A1(new_n1335_), .B0(new_n1438_), .Y(new_n3943_));
  AOI21X1  g3558(.A0(new_n3943_), .A1(new_n1440_), .B0(new_n1803_), .Y(new_n3944_));
  OAI21X1  g3559(.A0(new_n3944_), .A1(new_n712_), .B0(new_n714_), .Y(new_n3945_));
  AOI21X1  g3560(.A0(new_n3945_), .A1(new_n719_), .B0(new_n722_), .Y(new_n3946_));
  OAI21X1  g3561(.A0(new_n3946_), .A1(new_n727_), .B0(new_n729_), .Y(new_n3947_));
  AOI21X1  g3562(.A0(new_n3947_), .A1(new_n734_), .B0(new_n737_), .Y(new_n3948_));
  OAI21X1  g3563(.A0(new_n3948_), .A1(new_n742_), .B0(new_n744_), .Y(new_n3949_));
  AOI21X1  g3564(.A0(new_n3949_), .A1(new_n749_), .B0(new_n752_), .Y(new_n3950_));
  OAI21X1  g3565(.A0(new_n3950_), .A1(new_n757_), .B0(new_n759_), .Y(new_n3951_));
  AOI21X1  g3566(.A0(new_n3951_), .A1(new_n764_), .B0(new_n767_), .Y(new_n3952_));
  OAI21X1  g3567(.A0(new_n3952_), .A1(new_n772_), .B0(new_n774_), .Y(new_n3953_));
  AOI21X1  g3568(.A0(new_n3953_), .A1(new_n779_), .B0(new_n782_), .Y(new_n3954_));
  OAI21X1  g3569(.A0(new_n3954_), .A1(new_n787_), .B0(new_n789_), .Y(new_n3955_));
  AOI21X1  g3570(.A0(new_n3955_), .A1(new_n794_), .B0(new_n797_), .Y(new_n3956_));
  OAI21X1  g3571(.A0(new_n3956_), .A1(new_n802_), .B0(new_n804_), .Y(new_n3957_));
  AOI21X1  g3572(.A0(new_n3957_), .A1(new_n809_), .B0(new_n812_), .Y(new_n3958_));
  OAI21X1  g3573(.A0(new_n3958_), .A1(new_n817_), .B0(new_n819_), .Y(new_n3959_));
  AOI21X1  g3574(.A0(new_n3959_), .A1(new_n824_), .B0(new_n827_), .Y(new_n3960_));
  OAI21X1  g3575(.A0(new_n3960_), .A1(new_n832_), .B0(new_n834_), .Y(new_n3961_));
  OAI21X1  g3576(.A0(new_n1151_), .A1(\priority[57] ), .B0(\req[57] ), .Y(new_n3962_));
  AOI21X1  g3577(.A0(new_n3961_), .A1(new_n839_), .B0(new_n3962_), .Y(\grant[57] ));
  NOR2X1   g3578(.A(new_n1160_), .B(new_n848_), .Y(new_n3964_));
  OAI21X1  g3579(.A0(new_n3964_), .A1(new_n1477_), .B0(new_n856_), .Y(new_n3965_));
  AOI21X1  g3580(.A0(new_n3965_), .A1(new_n1475_), .B0(new_n1476_), .Y(new_n3966_));
  OAI21X1  g3581(.A0(new_n3966_), .A1(new_n1474_), .B0(new_n871_), .Y(new_n3967_));
  AOI21X1  g3582(.A0(new_n3967_), .A1(new_n1472_), .B0(new_n1473_), .Y(new_n3968_));
  OAI21X1  g3583(.A0(new_n3968_), .A1(new_n1471_), .B0(new_n886_), .Y(new_n3969_));
  AOI21X1  g3584(.A0(new_n3969_), .A1(new_n1469_), .B0(new_n1470_), .Y(new_n3970_));
  OAI21X1  g3585(.A0(new_n3970_), .A1(new_n1468_), .B0(new_n901_), .Y(new_n3971_));
  AOI21X1  g3586(.A0(new_n3971_), .A1(new_n1466_), .B0(new_n1467_), .Y(new_n3972_));
  OAI21X1  g3587(.A0(new_n3972_), .A1(new_n1465_), .B0(new_n916_), .Y(new_n3973_));
  AOI21X1  g3588(.A0(new_n3973_), .A1(new_n1463_), .B0(new_n1464_), .Y(new_n3974_));
  OAI21X1  g3589(.A0(new_n3974_), .A1(new_n1462_), .B0(new_n931_), .Y(new_n3975_));
  AOI21X1  g3590(.A0(new_n3975_), .A1(new_n1460_), .B0(new_n1461_), .Y(new_n3976_));
  OAI21X1  g3591(.A0(new_n3976_), .A1(new_n1459_), .B0(new_n946_), .Y(new_n3977_));
  AOI21X1  g3592(.A0(new_n3977_), .A1(new_n1457_), .B0(new_n1458_), .Y(new_n3978_));
  OAI21X1  g3593(.A0(new_n3978_), .A1(new_n1456_), .B0(new_n961_), .Y(new_n3979_));
  AOI21X1  g3594(.A0(new_n3979_), .A1(new_n1454_), .B0(new_n1455_), .Y(new_n3980_));
  OAI21X1  g3595(.A0(new_n3980_), .A1(new_n1453_), .B0(new_n976_), .Y(new_n3981_));
  AOI21X1  g3596(.A0(new_n3981_), .A1(new_n1451_), .B0(new_n1452_), .Y(new_n3982_));
  OAI21X1  g3597(.A0(new_n3982_), .A1(new_n1450_), .B0(new_n991_), .Y(new_n3983_));
  AOI21X1  g3598(.A0(new_n3983_), .A1(new_n1448_), .B0(new_n1449_), .Y(new_n3984_));
  OAI21X1  g3599(.A0(new_n3984_), .A1(new_n1447_), .B0(new_n1006_), .Y(new_n3985_));
  AOI21X1  g3600(.A0(new_n3985_), .A1(new_n1445_), .B0(new_n1446_), .Y(new_n3986_));
  OAI21X1  g3601(.A0(new_n3986_), .A1(new_n1444_), .B0(new_n1547_), .Y(new_n3987_));
  AOI21X1  g3602(.A0(new_n3987_), .A1(new_n1549_), .B0(new_n1848_), .Y(new_n3988_));
  OAI21X1  g3603(.A0(new_n3988_), .A1(new_n1026_), .B0(new_n1028_), .Y(new_n3989_));
  AOI21X1  g3604(.A0(new_n3989_), .A1(new_n1033_), .B0(new_n1036_), .Y(new_n3990_));
  OAI21X1  g3605(.A0(new_n3990_), .A1(new_n1041_), .B0(new_n1043_), .Y(new_n3991_));
  AOI21X1  g3606(.A0(new_n3991_), .A1(new_n1048_), .B0(new_n1051_), .Y(new_n3992_));
  OAI21X1  g3607(.A0(new_n3992_), .A1(new_n1056_), .B0(new_n1058_), .Y(new_n3993_));
  AOI21X1  g3608(.A0(new_n3993_), .A1(new_n1063_), .B0(new_n1066_), .Y(new_n3994_));
  OAI21X1  g3609(.A0(new_n3994_), .A1(new_n1071_), .B0(new_n1073_), .Y(new_n3995_));
  AOI21X1  g3610(.A0(new_n3995_), .A1(new_n1078_), .B0(new_n1081_), .Y(new_n3996_));
  OAI21X1  g3611(.A0(new_n3996_), .A1(new_n1086_), .B0(new_n1088_), .Y(new_n3997_));
  AOI21X1  g3612(.A0(new_n3997_), .A1(new_n1093_), .B0(new_n1096_), .Y(new_n3998_));
  OAI21X1  g3613(.A0(new_n3998_), .A1(new_n1101_), .B0(new_n1103_), .Y(new_n3999_));
  AOI21X1  g3614(.A0(new_n3999_), .A1(new_n1108_), .B0(new_n1111_), .Y(new_n4000_));
  OAI21X1  g3615(.A0(new_n4000_), .A1(new_n1116_), .B0(new_n1118_), .Y(new_n4001_));
  AOI21X1  g3616(.A0(new_n4001_), .A1(new_n1123_), .B0(new_n1126_), .Y(new_n4002_));
  OAI21X1  g3617(.A0(new_n4002_), .A1(new_n1131_), .B0(new_n1133_), .Y(new_n4003_));
  AOI21X1  g3618(.A0(new_n4003_), .A1(new_n1138_), .B0(new_n1141_), .Y(new_n4004_));
  OAI21X1  g3619(.A0(new_n4004_), .A1(new_n1146_), .B0(new_n1148_), .Y(new_n4005_));
  OAI21X1  g3620(.A0(new_n527_), .A1(\priority[58] ), .B0(\req[58] ), .Y(new_n4006_));
  AOI21X1  g3621(.A0(new_n4005_), .A1(new_n1153_), .B0(new_n4006_), .Y(\grant[58] ));
  NOR2X1   g3622(.A(new_n1162_), .B(new_n535_), .Y(new_n4008_));
  OAI21X1  g3623(.A0(new_n4008_), .A1(new_n1586_), .B0(new_n1170_), .Y(new_n4009_));
  AOI21X1  g3624(.A0(new_n4009_), .A1(new_n1584_), .B0(new_n1585_), .Y(new_n4010_));
  OAI21X1  g3625(.A0(new_n4010_), .A1(new_n1583_), .B0(new_n1185_), .Y(new_n4011_));
  AOI21X1  g3626(.A0(new_n4011_), .A1(new_n1581_), .B0(new_n1582_), .Y(new_n4012_));
  OAI21X1  g3627(.A0(new_n4012_), .A1(new_n1580_), .B0(new_n1200_), .Y(new_n4013_));
  AOI21X1  g3628(.A0(new_n4013_), .A1(new_n1578_), .B0(new_n1579_), .Y(new_n4014_));
  OAI21X1  g3629(.A0(new_n4014_), .A1(new_n1577_), .B0(new_n1215_), .Y(new_n4015_));
  AOI21X1  g3630(.A0(new_n4015_), .A1(new_n1575_), .B0(new_n1576_), .Y(new_n4016_));
  OAI21X1  g3631(.A0(new_n4016_), .A1(new_n1574_), .B0(new_n1230_), .Y(new_n4017_));
  AOI21X1  g3632(.A0(new_n4017_), .A1(new_n1572_), .B0(new_n1573_), .Y(new_n4018_));
  OAI21X1  g3633(.A0(new_n4018_), .A1(new_n1571_), .B0(new_n1245_), .Y(new_n4019_));
  AOI21X1  g3634(.A0(new_n4019_), .A1(new_n1569_), .B0(new_n1570_), .Y(new_n4020_));
  OAI21X1  g3635(.A0(new_n4020_), .A1(new_n1568_), .B0(new_n1260_), .Y(new_n4021_));
  AOI21X1  g3636(.A0(new_n4021_), .A1(new_n1566_), .B0(new_n1567_), .Y(new_n4022_));
  OAI21X1  g3637(.A0(new_n4022_), .A1(new_n1565_), .B0(new_n1275_), .Y(new_n4023_));
  AOI21X1  g3638(.A0(new_n4023_), .A1(new_n1563_), .B0(new_n1564_), .Y(new_n4024_));
  OAI21X1  g3639(.A0(new_n4024_), .A1(new_n1562_), .B0(new_n1290_), .Y(new_n4025_));
  AOI21X1  g3640(.A0(new_n4025_), .A1(new_n1560_), .B0(new_n1561_), .Y(new_n4026_));
  OAI21X1  g3641(.A0(new_n4026_), .A1(new_n1559_), .B0(new_n1305_), .Y(new_n4027_));
  AOI21X1  g3642(.A0(new_n4027_), .A1(new_n1557_), .B0(new_n1558_), .Y(new_n4028_));
  OAI21X1  g3643(.A0(new_n4028_), .A1(new_n1556_), .B0(new_n1320_), .Y(new_n4029_));
  AOI21X1  g3644(.A0(new_n4029_), .A1(new_n1554_), .B0(new_n1555_), .Y(new_n4030_));
  OAI21X1  g3645(.A0(new_n4030_), .A1(new_n1553_), .B0(new_n1656_), .Y(new_n4031_));
  AOI21X1  g3646(.A0(new_n4031_), .A1(new_n1552_), .B0(new_n1893_), .Y(new_n4032_));
  OAI21X1  g3647(.A0(new_n4032_), .A1(new_n1395_), .B0(new_n403_), .Y(new_n4033_));
  AOI21X1  g3648(.A0(new_n4033_), .A1(new_n1393_), .B0(new_n1394_), .Y(new_n4034_));
  OAI21X1  g3649(.A0(new_n4034_), .A1(new_n1392_), .B0(new_n418_), .Y(new_n4035_));
  AOI21X1  g3650(.A0(new_n4035_), .A1(new_n1390_), .B0(new_n1391_), .Y(new_n4036_));
  OAI21X1  g3651(.A0(new_n4036_), .A1(new_n1389_), .B0(new_n433_), .Y(new_n4037_));
  AOI21X1  g3652(.A0(new_n4037_), .A1(new_n1387_), .B0(new_n1388_), .Y(new_n4038_));
  OAI21X1  g3653(.A0(new_n4038_), .A1(new_n1386_), .B0(new_n448_), .Y(new_n4039_));
  AOI21X1  g3654(.A0(new_n4039_), .A1(new_n1384_), .B0(new_n1385_), .Y(new_n4040_));
  OAI21X1  g3655(.A0(new_n4040_), .A1(new_n1383_), .B0(new_n463_), .Y(new_n4041_));
  AOI21X1  g3656(.A0(new_n4041_), .A1(new_n1381_), .B0(new_n1382_), .Y(new_n4042_));
  OAI21X1  g3657(.A0(new_n4042_), .A1(new_n1380_), .B0(new_n478_), .Y(new_n4043_));
  AOI21X1  g3658(.A0(new_n4043_), .A1(new_n1378_), .B0(new_n1379_), .Y(new_n4044_));
  OAI21X1  g3659(.A0(new_n4044_), .A1(new_n1377_), .B0(new_n493_), .Y(new_n4045_));
  AOI21X1  g3660(.A0(new_n4045_), .A1(new_n1375_), .B0(new_n1376_), .Y(new_n4046_));
  OAI21X1  g3661(.A0(new_n4046_), .A1(new_n1374_), .B0(new_n508_), .Y(new_n4047_));
  AOI21X1  g3662(.A0(new_n4047_), .A1(new_n1372_), .B0(new_n1373_), .Y(new_n4048_));
  OAI21X1  g3663(.A0(new_n4048_), .A1(new_n1371_), .B0(new_n523_), .Y(new_n4049_));
  OAI21X1  g3664(.A0(new_n845_), .A1(\priority[59] ), .B0(\req[59] ), .Y(new_n4050_));
  AOI21X1  g3665(.A0(new_n4049_), .A1(new_n1369_), .B0(new_n4050_), .Y(\grant[59] ));
  NOR2X1   g3666(.A(new_n853_), .B(new_n537_), .Y(new_n4052_));
  OAI21X1  g3667(.A0(new_n4052_), .A1(new_n544_), .B0(new_n546_), .Y(new_n4053_));
  AOI21X1  g3668(.A0(new_n4053_), .A1(new_n551_), .B0(new_n554_), .Y(new_n4054_));
  OAI21X1  g3669(.A0(new_n4054_), .A1(new_n559_), .B0(new_n561_), .Y(new_n4055_));
  AOI21X1  g3670(.A0(new_n4055_), .A1(new_n566_), .B0(new_n569_), .Y(new_n4056_));
  OAI21X1  g3671(.A0(new_n4056_), .A1(new_n574_), .B0(new_n576_), .Y(new_n4057_));
  AOI21X1  g3672(.A0(new_n4057_), .A1(new_n581_), .B0(new_n584_), .Y(new_n4058_));
  OAI21X1  g3673(.A0(new_n4058_), .A1(new_n589_), .B0(new_n591_), .Y(new_n4059_));
  AOI21X1  g3674(.A0(new_n4059_), .A1(new_n596_), .B0(new_n599_), .Y(new_n4060_));
  OAI21X1  g3675(.A0(new_n4060_), .A1(new_n604_), .B0(new_n606_), .Y(new_n4061_));
  AOI21X1  g3676(.A0(new_n4061_), .A1(new_n611_), .B0(new_n614_), .Y(new_n4062_));
  OAI21X1  g3677(.A0(new_n4062_), .A1(new_n619_), .B0(new_n621_), .Y(new_n4063_));
  AOI21X1  g3678(.A0(new_n4063_), .A1(new_n626_), .B0(new_n629_), .Y(new_n4064_));
  OAI21X1  g3679(.A0(new_n4064_), .A1(new_n634_), .B0(new_n636_), .Y(new_n4065_));
  AOI21X1  g3680(.A0(new_n4065_), .A1(new_n641_), .B0(new_n644_), .Y(new_n4066_));
  OAI21X1  g3681(.A0(new_n4066_), .A1(new_n649_), .B0(new_n651_), .Y(new_n4067_));
  AOI21X1  g3682(.A0(new_n4067_), .A1(new_n656_), .B0(new_n659_), .Y(new_n4068_));
  OAI21X1  g3683(.A0(new_n4068_), .A1(new_n664_), .B0(new_n666_), .Y(new_n4069_));
  AOI21X1  g3684(.A0(new_n4069_), .A1(new_n671_), .B0(new_n674_), .Y(new_n4070_));
  OAI21X1  g3685(.A0(new_n4070_), .A1(new_n679_), .B0(new_n681_), .Y(new_n4071_));
  AOI21X1  g3686(.A0(new_n4071_), .A1(new_n686_), .B0(new_n689_), .Y(new_n4072_));
  OAI21X1  g3687(.A0(new_n4072_), .A1(new_n694_), .B0(new_n696_), .Y(new_n4073_));
  AOI21X1  g3688(.A0(new_n4073_), .A1(new_n701_), .B0(new_n1662_), .Y(new_n4074_));
  OAI21X1  g3689(.A0(new_n4074_), .A1(new_n1661_), .B0(new_n1705_), .Y(new_n4075_));
  AOI21X1  g3690(.A0(new_n4075_), .A1(new_n1660_), .B0(new_n1938_), .Y(new_n4076_));
  OAI21X1  g3691(.A0(new_n4076_), .A1(new_n1504_), .B0(new_n721_), .Y(new_n4077_));
  AOI21X1  g3692(.A0(new_n4077_), .A1(new_n1502_), .B0(new_n1503_), .Y(new_n4078_));
  OAI21X1  g3693(.A0(new_n4078_), .A1(new_n1501_), .B0(new_n736_), .Y(new_n4079_));
  AOI21X1  g3694(.A0(new_n4079_), .A1(new_n1499_), .B0(new_n1500_), .Y(new_n4080_));
  OAI21X1  g3695(.A0(new_n4080_), .A1(new_n1498_), .B0(new_n751_), .Y(new_n4081_));
  AOI21X1  g3696(.A0(new_n4081_), .A1(new_n1496_), .B0(new_n1497_), .Y(new_n4082_));
  OAI21X1  g3697(.A0(new_n4082_), .A1(new_n1495_), .B0(new_n766_), .Y(new_n4083_));
  AOI21X1  g3698(.A0(new_n4083_), .A1(new_n1493_), .B0(new_n1494_), .Y(new_n4084_));
  OAI21X1  g3699(.A0(new_n4084_), .A1(new_n1492_), .B0(new_n781_), .Y(new_n4085_));
  AOI21X1  g3700(.A0(new_n4085_), .A1(new_n1490_), .B0(new_n1491_), .Y(new_n4086_));
  OAI21X1  g3701(.A0(new_n4086_), .A1(new_n1489_), .B0(new_n796_), .Y(new_n4087_));
  AOI21X1  g3702(.A0(new_n4087_), .A1(new_n1487_), .B0(new_n1488_), .Y(new_n4088_));
  OAI21X1  g3703(.A0(new_n4088_), .A1(new_n1486_), .B0(new_n811_), .Y(new_n4089_));
  AOI21X1  g3704(.A0(new_n4089_), .A1(new_n1484_), .B0(new_n1485_), .Y(new_n4090_));
  OAI21X1  g3705(.A0(new_n4090_), .A1(new_n1483_), .B0(new_n826_), .Y(new_n4091_));
  AOI21X1  g3706(.A0(new_n4091_), .A1(new_n1481_), .B0(new_n1482_), .Y(new_n4092_));
  OAI21X1  g3707(.A0(new_n4092_), .A1(new_n1480_), .B0(new_n841_), .Y(new_n4093_));
  OAI21X1  g3708(.A0(new_n1159_), .A1(\priority[60] ), .B0(\req[60] ), .Y(new_n4094_));
  AOI21X1  g3709(.A0(new_n4093_), .A1(new_n1478_), .B0(new_n4094_), .Y(\grant[60] ));
  NOR2X1   g3710(.A(new_n1167_), .B(new_n855_), .Y(new_n4096_));
  OAI21X1  g3711(.A0(new_n4096_), .A1(new_n862_), .B0(new_n864_), .Y(new_n4097_));
  AOI21X1  g3712(.A0(new_n4097_), .A1(new_n869_), .B0(new_n872_), .Y(new_n4098_));
  OAI21X1  g3713(.A0(new_n4098_), .A1(new_n877_), .B0(new_n879_), .Y(new_n4099_));
  AOI21X1  g3714(.A0(new_n4099_), .A1(new_n884_), .B0(new_n887_), .Y(new_n4100_));
  OAI21X1  g3715(.A0(new_n4100_), .A1(new_n892_), .B0(new_n894_), .Y(new_n4101_));
  AOI21X1  g3716(.A0(new_n4101_), .A1(new_n899_), .B0(new_n902_), .Y(new_n4102_));
  OAI21X1  g3717(.A0(new_n4102_), .A1(new_n907_), .B0(new_n909_), .Y(new_n4103_));
  AOI21X1  g3718(.A0(new_n4103_), .A1(new_n914_), .B0(new_n917_), .Y(new_n4104_));
  OAI21X1  g3719(.A0(new_n4104_), .A1(new_n922_), .B0(new_n924_), .Y(new_n4105_));
  AOI21X1  g3720(.A0(new_n4105_), .A1(new_n929_), .B0(new_n932_), .Y(new_n4106_));
  OAI21X1  g3721(.A0(new_n4106_), .A1(new_n937_), .B0(new_n939_), .Y(new_n4107_));
  AOI21X1  g3722(.A0(new_n4107_), .A1(new_n944_), .B0(new_n947_), .Y(new_n4108_));
  OAI21X1  g3723(.A0(new_n4108_), .A1(new_n952_), .B0(new_n954_), .Y(new_n4109_));
  AOI21X1  g3724(.A0(new_n4109_), .A1(new_n959_), .B0(new_n962_), .Y(new_n4110_));
  OAI21X1  g3725(.A0(new_n4110_), .A1(new_n967_), .B0(new_n969_), .Y(new_n4111_));
  AOI21X1  g3726(.A0(new_n4111_), .A1(new_n974_), .B0(new_n977_), .Y(new_n4112_));
  OAI21X1  g3727(.A0(new_n4112_), .A1(new_n982_), .B0(new_n984_), .Y(new_n4113_));
  AOI21X1  g3728(.A0(new_n4113_), .A1(new_n989_), .B0(new_n992_), .Y(new_n4114_));
  OAI21X1  g3729(.A0(new_n4114_), .A1(new_n997_), .B0(new_n999_), .Y(new_n4115_));
  AOI21X1  g3730(.A0(new_n4115_), .A1(new_n1004_), .B0(new_n1007_), .Y(new_n4116_));
  OAI21X1  g3731(.A0(new_n4116_), .A1(new_n1012_), .B0(new_n1014_), .Y(new_n4117_));
  AOI21X1  g3732(.A0(new_n4117_), .A1(new_n1017_), .B0(new_n1711_), .Y(new_n4118_));
  OAI21X1  g3733(.A0(new_n4118_), .A1(new_n1710_), .B0(new_n1754_), .Y(new_n4119_));
  AOI21X1  g3734(.A0(new_n4119_), .A1(new_n1709_), .B0(new_n1983_), .Y(new_n4120_));
  OAI21X1  g3735(.A0(new_n4120_), .A1(new_n1613_), .B0(new_n1035_), .Y(new_n4121_));
  AOI21X1  g3736(.A0(new_n4121_), .A1(new_n1611_), .B0(new_n1612_), .Y(new_n4122_));
  OAI21X1  g3737(.A0(new_n4122_), .A1(new_n1610_), .B0(new_n1050_), .Y(new_n4123_));
  AOI21X1  g3738(.A0(new_n4123_), .A1(new_n1608_), .B0(new_n1609_), .Y(new_n4124_));
  OAI21X1  g3739(.A0(new_n4124_), .A1(new_n1607_), .B0(new_n1065_), .Y(new_n4125_));
  AOI21X1  g3740(.A0(new_n4125_), .A1(new_n1605_), .B0(new_n1606_), .Y(new_n4126_));
  OAI21X1  g3741(.A0(new_n4126_), .A1(new_n1604_), .B0(new_n1080_), .Y(new_n4127_));
  AOI21X1  g3742(.A0(new_n4127_), .A1(new_n1602_), .B0(new_n1603_), .Y(new_n4128_));
  OAI21X1  g3743(.A0(new_n4128_), .A1(new_n1601_), .B0(new_n1095_), .Y(new_n4129_));
  AOI21X1  g3744(.A0(new_n4129_), .A1(new_n1599_), .B0(new_n1600_), .Y(new_n4130_));
  OAI21X1  g3745(.A0(new_n4130_), .A1(new_n1598_), .B0(new_n1110_), .Y(new_n4131_));
  AOI21X1  g3746(.A0(new_n4131_), .A1(new_n1596_), .B0(new_n1597_), .Y(new_n4132_));
  OAI21X1  g3747(.A0(new_n4132_), .A1(new_n1595_), .B0(new_n1125_), .Y(new_n4133_));
  AOI21X1  g3748(.A0(new_n4133_), .A1(new_n1593_), .B0(new_n1594_), .Y(new_n4134_));
  OAI21X1  g3749(.A0(new_n4134_), .A1(new_n1592_), .B0(new_n1140_), .Y(new_n4135_));
  AOI21X1  g3750(.A0(new_n4135_), .A1(new_n1590_), .B0(new_n1591_), .Y(new_n4136_));
  OAI21X1  g3751(.A0(new_n4136_), .A1(new_n1589_), .B0(new_n1155_), .Y(new_n4137_));
  OAI21X1  g3752(.A0(new_n534_), .A1(\priority[61] ), .B0(\req[61] ), .Y(new_n4138_));
  AOI21X1  g3753(.A0(new_n4137_), .A1(new_n1587_), .B0(new_n4138_), .Y(\grant[61] ));
  NOR2X1   g3754(.A(new_n1169_), .B(new_n543_), .Y(new_n4140_));
  OAI21X1  g3755(.A0(new_n4140_), .A1(new_n1176_), .B0(new_n1178_), .Y(new_n4141_));
  AOI21X1  g3756(.A0(new_n4141_), .A1(new_n1183_), .B0(new_n1186_), .Y(new_n4142_));
  OAI21X1  g3757(.A0(new_n4142_), .A1(new_n1191_), .B0(new_n1193_), .Y(new_n4143_));
  AOI21X1  g3758(.A0(new_n4143_), .A1(new_n1198_), .B0(new_n1201_), .Y(new_n4144_));
  OAI21X1  g3759(.A0(new_n4144_), .A1(new_n1206_), .B0(new_n1208_), .Y(new_n4145_));
  AOI21X1  g3760(.A0(new_n4145_), .A1(new_n1213_), .B0(new_n1216_), .Y(new_n4146_));
  OAI21X1  g3761(.A0(new_n4146_), .A1(new_n1221_), .B0(new_n1223_), .Y(new_n4147_));
  AOI21X1  g3762(.A0(new_n4147_), .A1(new_n1228_), .B0(new_n1231_), .Y(new_n4148_));
  OAI21X1  g3763(.A0(new_n4148_), .A1(new_n1236_), .B0(new_n1238_), .Y(new_n4149_));
  AOI21X1  g3764(.A0(new_n4149_), .A1(new_n1243_), .B0(new_n1246_), .Y(new_n4150_));
  OAI21X1  g3765(.A0(new_n4150_), .A1(new_n1251_), .B0(new_n1253_), .Y(new_n4151_));
  AOI21X1  g3766(.A0(new_n4151_), .A1(new_n1258_), .B0(new_n1261_), .Y(new_n4152_));
  OAI21X1  g3767(.A0(new_n4152_), .A1(new_n1266_), .B0(new_n1268_), .Y(new_n4153_));
  AOI21X1  g3768(.A0(new_n4153_), .A1(new_n1273_), .B0(new_n1276_), .Y(new_n4154_));
  OAI21X1  g3769(.A0(new_n4154_), .A1(new_n1281_), .B0(new_n1283_), .Y(new_n4155_));
  AOI21X1  g3770(.A0(new_n4155_), .A1(new_n1288_), .B0(new_n1291_), .Y(new_n4156_));
  OAI21X1  g3771(.A0(new_n4156_), .A1(new_n1296_), .B0(new_n1298_), .Y(new_n4157_));
  AOI21X1  g3772(.A0(new_n4157_), .A1(new_n1303_), .B0(new_n1306_), .Y(new_n4158_));
  OAI21X1  g3773(.A0(new_n4158_), .A1(new_n1311_), .B0(new_n1313_), .Y(new_n4159_));
  AOI21X1  g3774(.A0(new_n4159_), .A1(new_n1318_), .B0(new_n1321_), .Y(new_n4160_));
  OAI21X1  g3775(.A0(new_n4160_), .A1(new_n1326_), .B0(new_n1328_), .Y(new_n4161_));
  AOI21X1  g3776(.A0(new_n4161_), .A1(new_n1331_), .B0(new_n1758_), .Y(new_n4162_));
  OAI21X1  g3777(.A0(new_n4162_), .A1(new_n394_), .B0(new_n396_), .Y(new_n4163_));
  AOI21X1  g3778(.A0(new_n4163_), .A1(new_n401_), .B0(new_n404_), .Y(new_n4164_));
  OAI21X1  g3779(.A0(new_n4164_), .A1(new_n409_), .B0(new_n411_), .Y(new_n4165_));
  AOI21X1  g3780(.A0(new_n4165_), .A1(new_n416_), .B0(new_n419_), .Y(new_n4166_));
  OAI21X1  g3781(.A0(new_n4166_), .A1(new_n424_), .B0(new_n426_), .Y(new_n4167_));
  AOI21X1  g3782(.A0(new_n4167_), .A1(new_n431_), .B0(new_n434_), .Y(new_n4168_));
  OAI21X1  g3783(.A0(new_n4168_), .A1(new_n439_), .B0(new_n441_), .Y(new_n4169_));
  AOI21X1  g3784(.A0(new_n4169_), .A1(new_n446_), .B0(new_n449_), .Y(new_n4170_));
  OAI21X1  g3785(.A0(new_n4170_), .A1(new_n454_), .B0(new_n456_), .Y(new_n4171_));
  AOI21X1  g3786(.A0(new_n4171_), .A1(new_n461_), .B0(new_n464_), .Y(new_n4172_));
  OAI21X1  g3787(.A0(new_n4172_), .A1(new_n469_), .B0(new_n471_), .Y(new_n4173_));
  AOI21X1  g3788(.A0(new_n4173_), .A1(new_n476_), .B0(new_n479_), .Y(new_n4174_));
  OAI21X1  g3789(.A0(new_n4174_), .A1(new_n484_), .B0(new_n486_), .Y(new_n4175_));
  AOI21X1  g3790(.A0(new_n4175_), .A1(new_n491_), .B0(new_n494_), .Y(new_n4176_));
  OAI21X1  g3791(.A0(new_n4176_), .A1(new_n499_), .B0(new_n501_), .Y(new_n4177_));
  AOI21X1  g3792(.A0(new_n4177_), .A1(new_n506_), .B0(new_n509_), .Y(new_n4178_));
  OAI21X1  g3793(.A0(new_n4178_), .A1(new_n514_), .B0(new_n516_), .Y(new_n4179_));
  AOI21X1  g3794(.A0(new_n4179_), .A1(new_n521_), .B0(new_n524_), .Y(new_n4180_));
  OAI21X1  g3795(.A0(new_n4180_), .A1(new_n529_), .B0(new_n531_), .Y(new_n4181_));
  OAI21X1  g3796(.A0(new_n852_), .A1(\priority[62] ), .B0(\req[62] ), .Y(new_n4182_));
  AOI21X1  g3797(.A0(new_n4181_), .A1(new_n536_), .B0(new_n4182_), .Y(\grant[62] ));
  NOR2X1   g3798(.A(new_n861_), .B(new_n545_), .Y(new_n4184_));
  OAI21X1  g3799(.A0(new_n4184_), .A1(new_n1365_), .B0(new_n553_), .Y(new_n4185_));
  AOI21X1  g3800(.A0(new_n4185_), .A1(new_n1363_), .B0(new_n1364_), .Y(new_n4186_));
  OAI21X1  g3801(.A0(new_n4186_), .A1(new_n1362_), .B0(new_n568_), .Y(new_n4187_));
  AOI21X1  g3802(.A0(new_n4187_), .A1(new_n1360_), .B0(new_n1361_), .Y(new_n4188_));
  OAI21X1  g3803(.A0(new_n4188_), .A1(new_n1359_), .B0(new_n583_), .Y(new_n4189_));
  AOI21X1  g3804(.A0(new_n4189_), .A1(new_n1357_), .B0(new_n1358_), .Y(new_n4190_));
  OAI21X1  g3805(.A0(new_n4190_), .A1(new_n1356_), .B0(new_n598_), .Y(new_n4191_));
  AOI21X1  g3806(.A0(new_n4191_), .A1(new_n1354_), .B0(new_n1355_), .Y(new_n4192_));
  OAI21X1  g3807(.A0(new_n4192_), .A1(new_n1353_), .B0(new_n613_), .Y(new_n4193_));
  AOI21X1  g3808(.A0(new_n4193_), .A1(new_n1351_), .B0(new_n1352_), .Y(new_n4194_));
  OAI21X1  g3809(.A0(new_n4194_), .A1(new_n1350_), .B0(new_n628_), .Y(new_n4195_));
  AOI21X1  g3810(.A0(new_n4195_), .A1(new_n1348_), .B0(new_n1349_), .Y(new_n4196_));
  OAI21X1  g3811(.A0(new_n4196_), .A1(new_n1347_), .B0(new_n643_), .Y(new_n4197_));
  AOI21X1  g3812(.A0(new_n4197_), .A1(new_n1345_), .B0(new_n1346_), .Y(new_n4198_));
  OAI21X1  g3813(.A0(new_n4198_), .A1(new_n1344_), .B0(new_n658_), .Y(new_n4199_));
  AOI21X1  g3814(.A0(new_n4199_), .A1(new_n1342_), .B0(new_n1343_), .Y(new_n4200_));
  OAI21X1  g3815(.A0(new_n4200_), .A1(new_n1341_), .B0(new_n673_), .Y(new_n4201_));
  AOI21X1  g3816(.A0(new_n4201_), .A1(new_n1339_), .B0(new_n1340_), .Y(new_n4202_));
  OAI21X1  g3817(.A0(new_n4202_), .A1(new_n1338_), .B0(new_n688_), .Y(new_n4203_));
  AOI21X1  g3818(.A0(new_n4203_), .A1(new_n1336_), .B0(new_n1337_), .Y(new_n4204_));
  OAI21X1  g3819(.A0(new_n4204_), .A1(new_n1335_), .B0(new_n1438_), .Y(new_n4205_));
  AOI21X1  g3820(.A0(new_n4205_), .A1(new_n1440_), .B0(new_n1803_), .Y(new_n4206_));
  OAI21X1  g3821(.A0(new_n4206_), .A1(new_n712_), .B0(new_n714_), .Y(new_n4207_));
  AOI21X1  g3822(.A0(new_n4207_), .A1(new_n719_), .B0(new_n722_), .Y(new_n4208_));
  OAI21X1  g3823(.A0(new_n4208_), .A1(new_n727_), .B0(new_n729_), .Y(new_n4209_));
  AOI21X1  g3824(.A0(new_n4209_), .A1(new_n734_), .B0(new_n737_), .Y(new_n4210_));
  OAI21X1  g3825(.A0(new_n4210_), .A1(new_n742_), .B0(new_n744_), .Y(new_n4211_));
  AOI21X1  g3826(.A0(new_n4211_), .A1(new_n749_), .B0(new_n752_), .Y(new_n4212_));
  OAI21X1  g3827(.A0(new_n4212_), .A1(new_n757_), .B0(new_n759_), .Y(new_n4213_));
  AOI21X1  g3828(.A0(new_n4213_), .A1(new_n764_), .B0(new_n767_), .Y(new_n4214_));
  OAI21X1  g3829(.A0(new_n4214_), .A1(new_n772_), .B0(new_n774_), .Y(new_n4215_));
  AOI21X1  g3830(.A0(new_n4215_), .A1(new_n779_), .B0(new_n782_), .Y(new_n4216_));
  OAI21X1  g3831(.A0(new_n4216_), .A1(new_n787_), .B0(new_n789_), .Y(new_n4217_));
  AOI21X1  g3832(.A0(new_n4217_), .A1(new_n794_), .B0(new_n797_), .Y(new_n4218_));
  OAI21X1  g3833(.A0(new_n4218_), .A1(new_n802_), .B0(new_n804_), .Y(new_n4219_));
  AOI21X1  g3834(.A0(new_n4219_), .A1(new_n809_), .B0(new_n812_), .Y(new_n4220_));
  OAI21X1  g3835(.A0(new_n4220_), .A1(new_n817_), .B0(new_n819_), .Y(new_n4221_));
  AOI21X1  g3836(.A0(new_n4221_), .A1(new_n824_), .B0(new_n827_), .Y(new_n4222_));
  OAI21X1  g3837(.A0(new_n4222_), .A1(new_n832_), .B0(new_n834_), .Y(new_n4223_));
  AOI21X1  g3838(.A0(new_n4223_), .A1(new_n839_), .B0(new_n842_), .Y(new_n4224_));
  OAI21X1  g3839(.A0(new_n4224_), .A1(new_n847_), .B0(new_n849_), .Y(new_n4225_));
  OAI21X1  g3840(.A0(new_n1166_), .A1(\priority[63] ), .B0(\req[63] ), .Y(new_n4226_));
  AOI21X1  g3841(.A0(new_n4225_), .A1(new_n854_), .B0(new_n4226_), .Y(\grant[63] ));
  NOR2X1   g3842(.A(new_n1175_), .B(new_n863_), .Y(new_n4228_));
  OAI21X1  g3843(.A0(new_n4228_), .A1(new_n1474_), .B0(new_n871_), .Y(new_n4229_));
  AOI21X1  g3844(.A0(new_n4229_), .A1(new_n1472_), .B0(new_n1473_), .Y(new_n4230_));
  OAI21X1  g3845(.A0(new_n4230_), .A1(new_n1471_), .B0(new_n886_), .Y(new_n4231_));
  AOI21X1  g3846(.A0(new_n4231_), .A1(new_n1469_), .B0(new_n1470_), .Y(new_n4232_));
  OAI21X1  g3847(.A0(new_n4232_), .A1(new_n1468_), .B0(new_n901_), .Y(new_n4233_));
  AOI21X1  g3848(.A0(new_n4233_), .A1(new_n1466_), .B0(new_n1467_), .Y(new_n4234_));
  OAI21X1  g3849(.A0(new_n4234_), .A1(new_n1465_), .B0(new_n916_), .Y(new_n4235_));
  AOI21X1  g3850(.A0(new_n4235_), .A1(new_n1463_), .B0(new_n1464_), .Y(new_n4236_));
  OAI21X1  g3851(.A0(new_n4236_), .A1(new_n1462_), .B0(new_n931_), .Y(new_n4237_));
  AOI21X1  g3852(.A0(new_n4237_), .A1(new_n1460_), .B0(new_n1461_), .Y(new_n4238_));
  OAI21X1  g3853(.A0(new_n4238_), .A1(new_n1459_), .B0(new_n946_), .Y(new_n4239_));
  AOI21X1  g3854(.A0(new_n4239_), .A1(new_n1457_), .B0(new_n1458_), .Y(new_n4240_));
  OAI21X1  g3855(.A0(new_n4240_), .A1(new_n1456_), .B0(new_n961_), .Y(new_n4241_));
  AOI21X1  g3856(.A0(new_n4241_), .A1(new_n1454_), .B0(new_n1455_), .Y(new_n4242_));
  OAI21X1  g3857(.A0(new_n4242_), .A1(new_n1453_), .B0(new_n976_), .Y(new_n4243_));
  AOI21X1  g3858(.A0(new_n4243_), .A1(new_n1451_), .B0(new_n1452_), .Y(new_n4244_));
  OAI21X1  g3859(.A0(new_n4244_), .A1(new_n1450_), .B0(new_n991_), .Y(new_n4245_));
  AOI21X1  g3860(.A0(new_n4245_), .A1(new_n1448_), .B0(new_n1449_), .Y(new_n4246_));
  OAI21X1  g3861(.A0(new_n4246_), .A1(new_n1447_), .B0(new_n1006_), .Y(new_n4247_));
  AOI21X1  g3862(.A0(new_n4247_), .A1(new_n1445_), .B0(new_n1446_), .Y(new_n4248_));
  OAI21X1  g3863(.A0(new_n4248_), .A1(new_n1444_), .B0(new_n1547_), .Y(new_n4249_));
  AOI21X1  g3864(.A0(new_n4249_), .A1(new_n1549_), .B0(new_n1848_), .Y(new_n4250_));
  OAI21X1  g3865(.A0(new_n4250_), .A1(new_n1026_), .B0(new_n1028_), .Y(new_n4251_));
  AOI21X1  g3866(.A0(new_n4251_), .A1(new_n1033_), .B0(new_n1036_), .Y(new_n4252_));
  OAI21X1  g3867(.A0(new_n4252_), .A1(new_n1041_), .B0(new_n1043_), .Y(new_n4253_));
  AOI21X1  g3868(.A0(new_n4253_), .A1(new_n1048_), .B0(new_n1051_), .Y(new_n4254_));
  OAI21X1  g3869(.A0(new_n4254_), .A1(new_n1056_), .B0(new_n1058_), .Y(new_n4255_));
  AOI21X1  g3870(.A0(new_n4255_), .A1(new_n1063_), .B0(new_n1066_), .Y(new_n4256_));
  OAI21X1  g3871(.A0(new_n4256_), .A1(new_n1071_), .B0(new_n1073_), .Y(new_n4257_));
  AOI21X1  g3872(.A0(new_n4257_), .A1(new_n1078_), .B0(new_n1081_), .Y(new_n4258_));
  OAI21X1  g3873(.A0(new_n4258_), .A1(new_n1086_), .B0(new_n1088_), .Y(new_n4259_));
  AOI21X1  g3874(.A0(new_n4259_), .A1(new_n1093_), .B0(new_n1096_), .Y(new_n4260_));
  OAI21X1  g3875(.A0(new_n4260_), .A1(new_n1101_), .B0(new_n1103_), .Y(new_n4261_));
  AOI21X1  g3876(.A0(new_n4261_), .A1(new_n1108_), .B0(new_n1111_), .Y(new_n4262_));
  OAI21X1  g3877(.A0(new_n4262_), .A1(new_n1116_), .B0(new_n1118_), .Y(new_n4263_));
  AOI21X1  g3878(.A0(new_n4263_), .A1(new_n1123_), .B0(new_n1126_), .Y(new_n4264_));
  OAI21X1  g3879(.A0(new_n4264_), .A1(new_n1131_), .B0(new_n1133_), .Y(new_n4265_));
  AOI21X1  g3880(.A0(new_n4265_), .A1(new_n1138_), .B0(new_n1141_), .Y(new_n4266_));
  OAI21X1  g3881(.A0(new_n4266_), .A1(new_n1146_), .B0(new_n1148_), .Y(new_n4267_));
  AOI21X1  g3882(.A0(new_n4267_), .A1(new_n1153_), .B0(new_n1156_), .Y(new_n4268_));
  OAI21X1  g3883(.A0(new_n4268_), .A1(new_n1161_), .B0(new_n1163_), .Y(new_n4269_));
  OAI21X1  g3884(.A0(new_n542_), .A1(\priority[64] ), .B0(\req[64] ), .Y(new_n4270_));
  AOI21X1  g3885(.A0(new_n4269_), .A1(new_n1168_), .B0(new_n4270_), .Y(\grant[64] ));
  NOR2X1   g3886(.A(new_n1177_), .B(new_n550_), .Y(new_n4272_));
  OAI21X1  g3887(.A0(new_n4272_), .A1(new_n1583_), .B0(new_n1185_), .Y(new_n4273_));
  AOI21X1  g3888(.A0(new_n4273_), .A1(new_n1581_), .B0(new_n1582_), .Y(new_n4274_));
  OAI21X1  g3889(.A0(new_n4274_), .A1(new_n1580_), .B0(new_n1200_), .Y(new_n4275_));
  AOI21X1  g3890(.A0(new_n4275_), .A1(new_n1578_), .B0(new_n1579_), .Y(new_n4276_));
  OAI21X1  g3891(.A0(new_n4276_), .A1(new_n1577_), .B0(new_n1215_), .Y(new_n4277_));
  AOI21X1  g3892(.A0(new_n4277_), .A1(new_n1575_), .B0(new_n1576_), .Y(new_n4278_));
  OAI21X1  g3893(.A0(new_n4278_), .A1(new_n1574_), .B0(new_n1230_), .Y(new_n4279_));
  AOI21X1  g3894(.A0(new_n4279_), .A1(new_n1572_), .B0(new_n1573_), .Y(new_n4280_));
  OAI21X1  g3895(.A0(new_n4280_), .A1(new_n1571_), .B0(new_n1245_), .Y(new_n4281_));
  AOI21X1  g3896(.A0(new_n4281_), .A1(new_n1569_), .B0(new_n1570_), .Y(new_n4282_));
  OAI21X1  g3897(.A0(new_n4282_), .A1(new_n1568_), .B0(new_n1260_), .Y(new_n4283_));
  AOI21X1  g3898(.A0(new_n4283_), .A1(new_n1566_), .B0(new_n1567_), .Y(new_n4284_));
  OAI21X1  g3899(.A0(new_n4284_), .A1(new_n1565_), .B0(new_n1275_), .Y(new_n4285_));
  AOI21X1  g3900(.A0(new_n4285_), .A1(new_n1563_), .B0(new_n1564_), .Y(new_n4286_));
  OAI21X1  g3901(.A0(new_n4286_), .A1(new_n1562_), .B0(new_n1290_), .Y(new_n4287_));
  AOI21X1  g3902(.A0(new_n4287_), .A1(new_n1560_), .B0(new_n1561_), .Y(new_n4288_));
  OAI21X1  g3903(.A0(new_n4288_), .A1(new_n1559_), .B0(new_n1305_), .Y(new_n4289_));
  AOI21X1  g3904(.A0(new_n4289_), .A1(new_n1557_), .B0(new_n1558_), .Y(new_n4290_));
  OAI21X1  g3905(.A0(new_n4290_), .A1(new_n1556_), .B0(new_n1320_), .Y(new_n4291_));
  AOI21X1  g3906(.A0(new_n4291_), .A1(new_n1554_), .B0(new_n1555_), .Y(new_n4292_));
  OAI21X1  g3907(.A0(new_n4292_), .A1(new_n1553_), .B0(new_n1656_), .Y(new_n4293_));
  AOI21X1  g3908(.A0(new_n4293_), .A1(new_n1552_), .B0(new_n1893_), .Y(new_n4294_));
  OAI21X1  g3909(.A0(new_n4294_), .A1(new_n1395_), .B0(new_n403_), .Y(new_n4295_));
  AOI21X1  g3910(.A0(new_n4295_), .A1(new_n1393_), .B0(new_n1394_), .Y(new_n4296_));
  OAI21X1  g3911(.A0(new_n4296_), .A1(new_n1392_), .B0(new_n418_), .Y(new_n4297_));
  AOI21X1  g3912(.A0(new_n4297_), .A1(new_n1390_), .B0(new_n1391_), .Y(new_n4298_));
  OAI21X1  g3913(.A0(new_n4298_), .A1(new_n1389_), .B0(new_n433_), .Y(new_n4299_));
  AOI21X1  g3914(.A0(new_n4299_), .A1(new_n1387_), .B0(new_n1388_), .Y(new_n4300_));
  OAI21X1  g3915(.A0(new_n4300_), .A1(new_n1386_), .B0(new_n448_), .Y(new_n4301_));
  AOI21X1  g3916(.A0(new_n4301_), .A1(new_n1384_), .B0(new_n1385_), .Y(new_n4302_));
  OAI21X1  g3917(.A0(new_n4302_), .A1(new_n1383_), .B0(new_n463_), .Y(new_n4303_));
  AOI21X1  g3918(.A0(new_n4303_), .A1(new_n1381_), .B0(new_n1382_), .Y(new_n4304_));
  OAI21X1  g3919(.A0(new_n4304_), .A1(new_n1380_), .B0(new_n478_), .Y(new_n4305_));
  AOI21X1  g3920(.A0(new_n4305_), .A1(new_n1378_), .B0(new_n1379_), .Y(new_n4306_));
  OAI21X1  g3921(.A0(new_n4306_), .A1(new_n1377_), .B0(new_n493_), .Y(new_n4307_));
  AOI21X1  g3922(.A0(new_n4307_), .A1(new_n1375_), .B0(new_n1376_), .Y(new_n4308_));
  OAI21X1  g3923(.A0(new_n4308_), .A1(new_n1374_), .B0(new_n508_), .Y(new_n4309_));
  AOI21X1  g3924(.A0(new_n4309_), .A1(new_n1372_), .B0(new_n1373_), .Y(new_n4310_));
  OAI21X1  g3925(.A0(new_n4310_), .A1(new_n1371_), .B0(new_n523_), .Y(new_n4311_));
  AOI21X1  g3926(.A0(new_n4311_), .A1(new_n1369_), .B0(new_n1370_), .Y(new_n4312_));
  OAI21X1  g3927(.A0(new_n4312_), .A1(new_n1368_), .B0(new_n538_), .Y(new_n4313_));
  OAI21X1  g3928(.A0(new_n860_), .A1(\priority[65] ), .B0(\req[65] ), .Y(new_n4314_));
  AOI21X1  g3929(.A0(new_n4313_), .A1(new_n1366_), .B0(new_n4314_), .Y(\grant[65] ));
  NOR2X1   g3930(.A(new_n868_), .B(new_n552_), .Y(new_n4316_));
  OAI21X1  g3931(.A0(new_n4316_), .A1(new_n559_), .B0(new_n561_), .Y(new_n4317_));
  AOI21X1  g3932(.A0(new_n4317_), .A1(new_n566_), .B0(new_n569_), .Y(new_n4318_));
  OAI21X1  g3933(.A0(new_n4318_), .A1(new_n574_), .B0(new_n576_), .Y(new_n4319_));
  AOI21X1  g3934(.A0(new_n4319_), .A1(new_n581_), .B0(new_n584_), .Y(new_n4320_));
  OAI21X1  g3935(.A0(new_n4320_), .A1(new_n589_), .B0(new_n591_), .Y(new_n4321_));
  AOI21X1  g3936(.A0(new_n4321_), .A1(new_n596_), .B0(new_n599_), .Y(new_n4322_));
  OAI21X1  g3937(.A0(new_n4322_), .A1(new_n604_), .B0(new_n606_), .Y(new_n4323_));
  AOI21X1  g3938(.A0(new_n4323_), .A1(new_n611_), .B0(new_n614_), .Y(new_n4324_));
  OAI21X1  g3939(.A0(new_n4324_), .A1(new_n619_), .B0(new_n621_), .Y(new_n4325_));
  AOI21X1  g3940(.A0(new_n4325_), .A1(new_n626_), .B0(new_n629_), .Y(new_n4326_));
  OAI21X1  g3941(.A0(new_n4326_), .A1(new_n634_), .B0(new_n636_), .Y(new_n4327_));
  AOI21X1  g3942(.A0(new_n4327_), .A1(new_n641_), .B0(new_n644_), .Y(new_n4328_));
  OAI21X1  g3943(.A0(new_n4328_), .A1(new_n649_), .B0(new_n651_), .Y(new_n4329_));
  AOI21X1  g3944(.A0(new_n4329_), .A1(new_n656_), .B0(new_n659_), .Y(new_n4330_));
  OAI21X1  g3945(.A0(new_n4330_), .A1(new_n664_), .B0(new_n666_), .Y(new_n4331_));
  AOI21X1  g3946(.A0(new_n4331_), .A1(new_n671_), .B0(new_n674_), .Y(new_n4332_));
  OAI21X1  g3947(.A0(new_n4332_), .A1(new_n679_), .B0(new_n681_), .Y(new_n4333_));
  AOI21X1  g3948(.A0(new_n4333_), .A1(new_n686_), .B0(new_n689_), .Y(new_n4334_));
  OAI21X1  g3949(.A0(new_n4334_), .A1(new_n694_), .B0(new_n696_), .Y(new_n4335_));
  AOI21X1  g3950(.A0(new_n4335_), .A1(new_n701_), .B0(new_n1662_), .Y(new_n4336_));
  OAI21X1  g3951(.A0(new_n4336_), .A1(new_n1661_), .B0(new_n1705_), .Y(new_n4337_));
  AOI21X1  g3952(.A0(new_n4337_), .A1(new_n1660_), .B0(new_n1938_), .Y(new_n4338_));
  OAI21X1  g3953(.A0(new_n4338_), .A1(new_n1504_), .B0(new_n721_), .Y(new_n4339_));
  AOI21X1  g3954(.A0(new_n4339_), .A1(new_n1502_), .B0(new_n1503_), .Y(new_n4340_));
  OAI21X1  g3955(.A0(new_n4340_), .A1(new_n1501_), .B0(new_n736_), .Y(new_n4341_));
  AOI21X1  g3956(.A0(new_n4341_), .A1(new_n1499_), .B0(new_n1500_), .Y(new_n4342_));
  OAI21X1  g3957(.A0(new_n4342_), .A1(new_n1498_), .B0(new_n751_), .Y(new_n4343_));
  AOI21X1  g3958(.A0(new_n4343_), .A1(new_n1496_), .B0(new_n1497_), .Y(new_n4344_));
  OAI21X1  g3959(.A0(new_n4344_), .A1(new_n1495_), .B0(new_n766_), .Y(new_n4345_));
  AOI21X1  g3960(.A0(new_n4345_), .A1(new_n1493_), .B0(new_n1494_), .Y(new_n4346_));
  OAI21X1  g3961(.A0(new_n4346_), .A1(new_n1492_), .B0(new_n781_), .Y(new_n4347_));
  AOI21X1  g3962(.A0(new_n4347_), .A1(new_n1490_), .B0(new_n1491_), .Y(new_n4348_));
  OAI21X1  g3963(.A0(new_n4348_), .A1(new_n1489_), .B0(new_n796_), .Y(new_n4349_));
  AOI21X1  g3964(.A0(new_n4349_), .A1(new_n1487_), .B0(new_n1488_), .Y(new_n4350_));
  OAI21X1  g3965(.A0(new_n4350_), .A1(new_n1486_), .B0(new_n811_), .Y(new_n4351_));
  AOI21X1  g3966(.A0(new_n4351_), .A1(new_n1484_), .B0(new_n1485_), .Y(new_n4352_));
  OAI21X1  g3967(.A0(new_n4352_), .A1(new_n1483_), .B0(new_n826_), .Y(new_n4353_));
  AOI21X1  g3968(.A0(new_n4353_), .A1(new_n1481_), .B0(new_n1482_), .Y(new_n4354_));
  OAI21X1  g3969(.A0(new_n4354_), .A1(new_n1480_), .B0(new_n841_), .Y(new_n4355_));
  AOI21X1  g3970(.A0(new_n4355_), .A1(new_n1478_), .B0(new_n1479_), .Y(new_n4356_));
  OAI21X1  g3971(.A0(new_n4356_), .A1(new_n1477_), .B0(new_n856_), .Y(new_n4357_));
  OAI21X1  g3972(.A0(new_n1174_), .A1(\priority[66] ), .B0(\req[66] ), .Y(new_n4358_));
  AOI21X1  g3973(.A0(new_n4357_), .A1(new_n1475_), .B0(new_n4358_), .Y(\grant[66] ));
  NOR2X1   g3974(.A(new_n1182_), .B(new_n870_), .Y(new_n4360_));
  OAI21X1  g3975(.A0(new_n4360_), .A1(new_n877_), .B0(new_n879_), .Y(new_n4361_));
  AOI21X1  g3976(.A0(new_n4361_), .A1(new_n884_), .B0(new_n887_), .Y(new_n4362_));
  OAI21X1  g3977(.A0(new_n4362_), .A1(new_n892_), .B0(new_n894_), .Y(new_n4363_));
  AOI21X1  g3978(.A0(new_n4363_), .A1(new_n899_), .B0(new_n902_), .Y(new_n4364_));
  OAI21X1  g3979(.A0(new_n4364_), .A1(new_n907_), .B0(new_n909_), .Y(new_n4365_));
  AOI21X1  g3980(.A0(new_n4365_), .A1(new_n914_), .B0(new_n917_), .Y(new_n4366_));
  OAI21X1  g3981(.A0(new_n4366_), .A1(new_n922_), .B0(new_n924_), .Y(new_n4367_));
  AOI21X1  g3982(.A0(new_n4367_), .A1(new_n929_), .B0(new_n932_), .Y(new_n4368_));
  OAI21X1  g3983(.A0(new_n4368_), .A1(new_n937_), .B0(new_n939_), .Y(new_n4369_));
  AOI21X1  g3984(.A0(new_n4369_), .A1(new_n944_), .B0(new_n947_), .Y(new_n4370_));
  OAI21X1  g3985(.A0(new_n4370_), .A1(new_n952_), .B0(new_n954_), .Y(new_n4371_));
  AOI21X1  g3986(.A0(new_n4371_), .A1(new_n959_), .B0(new_n962_), .Y(new_n4372_));
  OAI21X1  g3987(.A0(new_n4372_), .A1(new_n967_), .B0(new_n969_), .Y(new_n4373_));
  AOI21X1  g3988(.A0(new_n4373_), .A1(new_n974_), .B0(new_n977_), .Y(new_n4374_));
  OAI21X1  g3989(.A0(new_n4374_), .A1(new_n982_), .B0(new_n984_), .Y(new_n4375_));
  AOI21X1  g3990(.A0(new_n4375_), .A1(new_n989_), .B0(new_n992_), .Y(new_n4376_));
  OAI21X1  g3991(.A0(new_n4376_), .A1(new_n997_), .B0(new_n999_), .Y(new_n4377_));
  AOI21X1  g3992(.A0(new_n4377_), .A1(new_n1004_), .B0(new_n1007_), .Y(new_n4378_));
  OAI21X1  g3993(.A0(new_n4378_), .A1(new_n1012_), .B0(new_n1014_), .Y(new_n4379_));
  AOI21X1  g3994(.A0(new_n4379_), .A1(new_n1017_), .B0(new_n1711_), .Y(new_n4380_));
  OAI21X1  g3995(.A0(new_n4380_), .A1(new_n1710_), .B0(new_n1754_), .Y(new_n4381_));
  AOI21X1  g3996(.A0(new_n4381_), .A1(new_n1709_), .B0(new_n1983_), .Y(new_n4382_));
  OAI21X1  g3997(.A0(new_n4382_), .A1(new_n1613_), .B0(new_n1035_), .Y(new_n4383_));
  AOI21X1  g3998(.A0(new_n4383_), .A1(new_n1611_), .B0(new_n1612_), .Y(new_n4384_));
  OAI21X1  g3999(.A0(new_n4384_), .A1(new_n1610_), .B0(new_n1050_), .Y(new_n4385_));
  AOI21X1  g4000(.A0(new_n4385_), .A1(new_n1608_), .B0(new_n1609_), .Y(new_n4386_));
  OAI21X1  g4001(.A0(new_n4386_), .A1(new_n1607_), .B0(new_n1065_), .Y(new_n4387_));
  AOI21X1  g4002(.A0(new_n4387_), .A1(new_n1605_), .B0(new_n1606_), .Y(new_n4388_));
  OAI21X1  g4003(.A0(new_n4388_), .A1(new_n1604_), .B0(new_n1080_), .Y(new_n4389_));
  AOI21X1  g4004(.A0(new_n4389_), .A1(new_n1602_), .B0(new_n1603_), .Y(new_n4390_));
  OAI21X1  g4005(.A0(new_n4390_), .A1(new_n1601_), .B0(new_n1095_), .Y(new_n4391_));
  AOI21X1  g4006(.A0(new_n4391_), .A1(new_n1599_), .B0(new_n1600_), .Y(new_n4392_));
  OAI21X1  g4007(.A0(new_n4392_), .A1(new_n1598_), .B0(new_n1110_), .Y(new_n4393_));
  AOI21X1  g4008(.A0(new_n4393_), .A1(new_n1596_), .B0(new_n1597_), .Y(new_n4394_));
  OAI21X1  g4009(.A0(new_n4394_), .A1(new_n1595_), .B0(new_n1125_), .Y(new_n4395_));
  AOI21X1  g4010(.A0(new_n4395_), .A1(new_n1593_), .B0(new_n1594_), .Y(new_n4396_));
  OAI21X1  g4011(.A0(new_n4396_), .A1(new_n1592_), .B0(new_n1140_), .Y(new_n4397_));
  AOI21X1  g4012(.A0(new_n4397_), .A1(new_n1590_), .B0(new_n1591_), .Y(new_n4398_));
  OAI21X1  g4013(.A0(new_n4398_), .A1(new_n1589_), .B0(new_n1155_), .Y(new_n4399_));
  AOI21X1  g4014(.A0(new_n4399_), .A1(new_n1587_), .B0(new_n1588_), .Y(new_n4400_));
  OAI21X1  g4015(.A0(new_n4400_), .A1(new_n1586_), .B0(new_n1170_), .Y(new_n4401_));
  OAI21X1  g4016(.A0(new_n549_), .A1(\priority[67] ), .B0(\req[67] ), .Y(new_n4402_));
  AOI21X1  g4017(.A0(new_n4401_), .A1(new_n1584_), .B0(new_n4402_), .Y(\grant[67] ));
  NOR2X1   g4018(.A(new_n1184_), .B(new_n558_), .Y(new_n4404_));
  OAI21X1  g4019(.A0(new_n4404_), .A1(new_n1191_), .B0(new_n1193_), .Y(new_n4405_));
  AOI21X1  g4020(.A0(new_n4405_), .A1(new_n1198_), .B0(new_n1201_), .Y(new_n4406_));
  OAI21X1  g4021(.A0(new_n4406_), .A1(new_n1206_), .B0(new_n1208_), .Y(new_n4407_));
  AOI21X1  g4022(.A0(new_n4407_), .A1(new_n1213_), .B0(new_n1216_), .Y(new_n4408_));
  OAI21X1  g4023(.A0(new_n4408_), .A1(new_n1221_), .B0(new_n1223_), .Y(new_n4409_));
  AOI21X1  g4024(.A0(new_n4409_), .A1(new_n1228_), .B0(new_n1231_), .Y(new_n4410_));
  OAI21X1  g4025(.A0(new_n4410_), .A1(new_n1236_), .B0(new_n1238_), .Y(new_n4411_));
  AOI21X1  g4026(.A0(new_n4411_), .A1(new_n1243_), .B0(new_n1246_), .Y(new_n4412_));
  OAI21X1  g4027(.A0(new_n4412_), .A1(new_n1251_), .B0(new_n1253_), .Y(new_n4413_));
  AOI21X1  g4028(.A0(new_n4413_), .A1(new_n1258_), .B0(new_n1261_), .Y(new_n4414_));
  OAI21X1  g4029(.A0(new_n4414_), .A1(new_n1266_), .B0(new_n1268_), .Y(new_n4415_));
  AOI21X1  g4030(.A0(new_n4415_), .A1(new_n1273_), .B0(new_n1276_), .Y(new_n4416_));
  OAI21X1  g4031(.A0(new_n4416_), .A1(new_n1281_), .B0(new_n1283_), .Y(new_n4417_));
  AOI21X1  g4032(.A0(new_n4417_), .A1(new_n1288_), .B0(new_n1291_), .Y(new_n4418_));
  OAI21X1  g4033(.A0(new_n4418_), .A1(new_n1296_), .B0(new_n1298_), .Y(new_n4419_));
  AOI21X1  g4034(.A0(new_n4419_), .A1(new_n1303_), .B0(new_n1306_), .Y(new_n4420_));
  OAI21X1  g4035(.A0(new_n4420_), .A1(new_n1311_), .B0(new_n1313_), .Y(new_n4421_));
  AOI21X1  g4036(.A0(new_n4421_), .A1(new_n1318_), .B0(new_n1321_), .Y(new_n4422_));
  OAI21X1  g4037(.A0(new_n4422_), .A1(new_n1326_), .B0(new_n1328_), .Y(new_n4423_));
  AOI21X1  g4038(.A0(new_n4423_), .A1(new_n1331_), .B0(new_n1758_), .Y(new_n4424_));
  OAI21X1  g4039(.A0(new_n4424_), .A1(new_n394_), .B0(new_n396_), .Y(new_n4425_));
  AOI21X1  g4040(.A0(new_n4425_), .A1(new_n401_), .B0(new_n404_), .Y(new_n4426_));
  OAI21X1  g4041(.A0(new_n4426_), .A1(new_n409_), .B0(new_n411_), .Y(new_n4427_));
  AOI21X1  g4042(.A0(new_n4427_), .A1(new_n416_), .B0(new_n419_), .Y(new_n4428_));
  OAI21X1  g4043(.A0(new_n4428_), .A1(new_n424_), .B0(new_n426_), .Y(new_n4429_));
  AOI21X1  g4044(.A0(new_n4429_), .A1(new_n431_), .B0(new_n434_), .Y(new_n4430_));
  OAI21X1  g4045(.A0(new_n4430_), .A1(new_n439_), .B0(new_n441_), .Y(new_n4431_));
  AOI21X1  g4046(.A0(new_n4431_), .A1(new_n446_), .B0(new_n449_), .Y(new_n4432_));
  OAI21X1  g4047(.A0(new_n4432_), .A1(new_n454_), .B0(new_n456_), .Y(new_n4433_));
  AOI21X1  g4048(.A0(new_n4433_), .A1(new_n461_), .B0(new_n464_), .Y(new_n4434_));
  OAI21X1  g4049(.A0(new_n4434_), .A1(new_n469_), .B0(new_n471_), .Y(new_n4435_));
  AOI21X1  g4050(.A0(new_n4435_), .A1(new_n476_), .B0(new_n479_), .Y(new_n4436_));
  OAI21X1  g4051(.A0(new_n4436_), .A1(new_n484_), .B0(new_n486_), .Y(new_n4437_));
  AOI21X1  g4052(.A0(new_n4437_), .A1(new_n491_), .B0(new_n494_), .Y(new_n4438_));
  OAI21X1  g4053(.A0(new_n4438_), .A1(new_n499_), .B0(new_n501_), .Y(new_n4439_));
  AOI21X1  g4054(.A0(new_n4439_), .A1(new_n506_), .B0(new_n509_), .Y(new_n4440_));
  OAI21X1  g4055(.A0(new_n4440_), .A1(new_n514_), .B0(new_n516_), .Y(new_n4441_));
  AOI21X1  g4056(.A0(new_n4441_), .A1(new_n521_), .B0(new_n524_), .Y(new_n4442_));
  OAI21X1  g4057(.A0(new_n4442_), .A1(new_n529_), .B0(new_n531_), .Y(new_n4443_));
  AOI21X1  g4058(.A0(new_n4443_), .A1(new_n536_), .B0(new_n539_), .Y(new_n4444_));
  OAI21X1  g4059(.A0(new_n4444_), .A1(new_n544_), .B0(new_n546_), .Y(new_n4445_));
  OAI21X1  g4060(.A0(new_n867_), .A1(\priority[68] ), .B0(\req[68] ), .Y(new_n4446_));
  AOI21X1  g4061(.A0(new_n4445_), .A1(new_n551_), .B0(new_n4446_), .Y(\grant[68] ));
  NOR2X1   g4062(.A(new_n876_), .B(new_n560_), .Y(new_n4448_));
  OAI21X1  g4063(.A0(new_n4448_), .A1(new_n1362_), .B0(new_n568_), .Y(new_n4449_));
  AOI21X1  g4064(.A0(new_n4449_), .A1(new_n1360_), .B0(new_n1361_), .Y(new_n4450_));
  OAI21X1  g4065(.A0(new_n4450_), .A1(new_n1359_), .B0(new_n583_), .Y(new_n4451_));
  AOI21X1  g4066(.A0(new_n4451_), .A1(new_n1357_), .B0(new_n1358_), .Y(new_n4452_));
  OAI21X1  g4067(.A0(new_n4452_), .A1(new_n1356_), .B0(new_n598_), .Y(new_n4453_));
  AOI21X1  g4068(.A0(new_n4453_), .A1(new_n1354_), .B0(new_n1355_), .Y(new_n4454_));
  OAI21X1  g4069(.A0(new_n4454_), .A1(new_n1353_), .B0(new_n613_), .Y(new_n4455_));
  AOI21X1  g4070(.A0(new_n4455_), .A1(new_n1351_), .B0(new_n1352_), .Y(new_n4456_));
  OAI21X1  g4071(.A0(new_n4456_), .A1(new_n1350_), .B0(new_n628_), .Y(new_n4457_));
  AOI21X1  g4072(.A0(new_n4457_), .A1(new_n1348_), .B0(new_n1349_), .Y(new_n4458_));
  OAI21X1  g4073(.A0(new_n4458_), .A1(new_n1347_), .B0(new_n643_), .Y(new_n4459_));
  AOI21X1  g4074(.A0(new_n4459_), .A1(new_n1345_), .B0(new_n1346_), .Y(new_n4460_));
  OAI21X1  g4075(.A0(new_n4460_), .A1(new_n1344_), .B0(new_n658_), .Y(new_n4461_));
  AOI21X1  g4076(.A0(new_n4461_), .A1(new_n1342_), .B0(new_n1343_), .Y(new_n4462_));
  OAI21X1  g4077(.A0(new_n4462_), .A1(new_n1341_), .B0(new_n673_), .Y(new_n4463_));
  AOI21X1  g4078(.A0(new_n4463_), .A1(new_n1339_), .B0(new_n1340_), .Y(new_n4464_));
  OAI21X1  g4079(.A0(new_n4464_), .A1(new_n1338_), .B0(new_n688_), .Y(new_n4465_));
  AOI21X1  g4080(.A0(new_n4465_), .A1(new_n1336_), .B0(new_n1337_), .Y(new_n4466_));
  OAI21X1  g4081(.A0(new_n4466_), .A1(new_n1335_), .B0(new_n1438_), .Y(new_n4467_));
  AOI21X1  g4082(.A0(new_n4467_), .A1(new_n1440_), .B0(new_n1803_), .Y(new_n4468_));
  OAI21X1  g4083(.A0(new_n4468_), .A1(new_n712_), .B0(new_n714_), .Y(new_n4469_));
  AOI21X1  g4084(.A0(new_n4469_), .A1(new_n719_), .B0(new_n722_), .Y(new_n4470_));
  OAI21X1  g4085(.A0(new_n4470_), .A1(new_n727_), .B0(new_n729_), .Y(new_n4471_));
  AOI21X1  g4086(.A0(new_n4471_), .A1(new_n734_), .B0(new_n737_), .Y(new_n4472_));
  OAI21X1  g4087(.A0(new_n4472_), .A1(new_n742_), .B0(new_n744_), .Y(new_n4473_));
  AOI21X1  g4088(.A0(new_n4473_), .A1(new_n749_), .B0(new_n752_), .Y(new_n4474_));
  OAI21X1  g4089(.A0(new_n4474_), .A1(new_n757_), .B0(new_n759_), .Y(new_n4475_));
  AOI21X1  g4090(.A0(new_n4475_), .A1(new_n764_), .B0(new_n767_), .Y(new_n4476_));
  OAI21X1  g4091(.A0(new_n4476_), .A1(new_n772_), .B0(new_n774_), .Y(new_n4477_));
  AOI21X1  g4092(.A0(new_n4477_), .A1(new_n779_), .B0(new_n782_), .Y(new_n4478_));
  OAI21X1  g4093(.A0(new_n4478_), .A1(new_n787_), .B0(new_n789_), .Y(new_n4479_));
  AOI21X1  g4094(.A0(new_n4479_), .A1(new_n794_), .B0(new_n797_), .Y(new_n4480_));
  OAI21X1  g4095(.A0(new_n4480_), .A1(new_n802_), .B0(new_n804_), .Y(new_n4481_));
  AOI21X1  g4096(.A0(new_n4481_), .A1(new_n809_), .B0(new_n812_), .Y(new_n4482_));
  OAI21X1  g4097(.A0(new_n4482_), .A1(new_n817_), .B0(new_n819_), .Y(new_n4483_));
  AOI21X1  g4098(.A0(new_n4483_), .A1(new_n824_), .B0(new_n827_), .Y(new_n4484_));
  OAI21X1  g4099(.A0(new_n4484_), .A1(new_n832_), .B0(new_n834_), .Y(new_n4485_));
  AOI21X1  g4100(.A0(new_n4485_), .A1(new_n839_), .B0(new_n842_), .Y(new_n4486_));
  OAI21X1  g4101(.A0(new_n4486_), .A1(new_n847_), .B0(new_n849_), .Y(new_n4487_));
  AOI21X1  g4102(.A0(new_n4487_), .A1(new_n854_), .B0(new_n857_), .Y(new_n4488_));
  OAI21X1  g4103(.A0(new_n4488_), .A1(new_n862_), .B0(new_n864_), .Y(new_n4489_));
  OAI21X1  g4104(.A0(new_n1181_), .A1(\priority[69] ), .B0(\req[69] ), .Y(new_n4490_));
  AOI21X1  g4105(.A0(new_n4489_), .A1(new_n869_), .B0(new_n4490_), .Y(\grant[69] ));
  NOR2X1   g4106(.A(new_n1190_), .B(new_n878_), .Y(new_n4492_));
  OAI21X1  g4107(.A0(new_n4492_), .A1(new_n1471_), .B0(new_n886_), .Y(new_n4493_));
  AOI21X1  g4108(.A0(new_n4493_), .A1(new_n1469_), .B0(new_n1470_), .Y(new_n4494_));
  OAI21X1  g4109(.A0(new_n4494_), .A1(new_n1468_), .B0(new_n901_), .Y(new_n4495_));
  AOI21X1  g4110(.A0(new_n4495_), .A1(new_n1466_), .B0(new_n1467_), .Y(new_n4496_));
  OAI21X1  g4111(.A0(new_n4496_), .A1(new_n1465_), .B0(new_n916_), .Y(new_n4497_));
  AOI21X1  g4112(.A0(new_n4497_), .A1(new_n1463_), .B0(new_n1464_), .Y(new_n4498_));
  OAI21X1  g4113(.A0(new_n4498_), .A1(new_n1462_), .B0(new_n931_), .Y(new_n4499_));
  AOI21X1  g4114(.A0(new_n4499_), .A1(new_n1460_), .B0(new_n1461_), .Y(new_n4500_));
  OAI21X1  g4115(.A0(new_n4500_), .A1(new_n1459_), .B0(new_n946_), .Y(new_n4501_));
  AOI21X1  g4116(.A0(new_n4501_), .A1(new_n1457_), .B0(new_n1458_), .Y(new_n4502_));
  OAI21X1  g4117(.A0(new_n4502_), .A1(new_n1456_), .B0(new_n961_), .Y(new_n4503_));
  AOI21X1  g4118(.A0(new_n4503_), .A1(new_n1454_), .B0(new_n1455_), .Y(new_n4504_));
  OAI21X1  g4119(.A0(new_n4504_), .A1(new_n1453_), .B0(new_n976_), .Y(new_n4505_));
  AOI21X1  g4120(.A0(new_n4505_), .A1(new_n1451_), .B0(new_n1452_), .Y(new_n4506_));
  OAI21X1  g4121(.A0(new_n4506_), .A1(new_n1450_), .B0(new_n991_), .Y(new_n4507_));
  AOI21X1  g4122(.A0(new_n4507_), .A1(new_n1448_), .B0(new_n1449_), .Y(new_n4508_));
  OAI21X1  g4123(.A0(new_n4508_), .A1(new_n1447_), .B0(new_n1006_), .Y(new_n4509_));
  AOI21X1  g4124(.A0(new_n4509_), .A1(new_n1445_), .B0(new_n1446_), .Y(new_n4510_));
  OAI21X1  g4125(.A0(new_n4510_), .A1(new_n1444_), .B0(new_n1547_), .Y(new_n4511_));
  AOI21X1  g4126(.A0(new_n4511_), .A1(new_n1549_), .B0(new_n1848_), .Y(new_n4512_));
  OAI21X1  g4127(.A0(new_n4512_), .A1(new_n1026_), .B0(new_n1028_), .Y(new_n4513_));
  AOI21X1  g4128(.A0(new_n4513_), .A1(new_n1033_), .B0(new_n1036_), .Y(new_n4514_));
  OAI21X1  g4129(.A0(new_n4514_), .A1(new_n1041_), .B0(new_n1043_), .Y(new_n4515_));
  AOI21X1  g4130(.A0(new_n4515_), .A1(new_n1048_), .B0(new_n1051_), .Y(new_n4516_));
  OAI21X1  g4131(.A0(new_n4516_), .A1(new_n1056_), .B0(new_n1058_), .Y(new_n4517_));
  AOI21X1  g4132(.A0(new_n4517_), .A1(new_n1063_), .B0(new_n1066_), .Y(new_n4518_));
  OAI21X1  g4133(.A0(new_n4518_), .A1(new_n1071_), .B0(new_n1073_), .Y(new_n4519_));
  AOI21X1  g4134(.A0(new_n4519_), .A1(new_n1078_), .B0(new_n1081_), .Y(new_n4520_));
  OAI21X1  g4135(.A0(new_n4520_), .A1(new_n1086_), .B0(new_n1088_), .Y(new_n4521_));
  AOI21X1  g4136(.A0(new_n4521_), .A1(new_n1093_), .B0(new_n1096_), .Y(new_n4522_));
  OAI21X1  g4137(.A0(new_n4522_), .A1(new_n1101_), .B0(new_n1103_), .Y(new_n4523_));
  AOI21X1  g4138(.A0(new_n4523_), .A1(new_n1108_), .B0(new_n1111_), .Y(new_n4524_));
  OAI21X1  g4139(.A0(new_n4524_), .A1(new_n1116_), .B0(new_n1118_), .Y(new_n4525_));
  AOI21X1  g4140(.A0(new_n4525_), .A1(new_n1123_), .B0(new_n1126_), .Y(new_n4526_));
  OAI21X1  g4141(.A0(new_n4526_), .A1(new_n1131_), .B0(new_n1133_), .Y(new_n4527_));
  AOI21X1  g4142(.A0(new_n4527_), .A1(new_n1138_), .B0(new_n1141_), .Y(new_n4528_));
  OAI21X1  g4143(.A0(new_n4528_), .A1(new_n1146_), .B0(new_n1148_), .Y(new_n4529_));
  AOI21X1  g4144(.A0(new_n4529_), .A1(new_n1153_), .B0(new_n1156_), .Y(new_n4530_));
  OAI21X1  g4145(.A0(new_n4530_), .A1(new_n1161_), .B0(new_n1163_), .Y(new_n4531_));
  AOI21X1  g4146(.A0(new_n4531_), .A1(new_n1168_), .B0(new_n1171_), .Y(new_n4532_));
  OAI21X1  g4147(.A0(new_n4532_), .A1(new_n1176_), .B0(new_n1178_), .Y(new_n4533_));
  OAI21X1  g4148(.A0(new_n557_), .A1(\priority[70] ), .B0(\req[70] ), .Y(new_n4534_));
  AOI21X1  g4149(.A0(new_n4533_), .A1(new_n1183_), .B0(new_n4534_), .Y(\grant[70] ));
  NOR2X1   g4150(.A(new_n1192_), .B(new_n565_), .Y(new_n4536_));
  OAI21X1  g4151(.A0(new_n4536_), .A1(new_n1580_), .B0(new_n1200_), .Y(new_n4537_));
  AOI21X1  g4152(.A0(new_n4537_), .A1(new_n1578_), .B0(new_n1579_), .Y(new_n4538_));
  OAI21X1  g4153(.A0(new_n4538_), .A1(new_n1577_), .B0(new_n1215_), .Y(new_n4539_));
  AOI21X1  g4154(.A0(new_n4539_), .A1(new_n1575_), .B0(new_n1576_), .Y(new_n4540_));
  OAI21X1  g4155(.A0(new_n4540_), .A1(new_n1574_), .B0(new_n1230_), .Y(new_n4541_));
  AOI21X1  g4156(.A0(new_n4541_), .A1(new_n1572_), .B0(new_n1573_), .Y(new_n4542_));
  OAI21X1  g4157(.A0(new_n4542_), .A1(new_n1571_), .B0(new_n1245_), .Y(new_n4543_));
  AOI21X1  g4158(.A0(new_n4543_), .A1(new_n1569_), .B0(new_n1570_), .Y(new_n4544_));
  OAI21X1  g4159(.A0(new_n4544_), .A1(new_n1568_), .B0(new_n1260_), .Y(new_n4545_));
  AOI21X1  g4160(.A0(new_n4545_), .A1(new_n1566_), .B0(new_n1567_), .Y(new_n4546_));
  OAI21X1  g4161(.A0(new_n4546_), .A1(new_n1565_), .B0(new_n1275_), .Y(new_n4547_));
  AOI21X1  g4162(.A0(new_n4547_), .A1(new_n1563_), .B0(new_n1564_), .Y(new_n4548_));
  OAI21X1  g4163(.A0(new_n4548_), .A1(new_n1562_), .B0(new_n1290_), .Y(new_n4549_));
  AOI21X1  g4164(.A0(new_n4549_), .A1(new_n1560_), .B0(new_n1561_), .Y(new_n4550_));
  OAI21X1  g4165(.A0(new_n4550_), .A1(new_n1559_), .B0(new_n1305_), .Y(new_n4551_));
  AOI21X1  g4166(.A0(new_n4551_), .A1(new_n1557_), .B0(new_n1558_), .Y(new_n4552_));
  OAI21X1  g4167(.A0(new_n4552_), .A1(new_n1556_), .B0(new_n1320_), .Y(new_n4553_));
  AOI21X1  g4168(.A0(new_n4553_), .A1(new_n1554_), .B0(new_n1555_), .Y(new_n4554_));
  OAI21X1  g4169(.A0(new_n4554_), .A1(new_n1553_), .B0(new_n1656_), .Y(new_n4555_));
  AOI21X1  g4170(.A0(new_n4555_), .A1(new_n1552_), .B0(new_n1893_), .Y(new_n4556_));
  OAI21X1  g4171(.A0(new_n4556_), .A1(new_n1395_), .B0(new_n403_), .Y(new_n4557_));
  AOI21X1  g4172(.A0(new_n4557_), .A1(new_n1393_), .B0(new_n1394_), .Y(new_n4558_));
  OAI21X1  g4173(.A0(new_n4558_), .A1(new_n1392_), .B0(new_n418_), .Y(new_n4559_));
  AOI21X1  g4174(.A0(new_n4559_), .A1(new_n1390_), .B0(new_n1391_), .Y(new_n4560_));
  OAI21X1  g4175(.A0(new_n4560_), .A1(new_n1389_), .B0(new_n433_), .Y(new_n4561_));
  AOI21X1  g4176(.A0(new_n4561_), .A1(new_n1387_), .B0(new_n1388_), .Y(new_n4562_));
  OAI21X1  g4177(.A0(new_n4562_), .A1(new_n1386_), .B0(new_n448_), .Y(new_n4563_));
  AOI21X1  g4178(.A0(new_n4563_), .A1(new_n1384_), .B0(new_n1385_), .Y(new_n4564_));
  OAI21X1  g4179(.A0(new_n4564_), .A1(new_n1383_), .B0(new_n463_), .Y(new_n4565_));
  AOI21X1  g4180(.A0(new_n4565_), .A1(new_n1381_), .B0(new_n1382_), .Y(new_n4566_));
  OAI21X1  g4181(.A0(new_n4566_), .A1(new_n1380_), .B0(new_n478_), .Y(new_n4567_));
  AOI21X1  g4182(.A0(new_n4567_), .A1(new_n1378_), .B0(new_n1379_), .Y(new_n4568_));
  OAI21X1  g4183(.A0(new_n4568_), .A1(new_n1377_), .B0(new_n493_), .Y(new_n4569_));
  AOI21X1  g4184(.A0(new_n4569_), .A1(new_n1375_), .B0(new_n1376_), .Y(new_n4570_));
  OAI21X1  g4185(.A0(new_n4570_), .A1(new_n1374_), .B0(new_n508_), .Y(new_n4571_));
  AOI21X1  g4186(.A0(new_n4571_), .A1(new_n1372_), .B0(new_n1373_), .Y(new_n4572_));
  OAI21X1  g4187(.A0(new_n4572_), .A1(new_n1371_), .B0(new_n523_), .Y(new_n4573_));
  AOI21X1  g4188(.A0(new_n4573_), .A1(new_n1369_), .B0(new_n1370_), .Y(new_n4574_));
  OAI21X1  g4189(.A0(new_n4574_), .A1(new_n1368_), .B0(new_n538_), .Y(new_n4575_));
  AOI21X1  g4190(.A0(new_n4575_), .A1(new_n1366_), .B0(new_n1367_), .Y(new_n4576_));
  OAI21X1  g4191(.A0(new_n4576_), .A1(new_n1365_), .B0(new_n553_), .Y(new_n4577_));
  OAI21X1  g4192(.A0(new_n875_), .A1(\priority[71] ), .B0(\req[71] ), .Y(new_n4578_));
  AOI21X1  g4193(.A0(new_n4577_), .A1(new_n1363_), .B0(new_n4578_), .Y(\grant[71] ));
  NOR2X1   g4194(.A(new_n883_), .B(new_n567_), .Y(new_n4580_));
  OAI21X1  g4195(.A0(new_n4580_), .A1(new_n574_), .B0(new_n576_), .Y(new_n4581_));
  AOI21X1  g4196(.A0(new_n4581_), .A1(new_n581_), .B0(new_n584_), .Y(new_n4582_));
  OAI21X1  g4197(.A0(new_n4582_), .A1(new_n589_), .B0(new_n591_), .Y(new_n4583_));
  AOI21X1  g4198(.A0(new_n4583_), .A1(new_n596_), .B0(new_n599_), .Y(new_n4584_));
  OAI21X1  g4199(.A0(new_n4584_), .A1(new_n604_), .B0(new_n606_), .Y(new_n4585_));
  AOI21X1  g4200(.A0(new_n4585_), .A1(new_n611_), .B0(new_n614_), .Y(new_n4586_));
  OAI21X1  g4201(.A0(new_n4586_), .A1(new_n619_), .B0(new_n621_), .Y(new_n4587_));
  AOI21X1  g4202(.A0(new_n4587_), .A1(new_n626_), .B0(new_n629_), .Y(new_n4588_));
  OAI21X1  g4203(.A0(new_n4588_), .A1(new_n634_), .B0(new_n636_), .Y(new_n4589_));
  AOI21X1  g4204(.A0(new_n4589_), .A1(new_n641_), .B0(new_n644_), .Y(new_n4590_));
  OAI21X1  g4205(.A0(new_n4590_), .A1(new_n649_), .B0(new_n651_), .Y(new_n4591_));
  AOI21X1  g4206(.A0(new_n4591_), .A1(new_n656_), .B0(new_n659_), .Y(new_n4592_));
  OAI21X1  g4207(.A0(new_n4592_), .A1(new_n664_), .B0(new_n666_), .Y(new_n4593_));
  AOI21X1  g4208(.A0(new_n4593_), .A1(new_n671_), .B0(new_n674_), .Y(new_n4594_));
  OAI21X1  g4209(.A0(new_n4594_), .A1(new_n679_), .B0(new_n681_), .Y(new_n4595_));
  AOI21X1  g4210(.A0(new_n4595_), .A1(new_n686_), .B0(new_n689_), .Y(new_n4596_));
  OAI21X1  g4211(.A0(new_n4596_), .A1(new_n694_), .B0(new_n696_), .Y(new_n4597_));
  AOI21X1  g4212(.A0(new_n4597_), .A1(new_n701_), .B0(new_n1662_), .Y(new_n4598_));
  OAI21X1  g4213(.A0(new_n4598_), .A1(new_n1661_), .B0(new_n1705_), .Y(new_n4599_));
  AOI21X1  g4214(.A0(new_n4599_), .A1(new_n1660_), .B0(new_n1938_), .Y(new_n4600_));
  OAI21X1  g4215(.A0(new_n4600_), .A1(new_n1504_), .B0(new_n721_), .Y(new_n4601_));
  AOI21X1  g4216(.A0(new_n4601_), .A1(new_n1502_), .B0(new_n1503_), .Y(new_n4602_));
  OAI21X1  g4217(.A0(new_n4602_), .A1(new_n1501_), .B0(new_n736_), .Y(new_n4603_));
  AOI21X1  g4218(.A0(new_n4603_), .A1(new_n1499_), .B0(new_n1500_), .Y(new_n4604_));
  OAI21X1  g4219(.A0(new_n4604_), .A1(new_n1498_), .B0(new_n751_), .Y(new_n4605_));
  AOI21X1  g4220(.A0(new_n4605_), .A1(new_n1496_), .B0(new_n1497_), .Y(new_n4606_));
  OAI21X1  g4221(.A0(new_n4606_), .A1(new_n1495_), .B0(new_n766_), .Y(new_n4607_));
  AOI21X1  g4222(.A0(new_n4607_), .A1(new_n1493_), .B0(new_n1494_), .Y(new_n4608_));
  OAI21X1  g4223(.A0(new_n4608_), .A1(new_n1492_), .B0(new_n781_), .Y(new_n4609_));
  AOI21X1  g4224(.A0(new_n4609_), .A1(new_n1490_), .B0(new_n1491_), .Y(new_n4610_));
  OAI21X1  g4225(.A0(new_n4610_), .A1(new_n1489_), .B0(new_n796_), .Y(new_n4611_));
  AOI21X1  g4226(.A0(new_n4611_), .A1(new_n1487_), .B0(new_n1488_), .Y(new_n4612_));
  OAI21X1  g4227(.A0(new_n4612_), .A1(new_n1486_), .B0(new_n811_), .Y(new_n4613_));
  AOI21X1  g4228(.A0(new_n4613_), .A1(new_n1484_), .B0(new_n1485_), .Y(new_n4614_));
  OAI21X1  g4229(.A0(new_n4614_), .A1(new_n1483_), .B0(new_n826_), .Y(new_n4615_));
  AOI21X1  g4230(.A0(new_n4615_), .A1(new_n1481_), .B0(new_n1482_), .Y(new_n4616_));
  OAI21X1  g4231(.A0(new_n4616_), .A1(new_n1480_), .B0(new_n841_), .Y(new_n4617_));
  AOI21X1  g4232(.A0(new_n4617_), .A1(new_n1478_), .B0(new_n1479_), .Y(new_n4618_));
  OAI21X1  g4233(.A0(new_n4618_), .A1(new_n1477_), .B0(new_n856_), .Y(new_n4619_));
  AOI21X1  g4234(.A0(new_n4619_), .A1(new_n1475_), .B0(new_n1476_), .Y(new_n4620_));
  OAI21X1  g4235(.A0(new_n4620_), .A1(new_n1474_), .B0(new_n871_), .Y(new_n4621_));
  OAI21X1  g4236(.A0(new_n1189_), .A1(\priority[72] ), .B0(\req[72] ), .Y(new_n4622_));
  AOI21X1  g4237(.A0(new_n4621_), .A1(new_n1472_), .B0(new_n4622_), .Y(\grant[72] ));
  NOR2X1   g4238(.A(new_n1197_), .B(new_n885_), .Y(new_n4624_));
  OAI21X1  g4239(.A0(new_n4624_), .A1(new_n892_), .B0(new_n894_), .Y(new_n4625_));
  AOI21X1  g4240(.A0(new_n4625_), .A1(new_n899_), .B0(new_n902_), .Y(new_n4626_));
  OAI21X1  g4241(.A0(new_n4626_), .A1(new_n907_), .B0(new_n909_), .Y(new_n4627_));
  AOI21X1  g4242(.A0(new_n4627_), .A1(new_n914_), .B0(new_n917_), .Y(new_n4628_));
  OAI21X1  g4243(.A0(new_n4628_), .A1(new_n922_), .B0(new_n924_), .Y(new_n4629_));
  AOI21X1  g4244(.A0(new_n4629_), .A1(new_n929_), .B0(new_n932_), .Y(new_n4630_));
  OAI21X1  g4245(.A0(new_n4630_), .A1(new_n937_), .B0(new_n939_), .Y(new_n4631_));
  AOI21X1  g4246(.A0(new_n4631_), .A1(new_n944_), .B0(new_n947_), .Y(new_n4632_));
  OAI21X1  g4247(.A0(new_n4632_), .A1(new_n952_), .B0(new_n954_), .Y(new_n4633_));
  AOI21X1  g4248(.A0(new_n4633_), .A1(new_n959_), .B0(new_n962_), .Y(new_n4634_));
  OAI21X1  g4249(.A0(new_n4634_), .A1(new_n967_), .B0(new_n969_), .Y(new_n4635_));
  AOI21X1  g4250(.A0(new_n4635_), .A1(new_n974_), .B0(new_n977_), .Y(new_n4636_));
  OAI21X1  g4251(.A0(new_n4636_), .A1(new_n982_), .B0(new_n984_), .Y(new_n4637_));
  AOI21X1  g4252(.A0(new_n4637_), .A1(new_n989_), .B0(new_n992_), .Y(new_n4638_));
  OAI21X1  g4253(.A0(new_n4638_), .A1(new_n997_), .B0(new_n999_), .Y(new_n4639_));
  AOI21X1  g4254(.A0(new_n4639_), .A1(new_n1004_), .B0(new_n1007_), .Y(new_n4640_));
  OAI21X1  g4255(.A0(new_n4640_), .A1(new_n1012_), .B0(new_n1014_), .Y(new_n4641_));
  AOI21X1  g4256(.A0(new_n4641_), .A1(new_n1017_), .B0(new_n1711_), .Y(new_n4642_));
  OAI21X1  g4257(.A0(new_n4642_), .A1(new_n1710_), .B0(new_n1754_), .Y(new_n4643_));
  AOI21X1  g4258(.A0(new_n4643_), .A1(new_n1709_), .B0(new_n1983_), .Y(new_n4644_));
  OAI21X1  g4259(.A0(new_n4644_), .A1(new_n1613_), .B0(new_n1035_), .Y(new_n4645_));
  AOI21X1  g4260(.A0(new_n4645_), .A1(new_n1611_), .B0(new_n1612_), .Y(new_n4646_));
  OAI21X1  g4261(.A0(new_n4646_), .A1(new_n1610_), .B0(new_n1050_), .Y(new_n4647_));
  AOI21X1  g4262(.A0(new_n4647_), .A1(new_n1608_), .B0(new_n1609_), .Y(new_n4648_));
  OAI21X1  g4263(.A0(new_n4648_), .A1(new_n1607_), .B0(new_n1065_), .Y(new_n4649_));
  AOI21X1  g4264(.A0(new_n4649_), .A1(new_n1605_), .B0(new_n1606_), .Y(new_n4650_));
  OAI21X1  g4265(.A0(new_n4650_), .A1(new_n1604_), .B0(new_n1080_), .Y(new_n4651_));
  AOI21X1  g4266(.A0(new_n4651_), .A1(new_n1602_), .B0(new_n1603_), .Y(new_n4652_));
  OAI21X1  g4267(.A0(new_n4652_), .A1(new_n1601_), .B0(new_n1095_), .Y(new_n4653_));
  AOI21X1  g4268(.A0(new_n4653_), .A1(new_n1599_), .B0(new_n1600_), .Y(new_n4654_));
  OAI21X1  g4269(.A0(new_n4654_), .A1(new_n1598_), .B0(new_n1110_), .Y(new_n4655_));
  AOI21X1  g4270(.A0(new_n4655_), .A1(new_n1596_), .B0(new_n1597_), .Y(new_n4656_));
  OAI21X1  g4271(.A0(new_n4656_), .A1(new_n1595_), .B0(new_n1125_), .Y(new_n4657_));
  AOI21X1  g4272(.A0(new_n4657_), .A1(new_n1593_), .B0(new_n1594_), .Y(new_n4658_));
  OAI21X1  g4273(.A0(new_n4658_), .A1(new_n1592_), .B0(new_n1140_), .Y(new_n4659_));
  AOI21X1  g4274(.A0(new_n4659_), .A1(new_n1590_), .B0(new_n1591_), .Y(new_n4660_));
  OAI21X1  g4275(.A0(new_n4660_), .A1(new_n1589_), .B0(new_n1155_), .Y(new_n4661_));
  AOI21X1  g4276(.A0(new_n4661_), .A1(new_n1587_), .B0(new_n1588_), .Y(new_n4662_));
  OAI21X1  g4277(.A0(new_n4662_), .A1(new_n1586_), .B0(new_n1170_), .Y(new_n4663_));
  AOI21X1  g4278(.A0(new_n4663_), .A1(new_n1584_), .B0(new_n1585_), .Y(new_n4664_));
  OAI21X1  g4279(.A0(new_n4664_), .A1(new_n1583_), .B0(new_n1185_), .Y(new_n4665_));
  OAI21X1  g4280(.A0(new_n564_), .A1(\priority[73] ), .B0(\req[73] ), .Y(new_n4666_));
  AOI21X1  g4281(.A0(new_n4665_), .A1(new_n1581_), .B0(new_n4666_), .Y(\grant[73] ));
  NOR2X1   g4282(.A(new_n1199_), .B(new_n573_), .Y(new_n4668_));
  OAI21X1  g4283(.A0(new_n4668_), .A1(new_n1206_), .B0(new_n1208_), .Y(new_n4669_));
  AOI21X1  g4284(.A0(new_n4669_), .A1(new_n1213_), .B0(new_n1216_), .Y(new_n4670_));
  OAI21X1  g4285(.A0(new_n4670_), .A1(new_n1221_), .B0(new_n1223_), .Y(new_n4671_));
  AOI21X1  g4286(.A0(new_n4671_), .A1(new_n1228_), .B0(new_n1231_), .Y(new_n4672_));
  OAI21X1  g4287(.A0(new_n4672_), .A1(new_n1236_), .B0(new_n1238_), .Y(new_n4673_));
  AOI21X1  g4288(.A0(new_n4673_), .A1(new_n1243_), .B0(new_n1246_), .Y(new_n4674_));
  OAI21X1  g4289(.A0(new_n4674_), .A1(new_n1251_), .B0(new_n1253_), .Y(new_n4675_));
  AOI21X1  g4290(.A0(new_n4675_), .A1(new_n1258_), .B0(new_n1261_), .Y(new_n4676_));
  OAI21X1  g4291(.A0(new_n4676_), .A1(new_n1266_), .B0(new_n1268_), .Y(new_n4677_));
  AOI21X1  g4292(.A0(new_n4677_), .A1(new_n1273_), .B0(new_n1276_), .Y(new_n4678_));
  OAI21X1  g4293(.A0(new_n4678_), .A1(new_n1281_), .B0(new_n1283_), .Y(new_n4679_));
  AOI21X1  g4294(.A0(new_n4679_), .A1(new_n1288_), .B0(new_n1291_), .Y(new_n4680_));
  OAI21X1  g4295(.A0(new_n4680_), .A1(new_n1296_), .B0(new_n1298_), .Y(new_n4681_));
  AOI21X1  g4296(.A0(new_n4681_), .A1(new_n1303_), .B0(new_n1306_), .Y(new_n4682_));
  OAI21X1  g4297(.A0(new_n4682_), .A1(new_n1311_), .B0(new_n1313_), .Y(new_n4683_));
  AOI21X1  g4298(.A0(new_n4683_), .A1(new_n1318_), .B0(new_n1321_), .Y(new_n4684_));
  OAI21X1  g4299(.A0(new_n4684_), .A1(new_n1326_), .B0(new_n1328_), .Y(new_n4685_));
  AOI21X1  g4300(.A0(new_n4685_), .A1(new_n1331_), .B0(new_n1758_), .Y(new_n4686_));
  OAI21X1  g4301(.A0(new_n4686_), .A1(new_n394_), .B0(new_n396_), .Y(new_n4687_));
  AOI21X1  g4302(.A0(new_n4687_), .A1(new_n401_), .B0(new_n404_), .Y(new_n4688_));
  OAI21X1  g4303(.A0(new_n4688_), .A1(new_n409_), .B0(new_n411_), .Y(new_n4689_));
  AOI21X1  g4304(.A0(new_n4689_), .A1(new_n416_), .B0(new_n419_), .Y(new_n4690_));
  OAI21X1  g4305(.A0(new_n4690_), .A1(new_n424_), .B0(new_n426_), .Y(new_n4691_));
  AOI21X1  g4306(.A0(new_n4691_), .A1(new_n431_), .B0(new_n434_), .Y(new_n4692_));
  OAI21X1  g4307(.A0(new_n4692_), .A1(new_n439_), .B0(new_n441_), .Y(new_n4693_));
  AOI21X1  g4308(.A0(new_n4693_), .A1(new_n446_), .B0(new_n449_), .Y(new_n4694_));
  OAI21X1  g4309(.A0(new_n4694_), .A1(new_n454_), .B0(new_n456_), .Y(new_n4695_));
  AOI21X1  g4310(.A0(new_n4695_), .A1(new_n461_), .B0(new_n464_), .Y(new_n4696_));
  OAI21X1  g4311(.A0(new_n4696_), .A1(new_n469_), .B0(new_n471_), .Y(new_n4697_));
  AOI21X1  g4312(.A0(new_n4697_), .A1(new_n476_), .B0(new_n479_), .Y(new_n4698_));
  OAI21X1  g4313(.A0(new_n4698_), .A1(new_n484_), .B0(new_n486_), .Y(new_n4699_));
  AOI21X1  g4314(.A0(new_n4699_), .A1(new_n491_), .B0(new_n494_), .Y(new_n4700_));
  OAI21X1  g4315(.A0(new_n4700_), .A1(new_n499_), .B0(new_n501_), .Y(new_n4701_));
  AOI21X1  g4316(.A0(new_n4701_), .A1(new_n506_), .B0(new_n509_), .Y(new_n4702_));
  OAI21X1  g4317(.A0(new_n4702_), .A1(new_n514_), .B0(new_n516_), .Y(new_n4703_));
  AOI21X1  g4318(.A0(new_n4703_), .A1(new_n521_), .B0(new_n524_), .Y(new_n4704_));
  OAI21X1  g4319(.A0(new_n4704_), .A1(new_n529_), .B0(new_n531_), .Y(new_n4705_));
  AOI21X1  g4320(.A0(new_n4705_), .A1(new_n536_), .B0(new_n539_), .Y(new_n4706_));
  OAI21X1  g4321(.A0(new_n4706_), .A1(new_n544_), .B0(new_n546_), .Y(new_n4707_));
  AOI21X1  g4322(.A0(new_n4707_), .A1(new_n551_), .B0(new_n554_), .Y(new_n4708_));
  OAI21X1  g4323(.A0(new_n4708_), .A1(new_n559_), .B0(new_n561_), .Y(new_n4709_));
  OAI21X1  g4324(.A0(new_n882_), .A1(\priority[74] ), .B0(\req[74] ), .Y(new_n4710_));
  AOI21X1  g4325(.A0(new_n4709_), .A1(new_n566_), .B0(new_n4710_), .Y(\grant[74] ));
  NOR2X1   g4326(.A(new_n891_), .B(new_n575_), .Y(new_n4712_));
  OAI21X1  g4327(.A0(new_n4712_), .A1(new_n1359_), .B0(new_n583_), .Y(new_n4713_));
  AOI21X1  g4328(.A0(new_n4713_), .A1(new_n1357_), .B0(new_n1358_), .Y(new_n4714_));
  OAI21X1  g4329(.A0(new_n4714_), .A1(new_n1356_), .B0(new_n598_), .Y(new_n4715_));
  AOI21X1  g4330(.A0(new_n4715_), .A1(new_n1354_), .B0(new_n1355_), .Y(new_n4716_));
  OAI21X1  g4331(.A0(new_n4716_), .A1(new_n1353_), .B0(new_n613_), .Y(new_n4717_));
  AOI21X1  g4332(.A0(new_n4717_), .A1(new_n1351_), .B0(new_n1352_), .Y(new_n4718_));
  OAI21X1  g4333(.A0(new_n4718_), .A1(new_n1350_), .B0(new_n628_), .Y(new_n4719_));
  AOI21X1  g4334(.A0(new_n4719_), .A1(new_n1348_), .B0(new_n1349_), .Y(new_n4720_));
  OAI21X1  g4335(.A0(new_n4720_), .A1(new_n1347_), .B0(new_n643_), .Y(new_n4721_));
  AOI21X1  g4336(.A0(new_n4721_), .A1(new_n1345_), .B0(new_n1346_), .Y(new_n4722_));
  OAI21X1  g4337(.A0(new_n4722_), .A1(new_n1344_), .B0(new_n658_), .Y(new_n4723_));
  AOI21X1  g4338(.A0(new_n4723_), .A1(new_n1342_), .B0(new_n1343_), .Y(new_n4724_));
  OAI21X1  g4339(.A0(new_n4724_), .A1(new_n1341_), .B0(new_n673_), .Y(new_n4725_));
  AOI21X1  g4340(.A0(new_n4725_), .A1(new_n1339_), .B0(new_n1340_), .Y(new_n4726_));
  OAI21X1  g4341(.A0(new_n4726_), .A1(new_n1338_), .B0(new_n688_), .Y(new_n4727_));
  AOI21X1  g4342(.A0(new_n4727_), .A1(new_n1336_), .B0(new_n1337_), .Y(new_n4728_));
  OAI21X1  g4343(.A0(new_n4728_), .A1(new_n1335_), .B0(new_n1438_), .Y(new_n4729_));
  AOI21X1  g4344(.A0(new_n4729_), .A1(new_n1440_), .B0(new_n1803_), .Y(new_n4730_));
  OAI21X1  g4345(.A0(new_n4730_), .A1(new_n712_), .B0(new_n714_), .Y(new_n4731_));
  AOI21X1  g4346(.A0(new_n4731_), .A1(new_n719_), .B0(new_n722_), .Y(new_n4732_));
  OAI21X1  g4347(.A0(new_n4732_), .A1(new_n727_), .B0(new_n729_), .Y(new_n4733_));
  AOI21X1  g4348(.A0(new_n4733_), .A1(new_n734_), .B0(new_n737_), .Y(new_n4734_));
  OAI21X1  g4349(.A0(new_n4734_), .A1(new_n742_), .B0(new_n744_), .Y(new_n4735_));
  AOI21X1  g4350(.A0(new_n4735_), .A1(new_n749_), .B0(new_n752_), .Y(new_n4736_));
  OAI21X1  g4351(.A0(new_n4736_), .A1(new_n757_), .B0(new_n759_), .Y(new_n4737_));
  AOI21X1  g4352(.A0(new_n4737_), .A1(new_n764_), .B0(new_n767_), .Y(new_n4738_));
  OAI21X1  g4353(.A0(new_n4738_), .A1(new_n772_), .B0(new_n774_), .Y(new_n4739_));
  AOI21X1  g4354(.A0(new_n4739_), .A1(new_n779_), .B0(new_n782_), .Y(new_n4740_));
  OAI21X1  g4355(.A0(new_n4740_), .A1(new_n787_), .B0(new_n789_), .Y(new_n4741_));
  AOI21X1  g4356(.A0(new_n4741_), .A1(new_n794_), .B0(new_n797_), .Y(new_n4742_));
  OAI21X1  g4357(.A0(new_n4742_), .A1(new_n802_), .B0(new_n804_), .Y(new_n4743_));
  AOI21X1  g4358(.A0(new_n4743_), .A1(new_n809_), .B0(new_n812_), .Y(new_n4744_));
  OAI21X1  g4359(.A0(new_n4744_), .A1(new_n817_), .B0(new_n819_), .Y(new_n4745_));
  AOI21X1  g4360(.A0(new_n4745_), .A1(new_n824_), .B0(new_n827_), .Y(new_n4746_));
  OAI21X1  g4361(.A0(new_n4746_), .A1(new_n832_), .B0(new_n834_), .Y(new_n4747_));
  AOI21X1  g4362(.A0(new_n4747_), .A1(new_n839_), .B0(new_n842_), .Y(new_n4748_));
  OAI21X1  g4363(.A0(new_n4748_), .A1(new_n847_), .B0(new_n849_), .Y(new_n4749_));
  AOI21X1  g4364(.A0(new_n4749_), .A1(new_n854_), .B0(new_n857_), .Y(new_n4750_));
  OAI21X1  g4365(.A0(new_n4750_), .A1(new_n862_), .B0(new_n864_), .Y(new_n4751_));
  AOI21X1  g4366(.A0(new_n4751_), .A1(new_n869_), .B0(new_n872_), .Y(new_n4752_));
  OAI21X1  g4367(.A0(new_n4752_), .A1(new_n877_), .B0(new_n879_), .Y(new_n4753_));
  OAI21X1  g4368(.A0(new_n1196_), .A1(\priority[75] ), .B0(\req[75] ), .Y(new_n4754_));
  AOI21X1  g4369(.A0(new_n4753_), .A1(new_n884_), .B0(new_n4754_), .Y(\grant[75] ));
  NOR2X1   g4370(.A(new_n1205_), .B(new_n893_), .Y(new_n4756_));
  OAI21X1  g4371(.A0(new_n4756_), .A1(new_n1468_), .B0(new_n901_), .Y(new_n4757_));
  AOI21X1  g4372(.A0(new_n4757_), .A1(new_n1466_), .B0(new_n1467_), .Y(new_n4758_));
  OAI21X1  g4373(.A0(new_n4758_), .A1(new_n1465_), .B0(new_n916_), .Y(new_n4759_));
  AOI21X1  g4374(.A0(new_n4759_), .A1(new_n1463_), .B0(new_n1464_), .Y(new_n4760_));
  OAI21X1  g4375(.A0(new_n4760_), .A1(new_n1462_), .B0(new_n931_), .Y(new_n4761_));
  AOI21X1  g4376(.A0(new_n4761_), .A1(new_n1460_), .B0(new_n1461_), .Y(new_n4762_));
  OAI21X1  g4377(.A0(new_n4762_), .A1(new_n1459_), .B0(new_n946_), .Y(new_n4763_));
  AOI21X1  g4378(.A0(new_n4763_), .A1(new_n1457_), .B0(new_n1458_), .Y(new_n4764_));
  OAI21X1  g4379(.A0(new_n4764_), .A1(new_n1456_), .B0(new_n961_), .Y(new_n4765_));
  AOI21X1  g4380(.A0(new_n4765_), .A1(new_n1454_), .B0(new_n1455_), .Y(new_n4766_));
  OAI21X1  g4381(.A0(new_n4766_), .A1(new_n1453_), .B0(new_n976_), .Y(new_n4767_));
  AOI21X1  g4382(.A0(new_n4767_), .A1(new_n1451_), .B0(new_n1452_), .Y(new_n4768_));
  OAI21X1  g4383(.A0(new_n4768_), .A1(new_n1450_), .B0(new_n991_), .Y(new_n4769_));
  AOI21X1  g4384(.A0(new_n4769_), .A1(new_n1448_), .B0(new_n1449_), .Y(new_n4770_));
  OAI21X1  g4385(.A0(new_n4770_), .A1(new_n1447_), .B0(new_n1006_), .Y(new_n4771_));
  AOI21X1  g4386(.A0(new_n4771_), .A1(new_n1445_), .B0(new_n1446_), .Y(new_n4772_));
  OAI21X1  g4387(.A0(new_n4772_), .A1(new_n1444_), .B0(new_n1547_), .Y(new_n4773_));
  AOI21X1  g4388(.A0(new_n4773_), .A1(new_n1549_), .B0(new_n1848_), .Y(new_n4774_));
  OAI21X1  g4389(.A0(new_n4774_), .A1(new_n1026_), .B0(new_n1028_), .Y(new_n4775_));
  AOI21X1  g4390(.A0(new_n4775_), .A1(new_n1033_), .B0(new_n1036_), .Y(new_n4776_));
  OAI21X1  g4391(.A0(new_n4776_), .A1(new_n1041_), .B0(new_n1043_), .Y(new_n4777_));
  AOI21X1  g4392(.A0(new_n4777_), .A1(new_n1048_), .B0(new_n1051_), .Y(new_n4778_));
  OAI21X1  g4393(.A0(new_n4778_), .A1(new_n1056_), .B0(new_n1058_), .Y(new_n4779_));
  AOI21X1  g4394(.A0(new_n4779_), .A1(new_n1063_), .B0(new_n1066_), .Y(new_n4780_));
  OAI21X1  g4395(.A0(new_n4780_), .A1(new_n1071_), .B0(new_n1073_), .Y(new_n4781_));
  AOI21X1  g4396(.A0(new_n4781_), .A1(new_n1078_), .B0(new_n1081_), .Y(new_n4782_));
  OAI21X1  g4397(.A0(new_n4782_), .A1(new_n1086_), .B0(new_n1088_), .Y(new_n4783_));
  AOI21X1  g4398(.A0(new_n4783_), .A1(new_n1093_), .B0(new_n1096_), .Y(new_n4784_));
  OAI21X1  g4399(.A0(new_n4784_), .A1(new_n1101_), .B0(new_n1103_), .Y(new_n4785_));
  AOI21X1  g4400(.A0(new_n4785_), .A1(new_n1108_), .B0(new_n1111_), .Y(new_n4786_));
  OAI21X1  g4401(.A0(new_n4786_), .A1(new_n1116_), .B0(new_n1118_), .Y(new_n4787_));
  AOI21X1  g4402(.A0(new_n4787_), .A1(new_n1123_), .B0(new_n1126_), .Y(new_n4788_));
  OAI21X1  g4403(.A0(new_n4788_), .A1(new_n1131_), .B0(new_n1133_), .Y(new_n4789_));
  AOI21X1  g4404(.A0(new_n4789_), .A1(new_n1138_), .B0(new_n1141_), .Y(new_n4790_));
  OAI21X1  g4405(.A0(new_n4790_), .A1(new_n1146_), .B0(new_n1148_), .Y(new_n4791_));
  AOI21X1  g4406(.A0(new_n4791_), .A1(new_n1153_), .B0(new_n1156_), .Y(new_n4792_));
  OAI21X1  g4407(.A0(new_n4792_), .A1(new_n1161_), .B0(new_n1163_), .Y(new_n4793_));
  AOI21X1  g4408(.A0(new_n4793_), .A1(new_n1168_), .B0(new_n1171_), .Y(new_n4794_));
  OAI21X1  g4409(.A0(new_n4794_), .A1(new_n1176_), .B0(new_n1178_), .Y(new_n4795_));
  AOI21X1  g4410(.A0(new_n4795_), .A1(new_n1183_), .B0(new_n1186_), .Y(new_n4796_));
  OAI21X1  g4411(.A0(new_n4796_), .A1(new_n1191_), .B0(new_n1193_), .Y(new_n4797_));
  OAI21X1  g4412(.A0(new_n572_), .A1(\priority[76] ), .B0(\req[76] ), .Y(new_n4798_));
  AOI21X1  g4413(.A0(new_n4797_), .A1(new_n1198_), .B0(new_n4798_), .Y(\grant[76] ));
  NOR2X1   g4414(.A(new_n1207_), .B(new_n580_), .Y(new_n4800_));
  OAI21X1  g4415(.A0(new_n4800_), .A1(new_n1577_), .B0(new_n1215_), .Y(new_n4801_));
  AOI21X1  g4416(.A0(new_n4801_), .A1(new_n1575_), .B0(new_n1576_), .Y(new_n4802_));
  OAI21X1  g4417(.A0(new_n4802_), .A1(new_n1574_), .B0(new_n1230_), .Y(new_n4803_));
  AOI21X1  g4418(.A0(new_n4803_), .A1(new_n1572_), .B0(new_n1573_), .Y(new_n4804_));
  OAI21X1  g4419(.A0(new_n4804_), .A1(new_n1571_), .B0(new_n1245_), .Y(new_n4805_));
  AOI21X1  g4420(.A0(new_n4805_), .A1(new_n1569_), .B0(new_n1570_), .Y(new_n4806_));
  OAI21X1  g4421(.A0(new_n4806_), .A1(new_n1568_), .B0(new_n1260_), .Y(new_n4807_));
  AOI21X1  g4422(.A0(new_n4807_), .A1(new_n1566_), .B0(new_n1567_), .Y(new_n4808_));
  OAI21X1  g4423(.A0(new_n4808_), .A1(new_n1565_), .B0(new_n1275_), .Y(new_n4809_));
  AOI21X1  g4424(.A0(new_n4809_), .A1(new_n1563_), .B0(new_n1564_), .Y(new_n4810_));
  OAI21X1  g4425(.A0(new_n4810_), .A1(new_n1562_), .B0(new_n1290_), .Y(new_n4811_));
  AOI21X1  g4426(.A0(new_n4811_), .A1(new_n1560_), .B0(new_n1561_), .Y(new_n4812_));
  OAI21X1  g4427(.A0(new_n4812_), .A1(new_n1559_), .B0(new_n1305_), .Y(new_n4813_));
  AOI21X1  g4428(.A0(new_n4813_), .A1(new_n1557_), .B0(new_n1558_), .Y(new_n4814_));
  OAI21X1  g4429(.A0(new_n4814_), .A1(new_n1556_), .B0(new_n1320_), .Y(new_n4815_));
  AOI21X1  g4430(.A0(new_n4815_), .A1(new_n1554_), .B0(new_n1555_), .Y(new_n4816_));
  OAI21X1  g4431(.A0(new_n4816_), .A1(new_n1553_), .B0(new_n1656_), .Y(new_n4817_));
  AOI21X1  g4432(.A0(new_n4817_), .A1(new_n1552_), .B0(new_n1893_), .Y(new_n4818_));
  OAI21X1  g4433(.A0(new_n4818_), .A1(new_n1395_), .B0(new_n403_), .Y(new_n4819_));
  AOI21X1  g4434(.A0(new_n4819_), .A1(new_n1393_), .B0(new_n1394_), .Y(new_n4820_));
  OAI21X1  g4435(.A0(new_n4820_), .A1(new_n1392_), .B0(new_n418_), .Y(new_n4821_));
  AOI21X1  g4436(.A0(new_n4821_), .A1(new_n1390_), .B0(new_n1391_), .Y(new_n4822_));
  OAI21X1  g4437(.A0(new_n4822_), .A1(new_n1389_), .B0(new_n433_), .Y(new_n4823_));
  AOI21X1  g4438(.A0(new_n4823_), .A1(new_n1387_), .B0(new_n1388_), .Y(new_n4824_));
  OAI21X1  g4439(.A0(new_n4824_), .A1(new_n1386_), .B0(new_n448_), .Y(new_n4825_));
  AOI21X1  g4440(.A0(new_n4825_), .A1(new_n1384_), .B0(new_n1385_), .Y(new_n4826_));
  OAI21X1  g4441(.A0(new_n4826_), .A1(new_n1383_), .B0(new_n463_), .Y(new_n4827_));
  AOI21X1  g4442(.A0(new_n4827_), .A1(new_n1381_), .B0(new_n1382_), .Y(new_n4828_));
  OAI21X1  g4443(.A0(new_n4828_), .A1(new_n1380_), .B0(new_n478_), .Y(new_n4829_));
  AOI21X1  g4444(.A0(new_n4829_), .A1(new_n1378_), .B0(new_n1379_), .Y(new_n4830_));
  OAI21X1  g4445(.A0(new_n4830_), .A1(new_n1377_), .B0(new_n493_), .Y(new_n4831_));
  AOI21X1  g4446(.A0(new_n4831_), .A1(new_n1375_), .B0(new_n1376_), .Y(new_n4832_));
  OAI21X1  g4447(.A0(new_n4832_), .A1(new_n1374_), .B0(new_n508_), .Y(new_n4833_));
  AOI21X1  g4448(.A0(new_n4833_), .A1(new_n1372_), .B0(new_n1373_), .Y(new_n4834_));
  OAI21X1  g4449(.A0(new_n4834_), .A1(new_n1371_), .B0(new_n523_), .Y(new_n4835_));
  AOI21X1  g4450(.A0(new_n4835_), .A1(new_n1369_), .B0(new_n1370_), .Y(new_n4836_));
  OAI21X1  g4451(.A0(new_n4836_), .A1(new_n1368_), .B0(new_n538_), .Y(new_n4837_));
  AOI21X1  g4452(.A0(new_n4837_), .A1(new_n1366_), .B0(new_n1367_), .Y(new_n4838_));
  OAI21X1  g4453(.A0(new_n4838_), .A1(new_n1365_), .B0(new_n553_), .Y(new_n4839_));
  AOI21X1  g4454(.A0(new_n4839_), .A1(new_n1363_), .B0(new_n1364_), .Y(new_n4840_));
  OAI21X1  g4455(.A0(new_n4840_), .A1(new_n1362_), .B0(new_n568_), .Y(new_n4841_));
  OAI21X1  g4456(.A0(new_n890_), .A1(\priority[77] ), .B0(\req[77] ), .Y(new_n4842_));
  AOI21X1  g4457(.A0(new_n4841_), .A1(new_n1360_), .B0(new_n4842_), .Y(\grant[77] ));
  NOR2X1   g4458(.A(new_n898_), .B(new_n582_), .Y(new_n4844_));
  OAI21X1  g4459(.A0(new_n4844_), .A1(new_n589_), .B0(new_n591_), .Y(new_n4845_));
  AOI21X1  g4460(.A0(new_n4845_), .A1(new_n596_), .B0(new_n599_), .Y(new_n4846_));
  OAI21X1  g4461(.A0(new_n4846_), .A1(new_n604_), .B0(new_n606_), .Y(new_n4847_));
  AOI21X1  g4462(.A0(new_n4847_), .A1(new_n611_), .B0(new_n614_), .Y(new_n4848_));
  OAI21X1  g4463(.A0(new_n4848_), .A1(new_n619_), .B0(new_n621_), .Y(new_n4849_));
  AOI21X1  g4464(.A0(new_n4849_), .A1(new_n626_), .B0(new_n629_), .Y(new_n4850_));
  OAI21X1  g4465(.A0(new_n4850_), .A1(new_n634_), .B0(new_n636_), .Y(new_n4851_));
  AOI21X1  g4466(.A0(new_n4851_), .A1(new_n641_), .B0(new_n644_), .Y(new_n4852_));
  OAI21X1  g4467(.A0(new_n4852_), .A1(new_n649_), .B0(new_n651_), .Y(new_n4853_));
  AOI21X1  g4468(.A0(new_n4853_), .A1(new_n656_), .B0(new_n659_), .Y(new_n4854_));
  OAI21X1  g4469(.A0(new_n4854_), .A1(new_n664_), .B0(new_n666_), .Y(new_n4855_));
  AOI21X1  g4470(.A0(new_n4855_), .A1(new_n671_), .B0(new_n674_), .Y(new_n4856_));
  OAI21X1  g4471(.A0(new_n4856_), .A1(new_n679_), .B0(new_n681_), .Y(new_n4857_));
  AOI21X1  g4472(.A0(new_n4857_), .A1(new_n686_), .B0(new_n689_), .Y(new_n4858_));
  OAI21X1  g4473(.A0(new_n4858_), .A1(new_n694_), .B0(new_n696_), .Y(new_n4859_));
  AOI21X1  g4474(.A0(new_n4859_), .A1(new_n701_), .B0(new_n1662_), .Y(new_n4860_));
  OAI21X1  g4475(.A0(new_n4860_), .A1(new_n1661_), .B0(new_n1705_), .Y(new_n4861_));
  AOI21X1  g4476(.A0(new_n4861_), .A1(new_n1660_), .B0(new_n1938_), .Y(new_n4862_));
  OAI21X1  g4477(.A0(new_n4862_), .A1(new_n1504_), .B0(new_n721_), .Y(new_n4863_));
  AOI21X1  g4478(.A0(new_n4863_), .A1(new_n1502_), .B0(new_n1503_), .Y(new_n4864_));
  OAI21X1  g4479(.A0(new_n4864_), .A1(new_n1501_), .B0(new_n736_), .Y(new_n4865_));
  AOI21X1  g4480(.A0(new_n4865_), .A1(new_n1499_), .B0(new_n1500_), .Y(new_n4866_));
  OAI21X1  g4481(.A0(new_n4866_), .A1(new_n1498_), .B0(new_n751_), .Y(new_n4867_));
  AOI21X1  g4482(.A0(new_n4867_), .A1(new_n1496_), .B0(new_n1497_), .Y(new_n4868_));
  OAI21X1  g4483(.A0(new_n4868_), .A1(new_n1495_), .B0(new_n766_), .Y(new_n4869_));
  AOI21X1  g4484(.A0(new_n4869_), .A1(new_n1493_), .B0(new_n1494_), .Y(new_n4870_));
  OAI21X1  g4485(.A0(new_n4870_), .A1(new_n1492_), .B0(new_n781_), .Y(new_n4871_));
  AOI21X1  g4486(.A0(new_n4871_), .A1(new_n1490_), .B0(new_n1491_), .Y(new_n4872_));
  OAI21X1  g4487(.A0(new_n4872_), .A1(new_n1489_), .B0(new_n796_), .Y(new_n4873_));
  AOI21X1  g4488(.A0(new_n4873_), .A1(new_n1487_), .B0(new_n1488_), .Y(new_n4874_));
  OAI21X1  g4489(.A0(new_n4874_), .A1(new_n1486_), .B0(new_n811_), .Y(new_n4875_));
  AOI21X1  g4490(.A0(new_n4875_), .A1(new_n1484_), .B0(new_n1485_), .Y(new_n4876_));
  OAI21X1  g4491(.A0(new_n4876_), .A1(new_n1483_), .B0(new_n826_), .Y(new_n4877_));
  AOI21X1  g4492(.A0(new_n4877_), .A1(new_n1481_), .B0(new_n1482_), .Y(new_n4878_));
  OAI21X1  g4493(.A0(new_n4878_), .A1(new_n1480_), .B0(new_n841_), .Y(new_n4879_));
  AOI21X1  g4494(.A0(new_n4879_), .A1(new_n1478_), .B0(new_n1479_), .Y(new_n4880_));
  OAI21X1  g4495(.A0(new_n4880_), .A1(new_n1477_), .B0(new_n856_), .Y(new_n4881_));
  AOI21X1  g4496(.A0(new_n4881_), .A1(new_n1475_), .B0(new_n1476_), .Y(new_n4882_));
  OAI21X1  g4497(.A0(new_n4882_), .A1(new_n1474_), .B0(new_n871_), .Y(new_n4883_));
  AOI21X1  g4498(.A0(new_n4883_), .A1(new_n1472_), .B0(new_n1473_), .Y(new_n4884_));
  OAI21X1  g4499(.A0(new_n4884_), .A1(new_n1471_), .B0(new_n886_), .Y(new_n4885_));
  OAI21X1  g4500(.A0(new_n1204_), .A1(\priority[78] ), .B0(\req[78] ), .Y(new_n4886_));
  AOI21X1  g4501(.A0(new_n4885_), .A1(new_n1469_), .B0(new_n4886_), .Y(\grant[78] ));
  NOR2X1   g4502(.A(new_n1212_), .B(new_n900_), .Y(new_n4888_));
  OAI21X1  g4503(.A0(new_n4888_), .A1(new_n907_), .B0(new_n909_), .Y(new_n4889_));
  AOI21X1  g4504(.A0(new_n4889_), .A1(new_n914_), .B0(new_n917_), .Y(new_n4890_));
  OAI21X1  g4505(.A0(new_n4890_), .A1(new_n922_), .B0(new_n924_), .Y(new_n4891_));
  AOI21X1  g4506(.A0(new_n4891_), .A1(new_n929_), .B0(new_n932_), .Y(new_n4892_));
  OAI21X1  g4507(.A0(new_n4892_), .A1(new_n937_), .B0(new_n939_), .Y(new_n4893_));
  AOI21X1  g4508(.A0(new_n4893_), .A1(new_n944_), .B0(new_n947_), .Y(new_n4894_));
  OAI21X1  g4509(.A0(new_n4894_), .A1(new_n952_), .B0(new_n954_), .Y(new_n4895_));
  AOI21X1  g4510(.A0(new_n4895_), .A1(new_n959_), .B0(new_n962_), .Y(new_n4896_));
  OAI21X1  g4511(.A0(new_n4896_), .A1(new_n967_), .B0(new_n969_), .Y(new_n4897_));
  AOI21X1  g4512(.A0(new_n4897_), .A1(new_n974_), .B0(new_n977_), .Y(new_n4898_));
  OAI21X1  g4513(.A0(new_n4898_), .A1(new_n982_), .B0(new_n984_), .Y(new_n4899_));
  AOI21X1  g4514(.A0(new_n4899_), .A1(new_n989_), .B0(new_n992_), .Y(new_n4900_));
  OAI21X1  g4515(.A0(new_n4900_), .A1(new_n997_), .B0(new_n999_), .Y(new_n4901_));
  AOI21X1  g4516(.A0(new_n4901_), .A1(new_n1004_), .B0(new_n1007_), .Y(new_n4902_));
  OAI21X1  g4517(.A0(new_n4902_), .A1(new_n1012_), .B0(new_n1014_), .Y(new_n4903_));
  AOI21X1  g4518(.A0(new_n4903_), .A1(new_n1017_), .B0(new_n1711_), .Y(new_n4904_));
  OAI21X1  g4519(.A0(new_n4904_), .A1(new_n1710_), .B0(new_n1754_), .Y(new_n4905_));
  AOI21X1  g4520(.A0(new_n4905_), .A1(new_n1709_), .B0(new_n1983_), .Y(new_n4906_));
  OAI21X1  g4521(.A0(new_n4906_), .A1(new_n1613_), .B0(new_n1035_), .Y(new_n4907_));
  AOI21X1  g4522(.A0(new_n4907_), .A1(new_n1611_), .B0(new_n1612_), .Y(new_n4908_));
  OAI21X1  g4523(.A0(new_n4908_), .A1(new_n1610_), .B0(new_n1050_), .Y(new_n4909_));
  AOI21X1  g4524(.A0(new_n4909_), .A1(new_n1608_), .B0(new_n1609_), .Y(new_n4910_));
  OAI21X1  g4525(.A0(new_n4910_), .A1(new_n1607_), .B0(new_n1065_), .Y(new_n4911_));
  AOI21X1  g4526(.A0(new_n4911_), .A1(new_n1605_), .B0(new_n1606_), .Y(new_n4912_));
  OAI21X1  g4527(.A0(new_n4912_), .A1(new_n1604_), .B0(new_n1080_), .Y(new_n4913_));
  AOI21X1  g4528(.A0(new_n4913_), .A1(new_n1602_), .B0(new_n1603_), .Y(new_n4914_));
  OAI21X1  g4529(.A0(new_n4914_), .A1(new_n1601_), .B0(new_n1095_), .Y(new_n4915_));
  AOI21X1  g4530(.A0(new_n4915_), .A1(new_n1599_), .B0(new_n1600_), .Y(new_n4916_));
  OAI21X1  g4531(.A0(new_n4916_), .A1(new_n1598_), .B0(new_n1110_), .Y(new_n4917_));
  AOI21X1  g4532(.A0(new_n4917_), .A1(new_n1596_), .B0(new_n1597_), .Y(new_n4918_));
  OAI21X1  g4533(.A0(new_n4918_), .A1(new_n1595_), .B0(new_n1125_), .Y(new_n4919_));
  AOI21X1  g4534(.A0(new_n4919_), .A1(new_n1593_), .B0(new_n1594_), .Y(new_n4920_));
  OAI21X1  g4535(.A0(new_n4920_), .A1(new_n1592_), .B0(new_n1140_), .Y(new_n4921_));
  AOI21X1  g4536(.A0(new_n4921_), .A1(new_n1590_), .B0(new_n1591_), .Y(new_n4922_));
  OAI21X1  g4537(.A0(new_n4922_), .A1(new_n1589_), .B0(new_n1155_), .Y(new_n4923_));
  AOI21X1  g4538(.A0(new_n4923_), .A1(new_n1587_), .B0(new_n1588_), .Y(new_n4924_));
  OAI21X1  g4539(.A0(new_n4924_), .A1(new_n1586_), .B0(new_n1170_), .Y(new_n4925_));
  AOI21X1  g4540(.A0(new_n4925_), .A1(new_n1584_), .B0(new_n1585_), .Y(new_n4926_));
  OAI21X1  g4541(.A0(new_n4926_), .A1(new_n1583_), .B0(new_n1185_), .Y(new_n4927_));
  AOI21X1  g4542(.A0(new_n4927_), .A1(new_n1581_), .B0(new_n1582_), .Y(new_n4928_));
  OAI21X1  g4543(.A0(new_n4928_), .A1(new_n1580_), .B0(new_n1200_), .Y(new_n4929_));
  OAI21X1  g4544(.A0(new_n579_), .A1(\priority[79] ), .B0(\req[79] ), .Y(new_n4930_));
  AOI21X1  g4545(.A0(new_n4929_), .A1(new_n1578_), .B0(new_n4930_), .Y(\grant[79] ));
  NOR2X1   g4546(.A(new_n1214_), .B(new_n588_), .Y(new_n4932_));
  OAI21X1  g4547(.A0(new_n4932_), .A1(new_n1221_), .B0(new_n1223_), .Y(new_n4933_));
  AOI21X1  g4548(.A0(new_n4933_), .A1(new_n1228_), .B0(new_n1231_), .Y(new_n4934_));
  OAI21X1  g4549(.A0(new_n4934_), .A1(new_n1236_), .B0(new_n1238_), .Y(new_n4935_));
  AOI21X1  g4550(.A0(new_n4935_), .A1(new_n1243_), .B0(new_n1246_), .Y(new_n4936_));
  OAI21X1  g4551(.A0(new_n4936_), .A1(new_n1251_), .B0(new_n1253_), .Y(new_n4937_));
  AOI21X1  g4552(.A0(new_n4937_), .A1(new_n1258_), .B0(new_n1261_), .Y(new_n4938_));
  OAI21X1  g4553(.A0(new_n4938_), .A1(new_n1266_), .B0(new_n1268_), .Y(new_n4939_));
  AOI21X1  g4554(.A0(new_n4939_), .A1(new_n1273_), .B0(new_n1276_), .Y(new_n4940_));
  OAI21X1  g4555(.A0(new_n4940_), .A1(new_n1281_), .B0(new_n1283_), .Y(new_n4941_));
  AOI21X1  g4556(.A0(new_n4941_), .A1(new_n1288_), .B0(new_n1291_), .Y(new_n4942_));
  OAI21X1  g4557(.A0(new_n4942_), .A1(new_n1296_), .B0(new_n1298_), .Y(new_n4943_));
  AOI21X1  g4558(.A0(new_n4943_), .A1(new_n1303_), .B0(new_n1306_), .Y(new_n4944_));
  OAI21X1  g4559(.A0(new_n4944_), .A1(new_n1311_), .B0(new_n1313_), .Y(new_n4945_));
  AOI21X1  g4560(.A0(new_n4945_), .A1(new_n1318_), .B0(new_n1321_), .Y(new_n4946_));
  OAI21X1  g4561(.A0(new_n4946_), .A1(new_n1326_), .B0(new_n1328_), .Y(new_n4947_));
  AOI21X1  g4562(.A0(new_n4947_), .A1(new_n1331_), .B0(new_n1758_), .Y(new_n4948_));
  OAI21X1  g4563(.A0(new_n4948_), .A1(new_n394_), .B0(new_n396_), .Y(new_n4949_));
  AOI21X1  g4564(.A0(new_n4949_), .A1(new_n401_), .B0(new_n404_), .Y(new_n4950_));
  OAI21X1  g4565(.A0(new_n4950_), .A1(new_n409_), .B0(new_n411_), .Y(new_n4951_));
  AOI21X1  g4566(.A0(new_n4951_), .A1(new_n416_), .B0(new_n419_), .Y(new_n4952_));
  OAI21X1  g4567(.A0(new_n4952_), .A1(new_n424_), .B0(new_n426_), .Y(new_n4953_));
  AOI21X1  g4568(.A0(new_n4953_), .A1(new_n431_), .B0(new_n434_), .Y(new_n4954_));
  OAI21X1  g4569(.A0(new_n4954_), .A1(new_n439_), .B0(new_n441_), .Y(new_n4955_));
  AOI21X1  g4570(.A0(new_n4955_), .A1(new_n446_), .B0(new_n449_), .Y(new_n4956_));
  OAI21X1  g4571(.A0(new_n4956_), .A1(new_n454_), .B0(new_n456_), .Y(new_n4957_));
  AOI21X1  g4572(.A0(new_n4957_), .A1(new_n461_), .B0(new_n464_), .Y(new_n4958_));
  OAI21X1  g4573(.A0(new_n4958_), .A1(new_n469_), .B0(new_n471_), .Y(new_n4959_));
  AOI21X1  g4574(.A0(new_n4959_), .A1(new_n476_), .B0(new_n479_), .Y(new_n4960_));
  OAI21X1  g4575(.A0(new_n4960_), .A1(new_n484_), .B0(new_n486_), .Y(new_n4961_));
  AOI21X1  g4576(.A0(new_n4961_), .A1(new_n491_), .B0(new_n494_), .Y(new_n4962_));
  OAI21X1  g4577(.A0(new_n4962_), .A1(new_n499_), .B0(new_n501_), .Y(new_n4963_));
  AOI21X1  g4578(.A0(new_n4963_), .A1(new_n506_), .B0(new_n509_), .Y(new_n4964_));
  OAI21X1  g4579(.A0(new_n4964_), .A1(new_n514_), .B0(new_n516_), .Y(new_n4965_));
  AOI21X1  g4580(.A0(new_n4965_), .A1(new_n521_), .B0(new_n524_), .Y(new_n4966_));
  OAI21X1  g4581(.A0(new_n4966_), .A1(new_n529_), .B0(new_n531_), .Y(new_n4967_));
  AOI21X1  g4582(.A0(new_n4967_), .A1(new_n536_), .B0(new_n539_), .Y(new_n4968_));
  OAI21X1  g4583(.A0(new_n4968_), .A1(new_n544_), .B0(new_n546_), .Y(new_n4969_));
  AOI21X1  g4584(.A0(new_n4969_), .A1(new_n551_), .B0(new_n554_), .Y(new_n4970_));
  OAI21X1  g4585(.A0(new_n4970_), .A1(new_n559_), .B0(new_n561_), .Y(new_n4971_));
  AOI21X1  g4586(.A0(new_n4971_), .A1(new_n566_), .B0(new_n569_), .Y(new_n4972_));
  OAI21X1  g4587(.A0(new_n4972_), .A1(new_n574_), .B0(new_n576_), .Y(new_n4973_));
  OAI21X1  g4588(.A0(new_n897_), .A1(\priority[80] ), .B0(\req[80] ), .Y(new_n4974_));
  AOI21X1  g4589(.A0(new_n4973_), .A1(new_n581_), .B0(new_n4974_), .Y(\grant[80] ));
  NOR2X1   g4590(.A(new_n906_), .B(new_n590_), .Y(new_n4976_));
  OAI21X1  g4591(.A0(new_n4976_), .A1(new_n1356_), .B0(new_n598_), .Y(new_n4977_));
  AOI21X1  g4592(.A0(new_n4977_), .A1(new_n1354_), .B0(new_n1355_), .Y(new_n4978_));
  OAI21X1  g4593(.A0(new_n4978_), .A1(new_n1353_), .B0(new_n613_), .Y(new_n4979_));
  AOI21X1  g4594(.A0(new_n4979_), .A1(new_n1351_), .B0(new_n1352_), .Y(new_n4980_));
  OAI21X1  g4595(.A0(new_n4980_), .A1(new_n1350_), .B0(new_n628_), .Y(new_n4981_));
  AOI21X1  g4596(.A0(new_n4981_), .A1(new_n1348_), .B0(new_n1349_), .Y(new_n4982_));
  OAI21X1  g4597(.A0(new_n4982_), .A1(new_n1347_), .B0(new_n643_), .Y(new_n4983_));
  AOI21X1  g4598(.A0(new_n4983_), .A1(new_n1345_), .B0(new_n1346_), .Y(new_n4984_));
  OAI21X1  g4599(.A0(new_n4984_), .A1(new_n1344_), .B0(new_n658_), .Y(new_n4985_));
  AOI21X1  g4600(.A0(new_n4985_), .A1(new_n1342_), .B0(new_n1343_), .Y(new_n4986_));
  OAI21X1  g4601(.A0(new_n4986_), .A1(new_n1341_), .B0(new_n673_), .Y(new_n4987_));
  AOI21X1  g4602(.A0(new_n4987_), .A1(new_n1339_), .B0(new_n1340_), .Y(new_n4988_));
  OAI21X1  g4603(.A0(new_n4988_), .A1(new_n1338_), .B0(new_n688_), .Y(new_n4989_));
  AOI21X1  g4604(.A0(new_n4989_), .A1(new_n1336_), .B0(new_n1337_), .Y(new_n4990_));
  OAI21X1  g4605(.A0(new_n4990_), .A1(new_n1335_), .B0(new_n1438_), .Y(new_n4991_));
  AOI21X1  g4606(.A0(new_n4991_), .A1(new_n1440_), .B0(new_n1803_), .Y(new_n4992_));
  OAI21X1  g4607(.A0(new_n4992_), .A1(new_n712_), .B0(new_n714_), .Y(new_n4993_));
  AOI21X1  g4608(.A0(new_n4993_), .A1(new_n719_), .B0(new_n722_), .Y(new_n4994_));
  OAI21X1  g4609(.A0(new_n4994_), .A1(new_n727_), .B0(new_n729_), .Y(new_n4995_));
  AOI21X1  g4610(.A0(new_n4995_), .A1(new_n734_), .B0(new_n737_), .Y(new_n4996_));
  OAI21X1  g4611(.A0(new_n4996_), .A1(new_n742_), .B0(new_n744_), .Y(new_n4997_));
  AOI21X1  g4612(.A0(new_n4997_), .A1(new_n749_), .B0(new_n752_), .Y(new_n4998_));
  OAI21X1  g4613(.A0(new_n4998_), .A1(new_n757_), .B0(new_n759_), .Y(new_n4999_));
  AOI21X1  g4614(.A0(new_n4999_), .A1(new_n764_), .B0(new_n767_), .Y(new_n5000_));
  OAI21X1  g4615(.A0(new_n5000_), .A1(new_n772_), .B0(new_n774_), .Y(new_n5001_));
  AOI21X1  g4616(.A0(new_n5001_), .A1(new_n779_), .B0(new_n782_), .Y(new_n5002_));
  OAI21X1  g4617(.A0(new_n5002_), .A1(new_n787_), .B0(new_n789_), .Y(new_n5003_));
  AOI21X1  g4618(.A0(new_n5003_), .A1(new_n794_), .B0(new_n797_), .Y(new_n5004_));
  OAI21X1  g4619(.A0(new_n5004_), .A1(new_n802_), .B0(new_n804_), .Y(new_n5005_));
  AOI21X1  g4620(.A0(new_n5005_), .A1(new_n809_), .B0(new_n812_), .Y(new_n5006_));
  OAI21X1  g4621(.A0(new_n5006_), .A1(new_n817_), .B0(new_n819_), .Y(new_n5007_));
  AOI21X1  g4622(.A0(new_n5007_), .A1(new_n824_), .B0(new_n827_), .Y(new_n5008_));
  OAI21X1  g4623(.A0(new_n5008_), .A1(new_n832_), .B0(new_n834_), .Y(new_n5009_));
  AOI21X1  g4624(.A0(new_n5009_), .A1(new_n839_), .B0(new_n842_), .Y(new_n5010_));
  OAI21X1  g4625(.A0(new_n5010_), .A1(new_n847_), .B0(new_n849_), .Y(new_n5011_));
  AOI21X1  g4626(.A0(new_n5011_), .A1(new_n854_), .B0(new_n857_), .Y(new_n5012_));
  OAI21X1  g4627(.A0(new_n5012_), .A1(new_n862_), .B0(new_n864_), .Y(new_n5013_));
  AOI21X1  g4628(.A0(new_n5013_), .A1(new_n869_), .B0(new_n872_), .Y(new_n5014_));
  OAI21X1  g4629(.A0(new_n5014_), .A1(new_n877_), .B0(new_n879_), .Y(new_n5015_));
  AOI21X1  g4630(.A0(new_n5015_), .A1(new_n884_), .B0(new_n887_), .Y(new_n5016_));
  OAI21X1  g4631(.A0(new_n5016_), .A1(new_n892_), .B0(new_n894_), .Y(new_n5017_));
  OAI21X1  g4632(.A0(new_n1211_), .A1(\priority[81] ), .B0(\req[81] ), .Y(new_n5018_));
  AOI21X1  g4633(.A0(new_n5017_), .A1(new_n899_), .B0(new_n5018_), .Y(\grant[81] ));
  NOR2X1   g4634(.A(new_n1220_), .B(new_n908_), .Y(new_n5020_));
  OAI21X1  g4635(.A0(new_n5020_), .A1(new_n1465_), .B0(new_n916_), .Y(new_n5021_));
  AOI21X1  g4636(.A0(new_n5021_), .A1(new_n1463_), .B0(new_n1464_), .Y(new_n5022_));
  OAI21X1  g4637(.A0(new_n5022_), .A1(new_n1462_), .B0(new_n931_), .Y(new_n5023_));
  AOI21X1  g4638(.A0(new_n5023_), .A1(new_n1460_), .B0(new_n1461_), .Y(new_n5024_));
  OAI21X1  g4639(.A0(new_n5024_), .A1(new_n1459_), .B0(new_n946_), .Y(new_n5025_));
  AOI21X1  g4640(.A0(new_n5025_), .A1(new_n1457_), .B0(new_n1458_), .Y(new_n5026_));
  OAI21X1  g4641(.A0(new_n5026_), .A1(new_n1456_), .B0(new_n961_), .Y(new_n5027_));
  AOI21X1  g4642(.A0(new_n5027_), .A1(new_n1454_), .B0(new_n1455_), .Y(new_n5028_));
  OAI21X1  g4643(.A0(new_n5028_), .A1(new_n1453_), .B0(new_n976_), .Y(new_n5029_));
  AOI21X1  g4644(.A0(new_n5029_), .A1(new_n1451_), .B0(new_n1452_), .Y(new_n5030_));
  OAI21X1  g4645(.A0(new_n5030_), .A1(new_n1450_), .B0(new_n991_), .Y(new_n5031_));
  AOI21X1  g4646(.A0(new_n5031_), .A1(new_n1448_), .B0(new_n1449_), .Y(new_n5032_));
  OAI21X1  g4647(.A0(new_n5032_), .A1(new_n1447_), .B0(new_n1006_), .Y(new_n5033_));
  AOI21X1  g4648(.A0(new_n5033_), .A1(new_n1445_), .B0(new_n1446_), .Y(new_n5034_));
  OAI21X1  g4649(.A0(new_n5034_), .A1(new_n1444_), .B0(new_n1547_), .Y(new_n5035_));
  AOI21X1  g4650(.A0(new_n5035_), .A1(new_n1549_), .B0(new_n1848_), .Y(new_n5036_));
  OAI21X1  g4651(.A0(new_n5036_), .A1(new_n1026_), .B0(new_n1028_), .Y(new_n5037_));
  AOI21X1  g4652(.A0(new_n5037_), .A1(new_n1033_), .B0(new_n1036_), .Y(new_n5038_));
  OAI21X1  g4653(.A0(new_n5038_), .A1(new_n1041_), .B0(new_n1043_), .Y(new_n5039_));
  AOI21X1  g4654(.A0(new_n5039_), .A1(new_n1048_), .B0(new_n1051_), .Y(new_n5040_));
  OAI21X1  g4655(.A0(new_n5040_), .A1(new_n1056_), .B0(new_n1058_), .Y(new_n5041_));
  AOI21X1  g4656(.A0(new_n5041_), .A1(new_n1063_), .B0(new_n1066_), .Y(new_n5042_));
  OAI21X1  g4657(.A0(new_n5042_), .A1(new_n1071_), .B0(new_n1073_), .Y(new_n5043_));
  AOI21X1  g4658(.A0(new_n5043_), .A1(new_n1078_), .B0(new_n1081_), .Y(new_n5044_));
  OAI21X1  g4659(.A0(new_n5044_), .A1(new_n1086_), .B0(new_n1088_), .Y(new_n5045_));
  AOI21X1  g4660(.A0(new_n5045_), .A1(new_n1093_), .B0(new_n1096_), .Y(new_n5046_));
  OAI21X1  g4661(.A0(new_n5046_), .A1(new_n1101_), .B0(new_n1103_), .Y(new_n5047_));
  AOI21X1  g4662(.A0(new_n5047_), .A1(new_n1108_), .B0(new_n1111_), .Y(new_n5048_));
  OAI21X1  g4663(.A0(new_n5048_), .A1(new_n1116_), .B0(new_n1118_), .Y(new_n5049_));
  AOI21X1  g4664(.A0(new_n5049_), .A1(new_n1123_), .B0(new_n1126_), .Y(new_n5050_));
  OAI21X1  g4665(.A0(new_n5050_), .A1(new_n1131_), .B0(new_n1133_), .Y(new_n5051_));
  AOI21X1  g4666(.A0(new_n5051_), .A1(new_n1138_), .B0(new_n1141_), .Y(new_n5052_));
  OAI21X1  g4667(.A0(new_n5052_), .A1(new_n1146_), .B0(new_n1148_), .Y(new_n5053_));
  AOI21X1  g4668(.A0(new_n5053_), .A1(new_n1153_), .B0(new_n1156_), .Y(new_n5054_));
  OAI21X1  g4669(.A0(new_n5054_), .A1(new_n1161_), .B0(new_n1163_), .Y(new_n5055_));
  AOI21X1  g4670(.A0(new_n5055_), .A1(new_n1168_), .B0(new_n1171_), .Y(new_n5056_));
  OAI21X1  g4671(.A0(new_n5056_), .A1(new_n1176_), .B0(new_n1178_), .Y(new_n5057_));
  AOI21X1  g4672(.A0(new_n5057_), .A1(new_n1183_), .B0(new_n1186_), .Y(new_n5058_));
  OAI21X1  g4673(.A0(new_n5058_), .A1(new_n1191_), .B0(new_n1193_), .Y(new_n5059_));
  AOI21X1  g4674(.A0(new_n5059_), .A1(new_n1198_), .B0(new_n1201_), .Y(new_n5060_));
  OAI21X1  g4675(.A0(new_n5060_), .A1(new_n1206_), .B0(new_n1208_), .Y(new_n5061_));
  OAI21X1  g4676(.A0(new_n587_), .A1(\priority[82] ), .B0(\req[82] ), .Y(new_n5062_));
  AOI21X1  g4677(.A0(new_n5061_), .A1(new_n1213_), .B0(new_n5062_), .Y(\grant[82] ));
  NOR2X1   g4678(.A(new_n1222_), .B(new_n595_), .Y(new_n5064_));
  OAI21X1  g4679(.A0(new_n5064_), .A1(new_n1574_), .B0(new_n1230_), .Y(new_n5065_));
  AOI21X1  g4680(.A0(new_n5065_), .A1(new_n1572_), .B0(new_n1573_), .Y(new_n5066_));
  OAI21X1  g4681(.A0(new_n5066_), .A1(new_n1571_), .B0(new_n1245_), .Y(new_n5067_));
  AOI21X1  g4682(.A0(new_n5067_), .A1(new_n1569_), .B0(new_n1570_), .Y(new_n5068_));
  OAI21X1  g4683(.A0(new_n5068_), .A1(new_n1568_), .B0(new_n1260_), .Y(new_n5069_));
  AOI21X1  g4684(.A0(new_n5069_), .A1(new_n1566_), .B0(new_n1567_), .Y(new_n5070_));
  OAI21X1  g4685(.A0(new_n5070_), .A1(new_n1565_), .B0(new_n1275_), .Y(new_n5071_));
  AOI21X1  g4686(.A0(new_n5071_), .A1(new_n1563_), .B0(new_n1564_), .Y(new_n5072_));
  OAI21X1  g4687(.A0(new_n5072_), .A1(new_n1562_), .B0(new_n1290_), .Y(new_n5073_));
  AOI21X1  g4688(.A0(new_n5073_), .A1(new_n1560_), .B0(new_n1561_), .Y(new_n5074_));
  OAI21X1  g4689(.A0(new_n5074_), .A1(new_n1559_), .B0(new_n1305_), .Y(new_n5075_));
  AOI21X1  g4690(.A0(new_n5075_), .A1(new_n1557_), .B0(new_n1558_), .Y(new_n5076_));
  OAI21X1  g4691(.A0(new_n5076_), .A1(new_n1556_), .B0(new_n1320_), .Y(new_n5077_));
  AOI21X1  g4692(.A0(new_n5077_), .A1(new_n1554_), .B0(new_n1555_), .Y(new_n5078_));
  OAI21X1  g4693(.A0(new_n5078_), .A1(new_n1553_), .B0(new_n1656_), .Y(new_n5079_));
  AOI21X1  g4694(.A0(new_n5079_), .A1(new_n1552_), .B0(new_n1893_), .Y(new_n5080_));
  OAI21X1  g4695(.A0(new_n5080_), .A1(new_n1395_), .B0(new_n403_), .Y(new_n5081_));
  AOI21X1  g4696(.A0(new_n5081_), .A1(new_n1393_), .B0(new_n1394_), .Y(new_n5082_));
  OAI21X1  g4697(.A0(new_n5082_), .A1(new_n1392_), .B0(new_n418_), .Y(new_n5083_));
  AOI21X1  g4698(.A0(new_n5083_), .A1(new_n1390_), .B0(new_n1391_), .Y(new_n5084_));
  OAI21X1  g4699(.A0(new_n5084_), .A1(new_n1389_), .B0(new_n433_), .Y(new_n5085_));
  AOI21X1  g4700(.A0(new_n5085_), .A1(new_n1387_), .B0(new_n1388_), .Y(new_n5086_));
  OAI21X1  g4701(.A0(new_n5086_), .A1(new_n1386_), .B0(new_n448_), .Y(new_n5087_));
  AOI21X1  g4702(.A0(new_n5087_), .A1(new_n1384_), .B0(new_n1385_), .Y(new_n5088_));
  OAI21X1  g4703(.A0(new_n5088_), .A1(new_n1383_), .B0(new_n463_), .Y(new_n5089_));
  AOI21X1  g4704(.A0(new_n5089_), .A1(new_n1381_), .B0(new_n1382_), .Y(new_n5090_));
  OAI21X1  g4705(.A0(new_n5090_), .A1(new_n1380_), .B0(new_n478_), .Y(new_n5091_));
  AOI21X1  g4706(.A0(new_n5091_), .A1(new_n1378_), .B0(new_n1379_), .Y(new_n5092_));
  OAI21X1  g4707(.A0(new_n5092_), .A1(new_n1377_), .B0(new_n493_), .Y(new_n5093_));
  AOI21X1  g4708(.A0(new_n5093_), .A1(new_n1375_), .B0(new_n1376_), .Y(new_n5094_));
  OAI21X1  g4709(.A0(new_n5094_), .A1(new_n1374_), .B0(new_n508_), .Y(new_n5095_));
  AOI21X1  g4710(.A0(new_n5095_), .A1(new_n1372_), .B0(new_n1373_), .Y(new_n5096_));
  OAI21X1  g4711(.A0(new_n5096_), .A1(new_n1371_), .B0(new_n523_), .Y(new_n5097_));
  AOI21X1  g4712(.A0(new_n5097_), .A1(new_n1369_), .B0(new_n1370_), .Y(new_n5098_));
  OAI21X1  g4713(.A0(new_n5098_), .A1(new_n1368_), .B0(new_n538_), .Y(new_n5099_));
  AOI21X1  g4714(.A0(new_n5099_), .A1(new_n1366_), .B0(new_n1367_), .Y(new_n5100_));
  OAI21X1  g4715(.A0(new_n5100_), .A1(new_n1365_), .B0(new_n553_), .Y(new_n5101_));
  AOI21X1  g4716(.A0(new_n5101_), .A1(new_n1363_), .B0(new_n1364_), .Y(new_n5102_));
  OAI21X1  g4717(.A0(new_n5102_), .A1(new_n1362_), .B0(new_n568_), .Y(new_n5103_));
  AOI21X1  g4718(.A0(new_n5103_), .A1(new_n1360_), .B0(new_n1361_), .Y(new_n5104_));
  OAI21X1  g4719(.A0(new_n5104_), .A1(new_n1359_), .B0(new_n583_), .Y(new_n5105_));
  OAI21X1  g4720(.A0(new_n905_), .A1(\priority[83] ), .B0(\req[83] ), .Y(new_n5106_));
  AOI21X1  g4721(.A0(new_n5105_), .A1(new_n1357_), .B0(new_n5106_), .Y(\grant[83] ));
  NOR2X1   g4722(.A(new_n913_), .B(new_n597_), .Y(new_n5108_));
  OAI21X1  g4723(.A0(new_n5108_), .A1(new_n604_), .B0(new_n606_), .Y(new_n5109_));
  AOI21X1  g4724(.A0(new_n5109_), .A1(new_n611_), .B0(new_n614_), .Y(new_n5110_));
  OAI21X1  g4725(.A0(new_n5110_), .A1(new_n619_), .B0(new_n621_), .Y(new_n5111_));
  AOI21X1  g4726(.A0(new_n5111_), .A1(new_n626_), .B0(new_n629_), .Y(new_n5112_));
  OAI21X1  g4727(.A0(new_n5112_), .A1(new_n634_), .B0(new_n636_), .Y(new_n5113_));
  AOI21X1  g4728(.A0(new_n5113_), .A1(new_n641_), .B0(new_n644_), .Y(new_n5114_));
  OAI21X1  g4729(.A0(new_n5114_), .A1(new_n649_), .B0(new_n651_), .Y(new_n5115_));
  AOI21X1  g4730(.A0(new_n5115_), .A1(new_n656_), .B0(new_n659_), .Y(new_n5116_));
  OAI21X1  g4731(.A0(new_n5116_), .A1(new_n664_), .B0(new_n666_), .Y(new_n5117_));
  AOI21X1  g4732(.A0(new_n5117_), .A1(new_n671_), .B0(new_n674_), .Y(new_n5118_));
  OAI21X1  g4733(.A0(new_n5118_), .A1(new_n679_), .B0(new_n681_), .Y(new_n5119_));
  AOI21X1  g4734(.A0(new_n5119_), .A1(new_n686_), .B0(new_n689_), .Y(new_n5120_));
  OAI21X1  g4735(.A0(new_n5120_), .A1(new_n694_), .B0(new_n696_), .Y(new_n5121_));
  AOI21X1  g4736(.A0(new_n5121_), .A1(new_n701_), .B0(new_n1662_), .Y(new_n5122_));
  OAI21X1  g4737(.A0(new_n5122_), .A1(new_n1661_), .B0(new_n1705_), .Y(new_n5123_));
  AOI21X1  g4738(.A0(new_n5123_), .A1(new_n1660_), .B0(new_n1938_), .Y(new_n5124_));
  OAI21X1  g4739(.A0(new_n5124_), .A1(new_n1504_), .B0(new_n721_), .Y(new_n5125_));
  AOI21X1  g4740(.A0(new_n5125_), .A1(new_n1502_), .B0(new_n1503_), .Y(new_n5126_));
  OAI21X1  g4741(.A0(new_n5126_), .A1(new_n1501_), .B0(new_n736_), .Y(new_n5127_));
  AOI21X1  g4742(.A0(new_n5127_), .A1(new_n1499_), .B0(new_n1500_), .Y(new_n5128_));
  OAI21X1  g4743(.A0(new_n5128_), .A1(new_n1498_), .B0(new_n751_), .Y(new_n5129_));
  AOI21X1  g4744(.A0(new_n5129_), .A1(new_n1496_), .B0(new_n1497_), .Y(new_n5130_));
  OAI21X1  g4745(.A0(new_n5130_), .A1(new_n1495_), .B0(new_n766_), .Y(new_n5131_));
  AOI21X1  g4746(.A0(new_n5131_), .A1(new_n1493_), .B0(new_n1494_), .Y(new_n5132_));
  OAI21X1  g4747(.A0(new_n5132_), .A1(new_n1492_), .B0(new_n781_), .Y(new_n5133_));
  AOI21X1  g4748(.A0(new_n5133_), .A1(new_n1490_), .B0(new_n1491_), .Y(new_n5134_));
  OAI21X1  g4749(.A0(new_n5134_), .A1(new_n1489_), .B0(new_n796_), .Y(new_n5135_));
  AOI21X1  g4750(.A0(new_n5135_), .A1(new_n1487_), .B0(new_n1488_), .Y(new_n5136_));
  OAI21X1  g4751(.A0(new_n5136_), .A1(new_n1486_), .B0(new_n811_), .Y(new_n5137_));
  AOI21X1  g4752(.A0(new_n5137_), .A1(new_n1484_), .B0(new_n1485_), .Y(new_n5138_));
  OAI21X1  g4753(.A0(new_n5138_), .A1(new_n1483_), .B0(new_n826_), .Y(new_n5139_));
  AOI21X1  g4754(.A0(new_n5139_), .A1(new_n1481_), .B0(new_n1482_), .Y(new_n5140_));
  OAI21X1  g4755(.A0(new_n5140_), .A1(new_n1480_), .B0(new_n841_), .Y(new_n5141_));
  AOI21X1  g4756(.A0(new_n5141_), .A1(new_n1478_), .B0(new_n1479_), .Y(new_n5142_));
  OAI21X1  g4757(.A0(new_n5142_), .A1(new_n1477_), .B0(new_n856_), .Y(new_n5143_));
  AOI21X1  g4758(.A0(new_n5143_), .A1(new_n1475_), .B0(new_n1476_), .Y(new_n5144_));
  OAI21X1  g4759(.A0(new_n5144_), .A1(new_n1474_), .B0(new_n871_), .Y(new_n5145_));
  AOI21X1  g4760(.A0(new_n5145_), .A1(new_n1472_), .B0(new_n1473_), .Y(new_n5146_));
  OAI21X1  g4761(.A0(new_n5146_), .A1(new_n1471_), .B0(new_n886_), .Y(new_n5147_));
  AOI21X1  g4762(.A0(new_n5147_), .A1(new_n1469_), .B0(new_n1470_), .Y(new_n5148_));
  OAI21X1  g4763(.A0(new_n5148_), .A1(new_n1468_), .B0(new_n901_), .Y(new_n5149_));
  OAI21X1  g4764(.A0(new_n1219_), .A1(\priority[84] ), .B0(\req[84] ), .Y(new_n5150_));
  AOI21X1  g4765(.A0(new_n5149_), .A1(new_n1466_), .B0(new_n5150_), .Y(\grant[84] ));
  NOR2X1   g4766(.A(new_n1227_), .B(new_n915_), .Y(new_n5152_));
  OAI21X1  g4767(.A0(new_n5152_), .A1(new_n922_), .B0(new_n924_), .Y(new_n5153_));
  AOI21X1  g4768(.A0(new_n5153_), .A1(new_n929_), .B0(new_n932_), .Y(new_n5154_));
  OAI21X1  g4769(.A0(new_n5154_), .A1(new_n937_), .B0(new_n939_), .Y(new_n5155_));
  AOI21X1  g4770(.A0(new_n5155_), .A1(new_n944_), .B0(new_n947_), .Y(new_n5156_));
  OAI21X1  g4771(.A0(new_n5156_), .A1(new_n952_), .B0(new_n954_), .Y(new_n5157_));
  AOI21X1  g4772(.A0(new_n5157_), .A1(new_n959_), .B0(new_n962_), .Y(new_n5158_));
  OAI21X1  g4773(.A0(new_n5158_), .A1(new_n967_), .B0(new_n969_), .Y(new_n5159_));
  AOI21X1  g4774(.A0(new_n5159_), .A1(new_n974_), .B0(new_n977_), .Y(new_n5160_));
  OAI21X1  g4775(.A0(new_n5160_), .A1(new_n982_), .B0(new_n984_), .Y(new_n5161_));
  AOI21X1  g4776(.A0(new_n5161_), .A1(new_n989_), .B0(new_n992_), .Y(new_n5162_));
  OAI21X1  g4777(.A0(new_n5162_), .A1(new_n997_), .B0(new_n999_), .Y(new_n5163_));
  AOI21X1  g4778(.A0(new_n5163_), .A1(new_n1004_), .B0(new_n1007_), .Y(new_n5164_));
  OAI21X1  g4779(.A0(new_n5164_), .A1(new_n1012_), .B0(new_n1014_), .Y(new_n5165_));
  AOI21X1  g4780(.A0(new_n5165_), .A1(new_n1017_), .B0(new_n1711_), .Y(new_n5166_));
  OAI21X1  g4781(.A0(new_n5166_), .A1(new_n1710_), .B0(new_n1754_), .Y(new_n5167_));
  AOI21X1  g4782(.A0(new_n5167_), .A1(new_n1709_), .B0(new_n1983_), .Y(new_n5168_));
  OAI21X1  g4783(.A0(new_n5168_), .A1(new_n1613_), .B0(new_n1035_), .Y(new_n5169_));
  AOI21X1  g4784(.A0(new_n5169_), .A1(new_n1611_), .B0(new_n1612_), .Y(new_n5170_));
  OAI21X1  g4785(.A0(new_n5170_), .A1(new_n1610_), .B0(new_n1050_), .Y(new_n5171_));
  AOI21X1  g4786(.A0(new_n5171_), .A1(new_n1608_), .B0(new_n1609_), .Y(new_n5172_));
  OAI21X1  g4787(.A0(new_n5172_), .A1(new_n1607_), .B0(new_n1065_), .Y(new_n5173_));
  AOI21X1  g4788(.A0(new_n5173_), .A1(new_n1605_), .B0(new_n1606_), .Y(new_n5174_));
  OAI21X1  g4789(.A0(new_n5174_), .A1(new_n1604_), .B0(new_n1080_), .Y(new_n5175_));
  AOI21X1  g4790(.A0(new_n5175_), .A1(new_n1602_), .B0(new_n1603_), .Y(new_n5176_));
  OAI21X1  g4791(.A0(new_n5176_), .A1(new_n1601_), .B0(new_n1095_), .Y(new_n5177_));
  AOI21X1  g4792(.A0(new_n5177_), .A1(new_n1599_), .B0(new_n1600_), .Y(new_n5178_));
  OAI21X1  g4793(.A0(new_n5178_), .A1(new_n1598_), .B0(new_n1110_), .Y(new_n5179_));
  AOI21X1  g4794(.A0(new_n5179_), .A1(new_n1596_), .B0(new_n1597_), .Y(new_n5180_));
  OAI21X1  g4795(.A0(new_n5180_), .A1(new_n1595_), .B0(new_n1125_), .Y(new_n5181_));
  AOI21X1  g4796(.A0(new_n5181_), .A1(new_n1593_), .B0(new_n1594_), .Y(new_n5182_));
  OAI21X1  g4797(.A0(new_n5182_), .A1(new_n1592_), .B0(new_n1140_), .Y(new_n5183_));
  AOI21X1  g4798(.A0(new_n5183_), .A1(new_n1590_), .B0(new_n1591_), .Y(new_n5184_));
  OAI21X1  g4799(.A0(new_n5184_), .A1(new_n1589_), .B0(new_n1155_), .Y(new_n5185_));
  AOI21X1  g4800(.A0(new_n5185_), .A1(new_n1587_), .B0(new_n1588_), .Y(new_n5186_));
  OAI21X1  g4801(.A0(new_n5186_), .A1(new_n1586_), .B0(new_n1170_), .Y(new_n5187_));
  AOI21X1  g4802(.A0(new_n5187_), .A1(new_n1584_), .B0(new_n1585_), .Y(new_n5188_));
  OAI21X1  g4803(.A0(new_n5188_), .A1(new_n1583_), .B0(new_n1185_), .Y(new_n5189_));
  AOI21X1  g4804(.A0(new_n5189_), .A1(new_n1581_), .B0(new_n1582_), .Y(new_n5190_));
  OAI21X1  g4805(.A0(new_n5190_), .A1(new_n1580_), .B0(new_n1200_), .Y(new_n5191_));
  AOI21X1  g4806(.A0(new_n5191_), .A1(new_n1578_), .B0(new_n1579_), .Y(new_n5192_));
  OAI21X1  g4807(.A0(new_n5192_), .A1(new_n1577_), .B0(new_n1215_), .Y(new_n5193_));
  OAI21X1  g4808(.A0(new_n594_), .A1(\priority[85] ), .B0(\req[85] ), .Y(new_n5194_));
  AOI21X1  g4809(.A0(new_n5193_), .A1(new_n1575_), .B0(new_n5194_), .Y(\grant[85] ));
  NOR2X1   g4810(.A(new_n1229_), .B(new_n603_), .Y(new_n5196_));
  OAI21X1  g4811(.A0(new_n5196_), .A1(new_n1236_), .B0(new_n1238_), .Y(new_n5197_));
  AOI21X1  g4812(.A0(new_n5197_), .A1(new_n1243_), .B0(new_n1246_), .Y(new_n5198_));
  OAI21X1  g4813(.A0(new_n5198_), .A1(new_n1251_), .B0(new_n1253_), .Y(new_n5199_));
  AOI21X1  g4814(.A0(new_n5199_), .A1(new_n1258_), .B0(new_n1261_), .Y(new_n5200_));
  OAI21X1  g4815(.A0(new_n5200_), .A1(new_n1266_), .B0(new_n1268_), .Y(new_n5201_));
  AOI21X1  g4816(.A0(new_n5201_), .A1(new_n1273_), .B0(new_n1276_), .Y(new_n5202_));
  OAI21X1  g4817(.A0(new_n5202_), .A1(new_n1281_), .B0(new_n1283_), .Y(new_n5203_));
  AOI21X1  g4818(.A0(new_n5203_), .A1(new_n1288_), .B0(new_n1291_), .Y(new_n5204_));
  OAI21X1  g4819(.A0(new_n5204_), .A1(new_n1296_), .B0(new_n1298_), .Y(new_n5205_));
  AOI21X1  g4820(.A0(new_n5205_), .A1(new_n1303_), .B0(new_n1306_), .Y(new_n5206_));
  OAI21X1  g4821(.A0(new_n5206_), .A1(new_n1311_), .B0(new_n1313_), .Y(new_n5207_));
  AOI21X1  g4822(.A0(new_n5207_), .A1(new_n1318_), .B0(new_n1321_), .Y(new_n5208_));
  OAI21X1  g4823(.A0(new_n5208_), .A1(new_n1326_), .B0(new_n1328_), .Y(new_n5209_));
  AOI21X1  g4824(.A0(new_n5209_), .A1(new_n1331_), .B0(new_n1758_), .Y(new_n5210_));
  OAI21X1  g4825(.A0(new_n5210_), .A1(new_n394_), .B0(new_n396_), .Y(new_n5211_));
  AOI21X1  g4826(.A0(new_n5211_), .A1(new_n401_), .B0(new_n404_), .Y(new_n5212_));
  OAI21X1  g4827(.A0(new_n5212_), .A1(new_n409_), .B0(new_n411_), .Y(new_n5213_));
  AOI21X1  g4828(.A0(new_n5213_), .A1(new_n416_), .B0(new_n419_), .Y(new_n5214_));
  OAI21X1  g4829(.A0(new_n5214_), .A1(new_n424_), .B0(new_n426_), .Y(new_n5215_));
  AOI21X1  g4830(.A0(new_n5215_), .A1(new_n431_), .B0(new_n434_), .Y(new_n5216_));
  OAI21X1  g4831(.A0(new_n5216_), .A1(new_n439_), .B0(new_n441_), .Y(new_n5217_));
  AOI21X1  g4832(.A0(new_n5217_), .A1(new_n446_), .B0(new_n449_), .Y(new_n5218_));
  OAI21X1  g4833(.A0(new_n5218_), .A1(new_n454_), .B0(new_n456_), .Y(new_n5219_));
  AOI21X1  g4834(.A0(new_n5219_), .A1(new_n461_), .B0(new_n464_), .Y(new_n5220_));
  OAI21X1  g4835(.A0(new_n5220_), .A1(new_n469_), .B0(new_n471_), .Y(new_n5221_));
  AOI21X1  g4836(.A0(new_n5221_), .A1(new_n476_), .B0(new_n479_), .Y(new_n5222_));
  OAI21X1  g4837(.A0(new_n5222_), .A1(new_n484_), .B0(new_n486_), .Y(new_n5223_));
  AOI21X1  g4838(.A0(new_n5223_), .A1(new_n491_), .B0(new_n494_), .Y(new_n5224_));
  OAI21X1  g4839(.A0(new_n5224_), .A1(new_n499_), .B0(new_n501_), .Y(new_n5225_));
  AOI21X1  g4840(.A0(new_n5225_), .A1(new_n506_), .B0(new_n509_), .Y(new_n5226_));
  OAI21X1  g4841(.A0(new_n5226_), .A1(new_n514_), .B0(new_n516_), .Y(new_n5227_));
  AOI21X1  g4842(.A0(new_n5227_), .A1(new_n521_), .B0(new_n524_), .Y(new_n5228_));
  OAI21X1  g4843(.A0(new_n5228_), .A1(new_n529_), .B0(new_n531_), .Y(new_n5229_));
  AOI21X1  g4844(.A0(new_n5229_), .A1(new_n536_), .B0(new_n539_), .Y(new_n5230_));
  OAI21X1  g4845(.A0(new_n5230_), .A1(new_n544_), .B0(new_n546_), .Y(new_n5231_));
  AOI21X1  g4846(.A0(new_n5231_), .A1(new_n551_), .B0(new_n554_), .Y(new_n5232_));
  OAI21X1  g4847(.A0(new_n5232_), .A1(new_n559_), .B0(new_n561_), .Y(new_n5233_));
  AOI21X1  g4848(.A0(new_n5233_), .A1(new_n566_), .B0(new_n569_), .Y(new_n5234_));
  OAI21X1  g4849(.A0(new_n5234_), .A1(new_n574_), .B0(new_n576_), .Y(new_n5235_));
  AOI21X1  g4850(.A0(new_n5235_), .A1(new_n581_), .B0(new_n584_), .Y(new_n5236_));
  OAI21X1  g4851(.A0(new_n5236_), .A1(new_n589_), .B0(new_n591_), .Y(new_n5237_));
  OAI21X1  g4852(.A0(new_n912_), .A1(\priority[86] ), .B0(\req[86] ), .Y(new_n5238_));
  AOI21X1  g4853(.A0(new_n5237_), .A1(new_n596_), .B0(new_n5238_), .Y(\grant[86] ));
  NOR2X1   g4854(.A(new_n921_), .B(new_n605_), .Y(new_n5240_));
  OAI21X1  g4855(.A0(new_n5240_), .A1(new_n1353_), .B0(new_n613_), .Y(new_n5241_));
  AOI21X1  g4856(.A0(new_n5241_), .A1(new_n1351_), .B0(new_n1352_), .Y(new_n5242_));
  OAI21X1  g4857(.A0(new_n5242_), .A1(new_n1350_), .B0(new_n628_), .Y(new_n5243_));
  AOI21X1  g4858(.A0(new_n5243_), .A1(new_n1348_), .B0(new_n1349_), .Y(new_n5244_));
  OAI21X1  g4859(.A0(new_n5244_), .A1(new_n1347_), .B0(new_n643_), .Y(new_n5245_));
  AOI21X1  g4860(.A0(new_n5245_), .A1(new_n1345_), .B0(new_n1346_), .Y(new_n5246_));
  OAI21X1  g4861(.A0(new_n5246_), .A1(new_n1344_), .B0(new_n658_), .Y(new_n5247_));
  AOI21X1  g4862(.A0(new_n5247_), .A1(new_n1342_), .B0(new_n1343_), .Y(new_n5248_));
  OAI21X1  g4863(.A0(new_n5248_), .A1(new_n1341_), .B0(new_n673_), .Y(new_n5249_));
  AOI21X1  g4864(.A0(new_n5249_), .A1(new_n1339_), .B0(new_n1340_), .Y(new_n5250_));
  OAI21X1  g4865(.A0(new_n5250_), .A1(new_n1338_), .B0(new_n688_), .Y(new_n5251_));
  AOI21X1  g4866(.A0(new_n5251_), .A1(new_n1336_), .B0(new_n1337_), .Y(new_n5252_));
  OAI21X1  g4867(.A0(new_n5252_), .A1(new_n1335_), .B0(new_n1438_), .Y(new_n5253_));
  AOI21X1  g4868(.A0(new_n5253_), .A1(new_n1440_), .B0(new_n1803_), .Y(new_n5254_));
  OAI21X1  g4869(.A0(new_n5254_), .A1(new_n712_), .B0(new_n714_), .Y(new_n5255_));
  AOI21X1  g4870(.A0(new_n5255_), .A1(new_n719_), .B0(new_n722_), .Y(new_n5256_));
  OAI21X1  g4871(.A0(new_n5256_), .A1(new_n727_), .B0(new_n729_), .Y(new_n5257_));
  AOI21X1  g4872(.A0(new_n5257_), .A1(new_n734_), .B0(new_n737_), .Y(new_n5258_));
  OAI21X1  g4873(.A0(new_n5258_), .A1(new_n742_), .B0(new_n744_), .Y(new_n5259_));
  AOI21X1  g4874(.A0(new_n5259_), .A1(new_n749_), .B0(new_n752_), .Y(new_n5260_));
  OAI21X1  g4875(.A0(new_n5260_), .A1(new_n757_), .B0(new_n759_), .Y(new_n5261_));
  AOI21X1  g4876(.A0(new_n5261_), .A1(new_n764_), .B0(new_n767_), .Y(new_n5262_));
  OAI21X1  g4877(.A0(new_n5262_), .A1(new_n772_), .B0(new_n774_), .Y(new_n5263_));
  AOI21X1  g4878(.A0(new_n5263_), .A1(new_n779_), .B0(new_n782_), .Y(new_n5264_));
  OAI21X1  g4879(.A0(new_n5264_), .A1(new_n787_), .B0(new_n789_), .Y(new_n5265_));
  AOI21X1  g4880(.A0(new_n5265_), .A1(new_n794_), .B0(new_n797_), .Y(new_n5266_));
  OAI21X1  g4881(.A0(new_n5266_), .A1(new_n802_), .B0(new_n804_), .Y(new_n5267_));
  AOI21X1  g4882(.A0(new_n5267_), .A1(new_n809_), .B0(new_n812_), .Y(new_n5268_));
  OAI21X1  g4883(.A0(new_n5268_), .A1(new_n817_), .B0(new_n819_), .Y(new_n5269_));
  AOI21X1  g4884(.A0(new_n5269_), .A1(new_n824_), .B0(new_n827_), .Y(new_n5270_));
  OAI21X1  g4885(.A0(new_n5270_), .A1(new_n832_), .B0(new_n834_), .Y(new_n5271_));
  AOI21X1  g4886(.A0(new_n5271_), .A1(new_n839_), .B0(new_n842_), .Y(new_n5272_));
  OAI21X1  g4887(.A0(new_n5272_), .A1(new_n847_), .B0(new_n849_), .Y(new_n5273_));
  AOI21X1  g4888(.A0(new_n5273_), .A1(new_n854_), .B0(new_n857_), .Y(new_n5274_));
  OAI21X1  g4889(.A0(new_n5274_), .A1(new_n862_), .B0(new_n864_), .Y(new_n5275_));
  AOI21X1  g4890(.A0(new_n5275_), .A1(new_n869_), .B0(new_n872_), .Y(new_n5276_));
  OAI21X1  g4891(.A0(new_n5276_), .A1(new_n877_), .B0(new_n879_), .Y(new_n5277_));
  AOI21X1  g4892(.A0(new_n5277_), .A1(new_n884_), .B0(new_n887_), .Y(new_n5278_));
  OAI21X1  g4893(.A0(new_n5278_), .A1(new_n892_), .B0(new_n894_), .Y(new_n5279_));
  AOI21X1  g4894(.A0(new_n5279_), .A1(new_n899_), .B0(new_n902_), .Y(new_n5280_));
  OAI21X1  g4895(.A0(new_n5280_), .A1(new_n907_), .B0(new_n909_), .Y(new_n5281_));
  OAI21X1  g4896(.A0(new_n1226_), .A1(\priority[87] ), .B0(\req[87] ), .Y(new_n5282_));
  AOI21X1  g4897(.A0(new_n5281_), .A1(new_n914_), .B0(new_n5282_), .Y(\grant[87] ));
  NOR2X1   g4898(.A(new_n1235_), .B(new_n923_), .Y(new_n5284_));
  OAI21X1  g4899(.A0(new_n5284_), .A1(new_n1462_), .B0(new_n931_), .Y(new_n5285_));
  AOI21X1  g4900(.A0(new_n5285_), .A1(new_n1460_), .B0(new_n1461_), .Y(new_n5286_));
  OAI21X1  g4901(.A0(new_n5286_), .A1(new_n1459_), .B0(new_n946_), .Y(new_n5287_));
  AOI21X1  g4902(.A0(new_n5287_), .A1(new_n1457_), .B0(new_n1458_), .Y(new_n5288_));
  OAI21X1  g4903(.A0(new_n5288_), .A1(new_n1456_), .B0(new_n961_), .Y(new_n5289_));
  AOI21X1  g4904(.A0(new_n5289_), .A1(new_n1454_), .B0(new_n1455_), .Y(new_n5290_));
  OAI21X1  g4905(.A0(new_n5290_), .A1(new_n1453_), .B0(new_n976_), .Y(new_n5291_));
  AOI21X1  g4906(.A0(new_n5291_), .A1(new_n1451_), .B0(new_n1452_), .Y(new_n5292_));
  OAI21X1  g4907(.A0(new_n5292_), .A1(new_n1450_), .B0(new_n991_), .Y(new_n5293_));
  AOI21X1  g4908(.A0(new_n5293_), .A1(new_n1448_), .B0(new_n1449_), .Y(new_n5294_));
  OAI21X1  g4909(.A0(new_n5294_), .A1(new_n1447_), .B0(new_n1006_), .Y(new_n5295_));
  AOI21X1  g4910(.A0(new_n5295_), .A1(new_n1445_), .B0(new_n1446_), .Y(new_n5296_));
  OAI21X1  g4911(.A0(new_n5296_), .A1(new_n1444_), .B0(new_n1547_), .Y(new_n5297_));
  AOI21X1  g4912(.A0(new_n5297_), .A1(new_n1549_), .B0(new_n1848_), .Y(new_n5298_));
  OAI21X1  g4913(.A0(new_n5298_), .A1(new_n1026_), .B0(new_n1028_), .Y(new_n5299_));
  AOI21X1  g4914(.A0(new_n5299_), .A1(new_n1033_), .B0(new_n1036_), .Y(new_n5300_));
  OAI21X1  g4915(.A0(new_n5300_), .A1(new_n1041_), .B0(new_n1043_), .Y(new_n5301_));
  AOI21X1  g4916(.A0(new_n5301_), .A1(new_n1048_), .B0(new_n1051_), .Y(new_n5302_));
  OAI21X1  g4917(.A0(new_n5302_), .A1(new_n1056_), .B0(new_n1058_), .Y(new_n5303_));
  AOI21X1  g4918(.A0(new_n5303_), .A1(new_n1063_), .B0(new_n1066_), .Y(new_n5304_));
  OAI21X1  g4919(.A0(new_n5304_), .A1(new_n1071_), .B0(new_n1073_), .Y(new_n5305_));
  AOI21X1  g4920(.A0(new_n5305_), .A1(new_n1078_), .B0(new_n1081_), .Y(new_n5306_));
  OAI21X1  g4921(.A0(new_n5306_), .A1(new_n1086_), .B0(new_n1088_), .Y(new_n5307_));
  AOI21X1  g4922(.A0(new_n5307_), .A1(new_n1093_), .B0(new_n1096_), .Y(new_n5308_));
  OAI21X1  g4923(.A0(new_n5308_), .A1(new_n1101_), .B0(new_n1103_), .Y(new_n5309_));
  AOI21X1  g4924(.A0(new_n5309_), .A1(new_n1108_), .B0(new_n1111_), .Y(new_n5310_));
  OAI21X1  g4925(.A0(new_n5310_), .A1(new_n1116_), .B0(new_n1118_), .Y(new_n5311_));
  AOI21X1  g4926(.A0(new_n5311_), .A1(new_n1123_), .B0(new_n1126_), .Y(new_n5312_));
  OAI21X1  g4927(.A0(new_n5312_), .A1(new_n1131_), .B0(new_n1133_), .Y(new_n5313_));
  AOI21X1  g4928(.A0(new_n5313_), .A1(new_n1138_), .B0(new_n1141_), .Y(new_n5314_));
  OAI21X1  g4929(.A0(new_n5314_), .A1(new_n1146_), .B0(new_n1148_), .Y(new_n5315_));
  AOI21X1  g4930(.A0(new_n5315_), .A1(new_n1153_), .B0(new_n1156_), .Y(new_n5316_));
  OAI21X1  g4931(.A0(new_n5316_), .A1(new_n1161_), .B0(new_n1163_), .Y(new_n5317_));
  AOI21X1  g4932(.A0(new_n5317_), .A1(new_n1168_), .B0(new_n1171_), .Y(new_n5318_));
  OAI21X1  g4933(.A0(new_n5318_), .A1(new_n1176_), .B0(new_n1178_), .Y(new_n5319_));
  AOI21X1  g4934(.A0(new_n5319_), .A1(new_n1183_), .B0(new_n1186_), .Y(new_n5320_));
  OAI21X1  g4935(.A0(new_n5320_), .A1(new_n1191_), .B0(new_n1193_), .Y(new_n5321_));
  AOI21X1  g4936(.A0(new_n5321_), .A1(new_n1198_), .B0(new_n1201_), .Y(new_n5322_));
  OAI21X1  g4937(.A0(new_n5322_), .A1(new_n1206_), .B0(new_n1208_), .Y(new_n5323_));
  AOI21X1  g4938(.A0(new_n5323_), .A1(new_n1213_), .B0(new_n1216_), .Y(new_n5324_));
  OAI21X1  g4939(.A0(new_n5324_), .A1(new_n1221_), .B0(new_n1223_), .Y(new_n5325_));
  OAI21X1  g4940(.A0(new_n602_), .A1(\priority[88] ), .B0(\req[88] ), .Y(new_n5326_));
  AOI21X1  g4941(.A0(new_n5325_), .A1(new_n1228_), .B0(new_n5326_), .Y(\grant[88] ));
  NOR2X1   g4942(.A(new_n1237_), .B(new_n610_), .Y(new_n5328_));
  OAI21X1  g4943(.A0(new_n5328_), .A1(new_n1571_), .B0(new_n1245_), .Y(new_n5329_));
  AOI21X1  g4944(.A0(new_n5329_), .A1(new_n1569_), .B0(new_n1570_), .Y(new_n5330_));
  OAI21X1  g4945(.A0(new_n5330_), .A1(new_n1568_), .B0(new_n1260_), .Y(new_n5331_));
  AOI21X1  g4946(.A0(new_n5331_), .A1(new_n1566_), .B0(new_n1567_), .Y(new_n5332_));
  OAI21X1  g4947(.A0(new_n5332_), .A1(new_n1565_), .B0(new_n1275_), .Y(new_n5333_));
  AOI21X1  g4948(.A0(new_n5333_), .A1(new_n1563_), .B0(new_n1564_), .Y(new_n5334_));
  OAI21X1  g4949(.A0(new_n5334_), .A1(new_n1562_), .B0(new_n1290_), .Y(new_n5335_));
  AOI21X1  g4950(.A0(new_n5335_), .A1(new_n1560_), .B0(new_n1561_), .Y(new_n5336_));
  OAI21X1  g4951(.A0(new_n5336_), .A1(new_n1559_), .B0(new_n1305_), .Y(new_n5337_));
  AOI21X1  g4952(.A0(new_n5337_), .A1(new_n1557_), .B0(new_n1558_), .Y(new_n5338_));
  OAI21X1  g4953(.A0(new_n5338_), .A1(new_n1556_), .B0(new_n1320_), .Y(new_n5339_));
  AOI21X1  g4954(.A0(new_n5339_), .A1(new_n1554_), .B0(new_n1555_), .Y(new_n5340_));
  OAI21X1  g4955(.A0(new_n5340_), .A1(new_n1553_), .B0(new_n1656_), .Y(new_n5341_));
  AOI21X1  g4956(.A0(new_n5341_), .A1(new_n1552_), .B0(new_n1893_), .Y(new_n5342_));
  OAI21X1  g4957(.A0(new_n5342_), .A1(new_n1395_), .B0(new_n403_), .Y(new_n5343_));
  AOI21X1  g4958(.A0(new_n5343_), .A1(new_n1393_), .B0(new_n1394_), .Y(new_n5344_));
  OAI21X1  g4959(.A0(new_n5344_), .A1(new_n1392_), .B0(new_n418_), .Y(new_n5345_));
  AOI21X1  g4960(.A0(new_n5345_), .A1(new_n1390_), .B0(new_n1391_), .Y(new_n5346_));
  OAI21X1  g4961(.A0(new_n5346_), .A1(new_n1389_), .B0(new_n433_), .Y(new_n5347_));
  AOI21X1  g4962(.A0(new_n5347_), .A1(new_n1387_), .B0(new_n1388_), .Y(new_n5348_));
  OAI21X1  g4963(.A0(new_n5348_), .A1(new_n1386_), .B0(new_n448_), .Y(new_n5349_));
  AOI21X1  g4964(.A0(new_n5349_), .A1(new_n1384_), .B0(new_n1385_), .Y(new_n5350_));
  OAI21X1  g4965(.A0(new_n5350_), .A1(new_n1383_), .B0(new_n463_), .Y(new_n5351_));
  AOI21X1  g4966(.A0(new_n5351_), .A1(new_n1381_), .B0(new_n1382_), .Y(new_n5352_));
  OAI21X1  g4967(.A0(new_n5352_), .A1(new_n1380_), .B0(new_n478_), .Y(new_n5353_));
  AOI21X1  g4968(.A0(new_n5353_), .A1(new_n1378_), .B0(new_n1379_), .Y(new_n5354_));
  OAI21X1  g4969(.A0(new_n5354_), .A1(new_n1377_), .B0(new_n493_), .Y(new_n5355_));
  AOI21X1  g4970(.A0(new_n5355_), .A1(new_n1375_), .B0(new_n1376_), .Y(new_n5356_));
  OAI21X1  g4971(.A0(new_n5356_), .A1(new_n1374_), .B0(new_n508_), .Y(new_n5357_));
  AOI21X1  g4972(.A0(new_n5357_), .A1(new_n1372_), .B0(new_n1373_), .Y(new_n5358_));
  OAI21X1  g4973(.A0(new_n5358_), .A1(new_n1371_), .B0(new_n523_), .Y(new_n5359_));
  AOI21X1  g4974(.A0(new_n5359_), .A1(new_n1369_), .B0(new_n1370_), .Y(new_n5360_));
  OAI21X1  g4975(.A0(new_n5360_), .A1(new_n1368_), .B0(new_n538_), .Y(new_n5361_));
  AOI21X1  g4976(.A0(new_n5361_), .A1(new_n1366_), .B0(new_n1367_), .Y(new_n5362_));
  OAI21X1  g4977(.A0(new_n5362_), .A1(new_n1365_), .B0(new_n553_), .Y(new_n5363_));
  AOI21X1  g4978(.A0(new_n5363_), .A1(new_n1363_), .B0(new_n1364_), .Y(new_n5364_));
  OAI21X1  g4979(.A0(new_n5364_), .A1(new_n1362_), .B0(new_n568_), .Y(new_n5365_));
  AOI21X1  g4980(.A0(new_n5365_), .A1(new_n1360_), .B0(new_n1361_), .Y(new_n5366_));
  OAI21X1  g4981(.A0(new_n5366_), .A1(new_n1359_), .B0(new_n583_), .Y(new_n5367_));
  AOI21X1  g4982(.A0(new_n5367_), .A1(new_n1357_), .B0(new_n1358_), .Y(new_n5368_));
  OAI21X1  g4983(.A0(new_n5368_), .A1(new_n1356_), .B0(new_n598_), .Y(new_n5369_));
  OAI21X1  g4984(.A0(new_n920_), .A1(\priority[89] ), .B0(\req[89] ), .Y(new_n5370_));
  AOI21X1  g4985(.A0(new_n5369_), .A1(new_n1354_), .B0(new_n5370_), .Y(\grant[89] ));
  NOR2X1   g4986(.A(new_n928_), .B(new_n612_), .Y(new_n5372_));
  OAI21X1  g4987(.A0(new_n5372_), .A1(new_n619_), .B0(new_n621_), .Y(new_n5373_));
  AOI21X1  g4988(.A0(new_n5373_), .A1(new_n626_), .B0(new_n629_), .Y(new_n5374_));
  OAI21X1  g4989(.A0(new_n5374_), .A1(new_n634_), .B0(new_n636_), .Y(new_n5375_));
  AOI21X1  g4990(.A0(new_n5375_), .A1(new_n641_), .B0(new_n644_), .Y(new_n5376_));
  OAI21X1  g4991(.A0(new_n5376_), .A1(new_n649_), .B0(new_n651_), .Y(new_n5377_));
  AOI21X1  g4992(.A0(new_n5377_), .A1(new_n656_), .B0(new_n659_), .Y(new_n5378_));
  OAI21X1  g4993(.A0(new_n5378_), .A1(new_n664_), .B0(new_n666_), .Y(new_n5379_));
  AOI21X1  g4994(.A0(new_n5379_), .A1(new_n671_), .B0(new_n674_), .Y(new_n5380_));
  OAI21X1  g4995(.A0(new_n5380_), .A1(new_n679_), .B0(new_n681_), .Y(new_n5381_));
  AOI21X1  g4996(.A0(new_n5381_), .A1(new_n686_), .B0(new_n689_), .Y(new_n5382_));
  OAI21X1  g4997(.A0(new_n5382_), .A1(new_n694_), .B0(new_n696_), .Y(new_n5383_));
  AOI21X1  g4998(.A0(new_n5383_), .A1(new_n701_), .B0(new_n1662_), .Y(new_n5384_));
  OAI21X1  g4999(.A0(new_n5384_), .A1(new_n1661_), .B0(new_n1705_), .Y(new_n5385_));
  AOI21X1  g5000(.A0(new_n5385_), .A1(new_n1660_), .B0(new_n1938_), .Y(new_n5386_));
  OAI21X1  g5001(.A0(new_n5386_), .A1(new_n1504_), .B0(new_n721_), .Y(new_n5387_));
  AOI21X1  g5002(.A0(new_n5387_), .A1(new_n1502_), .B0(new_n1503_), .Y(new_n5388_));
  OAI21X1  g5003(.A0(new_n5388_), .A1(new_n1501_), .B0(new_n736_), .Y(new_n5389_));
  AOI21X1  g5004(.A0(new_n5389_), .A1(new_n1499_), .B0(new_n1500_), .Y(new_n5390_));
  OAI21X1  g5005(.A0(new_n5390_), .A1(new_n1498_), .B0(new_n751_), .Y(new_n5391_));
  AOI21X1  g5006(.A0(new_n5391_), .A1(new_n1496_), .B0(new_n1497_), .Y(new_n5392_));
  OAI21X1  g5007(.A0(new_n5392_), .A1(new_n1495_), .B0(new_n766_), .Y(new_n5393_));
  AOI21X1  g5008(.A0(new_n5393_), .A1(new_n1493_), .B0(new_n1494_), .Y(new_n5394_));
  OAI21X1  g5009(.A0(new_n5394_), .A1(new_n1492_), .B0(new_n781_), .Y(new_n5395_));
  AOI21X1  g5010(.A0(new_n5395_), .A1(new_n1490_), .B0(new_n1491_), .Y(new_n5396_));
  OAI21X1  g5011(.A0(new_n5396_), .A1(new_n1489_), .B0(new_n796_), .Y(new_n5397_));
  AOI21X1  g5012(.A0(new_n5397_), .A1(new_n1487_), .B0(new_n1488_), .Y(new_n5398_));
  OAI21X1  g5013(.A0(new_n5398_), .A1(new_n1486_), .B0(new_n811_), .Y(new_n5399_));
  AOI21X1  g5014(.A0(new_n5399_), .A1(new_n1484_), .B0(new_n1485_), .Y(new_n5400_));
  OAI21X1  g5015(.A0(new_n5400_), .A1(new_n1483_), .B0(new_n826_), .Y(new_n5401_));
  AOI21X1  g5016(.A0(new_n5401_), .A1(new_n1481_), .B0(new_n1482_), .Y(new_n5402_));
  OAI21X1  g5017(.A0(new_n5402_), .A1(new_n1480_), .B0(new_n841_), .Y(new_n5403_));
  AOI21X1  g5018(.A0(new_n5403_), .A1(new_n1478_), .B0(new_n1479_), .Y(new_n5404_));
  OAI21X1  g5019(.A0(new_n5404_), .A1(new_n1477_), .B0(new_n856_), .Y(new_n5405_));
  AOI21X1  g5020(.A0(new_n5405_), .A1(new_n1475_), .B0(new_n1476_), .Y(new_n5406_));
  OAI21X1  g5021(.A0(new_n5406_), .A1(new_n1474_), .B0(new_n871_), .Y(new_n5407_));
  AOI21X1  g5022(.A0(new_n5407_), .A1(new_n1472_), .B0(new_n1473_), .Y(new_n5408_));
  OAI21X1  g5023(.A0(new_n5408_), .A1(new_n1471_), .B0(new_n886_), .Y(new_n5409_));
  AOI21X1  g5024(.A0(new_n5409_), .A1(new_n1469_), .B0(new_n1470_), .Y(new_n5410_));
  OAI21X1  g5025(.A0(new_n5410_), .A1(new_n1468_), .B0(new_n901_), .Y(new_n5411_));
  AOI21X1  g5026(.A0(new_n5411_), .A1(new_n1466_), .B0(new_n1467_), .Y(new_n5412_));
  OAI21X1  g5027(.A0(new_n5412_), .A1(new_n1465_), .B0(new_n916_), .Y(new_n5413_));
  OAI21X1  g5028(.A0(new_n1234_), .A1(\priority[90] ), .B0(\req[90] ), .Y(new_n5414_));
  AOI21X1  g5029(.A0(new_n5413_), .A1(new_n1463_), .B0(new_n5414_), .Y(\grant[90] ));
  NOR2X1   g5030(.A(new_n1242_), .B(new_n930_), .Y(new_n5416_));
  OAI21X1  g5031(.A0(new_n5416_), .A1(new_n937_), .B0(new_n939_), .Y(new_n5417_));
  AOI21X1  g5032(.A0(new_n5417_), .A1(new_n944_), .B0(new_n947_), .Y(new_n5418_));
  OAI21X1  g5033(.A0(new_n5418_), .A1(new_n952_), .B0(new_n954_), .Y(new_n5419_));
  AOI21X1  g5034(.A0(new_n5419_), .A1(new_n959_), .B0(new_n962_), .Y(new_n5420_));
  OAI21X1  g5035(.A0(new_n5420_), .A1(new_n967_), .B0(new_n969_), .Y(new_n5421_));
  AOI21X1  g5036(.A0(new_n5421_), .A1(new_n974_), .B0(new_n977_), .Y(new_n5422_));
  OAI21X1  g5037(.A0(new_n5422_), .A1(new_n982_), .B0(new_n984_), .Y(new_n5423_));
  AOI21X1  g5038(.A0(new_n5423_), .A1(new_n989_), .B0(new_n992_), .Y(new_n5424_));
  OAI21X1  g5039(.A0(new_n5424_), .A1(new_n997_), .B0(new_n999_), .Y(new_n5425_));
  AOI21X1  g5040(.A0(new_n5425_), .A1(new_n1004_), .B0(new_n1007_), .Y(new_n5426_));
  OAI21X1  g5041(.A0(new_n5426_), .A1(new_n1012_), .B0(new_n1014_), .Y(new_n5427_));
  AOI21X1  g5042(.A0(new_n5427_), .A1(new_n1017_), .B0(new_n1711_), .Y(new_n5428_));
  OAI21X1  g5043(.A0(new_n5428_), .A1(new_n1710_), .B0(new_n1754_), .Y(new_n5429_));
  AOI21X1  g5044(.A0(new_n5429_), .A1(new_n1709_), .B0(new_n1983_), .Y(new_n5430_));
  OAI21X1  g5045(.A0(new_n5430_), .A1(new_n1613_), .B0(new_n1035_), .Y(new_n5431_));
  AOI21X1  g5046(.A0(new_n5431_), .A1(new_n1611_), .B0(new_n1612_), .Y(new_n5432_));
  OAI21X1  g5047(.A0(new_n5432_), .A1(new_n1610_), .B0(new_n1050_), .Y(new_n5433_));
  AOI21X1  g5048(.A0(new_n5433_), .A1(new_n1608_), .B0(new_n1609_), .Y(new_n5434_));
  OAI21X1  g5049(.A0(new_n5434_), .A1(new_n1607_), .B0(new_n1065_), .Y(new_n5435_));
  AOI21X1  g5050(.A0(new_n5435_), .A1(new_n1605_), .B0(new_n1606_), .Y(new_n5436_));
  OAI21X1  g5051(.A0(new_n5436_), .A1(new_n1604_), .B0(new_n1080_), .Y(new_n5437_));
  AOI21X1  g5052(.A0(new_n5437_), .A1(new_n1602_), .B0(new_n1603_), .Y(new_n5438_));
  OAI21X1  g5053(.A0(new_n5438_), .A1(new_n1601_), .B0(new_n1095_), .Y(new_n5439_));
  AOI21X1  g5054(.A0(new_n5439_), .A1(new_n1599_), .B0(new_n1600_), .Y(new_n5440_));
  OAI21X1  g5055(.A0(new_n5440_), .A1(new_n1598_), .B0(new_n1110_), .Y(new_n5441_));
  AOI21X1  g5056(.A0(new_n5441_), .A1(new_n1596_), .B0(new_n1597_), .Y(new_n5442_));
  OAI21X1  g5057(.A0(new_n5442_), .A1(new_n1595_), .B0(new_n1125_), .Y(new_n5443_));
  AOI21X1  g5058(.A0(new_n5443_), .A1(new_n1593_), .B0(new_n1594_), .Y(new_n5444_));
  OAI21X1  g5059(.A0(new_n5444_), .A1(new_n1592_), .B0(new_n1140_), .Y(new_n5445_));
  AOI21X1  g5060(.A0(new_n5445_), .A1(new_n1590_), .B0(new_n1591_), .Y(new_n5446_));
  OAI21X1  g5061(.A0(new_n5446_), .A1(new_n1589_), .B0(new_n1155_), .Y(new_n5447_));
  AOI21X1  g5062(.A0(new_n5447_), .A1(new_n1587_), .B0(new_n1588_), .Y(new_n5448_));
  OAI21X1  g5063(.A0(new_n5448_), .A1(new_n1586_), .B0(new_n1170_), .Y(new_n5449_));
  AOI21X1  g5064(.A0(new_n5449_), .A1(new_n1584_), .B0(new_n1585_), .Y(new_n5450_));
  OAI21X1  g5065(.A0(new_n5450_), .A1(new_n1583_), .B0(new_n1185_), .Y(new_n5451_));
  AOI21X1  g5066(.A0(new_n5451_), .A1(new_n1581_), .B0(new_n1582_), .Y(new_n5452_));
  OAI21X1  g5067(.A0(new_n5452_), .A1(new_n1580_), .B0(new_n1200_), .Y(new_n5453_));
  AOI21X1  g5068(.A0(new_n5453_), .A1(new_n1578_), .B0(new_n1579_), .Y(new_n5454_));
  OAI21X1  g5069(.A0(new_n5454_), .A1(new_n1577_), .B0(new_n1215_), .Y(new_n5455_));
  AOI21X1  g5070(.A0(new_n5455_), .A1(new_n1575_), .B0(new_n1576_), .Y(new_n5456_));
  OAI21X1  g5071(.A0(new_n5456_), .A1(new_n1574_), .B0(new_n1230_), .Y(new_n5457_));
  OAI21X1  g5072(.A0(new_n609_), .A1(\priority[91] ), .B0(\req[91] ), .Y(new_n5458_));
  AOI21X1  g5073(.A0(new_n5457_), .A1(new_n1572_), .B0(new_n5458_), .Y(\grant[91] ));
  NOR2X1   g5074(.A(new_n1244_), .B(new_n618_), .Y(new_n5460_));
  OAI21X1  g5075(.A0(new_n5460_), .A1(new_n1251_), .B0(new_n1253_), .Y(new_n5461_));
  AOI21X1  g5076(.A0(new_n5461_), .A1(new_n1258_), .B0(new_n1261_), .Y(new_n5462_));
  OAI21X1  g5077(.A0(new_n5462_), .A1(new_n1266_), .B0(new_n1268_), .Y(new_n5463_));
  AOI21X1  g5078(.A0(new_n5463_), .A1(new_n1273_), .B0(new_n1276_), .Y(new_n5464_));
  OAI21X1  g5079(.A0(new_n5464_), .A1(new_n1281_), .B0(new_n1283_), .Y(new_n5465_));
  AOI21X1  g5080(.A0(new_n5465_), .A1(new_n1288_), .B0(new_n1291_), .Y(new_n5466_));
  OAI21X1  g5081(.A0(new_n5466_), .A1(new_n1296_), .B0(new_n1298_), .Y(new_n5467_));
  AOI21X1  g5082(.A0(new_n5467_), .A1(new_n1303_), .B0(new_n1306_), .Y(new_n5468_));
  OAI21X1  g5083(.A0(new_n5468_), .A1(new_n1311_), .B0(new_n1313_), .Y(new_n5469_));
  AOI21X1  g5084(.A0(new_n5469_), .A1(new_n1318_), .B0(new_n1321_), .Y(new_n5470_));
  OAI21X1  g5085(.A0(new_n5470_), .A1(new_n1326_), .B0(new_n1328_), .Y(new_n5471_));
  AOI21X1  g5086(.A0(new_n5471_), .A1(new_n1331_), .B0(new_n1758_), .Y(new_n5472_));
  OAI21X1  g5087(.A0(new_n5472_), .A1(new_n394_), .B0(new_n396_), .Y(new_n5473_));
  AOI21X1  g5088(.A0(new_n5473_), .A1(new_n401_), .B0(new_n404_), .Y(new_n5474_));
  OAI21X1  g5089(.A0(new_n5474_), .A1(new_n409_), .B0(new_n411_), .Y(new_n5475_));
  AOI21X1  g5090(.A0(new_n5475_), .A1(new_n416_), .B0(new_n419_), .Y(new_n5476_));
  OAI21X1  g5091(.A0(new_n5476_), .A1(new_n424_), .B0(new_n426_), .Y(new_n5477_));
  AOI21X1  g5092(.A0(new_n5477_), .A1(new_n431_), .B0(new_n434_), .Y(new_n5478_));
  OAI21X1  g5093(.A0(new_n5478_), .A1(new_n439_), .B0(new_n441_), .Y(new_n5479_));
  AOI21X1  g5094(.A0(new_n5479_), .A1(new_n446_), .B0(new_n449_), .Y(new_n5480_));
  OAI21X1  g5095(.A0(new_n5480_), .A1(new_n454_), .B0(new_n456_), .Y(new_n5481_));
  AOI21X1  g5096(.A0(new_n5481_), .A1(new_n461_), .B0(new_n464_), .Y(new_n5482_));
  OAI21X1  g5097(.A0(new_n5482_), .A1(new_n469_), .B0(new_n471_), .Y(new_n5483_));
  AOI21X1  g5098(.A0(new_n5483_), .A1(new_n476_), .B0(new_n479_), .Y(new_n5484_));
  OAI21X1  g5099(.A0(new_n5484_), .A1(new_n484_), .B0(new_n486_), .Y(new_n5485_));
  AOI21X1  g5100(.A0(new_n5485_), .A1(new_n491_), .B0(new_n494_), .Y(new_n5486_));
  OAI21X1  g5101(.A0(new_n5486_), .A1(new_n499_), .B0(new_n501_), .Y(new_n5487_));
  AOI21X1  g5102(.A0(new_n5487_), .A1(new_n506_), .B0(new_n509_), .Y(new_n5488_));
  OAI21X1  g5103(.A0(new_n5488_), .A1(new_n514_), .B0(new_n516_), .Y(new_n5489_));
  AOI21X1  g5104(.A0(new_n5489_), .A1(new_n521_), .B0(new_n524_), .Y(new_n5490_));
  OAI21X1  g5105(.A0(new_n5490_), .A1(new_n529_), .B0(new_n531_), .Y(new_n5491_));
  AOI21X1  g5106(.A0(new_n5491_), .A1(new_n536_), .B0(new_n539_), .Y(new_n5492_));
  OAI21X1  g5107(.A0(new_n5492_), .A1(new_n544_), .B0(new_n546_), .Y(new_n5493_));
  AOI21X1  g5108(.A0(new_n5493_), .A1(new_n551_), .B0(new_n554_), .Y(new_n5494_));
  OAI21X1  g5109(.A0(new_n5494_), .A1(new_n559_), .B0(new_n561_), .Y(new_n5495_));
  AOI21X1  g5110(.A0(new_n5495_), .A1(new_n566_), .B0(new_n569_), .Y(new_n5496_));
  OAI21X1  g5111(.A0(new_n5496_), .A1(new_n574_), .B0(new_n576_), .Y(new_n5497_));
  AOI21X1  g5112(.A0(new_n5497_), .A1(new_n581_), .B0(new_n584_), .Y(new_n5498_));
  OAI21X1  g5113(.A0(new_n5498_), .A1(new_n589_), .B0(new_n591_), .Y(new_n5499_));
  AOI21X1  g5114(.A0(new_n5499_), .A1(new_n596_), .B0(new_n599_), .Y(new_n5500_));
  OAI21X1  g5115(.A0(new_n5500_), .A1(new_n604_), .B0(new_n606_), .Y(new_n5501_));
  OAI21X1  g5116(.A0(new_n927_), .A1(\priority[92] ), .B0(\req[92] ), .Y(new_n5502_));
  AOI21X1  g5117(.A0(new_n5501_), .A1(new_n611_), .B0(new_n5502_), .Y(\grant[92] ));
  NOR2X1   g5118(.A(new_n936_), .B(new_n620_), .Y(new_n5504_));
  OAI21X1  g5119(.A0(new_n5504_), .A1(new_n1350_), .B0(new_n628_), .Y(new_n5505_));
  AOI21X1  g5120(.A0(new_n5505_), .A1(new_n1348_), .B0(new_n1349_), .Y(new_n5506_));
  OAI21X1  g5121(.A0(new_n5506_), .A1(new_n1347_), .B0(new_n643_), .Y(new_n5507_));
  AOI21X1  g5122(.A0(new_n5507_), .A1(new_n1345_), .B0(new_n1346_), .Y(new_n5508_));
  OAI21X1  g5123(.A0(new_n5508_), .A1(new_n1344_), .B0(new_n658_), .Y(new_n5509_));
  AOI21X1  g5124(.A0(new_n5509_), .A1(new_n1342_), .B0(new_n1343_), .Y(new_n5510_));
  OAI21X1  g5125(.A0(new_n5510_), .A1(new_n1341_), .B0(new_n673_), .Y(new_n5511_));
  AOI21X1  g5126(.A0(new_n5511_), .A1(new_n1339_), .B0(new_n1340_), .Y(new_n5512_));
  OAI21X1  g5127(.A0(new_n5512_), .A1(new_n1338_), .B0(new_n688_), .Y(new_n5513_));
  AOI21X1  g5128(.A0(new_n5513_), .A1(new_n1336_), .B0(new_n1337_), .Y(new_n5514_));
  OAI21X1  g5129(.A0(new_n5514_), .A1(new_n1335_), .B0(new_n1438_), .Y(new_n5515_));
  AOI21X1  g5130(.A0(new_n5515_), .A1(new_n1440_), .B0(new_n1803_), .Y(new_n5516_));
  OAI21X1  g5131(.A0(new_n5516_), .A1(new_n712_), .B0(new_n714_), .Y(new_n5517_));
  AOI21X1  g5132(.A0(new_n5517_), .A1(new_n719_), .B0(new_n722_), .Y(new_n5518_));
  OAI21X1  g5133(.A0(new_n5518_), .A1(new_n727_), .B0(new_n729_), .Y(new_n5519_));
  AOI21X1  g5134(.A0(new_n5519_), .A1(new_n734_), .B0(new_n737_), .Y(new_n5520_));
  OAI21X1  g5135(.A0(new_n5520_), .A1(new_n742_), .B0(new_n744_), .Y(new_n5521_));
  AOI21X1  g5136(.A0(new_n5521_), .A1(new_n749_), .B0(new_n752_), .Y(new_n5522_));
  OAI21X1  g5137(.A0(new_n5522_), .A1(new_n757_), .B0(new_n759_), .Y(new_n5523_));
  AOI21X1  g5138(.A0(new_n5523_), .A1(new_n764_), .B0(new_n767_), .Y(new_n5524_));
  OAI21X1  g5139(.A0(new_n5524_), .A1(new_n772_), .B0(new_n774_), .Y(new_n5525_));
  AOI21X1  g5140(.A0(new_n5525_), .A1(new_n779_), .B0(new_n782_), .Y(new_n5526_));
  OAI21X1  g5141(.A0(new_n5526_), .A1(new_n787_), .B0(new_n789_), .Y(new_n5527_));
  AOI21X1  g5142(.A0(new_n5527_), .A1(new_n794_), .B0(new_n797_), .Y(new_n5528_));
  OAI21X1  g5143(.A0(new_n5528_), .A1(new_n802_), .B0(new_n804_), .Y(new_n5529_));
  AOI21X1  g5144(.A0(new_n5529_), .A1(new_n809_), .B0(new_n812_), .Y(new_n5530_));
  OAI21X1  g5145(.A0(new_n5530_), .A1(new_n817_), .B0(new_n819_), .Y(new_n5531_));
  AOI21X1  g5146(.A0(new_n5531_), .A1(new_n824_), .B0(new_n827_), .Y(new_n5532_));
  OAI21X1  g5147(.A0(new_n5532_), .A1(new_n832_), .B0(new_n834_), .Y(new_n5533_));
  AOI21X1  g5148(.A0(new_n5533_), .A1(new_n839_), .B0(new_n842_), .Y(new_n5534_));
  OAI21X1  g5149(.A0(new_n5534_), .A1(new_n847_), .B0(new_n849_), .Y(new_n5535_));
  AOI21X1  g5150(.A0(new_n5535_), .A1(new_n854_), .B0(new_n857_), .Y(new_n5536_));
  OAI21X1  g5151(.A0(new_n5536_), .A1(new_n862_), .B0(new_n864_), .Y(new_n5537_));
  AOI21X1  g5152(.A0(new_n5537_), .A1(new_n869_), .B0(new_n872_), .Y(new_n5538_));
  OAI21X1  g5153(.A0(new_n5538_), .A1(new_n877_), .B0(new_n879_), .Y(new_n5539_));
  AOI21X1  g5154(.A0(new_n5539_), .A1(new_n884_), .B0(new_n887_), .Y(new_n5540_));
  OAI21X1  g5155(.A0(new_n5540_), .A1(new_n892_), .B0(new_n894_), .Y(new_n5541_));
  AOI21X1  g5156(.A0(new_n5541_), .A1(new_n899_), .B0(new_n902_), .Y(new_n5542_));
  OAI21X1  g5157(.A0(new_n5542_), .A1(new_n907_), .B0(new_n909_), .Y(new_n5543_));
  AOI21X1  g5158(.A0(new_n5543_), .A1(new_n914_), .B0(new_n917_), .Y(new_n5544_));
  OAI21X1  g5159(.A0(new_n5544_), .A1(new_n922_), .B0(new_n924_), .Y(new_n5545_));
  OAI21X1  g5160(.A0(new_n1241_), .A1(\priority[93] ), .B0(\req[93] ), .Y(new_n5546_));
  AOI21X1  g5161(.A0(new_n5545_), .A1(new_n929_), .B0(new_n5546_), .Y(\grant[93] ));
  NOR2X1   g5162(.A(new_n1250_), .B(new_n938_), .Y(new_n5548_));
  OAI21X1  g5163(.A0(new_n5548_), .A1(new_n1459_), .B0(new_n946_), .Y(new_n5549_));
  AOI21X1  g5164(.A0(new_n5549_), .A1(new_n1457_), .B0(new_n1458_), .Y(new_n5550_));
  OAI21X1  g5165(.A0(new_n5550_), .A1(new_n1456_), .B0(new_n961_), .Y(new_n5551_));
  AOI21X1  g5166(.A0(new_n5551_), .A1(new_n1454_), .B0(new_n1455_), .Y(new_n5552_));
  OAI21X1  g5167(.A0(new_n5552_), .A1(new_n1453_), .B0(new_n976_), .Y(new_n5553_));
  AOI21X1  g5168(.A0(new_n5553_), .A1(new_n1451_), .B0(new_n1452_), .Y(new_n5554_));
  OAI21X1  g5169(.A0(new_n5554_), .A1(new_n1450_), .B0(new_n991_), .Y(new_n5555_));
  AOI21X1  g5170(.A0(new_n5555_), .A1(new_n1448_), .B0(new_n1449_), .Y(new_n5556_));
  OAI21X1  g5171(.A0(new_n5556_), .A1(new_n1447_), .B0(new_n1006_), .Y(new_n5557_));
  AOI21X1  g5172(.A0(new_n5557_), .A1(new_n1445_), .B0(new_n1446_), .Y(new_n5558_));
  OAI21X1  g5173(.A0(new_n5558_), .A1(new_n1444_), .B0(new_n1547_), .Y(new_n5559_));
  AOI21X1  g5174(.A0(new_n5559_), .A1(new_n1549_), .B0(new_n1848_), .Y(new_n5560_));
  OAI21X1  g5175(.A0(new_n5560_), .A1(new_n1026_), .B0(new_n1028_), .Y(new_n5561_));
  AOI21X1  g5176(.A0(new_n5561_), .A1(new_n1033_), .B0(new_n1036_), .Y(new_n5562_));
  OAI21X1  g5177(.A0(new_n5562_), .A1(new_n1041_), .B0(new_n1043_), .Y(new_n5563_));
  AOI21X1  g5178(.A0(new_n5563_), .A1(new_n1048_), .B0(new_n1051_), .Y(new_n5564_));
  OAI21X1  g5179(.A0(new_n5564_), .A1(new_n1056_), .B0(new_n1058_), .Y(new_n5565_));
  AOI21X1  g5180(.A0(new_n5565_), .A1(new_n1063_), .B0(new_n1066_), .Y(new_n5566_));
  OAI21X1  g5181(.A0(new_n5566_), .A1(new_n1071_), .B0(new_n1073_), .Y(new_n5567_));
  AOI21X1  g5182(.A0(new_n5567_), .A1(new_n1078_), .B0(new_n1081_), .Y(new_n5568_));
  OAI21X1  g5183(.A0(new_n5568_), .A1(new_n1086_), .B0(new_n1088_), .Y(new_n5569_));
  AOI21X1  g5184(.A0(new_n5569_), .A1(new_n1093_), .B0(new_n1096_), .Y(new_n5570_));
  OAI21X1  g5185(.A0(new_n5570_), .A1(new_n1101_), .B0(new_n1103_), .Y(new_n5571_));
  AOI21X1  g5186(.A0(new_n5571_), .A1(new_n1108_), .B0(new_n1111_), .Y(new_n5572_));
  OAI21X1  g5187(.A0(new_n5572_), .A1(new_n1116_), .B0(new_n1118_), .Y(new_n5573_));
  AOI21X1  g5188(.A0(new_n5573_), .A1(new_n1123_), .B0(new_n1126_), .Y(new_n5574_));
  OAI21X1  g5189(.A0(new_n5574_), .A1(new_n1131_), .B0(new_n1133_), .Y(new_n5575_));
  AOI21X1  g5190(.A0(new_n5575_), .A1(new_n1138_), .B0(new_n1141_), .Y(new_n5576_));
  OAI21X1  g5191(.A0(new_n5576_), .A1(new_n1146_), .B0(new_n1148_), .Y(new_n5577_));
  AOI21X1  g5192(.A0(new_n5577_), .A1(new_n1153_), .B0(new_n1156_), .Y(new_n5578_));
  OAI21X1  g5193(.A0(new_n5578_), .A1(new_n1161_), .B0(new_n1163_), .Y(new_n5579_));
  AOI21X1  g5194(.A0(new_n5579_), .A1(new_n1168_), .B0(new_n1171_), .Y(new_n5580_));
  OAI21X1  g5195(.A0(new_n5580_), .A1(new_n1176_), .B0(new_n1178_), .Y(new_n5581_));
  AOI21X1  g5196(.A0(new_n5581_), .A1(new_n1183_), .B0(new_n1186_), .Y(new_n5582_));
  OAI21X1  g5197(.A0(new_n5582_), .A1(new_n1191_), .B0(new_n1193_), .Y(new_n5583_));
  AOI21X1  g5198(.A0(new_n5583_), .A1(new_n1198_), .B0(new_n1201_), .Y(new_n5584_));
  OAI21X1  g5199(.A0(new_n5584_), .A1(new_n1206_), .B0(new_n1208_), .Y(new_n5585_));
  AOI21X1  g5200(.A0(new_n5585_), .A1(new_n1213_), .B0(new_n1216_), .Y(new_n5586_));
  OAI21X1  g5201(.A0(new_n5586_), .A1(new_n1221_), .B0(new_n1223_), .Y(new_n5587_));
  AOI21X1  g5202(.A0(new_n5587_), .A1(new_n1228_), .B0(new_n1231_), .Y(new_n5588_));
  OAI21X1  g5203(.A0(new_n5588_), .A1(new_n1236_), .B0(new_n1238_), .Y(new_n5589_));
  OAI21X1  g5204(.A0(new_n617_), .A1(\priority[94] ), .B0(\req[94] ), .Y(new_n5590_));
  AOI21X1  g5205(.A0(new_n5589_), .A1(new_n1243_), .B0(new_n5590_), .Y(\grant[94] ));
  NOR2X1   g5206(.A(new_n1252_), .B(new_n625_), .Y(new_n5592_));
  OAI21X1  g5207(.A0(new_n5592_), .A1(new_n1568_), .B0(new_n1260_), .Y(new_n5593_));
  AOI21X1  g5208(.A0(new_n5593_), .A1(new_n1566_), .B0(new_n1567_), .Y(new_n5594_));
  OAI21X1  g5209(.A0(new_n5594_), .A1(new_n1565_), .B0(new_n1275_), .Y(new_n5595_));
  AOI21X1  g5210(.A0(new_n5595_), .A1(new_n1563_), .B0(new_n1564_), .Y(new_n5596_));
  OAI21X1  g5211(.A0(new_n5596_), .A1(new_n1562_), .B0(new_n1290_), .Y(new_n5597_));
  AOI21X1  g5212(.A0(new_n5597_), .A1(new_n1560_), .B0(new_n1561_), .Y(new_n5598_));
  OAI21X1  g5213(.A0(new_n5598_), .A1(new_n1559_), .B0(new_n1305_), .Y(new_n5599_));
  AOI21X1  g5214(.A0(new_n5599_), .A1(new_n1557_), .B0(new_n1558_), .Y(new_n5600_));
  OAI21X1  g5215(.A0(new_n5600_), .A1(new_n1556_), .B0(new_n1320_), .Y(new_n5601_));
  AOI21X1  g5216(.A0(new_n5601_), .A1(new_n1554_), .B0(new_n1555_), .Y(new_n5602_));
  OAI21X1  g5217(.A0(new_n5602_), .A1(new_n1553_), .B0(new_n1656_), .Y(new_n5603_));
  AOI21X1  g5218(.A0(new_n5603_), .A1(new_n1552_), .B0(new_n1893_), .Y(new_n5604_));
  OAI21X1  g5219(.A0(new_n5604_), .A1(new_n1395_), .B0(new_n403_), .Y(new_n5605_));
  AOI21X1  g5220(.A0(new_n5605_), .A1(new_n1393_), .B0(new_n1394_), .Y(new_n5606_));
  OAI21X1  g5221(.A0(new_n5606_), .A1(new_n1392_), .B0(new_n418_), .Y(new_n5607_));
  AOI21X1  g5222(.A0(new_n5607_), .A1(new_n1390_), .B0(new_n1391_), .Y(new_n5608_));
  OAI21X1  g5223(.A0(new_n5608_), .A1(new_n1389_), .B0(new_n433_), .Y(new_n5609_));
  AOI21X1  g5224(.A0(new_n5609_), .A1(new_n1387_), .B0(new_n1388_), .Y(new_n5610_));
  OAI21X1  g5225(.A0(new_n5610_), .A1(new_n1386_), .B0(new_n448_), .Y(new_n5611_));
  AOI21X1  g5226(.A0(new_n5611_), .A1(new_n1384_), .B0(new_n1385_), .Y(new_n5612_));
  OAI21X1  g5227(.A0(new_n5612_), .A1(new_n1383_), .B0(new_n463_), .Y(new_n5613_));
  AOI21X1  g5228(.A0(new_n5613_), .A1(new_n1381_), .B0(new_n1382_), .Y(new_n5614_));
  OAI21X1  g5229(.A0(new_n5614_), .A1(new_n1380_), .B0(new_n478_), .Y(new_n5615_));
  AOI21X1  g5230(.A0(new_n5615_), .A1(new_n1378_), .B0(new_n1379_), .Y(new_n5616_));
  OAI21X1  g5231(.A0(new_n5616_), .A1(new_n1377_), .B0(new_n493_), .Y(new_n5617_));
  AOI21X1  g5232(.A0(new_n5617_), .A1(new_n1375_), .B0(new_n1376_), .Y(new_n5618_));
  OAI21X1  g5233(.A0(new_n5618_), .A1(new_n1374_), .B0(new_n508_), .Y(new_n5619_));
  AOI21X1  g5234(.A0(new_n5619_), .A1(new_n1372_), .B0(new_n1373_), .Y(new_n5620_));
  OAI21X1  g5235(.A0(new_n5620_), .A1(new_n1371_), .B0(new_n523_), .Y(new_n5621_));
  AOI21X1  g5236(.A0(new_n5621_), .A1(new_n1369_), .B0(new_n1370_), .Y(new_n5622_));
  OAI21X1  g5237(.A0(new_n5622_), .A1(new_n1368_), .B0(new_n538_), .Y(new_n5623_));
  AOI21X1  g5238(.A0(new_n5623_), .A1(new_n1366_), .B0(new_n1367_), .Y(new_n5624_));
  OAI21X1  g5239(.A0(new_n5624_), .A1(new_n1365_), .B0(new_n553_), .Y(new_n5625_));
  AOI21X1  g5240(.A0(new_n5625_), .A1(new_n1363_), .B0(new_n1364_), .Y(new_n5626_));
  OAI21X1  g5241(.A0(new_n5626_), .A1(new_n1362_), .B0(new_n568_), .Y(new_n5627_));
  AOI21X1  g5242(.A0(new_n5627_), .A1(new_n1360_), .B0(new_n1361_), .Y(new_n5628_));
  OAI21X1  g5243(.A0(new_n5628_), .A1(new_n1359_), .B0(new_n583_), .Y(new_n5629_));
  AOI21X1  g5244(.A0(new_n5629_), .A1(new_n1357_), .B0(new_n1358_), .Y(new_n5630_));
  OAI21X1  g5245(.A0(new_n5630_), .A1(new_n1356_), .B0(new_n598_), .Y(new_n5631_));
  AOI21X1  g5246(.A0(new_n5631_), .A1(new_n1354_), .B0(new_n1355_), .Y(new_n5632_));
  OAI21X1  g5247(.A0(new_n5632_), .A1(new_n1353_), .B0(new_n613_), .Y(new_n5633_));
  OAI21X1  g5248(.A0(new_n935_), .A1(\priority[95] ), .B0(\req[95] ), .Y(new_n5634_));
  AOI21X1  g5249(.A0(new_n5633_), .A1(new_n1351_), .B0(new_n5634_), .Y(\grant[95] ));
  NOR2X1   g5250(.A(new_n943_), .B(new_n627_), .Y(new_n5636_));
  OAI21X1  g5251(.A0(new_n5636_), .A1(new_n634_), .B0(new_n636_), .Y(new_n5637_));
  AOI21X1  g5252(.A0(new_n5637_), .A1(new_n641_), .B0(new_n644_), .Y(new_n5638_));
  OAI21X1  g5253(.A0(new_n5638_), .A1(new_n649_), .B0(new_n651_), .Y(new_n5639_));
  AOI21X1  g5254(.A0(new_n5639_), .A1(new_n656_), .B0(new_n659_), .Y(new_n5640_));
  OAI21X1  g5255(.A0(new_n5640_), .A1(new_n664_), .B0(new_n666_), .Y(new_n5641_));
  AOI21X1  g5256(.A0(new_n5641_), .A1(new_n671_), .B0(new_n674_), .Y(new_n5642_));
  OAI21X1  g5257(.A0(new_n5642_), .A1(new_n679_), .B0(new_n681_), .Y(new_n5643_));
  AOI21X1  g5258(.A0(new_n5643_), .A1(new_n686_), .B0(new_n689_), .Y(new_n5644_));
  OAI21X1  g5259(.A0(new_n5644_), .A1(new_n694_), .B0(new_n696_), .Y(new_n5645_));
  AOI21X1  g5260(.A0(new_n5645_), .A1(new_n701_), .B0(new_n1662_), .Y(new_n5646_));
  OAI21X1  g5261(.A0(new_n5646_), .A1(new_n1661_), .B0(new_n1705_), .Y(new_n5647_));
  AOI21X1  g5262(.A0(new_n5647_), .A1(new_n1660_), .B0(new_n1938_), .Y(new_n5648_));
  OAI21X1  g5263(.A0(new_n5648_), .A1(new_n1504_), .B0(new_n721_), .Y(new_n5649_));
  AOI21X1  g5264(.A0(new_n5649_), .A1(new_n1502_), .B0(new_n1503_), .Y(new_n5650_));
  OAI21X1  g5265(.A0(new_n5650_), .A1(new_n1501_), .B0(new_n736_), .Y(new_n5651_));
  AOI21X1  g5266(.A0(new_n5651_), .A1(new_n1499_), .B0(new_n1500_), .Y(new_n5652_));
  OAI21X1  g5267(.A0(new_n5652_), .A1(new_n1498_), .B0(new_n751_), .Y(new_n5653_));
  AOI21X1  g5268(.A0(new_n5653_), .A1(new_n1496_), .B0(new_n1497_), .Y(new_n5654_));
  OAI21X1  g5269(.A0(new_n5654_), .A1(new_n1495_), .B0(new_n766_), .Y(new_n5655_));
  AOI21X1  g5270(.A0(new_n5655_), .A1(new_n1493_), .B0(new_n1494_), .Y(new_n5656_));
  OAI21X1  g5271(.A0(new_n5656_), .A1(new_n1492_), .B0(new_n781_), .Y(new_n5657_));
  AOI21X1  g5272(.A0(new_n5657_), .A1(new_n1490_), .B0(new_n1491_), .Y(new_n5658_));
  OAI21X1  g5273(.A0(new_n5658_), .A1(new_n1489_), .B0(new_n796_), .Y(new_n5659_));
  AOI21X1  g5274(.A0(new_n5659_), .A1(new_n1487_), .B0(new_n1488_), .Y(new_n5660_));
  OAI21X1  g5275(.A0(new_n5660_), .A1(new_n1486_), .B0(new_n811_), .Y(new_n5661_));
  AOI21X1  g5276(.A0(new_n5661_), .A1(new_n1484_), .B0(new_n1485_), .Y(new_n5662_));
  OAI21X1  g5277(.A0(new_n5662_), .A1(new_n1483_), .B0(new_n826_), .Y(new_n5663_));
  AOI21X1  g5278(.A0(new_n5663_), .A1(new_n1481_), .B0(new_n1482_), .Y(new_n5664_));
  OAI21X1  g5279(.A0(new_n5664_), .A1(new_n1480_), .B0(new_n841_), .Y(new_n5665_));
  AOI21X1  g5280(.A0(new_n5665_), .A1(new_n1478_), .B0(new_n1479_), .Y(new_n5666_));
  OAI21X1  g5281(.A0(new_n5666_), .A1(new_n1477_), .B0(new_n856_), .Y(new_n5667_));
  AOI21X1  g5282(.A0(new_n5667_), .A1(new_n1475_), .B0(new_n1476_), .Y(new_n5668_));
  OAI21X1  g5283(.A0(new_n5668_), .A1(new_n1474_), .B0(new_n871_), .Y(new_n5669_));
  AOI21X1  g5284(.A0(new_n5669_), .A1(new_n1472_), .B0(new_n1473_), .Y(new_n5670_));
  OAI21X1  g5285(.A0(new_n5670_), .A1(new_n1471_), .B0(new_n886_), .Y(new_n5671_));
  AOI21X1  g5286(.A0(new_n5671_), .A1(new_n1469_), .B0(new_n1470_), .Y(new_n5672_));
  OAI21X1  g5287(.A0(new_n5672_), .A1(new_n1468_), .B0(new_n901_), .Y(new_n5673_));
  AOI21X1  g5288(.A0(new_n5673_), .A1(new_n1466_), .B0(new_n1467_), .Y(new_n5674_));
  OAI21X1  g5289(.A0(new_n5674_), .A1(new_n1465_), .B0(new_n916_), .Y(new_n5675_));
  AOI21X1  g5290(.A0(new_n5675_), .A1(new_n1463_), .B0(new_n1464_), .Y(new_n5676_));
  OAI21X1  g5291(.A0(new_n5676_), .A1(new_n1462_), .B0(new_n931_), .Y(new_n5677_));
  OAI21X1  g5292(.A0(new_n1249_), .A1(\priority[96] ), .B0(\req[96] ), .Y(new_n5678_));
  AOI21X1  g5293(.A0(new_n5677_), .A1(new_n1460_), .B0(new_n5678_), .Y(\grant[96] ));
  NOR2X1   g5294(.A(new_n1257_), .B(new_n945_), .Y(new_n5680_));
  OAI21X1  g5295(.A0(new_n5680_), .A1(new_n952_), .B0(new_n954_), .Y(new_n5681_));
  AOI21X1  g5296(.A0(new_n5681_), .A1(new_n959_), .B0(new_n962_), .Y(new_n5682_));
  OAI21X1  g5297(.A0(new_n5682_), .A1(new_n967_), .B0(new_n969_), .Y(new_n5683_));
  AOI21X1  g5298(.A0(new_n5683_), .A1(new_n974_), .B0(new_n977_), .Y(new_n5684_));
  OAI21X1  g5299(.A0(new_n5684_), .A1(new_n982_), .B0(new_n984_), .Y(new_n5685_));
  AOI21X1  g5300(.A0(new_n5685_), .A1(new_n989_), .B0(new_n992_), .Y(new_n5686_));
  OAI21X1  g5301(.A0(new_n5686_), .A1(new_n997_), .B0(new_n999_), .Y(new_n5687_));
  AOI21X1  g5302(.A0(new_n5687_), .A1(new_n1004_), .B0(new_n1007_), .Y(new_n5688_));
  OAI21X1  g5303(.A0(new_n5688_), .A1(new_n1012_), .B0(new_n1014_), .Y(new_n5689_));
  AOI21X1  g5304(.A0(new_n5689_), .A1(new_n1017_), .B0(new_n1711_), .Y(new_n5690_));
  OAI21X1  g5305(.A0(new_n5690_), .A1(new_n1710_), .B0(new_n1754_), .Y(new_n5691_));
  AOI21X1  g5306(.A0(new_n5691_), .A1(new_n1709_), .B0(new_n1983_), .Y(new_n5692_));
  OAI21X1  g5307(.A0(new_n5692_), .A1(new_n1613_), .B0(new_n1035_), .Y(new_n5693_));
  AOI21X1  g5308(.A0(new_n5693_), .A1(new_n1611_), .B0(new_n1612_), .Y(new_n5694_));
  OAI21X1  g5309(.A0(new_n5694_), .A1(new_n1610_), .B0(new_n1050_), .Y(new_n5695_));
  AOI21X1  g5310(.A0(new_n5695_), .A1(new_n1608_), .B0(new_n1609_), .Y(new_n5696_));
  OAI21X1  g5311(.A0(new_n5696_), .A1(new_n1607_), .B0(new_n1065_), .Y(new_n5697_));
  AOI21X1  g5312(.A0(new_n5697_), .A1(new_n1605_), .B0(new_n1606_), .Y(new_n5698_));
  OAI21X1  g5313(.A0(new_n5698_), .A1(new_n1604_), .B0(new_n1080_), .Y(new_n5699_));
  AOI21X1  g5314(.A0(new_n5699_), .A1(new_n1602_), .B0(new_n1603_), .Y(new_n5700_));
  OAI21X1  g5315(.A0(new_n5700_), .A1(new_n1601_), .B0(new_n1095_), .Y(new_n5701_));
  AOI21X1  g5316(.A0(new_n5701_), .A1(new_n1599_), .B0(new_n1600_), .Y(new_n5702_));
  OAI21X1  g5317(.A0(new_n5702_), .A1(new_n1598_), .B0(new_n1110_), .Y(new_n5703_));
  AOI21X1  g5318(.A0(new_n5703_), .A1(new_n1596_), .B0(new_n1597_), .Y(new_n5704_));
  OAI21X1  g5319(.A0(new_n5704_), .A1(new_n1595_), .B0(new_n1125_), .Y(new_n5705_));
  AOI21X1  g5320(.A0(new_n5705_), .A1(new_n1593_), .B0(new_n1594_), .Y(new_n5706_));
  OAI21X1  g5321(.A0(new_n5706_), .A1(new_n1592_), .B0(new_n1140_), .Y(new_n5707_));
  AOI21X1  g5322(.A0(new_n5707_), .A1(new_n1590_), .B0(new_n1591_), .Y(new_n5708_));
  OAI21X1  g5323(.A0(new_n5708_), .A1(new_n1589_), .B0(new_n1155_), .Y(new_n5709_));
  AOI21X1  g5324(.A0(new_n5709_), .A1(new_n1587_), .B0(new_n1588_), .Y(new_n5710_));
  OAI21X1  g5325(.A0(new_n5710_), .A1(new_n1586_), .B0(new_n1170_), .Y(new_n5711_));
  AOI21X1  g5326(.A0(new_n5711_), .A1(new_n1584_), .B0(new_n1585_), .Y(new_n5712_));
  OAI21X1  g5327(.A0(new_n5712_), .A1(new_n1583_), .B0(new_n1185_), .Y(new_n5713_));
  AOI21X1  g5328(.A0(new_n5713_), .A1(new_n1581_), .B0(new_n1582_), .Y(new_n5714_));
  OAI21X1  g5329(.A0(new_n5714_), .A1(new_n1580_), .B0(new_n1200_), .Y(new_n5715_));
  AOI21X1  g5330(.A0(new_n5715_), .A1(new_n1578_), .B0(new_n1579_), .Y(new_n5716_));
  OAI21X1  g5331(.A0(new_n5716_), .A1(new_n1577_), .B0(new_n1215_), .Y(new_n5717_));
  AOI21X1  g5332(.A0(new_n5717_), .A1(new_n1575_), .B0(new_n1576_), .Y(new_n5718_));
  OAI21X1  g5333(.A0(new_n5718_), .A1(new_n1574_), .B0(new_n1230_), .Y(new_n5719_));
  AOI21X1  g5334(.A0(new_n5719_), .A1(new_n1572_), .B0(new_n1573_), .Y(new_n5720_));
  OAI21X1  g5335(.A0(new_n5720_), .A1(new_n1571_), .B0(new_n1245_), .Y(new_n5721_));
  OAI21X1  g5336(.A0(new_n624_), .A1(\priority[97] ), .B0(\req[97] ), .Y(new_n5722_));
  AOI21X1  g5337(.A0(new_n5721_), .A1(new_n1569_), .B0(new_n5722_), .Y(\grant[97] ));
  NOR2X1   g5338(.A(new_n1259_), .B(new_n633_), .Y(new_n5724_));
  OAI21X1  g5339(.A0(new_n5724_), .A1(new_n1266_), .B0(new_n1268_), .Y(new_n5725_));
  AOI21X1  g5340(.A0(new_n5725_), .A1(new_n1273_), .B0(new_n1276_), .Y(new_n5726_));
  OAI21X1  g5341(.A0(new_n5726_), .A1(new_n1281_), .B0(new_n1283_), .Y(new_n5727_));
  AOI21X1  g5342(.A0(new_n5727_), .A1(new_n1288_), .B0(new_n1291_), .Y(new_n5728_));
  OAI21X1  g5343(.A0(new_n5728_), .A1(new_n1296_), .B0(new_n1298_), .Y(new_n5729_));
  AOI21X1  g5344(.A0(new_n5729_), .A1(new_n1303_), .B0(new_n1306_), .Y(new_n5730_));
  OAI21X1  g5345(.A0(new_n5730_), .A1(new_n1311_), .B0(new_n1313_), .Y(new_n5731_));
  AOI21X1  g5346(.A0(new_n5731_), .A1(new_n1318_), .B0(new_n1321_), .Y(new_n5732_));
  OAI21X1  g5347(.A0(new_n5732_), .A1(new_n1326_), .B0(new_n1328_), .Y(new_n5733_));
  AOI21X1  g5348(.A0(new_n5733_), .A1(new_n1331_), .B0(new_n1758_), .Y(new_n5734_));
  OAI21X1  g5349(.A0(new_n5734_), .A1(new_n394_), .B0(new_n396_), .Y(new_n5735_));
  AOI21X1  g5350(.A0(new_n5735_), .A1(new_n401_), .B0(new_n404_), .Y(new_n5736_));
  OAI21X1  g5351(.A0(new_n5736_), .A1(new_n409_), .B0(new_n411_), .Y(new_n5737_));
  AOI21X1  g5352(.A0(new_n5737_), .A1(new_n416_), .B0(new_n419_), .Y(new_n5738_));
  OAI21X1  g5353(.A0(new_n5738_), .A1(new_n424_), .B0(new_n426_), .Y(new_n5739_));
  AOI21X1  g5354(.A0(new_n5739_), .A1(new_n431_), .B0(new_n434_), .Y(new_n5740_));
  OAI21X1  g5355(.A0(new_n5740_), .A1(new_n439_), .B0(new_n441_), .Y(new_n5741_));
  AOI21X1  g5356(.A0(new_n5741_), .A1(new_n446_), .B0(new_n449_), .Y(new_n5742_));
  OAI21X1  g5357(.A0(new_n5742_), .A1(new_n454_), .B0(new_n456_), .Y(new_n5743_));
  AOI21X1  g5358(.A0(new_n5743_), .A1(new_n461_), .B0(new_n464_), .Y(new_n5744_));
  OAI21X1  g5359(.A0(new_n5744_), .A1(new_n469_), .B0(new_n471_), .Y(new_n5745_));
  AOI21X1  g5360(.A0(new_n5745_), .A1(new_n476_), .B0(new_n479_), .Y(new_n5746_));
  OAI21X1  g5361(.A0(new_n5746_), .A1(new_n484_), .B0(new_n486_), .Y(new_n5747_));
  AOI21X1  g5362(.A0(new_n5747_), .A1(new_n491_), .B0(new_n494_), .Y(new_n5748_));
  OAI21X1  g5363(.A0(new_n5748_), .A1(new_n499_), .B0(new_n501_), .Y(new_n5749_));
  AOI21X1  g5364(.A0(new_n5749_), .A1(new_n506_), .B0(new_n509_), .Y(new_n5750_));
  OAI21X1  g5365(.A0(new_n5750_), .A1(new_n514_), .B0(new_n516_), .Y(new_n5751_));
  AOI21X1  g5366(.A0(new_n5751_), .A1(new_n521_), .B0(new_n524_), .Y(new_n5752_));
  OAI21X1  g5367(.A0(new_n5752_), .A1(new_n529_), .B0(new_n531_), .Y(new_n5753_));
  AOI21X1  g5368(.A0(new_n5753_), .A1(new_n536_), .B0(new_n539_), .Y(new_n5754_));
  OAI21X1  g5369(.A0(new_n5754_), .A1(new_n544_), .B0(new_n546_), .Y(new_n5755_));
  AOI21X1  g5370(.A0(new_n5755_), .A1(new_n551_), .B0(new_n554_), .Y(new_n5756_));
  OAI21X1  g5371(.A0(new_n5756_), .A1(new_n559_), .B0(new_n561_), .Y(new_n5757_));
  AOI21X1  g5372(.A0(new_n5757_), .A1(new_n566_), .B0(new_n569_), .Y(new_n5758_));
  OAI21X1  g5373(.A0(new_n5758_), .A1(new_n574_), .B0(new_n576_), .Y(new_n5759_));
  AOI21X1  g5374(.A0(new_n5759_), .A1(new_n581_), .B0(new_n584_), .Y(new_n5760_));
  OAI21X1  g5375(.A0(new_n5760_), .A1(new_n589_), .B0(new_n591_), .Y(new_n5761_));
  AOI21X1  g5376(.A0(new_n5761_), .A1(new_n596_), .B0(new_n599_), .Y(new_n5762_));
  OAI21X1  g5377(.A0(new_n5762_), .A1(new_n604_), .B0(new_n606_), .Y(new_n5763_));
  AOI21X1  g5378(.A0(new_n5763_), .A1(new_n611_), .B0(new_n614_), .Y(new_n5764_));
  OAI21X1  g5379(.A0(new_n5764_), .A1(new_n619_), .B0(new_n621_), .Y(new_n5765_));
  OAI21X1  g5380(.A0(new_n942_), .A1(\priority[98] ), .B0(\req[98] ), .Y(new_n5766_));
  AOI21X1  g5381(.A0(new_n5765_), .A1(new_n626_), .B0(new_n5766_), .Y(\grant[98] ));
  NOR2X1   g5382(.A(new_n951_), .B(new_n635_), .Y(new_n5768_));
  OAI21X1  g5383(.A0(new_n5768_), .A1(new_n1347_), .B0(new_n643_), .Y(new_n5769_));
  AOI21X1  g5384(.A0(new_n5769_), .A1(new_n1345_), .B0(new_n1346_), .Y(new_n5770_));
  OAI21X1  g5385(.A0(new_n5770_), .A1(new_n1344_), .B0(new_n658_), .Y(new_n5771_));
  AOI21X1  g5386(.A0(new_n5771_), .A1(new_n1342_), .B0(new_n1343_), .Y(new_n5772_));
  OAI21X1  g5387(.A0(new_n5772_), .A1(new_n1341_), .B0(new_n673_), .Y(new_n5773_));
  AOI21X1  g5388(.A0(new_n5773_), .A1(new_n1339_), .B0(new_n1340_), .Y(new_n5774_));
  OAI21X1  g5389(.A0(new_n5774_), .A1(new_n1338_), .B0(new_n688_), .Y(new_n5775_));
  AOI21X1  g5390(.A0(new_n5775_), .A1(new_n1336_), .B0(new_n1337_), .Y(new_n5776_));
  OAI21X1  g5391(.A0(new_n5776_), .A1(new_n1335_), .B0(new_n1438_), .Y(new_n5777_));
  AOI21X1  g5392(.A0(new_n5777_), .A1(new_n1440_), .B0(new_n1803_), .Y(new_n5778_));
  OAI21X1  g5393(.A0(new_n5778_), .A1(new_n712_), .B0(new_n714_), .Y(new_n5779_));
  AOI21X1  g5394(.A0(new_n5779_), .A1(new_n719_), .B0(new_n722_), .Y(new_n5780_));
  OAI21X1  g5395(.A0(new_n5780_), .A1(new_n727_), .B0(new_n729_), .Y(new_n5781_));
  AOI21X1  g5396(.A0(new_n5781_), .A1(new_n734_), .B0(new_n737_), .Y(new_n5782_));
  OAI21X1  g5397(.A0(new_n5782_), .A1(new_n742_), .B0(new_n744_), .Y(new_n5783_));
  AOI21X1  g5398(.A0(new_n5783_), .A1(new_n749_), .B0(new_n752_), .Y(new_n5784_));
  OAI21X1  g5399(.A0(new_n5784_), .A1(new_n757_), .B0(new_n759_), .Y(new_n5785_));
  AOI21X1  g5400(.A0(new_n5785_), .A1(new_n764_), .B0(new_n767_), .Y(new_n5786_));
  OAI21X1  g5401(.A0(new_n5786_), .A1(new_n772_), .B0(new_n774_), .Y(new_n5787_));
  AOI21X1  g5402(.A0(new_n5787_), .A1(new_n779_), .B0(new_n782_), .Y(new_n5788_));
  OAI21X1  g5403(.A0(new_n5788_), .A1(new_n787_), .B0(new_n789_), .Y(new_n5789_));
  AOI21X1  g5404(.A0(new_n5789_), .A1(new_n794_), .B0(new_n797_), .Y(new_n5790_));
  OAI21X1  g5405(.A0(new_n5790_), .A1(new_n802_), .B0(new_n804_), .Y(new_n5791_));
  AOI21X1  g5406(.A0(new_n5791_), .A1(new_n809_), .B0(new_n812_), .Y(new_n5792_));
  OAI21X1  g5407(.A0(new_n5792_), .A1(new_n817_), .B0(new_n819_), .Y(new_n5793_));
  AOI21X1  g5408(.A0(new_n5793_), .A1(new_n824_), .B0(new_n827_), .Y(new_n5794_));
  OAI21X1  g5409(.A0(new_n5794_), .A1(new_n832_), .B0(new_n834_), .Y(new_n5795_));
  AOI21X1  g5410(.A0(new_n5795_), .A1(new_n839_), .B0(new_n842_), .Y(new_n5796_));
  OAI21X1  g5411(.A0(new_n5796_), .A1(new_n847_), .B0(new_n849_), .Y(new_n5797_));
  AOI21X1  g5412(.A0(new_n5797_), .A1(new_n854_), .B0(new_n857_), .Y(new_n5798_));
  OAI21X1  g5413(.A0(new_n5798_), .A1(new_n862_), .B0(new_n864_), .Y(new_n5799_));
  AOI21X1  g5414(.A0(new_n5799_), .A1(new_n869_), .B0(new_n872_), .Y(new_n5800_));
  OAI21X1  g5415(.A0(new_n5800_), .A1(new_n877_), .B0(new_n879_), .Y(new_n5801_));
  AOI21X1  g5416(.A0(new_n5801_), .A1(new_n884_), .B0(new_n887_), .Y(new_n5802_));
  OAI21X1  g5417(.A0(new_n5802_), .A1(new_n892_), .B0(new_n894_), .Y(new_n5803_));
  AOI21X1  g5418(.A0(new_n5803_), .A1(new_n899_), .B0(new_n902_), .Y(new_n5804_));
  OAI21X1  g5419(.A0(new_n5804_), .A1(new_n907_), .B0(new_n909_), .Y(new_n5805_));
  AOI21X1  g5420(.A0(new_n5805_), .A1(new_n914_), .B0(new_n917_), .Y(new_n5806_));
  OAI21X1  g5421(.A0(new_n5806_), .A1(new_n922_), .B0(new_n924_), .Y(new_n5807_));
  AOI21X1  g5422(.A0(new_n5807_), .A1(new_n929_), .B0(new_n932_), .Y(new_n5808_));
  OAI21X1  g5423(.A0(new_n5808_), .A1(new_n937_), .B0(new_n939_), .Y(new_n5809_));
  OAI21X1  g5424(.A0(new_n1256_), .A1(\priority[99] ), .B0(\req[99] ), .Y(new_n5810_));
  AOI21X1  g5425(.A0(new_n5809_), .A1(new_n944_), .B0(new_n5810_), .Y(\grant[99] ));
  NOR2X1   g5426(.A(new_n1265_), .B(new_n953_), .Y(new_n5812_));
  OAI21X1  g5427(.A0(new_n5812_), .A1(new_n1456_), .B0(new_n961_), .Y(new_n5813_));
  AOI21X1  g5428(.A0(new_n5813_), .A1(new_n1454_), .B0(new_n1455_), .Y(new_n5814_));
  OAI21X1  g5429(.A0(new_n5814_), .A1(new_n1453_), .B0(new_n976_), .Y(new_n5815_));
  AOI21X1  g5430(.A0(new_n5815_), .A1(new_n1451_), .B0(new_n1452_), .Y(new_n5816_));
  OAI21X1  g5431(.A0(new_n5816_), .A1(new_n1450_), .B0(new_n991_), .Y(new_n5817_));
  AOI21X1  g5432(.A0(new_n5817_), .A1(new_n1448_), .B0(new_n1449_), .Y(new_n5818_));
  OAI21X1  g5433(.A0(new_n5818_), .A1(new_n1447_), .B0(new_n1006_), .Y(new_n5819_));
  AOI21X1  g5434(.A0(new_n5819_), .A1(new_n1445_), .B0(new_n1446_), .Y(new_n5820_));
  OAI21X1  g5435(.A0(new_n5820_), .A1(new_n1444_), .B0(new_n1547_), .Y(new_n5821_));
  AOI21X1  g5436(.A0(new_n5821_), .A1(new_n1549_), .B0(new_n1848_), .Y(new_n5822_));
  OAI21X1  g5437(.A0(new_n5822_), .A1(new_n1026_), .B0(new_n1028_), .Y(new_n5823_));
  AOI21X1  g5438(.A0(new_n5823_), .A1(new_n1033_), .B0(new_n1036_), .Y(new_n5824_));
  OAI21X1  g5439(.A0(new_n5824_), .A1(new_n1041_), .B0(new_n1043_), .Y(new_n5825_));
  AOI21X1  g5440(.A0(new_n5825_), .A1(new_n1048_), .B0(new_n1051_), .Y(new_n5826_));
  OAI21X1  g5441(.A0(new_n5826_), .A1(new_n1056_), .B0(new_n1058_), .Y(new_n5827_));
  AOI21X1  g5442(.A0(new_n5827_), .A1(new_n1063_), .B0(new_n1066_), .Y(new_n5828_));
  OAI21X1  g5443(.A0(new_n5828_), .A1(new_n1071_), .B0(new_n1073_), .Y(new_n5829_));
  AOI21X1  g5444(.A0(new_n5829_), .A1(new_n1078_), .B0(new_n1081_), .Y(new_n5830_));
  OAI21X1  g5445(.A0(new_n5830_), .A1(new_n1086_), .B0(new_n1088_), .Y(new_n5831_));
  AOI21X1  g5446(.A0(new_n5831_), .A1(new_n1093_), .B0(new_n1096_), .Y(new_n5832_));
  OAI21X1  g5447(.A0(new_n5832_), .A1(new_n1101_), .B0(new_n1103_), .Y(new_n5833_));
  AOI21X1  g5448(.A0(new_n5833_), .A1(new_n1108_), .B0(new_n1111_), .Y(new_n5834_));
  OAI21X1  g5449(.A0(new_n5834_), .A1(new_n1116_), .B0(new_n1118_), .Y(new_n5835_));
  AOI21X1  g5450(.A0(new_n5835_), .A1(new_n1123_), .B0(new_n1126_), .Y(new_n5836_));
  OAI21X1  g5451(.A0(new_n5836_), .A1(new_n1131_), .B0(new_n1133_), .Y(new_n5837_));
  AOI21X1  g5452(.A0(new_n5837_), .A1(new_n1138_), .B0(new_n1141_), .Y(new_n5838_));
  OAI21X1  g5453(.A0(new_n5838_), .A1(new_n1146_), .B0(new_n1148_), .Y(new_n5839_));
  AOI21X1  g5454(.A0(new_n5839_), .A1(new_n1153_), .B0(new_n1156_), .Y(new_n5840_));
  OAI21X1  g5455(.A0(new_n5840_), .A1(new_n1161_), .B0(new_n1163_), .Y(new_n5841_));
  AOI21X1  g5456(.A0(new_n5841_), .A1(new_n1168_), .B0(new_n1171_), .Y(new_n5842_));
  OAI21X1  g5457(.A0(new_n5842_), .A1(new_n1176_), .B0(new_n1178_), .Y(new_n5843_));
  AOI21X1  g5458(.A0(new_n5843_), .A1(new_n1183_), .B0(new_n1186_), .Y(new_n5844_));
  OAI21X1  g5459(.A0(new_n5844_), .A1(new_n1191_), .B0(new_n1193_), .Y(new_n5845_));
  AOI21X1  g5460(.A0(new_n5845_), .A1(new_n1198_), .B0(new_n1201_), .Y(new_n5846_));
  OAI21X1  g5461(.A0(new_n5846_), .A1(new_n1206_), .B0(new_n1208_), .Y(new_n5847_));
  AOI21X1  g5462(.A0(new_n5847_), .A1(new_n1213_), .B0(new_n1216_), .Y(new_n5848_));
  OAI21X1  g5463(.A0(new_n5848_), .A1(new_n1221_), .B0(new_n1223_), .Y(new_n5849_));
  AOI21X1  g5464(.A0(new_n5849_), .A1(new_n1228_), .B0(new_n1231_), .Y(new_n5850_));
  OAI21X1  g5465(.A0(new_n5850_), .A1(new_n1236_), .B0(new_n1238_), .Y(new_n5851_));
  AOI21X1  g5466(.A0(new_n5851_), .A1(new_n1243_), .B0(new_n1246_), .Y(new_n5852_));
  OAI21X1  g5467(.A0(new_n5852_), .A1(new_n1251_), .B0(new_n1253_), .Y(new_n5853_));
  OAI21X1  g5468(.A0(new_n632_), .A1(\priority[100] ), .B0(\req[100] ), .Y(new_n5854_));
  AOI21X1  g5469(.A0(new_n5853_), .A1(new_n1258_), .B0(new_n5854_), .Y(\grant[100] ));
  NOR2X1   g5470(.A(new_n1267_), .B(new_n640_), .Y(new_n5856_));
  OAI21X1  g5471(.A0(new_n5856_), .A1(new_n1565_), .B0(new_n1275_), .Y(new_n5857_));
  AOI21X1  g5472(.A0(new_n5857_), .A1(new_n1563_), .B0(new_n1564_), .Y(new_n5858_));
  OAI21X1  g5473(.A0(new_n5858_), .A1(new_n1562_), .B0(new_n1290_), .Y(new_n5859_));
  AOI21X1  g5474(.A0(new_n5859_), .A1(new_n1560_), .B0(new_n1561_), .Y(new_n5860_));
  OAI21X1  g5475(.A0(new_n5860_), .A1(new_n1559_), .B0(new_n1305_), .Y(new_n5861_));
  AOI21X1  g5476(.A0(new_n5861_), .A1(new_n1557_), .B0(new_n1558_), .Y(new_n5862_));
  OAI21X1  g5477(.A0(new_n5862_), .A1(new_n1556_), .B0(new_n1320_), .Y(new_n5863_));
  AOI21X1  g5478(.A0(new_n5863_), .A1(new_n1554_), .B0(new_n1555_), .Y(new_n5864_));
  OAI21X1  g5479(.A0(new_n5864_), .A1(new_n1553_), .B0(new_n1656_), .Y(new_n5865_));
  AOI21X1  g5480(.A0(new_n5865_), .A1(new_n1552_), .B0(new_n1893_), .Y(new_n5866_));
  OAI21X1  g5481(.A0(new_n5866_), .A1(new_n1395_), .B0(new_n403_), .Y(new_n5867_));
  AOI21X1  g5482(.A0(new_n5867_), .A1(new_n1393_), .B0(new_n1394_), .Y(new_n5868_));
  OAI21X1  g5483(.A0(new_n5868_), .A1(new_n1392_), .B0(new_n418_), .Y(new_n5869_));
  AOI21X1  g5484(.A0(new_n5869_), .A1(new_n1390_), .B0(new_n1391_), .Y(new_n5870_));
  OAI21X1  g5485(.A0(new_n5870_), .A1(new_n1389_), .B0(new_n433_), .Y(new_n5871_));
  AOI21X1  g5486(.A0(new_n5871_), .A1(new_n1387_), .B0(new_n1388_), .Y(new_n5872_));
  OAI21X1  g5487(.A0(new_n5872_), .A1(new_n1386_), .B0(new_n448_), .Y(new_n5873_));
  AOI21X1  g5488(.A0(new_n5873_), .A1(new_n1384_), .B0(new_n1385_), .Y(new_n5874_));
  OAI21X1  g5489(.A0(new_n5874_), .A1(new_n1383_), .B0(new_n463_), .Y(new_n5875_));
  AOI21X1  g5490(.A0(new_n5875_), .A1(new_n1381_), .B0(new_n1382_), .Y(new_n5876_));
  OAI21X1  g5491(.A0(new_n5876_), .A1(new_n1380_), .B0(new_n478_), .Y(new_n5877_));
  AOI21X1  g5492(.A0(new_n5877_), .A1(new_n1378_), .B0(new_n1379_), .Y(new_n5878_));
  OAI21X1  g5493(.A0(new_n5878_), .A1(new_n1377_), .B0(new_n493_), .Y(new_n5879_));
  AOI21X1  g5494(.A0(new_n5879_), .A1(new_n1375_), .B0(new_n1376_), .Y(new_n5880_));
  OAI21X1  g5495(.A0(new_n5880_), .A1(new_n1374_), .B0(new_n508_), .Y(new_n5881_));
  AOI21X1  g5496(.A0(new_n5881_), .A1(new_n1372_), .B0(new_n1373_), .Y(new_n5882_));
  OAI21X1  g5497(.A0(new_n5882_), .A1(new_n1371_), .B0(new_n523_), .Y(new_n5883_));
  AOI21X1  g5498(.A0(new_n5883_), .A1(new_n1369_), .B0(new_n1370_), .Y(new_n5884_));
  OAI21X1  g5499(.A0(new_n5884_), .A1(new_n1368_), .B0(new_n538_), .Y(new_n5885_));
  AOI21X1  g5500(.A0(new_n5885_), .A1(new_n1366_), .B0(new_n1367_), .Y(new_n5886_));
  OAI21X1  g5501(.A0(new_n5886_), .A1(new_n1365_), .B0(new_n553_), .Y(new_n5887_));
  AOI21X1  g5502(.A0(new_n5887_), .A1(new_n1363_), .B0(new_n1364_), .Y(new_n5888_));
  OAI21X1  g5503(.A0(new_n5888_), .A1(new_n1362_), .B0(new_n568_), .Y(new_n5889_));
  AOI21X1  g5504(.A0(new_n5889_), .A1(new_n1360_), .B0(new_n1361_), .Y(new_n5890_));
  OAI21X1  g5505(.A0(new_n5890_), .A1(new_n1359_), .B0(new_n583_), .Y(new_n5891_));
  AOI21X1  g5506(.A0(new_n5891_), .A1(new_n1357_), .B0(new_n1358_), .Y(new_n5892_));
  OAI21X1  g5507(.A0(new_n5892_), .A1(new_n1356_), .B0(new_n598_), .Y(new_n5893_));
  AOI21X1  g5508(.A0(new_n5893_), .A1(new_n1354_), .B0(new_n1355_), .Y(new_n5894_));
  OAI21X1  g5509(.A0(new_n5894_), .A1(new_n1353_), .B0(new_n613_), .Y(new_n5895_));
  AOI21X1  g5510(.A0(new_n5895_), .A1(new_n1351_), .B0(new_n1352_), .Y(new_n5896_));
  OAI21X1  g5511(.A0(new_n5896_), .A1(new_n1350_), .B0(new_n628_), .Y(new_n5897_));
  OAI21X1  g5512(.A0(new_n950_), .A1(\priority[101] ), .B0(\req[101] ), .Y(new_n5898_));
  AOI21X1  g5513(.A0(new_n5897_), .A1(new_n1348_), .B0(new_n5898_), .Y(\grant[101] ));
  NOR2X1   g5514(.A(new_n958_), .B(new_n642_), .Y(new_n5900_));
  OAI21X1  g5515(.A0(new_n5900_), .A1(new_n649_), .B0(new_n651_), .Y(new_n5901_));
  AOI21X1  g5516(.A0(new_n5901_), .A1(new_n656_), .B0(new_n659_), .Y(new_n5902_));
  OAI21X1  g5517(.A0(new_n5902_), .A1(new_n664_), .B0(new_n666_), .Y(new_n5903_));
  AOI21X1  g5518(.A0(new_n5903_), .A1(new_n671_), .B0(new_n674_), .Y(new_n5904_));
  OAI21X1  g5519(.A0(new_n5904_), .A1(new_n679_), .B0(new_n681_), .Y(new_n5905_));
  AOI21X1  g5520(.A0(new_n5905_), .A1(new_n686_), .B0(new_n689_), .Y(new_n5906_));
  OAI21X1  g5521(.A0(new_n5906_), .A1(new_n694_), .B0(new_n696_), .Y(new_n5907_));
  AOI21X1  g5522(.A0(new_n5907_), .A1(new_n701_), .B0(new_n1662_), .Y(new_n5908_));
  OAI21X1  g5523(.A0(new_n5908_), .A1(new_n1661_), .B0(new_n1705_), .Y(new_n5909_));
  AOI21X1  g5524(.A0(new_n5909_), .A1(new_n1660_), .B0(new_n1938_), .Y(new_n5910_));
  OAI21X1  g5525(.A0(new_n5910_), .A1(new_n1504_), .B0(new_n721_), .Y(new_n5911_));
  AOI21X1  g5526(.A0(new_n5911_), .A1(new_n1502_), .B0(new_n1503_), .Y(new_n5912_));
  OAI21X1  g5527(.A0(new_n5912_), .A1(new_n1501_), .B0(new_n736_), .Y(new_n5913_));
  AOI21X1  g5528(.A0(new_n5913_), .A1(new_n1499_), .B0(new_n1500_), .Y(new_n5914_));
  OAI21X1  g5529(.A0(new_n5914_), .A1(new_n1498_), .B0(new_n751_), .Y(new_n5915_));
  AOI21X1  g5530(.A0(new_n5915_), .A1(new_n1496_), .B0(new_n1497_), .Y(new_n5916_));
  OAI21X1  g5531(.A0(new_n5916_), .A1(new_n1495_), .B0(new_n766_), .Y(new_n5917_));
  AOI21X1  g5532(.A0(new_n5917_), .A1(new_n1493_), .B0(new_n1494_), .Y(new_n5918_));
  OAI21X1  g5533(.A0(new_n5918_), .A1(new_n1492_), .B0(new_n781_), .Y(new_n5919_));
  AOI21X1  g5534(.A0(new_n5919_), .A1(new_n1490_), .B0(new_n1491_), .Y(new_n5920_));
  OAI21X1  g5535(.A0(new_n5920_), .A1(new_n1489_), .B0(new_n796_), .Y(new_n5921_));
  AOI21X1  g5536(.A0(new_n5921_), .A1(new_n1487_), .B0(new_n1488_), .Y(new_n5922_));
  OAI21X1  g5537(.A0(new_n5922_), .A1(new_n1486_), .B0(new_n811_), .Y(new_n5923_));
  AOI21X1  g5538(.A0(new_n5923_), .A1(new_n1484_), .B0(new_n1485_), .Y(new_n5924_));
  OAI21X1  g5539(.A0(new_n5924_), .A1(new_n1483_), .B0(new_n826_), .Y(new_n5925_));
  AOI21X1  g5540(.A0(new_n5925_), .A1(new_n1481_), .B0(new_n1482_), .Y(new_n5926_));
  OAI21X1  g5541(.A0(new_n5926_), .A1(new_n1480_), .B0(new_n841_), .Y(new_n5927_));
  AOI21X1  g5542(.A0(new_n5927_), .A1(new_n1478_), .B0(new_n1479_), .Y(new_n5928_));
  OAI21X1  g5543(.A0(new_n5928_), .A1(new_n1477_), .B0(new_n856_), .Y(new_n5929_));
  AOI21X1  g5544(.A0(new_n5929_), .A1(new_n1475_), .B0(new_n1476_), .Y(new_n5930_));
  OAI21X1  g5545(.A0(new_n5930_), .A1(new_n1474_), .B0(new_n871_), .Y(new_n5931_));
  AOI21X1  g5546(.A0(new_n5931_), .A1(new_n1472_), .B0(new_n1473_), .Y(new_n5932_));
  OAI21X1  g5547(.A0(new_n5932_), .A1(new_n1471_), .B0(new_n886_), .Y(new_n5933_));
  AOI21X1  g5548(.A0(new_n5933_), .A1(new_n1469_), .B0(new_n1470_), .Y(new_n5934_));
  OAI21X1  g5549(.A0(new_n5934_), .A1(new_n1468_), .B0(new_n901_), .Y(new_n5935_));
  AOI21X1  g5550(.A0(new_n5935_), .A1(new_n1466_), .B0(new_n1467_), .Y(new_n5936_));
  OAI21X1  g5551(.A0(new_n5936_), .A1(new_n1465_), .B0(new_n916_), .Y(new_n5937_));
  AOI21X1  g5552(.A0(new_n5937_), .A1(new_n1463_), .B0(new_n1464_), .Y(new_n5938_));
  OAI21X1  g5553(.A0(new_n5938_), .A1(new_n1462_), .B0(new_n931_), .Y(new_n5939_));
  AOI21X1  g5554(.A0(new_n5939_), .A1(new_n1460_), .B0(new_n1461_), .Y(new_n5940_));
  OAI21X1  g5555(.A0(new_n5940_), .A1(new_n1459_), .B0(new_n946_), .Y(new_n5941_));
  OAI21X1  g5556(.A0(new_n1264_), .A1(\priority[102] ), .B0(\req[102] ), .Y(new_n5942_));
  AOI21X1  g5557(.A0(new_n5941_), .A1(new_n1457_), .B0(new_n5942_), .Y(\grant[102] ));
  NOR2X1   g5558(.A(new_n1272_), .B(new_n960_), .Y(new_n5944_));
  OAI21X1  g5559(.A0(new_n5944_), .A1(new_n967_), .B0(new_n969_), .Y(new_n5945_));
  AOI21X1  g5560(.A0(new_n5945_), .A1(new_n974_), .B0(new_n977_), .Y(new_n5946_));
  OAI21X1  g5561(.A0(new_n5946_), .A1(new_n982_), .B0(new_n984_), .Y(new_n5947_));
  AOI21X1  g5562(.A0(new_n5947_), .A1(new_n989_), .B0(new_n992_), .Y(new_n5948_));
  OAI21X1  g5563(.A0(new_n5948_), .A1(new_n997_), .B0(new_n999_), .Y(new_n5949_));
  AOI21X1  g5564(.A0(new_n5949_), .A1(new_n1004_), .B0(new_n1007_), .Y(new_n5950_));
  OAI21X1  g5565(.A0(new_n5950_), .A1(new_n1012_), .B0(new_n1014_), .Y(new_n5951_));
  AOI21X1  g5566(.A0(new_n5951_), .A1(new_n1017_), .B0(new_n1711_), .Y(new_n5952_));
  OAI21X1  g5567(.A0(new_n5952_), .A1(new_n1710_), .B0(new_n1754_), .Y(new_n5953_));
  AOI21X1  g5568(.A0(new_n5953_), .A1(new_n1709_), .B0(new_n1983_), .Y(new_n5954_));
  OAI21X1  g5569(.A0(new_n5954_), .A1(new_n1613_), .B0(new_n1035_), .Y(new_n5955_));
  AOI21X1  g5570(.A0(new_n5955_), .A1(new_n1611_), .B0(new_n1612_), .Y(new_n5956_));
  OAI21X1  g5571(.A0(new_n5956_), .A1(new_n1610_), .B0(new_n1050_), .Y(new_n5957_));
  AOI21X1  g5572(.A0(new_n5957_), .A1(new_n1608_), .B0(new_n1609_), .Y(new_n5958_));
  OAI21X1  g5573(.A0(new_n5958_), .A1(new_n1607_), .B0(new_n1065_), .Y(new_n5959_));
  AOI21X1  g5574(.A0(new_n5959_), .A1(new_n1605_), .B0(new_n1606_), .Y(new_n5960_));
  OAI21X1  g5575(.A0(new_n5960_), .A1(new_n1604_), .B0(new_n1080_), .Y(new_n5961_));
  AOI21X1  g5576(.A0(new_n5961_), .A1(new_n1602_), .B0(new_n1603_), .Y(new_n5962_));
  OAI21X1  g5577(.A0(new_n5962_), .A1(new_n1601_), .B0(new_n1095_), .Y(new_n5963_));
  AOI21X1  g5578(.A0(new_n5963_), .A1(new_n1599_), .B0(new_n1600_), .Y(new_n5964_));
  OAI21X1  g5579(.A0(new_n5964_), .A1(new_n1598_), .B0(new_n1110_), .Y(new_n5965_));
  AOI21X1  g5580(.A0(new_n5965_), .A1(new_n1596_), .B0(new_n1597_), .Y(new_n5966_));
  OAI21X1  g5581(.A0(new_n5966_), .A1(new_n1595_), .B0(new_n1125_), .Y(new_n5967_));
  AOI21X1  g5582(.A0(new_n5967_), .A1(new_n1593_), .B0(new_n1594_), .Y(new_n5968_));
  OAI21X1  g5583(.A0(new_n5968_), .A1(new_n1592_), .B0(new_n1140_), .Y(new_n5969_));
  AOI21X1  g5584(.A0(new_n5969_), .A1(new_n1590_), .B0(new_n1591_), .Y(new_n5970_));
  OAI21X1  g5585(.A0(new_n5970_), .A1(new_n1589_), .B0(new_n1155_), .Y(new_n5971_));
  AOI21X1  g5586(.A0(new_n5971_), .A1(new_n1587_), .B0(new_n1588_), .Y(new_n5972_));
  OAI21X1  g5587(.A0(new_n5972_), .A1(new_n1586_), .B0(new_n1170_), .Y(new_n5973_));
  AOI21X1  g5588(.A0(new_n5973_), .A1(new_n1584_), .B0(new_n1585_), .Y(new_n5974_));
  OAI21X1  g5589(.A0(new_n5974_), .A1(new_n1583_), .B0(new_n1185_), .Y(new_n5975_));
  AOI21X1  g5590(.A0(new_n5975_), .A1(new_n1581_), .B0(new_n1582_), .Y(new_n5976_));
  OAI21X1  g5591(.A0(new_n5976_), .A1(new_n1580_), .B0(new_n1200_), .Y(new_n5977_));
  AOI21X1  g5592(.A0(new_n5977_), .A1(new_n1578_), .B0(new_n1579_), .Y(new_n5978_));
  OAI21X1  g5593(.A0(new_n5978_), .A1(new_n1577_), .B0(new_n1215_), .Y(new_n5979_));
  AOI21X1  g5594(.A0(new_n5979_), .A1(new_n1575_), .B0(new_n1576_), .Y(new_n5980_));
  OAI21X1  g5595(.A0(new_n5980_), .A1(new_n1574_), .B0(new_n1230_), .Y(new_n5981_));
  AOI21X1  g5596(.A0(new_n5981_), .A1(new_n1572_), .B0(new_n1573_), .Y(new_n5982_));
  OAI21X1  g5597(.A0(new_n5982_), .A1(new_n1571_), .B0(new_n1245_), .Y(new_n5983_));
  AOI21X1  g5598(.A0(new_n5983_), .A1(new_n1569_), .B0(new_n1570_), .Y(new_n5984_));
  OAI21X1  g5599(.A0(new_n5984_), .A1(new_n1568_), .B0(new_n1260_), .Y(new_n5985_));
  OAI21X1  g5600(.A0(new_n639_), .A1(\priority[103] ), .B0(\req[103] ), .Y(new_n5986_));
  AOI21X1  g5601(.A0(new_n5985_), .A1(new_n1566_), .B0(new_n5986_), .Y(\grant[103] ));
  NOR2X1   g5602(.A(new_n1274_), .B(new_n648_), .Y(new_n5988_));
  OAI21X1  g5603(.A0(new_n5988_), .A1(new_n1281_), .B0(new_n1283_), .Y(new_n5989_));
  AOI21X1  g5604(.A0(new_n5989_), .A1(new_n1288_), .B0(new_n1291_), .Y(new_n5990_));
  OAI21X1  g5605(.A0(new_n5990_), .A1(new_n1296_), .B0(new_n1298_), .Y(new_n5991_));
  AOI21X1  g5606(.A0(new_n5991_), .A1(new_n1303_), .B0(new_n1306_), .Y(new_n5992_));
  OAI21X1  g5607(.A0(new_n5992_), .A1(new_n1311_), .B0(new_n1313_), .Y(new_n5993_));
  AOI21X1  g5608(.A0(new_n5993_), .A1(new_n1318_), .B0(new_n1321_), .Y(new_n5994_));
  OAI21X1  g5609(.A0(new_n5994_), .A1(new_n1326_), .B0(new_n1328_), .Y(new_n5995_));
  AOI21X1  g5610(.A0(new_n5995_), .A1(new_n1331_), .B0(new_n1758_), .Y(new_n5996_));
  OAI21X1  g5611(.A0(new_n5996_), .A1(new_n394_), .B0(new_n396_), .Y(new_n5997_));
  AOI21X1  g5612(.A0(new_n5997_), .A1(new_n401_), .B0(new_n404_), .Y(new_n5998_));
  OAI21X1  g5613(.A0(new_n5998_), .A1(new_n409_), .B0(new_n411_), .Y(new_n5999_));
  AOI21X1  g5614(.A0(new_n5999_), .A1(new_n416_), .B0(new_n419_), .Y(new_n6000_));
  OAI21X1  g5615(.A0(new_n6000_), .A1(new_n424_), .B0(new_n426_), .Y(new_n6001_));
  AOI21X1  g5616(.A0(new_n6001_), .A1(new_n431_), .B0(new_n434_), .Y(new_n6002_));
  OAI21X1  g5617(.A0(new_n6002_), .A1(new_n439_), .B0(new_n441_), .Y(new_n6003_));
  AOI21X1  g5618(.A0(new_n6003_), .A1(new_n446_), .B0(new_n449_), .Y(new_n6004_));
  OAI21X1  g5619(.A0(new_n6004_), .A1(new_n454_), .B0(new_n456_), .Y(new_n6005_));
  AOI21X1  g5620(.A0(new_n6005_), .A1(new_n461_), .B0(new_n464_), .Y(new_n6006_));
  OAI21X1  g5621(.A0(new_n6006_), .A1(new_n469_), .B0(new_n471_), .Y(new_n6007_));
  AOI21X1  g5622(.A0(new_n6007_), .A1(new_n476_), .B0(new_n479_), .Y(new_n6008_));
  OAI21X1  g5623(.A0(new_n6008_), .A1(new_n484_), .B0(new_n486_), .Y(new_n6009_));
  AOI21X1  g5624(.A0(new_n6009_), .A1(new_n491_), .B0(new_n494_), .Y(new_n6010_));
  OAI21X1  g5625(.A0(new_n6010_), .A1(new_n499_), .B0(new_n501_), .Y(new_n6011_));
  AOI21X1  g5626(.A0(new_n6011_), .A1(new_n506_), .B0(new_n509_), .Y(new_n6012_));
  OAI21X1  g5627(.A0(new_n6012_), .A1(new_n514_), .B0(new_n516_), .Y(new_n6013_));
  AOI21X1  g5628(.A0(new_n6013_), .A1(new_n521_), .B0(new_n524_), .Y(new_n6014_));
  OAI21X1  g5629(.A0(new_n6014_), .A1(new_n529_), .B0(new_n531_), .Y(new_n6015_));
  AOI21X1  g5630(.A0(new_n6015_), .A1(new_n536_), .B0(new_n539_), .Y(new_n6016_));
  OAI21X1  g5631(.A0(new_n6016_), .A1(new_n544_), .B0(new_n546_), .Y(new_n6017_));
  AOI21X1  g5632(.A0(new_n6017_), .A1(new_n551_), .B0(new_n554_), .Y(new_n6018_));
  OAI21X1  g5633(.A0(new_n6018_), .A1(new_n559_), .B0(new_n561_), .Y(new_n6019_));
  AOI21X1  g5634(.A0(new_n6019_), .A1(new_n566_), .B0(new_n569_), .Y(new_n6020_));
  OAI21X1  g5635(.A0(new_n6020_), .A1(new_n574_), .B0(new_n576_), .Y(new_n6021_));
  AOI21X1  g5636(.A0(new_n6021_), .A1(new_n581_), .B0(new_n584_), .Y(new_n6022_));
  OAI21X1  g5637(.A0(new_n6022_), .A1(new_n589_), .B0(new_n591_), .Y(new_n6023_));
  AOI21X1  g5638(.A0(new_n6023_), .A1(new_n596_), .B0(new_n599_), .Y(new_n6024_));
  OAI21X1  g5639(.A0(new_n6024_), .A1(new_n604_), .B0(new_n606_), .Y(new_n6025_));
  AOI21X1  g5640(.A0(new_n6025_), .A1(new_n611_), .B0(new_n614_), .Y(new_n6026_));
  OAI21X1  g5641(.A0(new_n6026_), .A1(new_n619_), .B0(new_n621_), .Y(new_n6027_));
  AOI21X1  g5642(.A0(new_n6027_), .A1(new_n626_), .B0(new_n629_), .Y(new_n6028_));
  OAI21X1  g5643(.A0(new_n6028_), .A1(new_n634_), .B0(new_n636_), .Y(new_n6029_));
  OAI21X1  g5644(.A0(new_n957_), .A1(\priority[104] ), .B0(\req[104] ), .Y(new_n6030_));
  AOI21X1  g5645(.A0(new_n6029_), .A1(new_n641_), .B0(new_n6030_), .Y(\grant[104] ));
  NOR2X1   g5646(.A(new_n966_), .B(new_n650_), .Y(new_n6032_));
  OAI21X1  g5647(.A0(new_n6032_), .A1(new_n1344_), .B0(new_n658_), .Y(new_n6033_));
  AOI21X1  g5648(.A0(new_n6033_), .A1(new_n1342_), .B0(new_n1343_), .Y(new_n6034_));
  OAI21X1  g5649(.A0(new_n6034_), .A1(new_n1341_), .B0(new_n673_), .Y(new_n6035_));
  AOI21X1  g5650(.A0(new_n6035_), .A1(new_n1339_), .B0(new_n1340_), .Y(new_n6036_));
  OAI21X1  g5651(.A0(new_n6036_), .A1(new_n1338_), .B0(new_n688_), .Y(new_n6037_));
  AOI21X1  g5652(.A0(new_n6037_), .A1(new_n1336_), .B0(new_n1337_), .Y(new_n6038_));
  OAI21X1  g5653(.A0(new_n6038_), .A1(new_n1335_), .B0(new_n1438_), .Y(new_n6039_));
  AOI21X1  g5654(.A0(new_n6039_), .A1(new_n1440_), .B0(new_n1803_), .Y(new_n6040_));
  OAI21X1  g5655(.A0(new_n6040_), .A1(new_n712_), .B0(new_n714_), .Y(new_n6041_));
  AOI21X1  g5656(.A0(new_n6041_), .A1(new_n719_), .B0(new_n722_), .Y(new_n6042_));
  OAI21X1  g5657(.A0(new_n6042_), .A1(new_n727_), .B0(new_n729_), .Y(new_n6043_));
  AOI21X1  g5658(.A0(new_n6043_), .A1(new_n734_), .B0(new_n737_), .Y(new_n6044_));
  OAI21X1  g5659(.A0(new_n6044_), .A1(new_n742_), .B0(new_n744_), .Y(new_n6045_));
  AOI21X1  g5660(.A0(new_n6045_), .A1(new_n749_), .B0(new_n752_), .Y(new_n6046_));
  OAI21X1  g5661(.A0(new_n6046_), .A1(new_n757_), .B0(new_n759_), .Y(new_n6047_));
  AOI21X1  g5662(.A0(new_n6047_), .A1(new_n764_), .B0(new_n767_), .Y(new_n6048_));
  OAI21X1  g5663(.A0(new_n6048_), .A1(new_n772_), .B0(new_n774_), .Y(new_n6049_));
  AOI21X1  g5664(.A0(new_n6049_), .A1(new_n779_), .B0(new_n782_), .Y(new_n6050_));
  OAI21X1  g5665(.A0(new_n6050_), .A1(new_n787_), .B0(new_n789_), .Y(new_n6051_));
  AOI21X1  g5666(.A0(new_n6051_), .A1(new_n794_), .B0(new_n797_), .Y(new_n6052_));
  OAI21X1  g5667(.A0(new_n6052_), .A1(new_n802_), .B0(new_n804_), .Y(new_n6053_));
  AOI21X1  g5668(.A0(new_n6053_), .A1(new_n809_), .B0(new_n812_), .Y(new_n6054_));
  OAI21X1  g5669(.A0(new_n6054_), .A1(new_n817_), .B0(new_n819_), .Y(new_n6055_));
  AOI21X1  g5670(.A0(new_n6055_), .A1(new_n824_), .B0(new_n827_), .Y(new_n6056_));
  OAI21X1  g5671(.A0(new_n6056_), .A1(new_n832_), .B0(new_n834_), .Y(new_n6057_));
  AOI21X1  g5672(.A0(new_n6057_), .A1(new_n839_), .B0(new_n842_), .Y(new_n6058_));
  OAI21X1  g5673(.A0(new_n6058_), .A1(new_n847_), .B0(new_n849_), .Y(new_n6059_));
  AOI21X1  g5674(.A0(new_n6059_), .A1(new_n854_), .B0(new_n857_), .Y(new_n6060_));
  OAI21X1  g5675(.A0(new_n6060_), .A1(new_n862_), .B0(new_n864_), .Y(new_n6061_));
  AOI21X1  g5676(.A0(new_n6061_), .A1(new_n869_), .B0(new_n872_), .Y(new_n6062_));
  OAI21X1  g5677(.A0(new_n6062_), .A1(new_n877_), .B0(new_n879_), .Y(new_n6063_));
  AOI21X1  g5678(.A0(new_n6063_), .A1(new_n884_), .B0(new_n887_), .Y(new_n6064_));
  OAI21X1  g5679(.A0(new_n6064_), .A1(new_n892_), .B0(new_n894_), .Y(new_n6065_));
  AOI21X1  g5680(.A0(new_n6065_), .A1(new_n899_), .B0(new_n902_), .Y(new_n6066_));
  OAI21X1  g5681(.A0(new_n6066_), .A1(new_n907_), .B0(new_n909_), .Y(new_n6067_));
  AOI21X1  g5682(.A0(new_n6067_), .A1(new_n914_), .B0(new_n917_), .Y(new_n6068_));
  OAI21X1  g5683(.A0(new_n6068_), .A1(new_n922_), .B0(new_n924_), .Y(new_n6069_));
  AOI21X1  g5684(.A0(new_n6069_), .A1(new_n929_), .B0(new_n932_), .Y(new_n6070_));
  OAI21X1  g5685(.A0(new_n6070_), .A1(new_n937_), .B0(new_n939_), .Y(new_n6071_));
  AOI21X1  g5686(.A0(new_n6071_), .A1(new_n944_), .B0(new_n947_), .Y(new_n6072_));
  OAI21X1  g5687(.A0(new_n6072_), .A1(new_n952_), .B0(new_n954_), .Y(new_n6073_));
  OAI21X1  g5688(.A0(new_n1271_), .A1(\priority[105] ), .B0(\req[105] ), .Y(new_n6074_));
  AOI21X1  g5689(.A0(new_n6073_), .A1(new_n959_), .B0(new_n6074_), .Y(\grant[105] ));
  NOR2X1   g5690(.A(new_n1280_), .B(new_n968_), .Y(new_n6076_));
  OAI21X1  g5691(.A0(new_n6076_), .A1(new_n1453_), .B0(new_n976_), .Y(new_n6077_));
  AOI21X1  g5692(.A0(new_n6077_), .A1(new_n1451_), .B0(new_n1452_), .Y(new_n6078_));
  OAI21X1  g5693(.A0(new_n6078_), .A1(new_n1450_), .B0(new_n991_), .Y(new_n6079_));
  AOI21X1  g5694(.A0(new_n6079_), .A1(new_n1448_), .B0(new_n1449_), .Y(new_n6080_));
  OAI21X1  g5695(.A0(new_n6080_), .A1(new_n1447_), .B0(new_n1006_), .Y(new_n6081_));
  AOI21X1  g5696(.A0(new_n6081_), .A1(new_n1445_), .B0(new_n1446_), .Y(new_n6082_));
  OAI21X1  g5697(.A0(new_n6082_), .A1(new_n1444_), .B0(new_n1547_), .Y(new_n6083_));
  AOI21X1  g5698(.A0(new_n6083_), .A1(new_n1549_), .B0(new_n1848_), .Y(new_n6084_));
  OAI21X1  g5699(.A0(new_n6084_), .A1(new_n1026_), .B0(new_n1028_), .Y(new_n6085_));
  AOI21X1  g5700(.A0(new_n6085_), .A1(new_n1033_), .B0(new_n1036_), .Y(new_n6086_));
  OAI21X1  g5701(.A0(new_n6086_), .A1(new_n1041_), .B0(new_n1043_), .Y(new_n6087_));
  AOI21X1  g5702(.A0(new_n6087_), .A1(new_n1048_), .B0(new_n1051_), .Y(new_n6088_));
  OAI21X1  g5703(.A0(new_n6088_), .A1(new_n1056_), .B0(new_n1058_), .Y(new_n6089_));
  AOI21X1  g5704(.A0(new_n6089_), .A1(new_n1063_), .B0(new_n1066_), .Y(new_n6090_));
  OAI21X1  g5705(.A0(new_n6090_), .A1(new_n1071_), .B0(new_n1073_), .Y(new_n6091_));
  AOI21X1  g5706(.A0(new_n6091_), .A1(new_n1078_), .B0(new_n1081_), .Y(new_n6092_));
  OAI21X1  g5707(.A0(new_n6092_), .A1(new_n1086_), .B0(new_n1088_), .Y(new_n6093_));
  AOI21X1  g5708(.A0(new_n6093_), .A1(new_n1093_), .B0(new_n1096_), .Y(new_n6094_));
  OAI21X1  g5709(.A0(new_n6094_), .A1(new_n1101_), .B0(new_n1103_), .Y(new_n6095_));
  AOI21X1  g5710(.A0(new_n6095_), .A1(new_n1108_), .B0(new_n1111_), .Y(new_n6096_));
  OAI21X1  g5711(.A0(new_n6096_), .A1(new_n1116_), .B0(new_n1118_), .Y(new_n6097_));
  AOI21X1  g5712(.A0(new_n6097_), .A1(new_n1123_), .B0(new_n1126_), .Y(new_n6098_));
  OAI21X1  g5713(.A0(new_n6098_), .A1(new_n1131_), .B0(new_n1133_), .Y(new_n6099_));
  AOI21X1  g5714(.A0(new_n6099_), .A1(new_n1138_), .B0(new_n1141_), .Y(new_n6100_));
  OAI21X1  g5715(.A0(new_n6100_), .A1(new_n1146_), .B0(new_n1148_), .Y(new_n6101_));
  AOI21X1  g5716(.A0(new_n6101_), .A1(new_n1153_), .B0(new_n1156_), .Y(new_n6102_));
  OAI21X1  g5717(.A0(new_n6102_), .A1(new_n1161_), .B0(new_n1163_), .Y(new_n6103_));
  AOI21X1  g5718(.A0(new_n6103_), .A1(new_n1168_), .B0(new_n1171_), .Y(new_n6104_));
  OAI21X1  g5719(.A0(new_n6104_), .A1(new_n1176_), .B0(new_n1178_), .Y(new_n6105_));
  AOI21X1  g5720(.A0(new_n6105_), .A1(new_n1183_), .B0(new_n1186_), .Y(new_n6106_));
  OAI21X1  g5721(.A0(new_n6106_), .A1(new_n1191_), .B0(new_n1193_), .Y(new_n6107_));
  AOI21X1  g5722(.A0(new_n6107_), .A1(new_n1198_), .B0(new_n1201_), .Y(new_n6108_));
  OAI21X1  g5723(.A0(new_n6108_), .A1(new_n1206_), .B0(new_n1208_), .Y(new_n6109_));
  AOI21X1  g5724(.A0(new_n6109_), .A1(new_n1213_), .B0(new_n1216_), .Y(new_n6110_));
  OAI21X1  g5725(.A0(new_n6110_), .A1(new_n1221_), .B0(new_n1223_), .Y(new_n6111_));
  AOI21X1  g5726(.A0(new_n6111_), .A1(new_n1228_), .B0(new_n1231_), .Y(new_n6112_));
  OAI21X1  g5727(.A0(new_n6112_), .A1(new_n1236_), .B0(new_n1238_), .Y(new_n6113_));
  AOI21X1  g5728(.A0(new_n6113_), .A1(new_n1243_), .B0(new_n1246_), .Y(new_n6114_));
  OAI21X1  g5729(.A0(new_n6114_), .A1(new_n1251_), .B0(new_n1253_), .Y(new_n6115_));
  AOI21X1  g5730(.A0(new_n6115_), .A1(new_n1258_), .B0(new_n1261_), .Y(new_n6116_));
  OAI21X1  g5731(.A0(new_n6116_), .A1(new_n1266_), .B0(new_n1268_), .Y(new_n6117_));
  OAI21X1  g5732(.A0(new_n647_), .A1(\priority[106] ), .B0(\req[106] ), .Y(new_n6118_));
  AOI21X1  g5733(.A0(new_n6117_), .A1(new_n1273_), .B0(new_n6118_), .Y(\grant[106] ));
  NOR2X1   g5734(.A(new_n1282_), .B(new_n655_), .Y(new_n6120_));
  OAI21X1  g5735(.A0(new_n6120_), .A1(new_n1562_), .B0(new_n1290_), .Y(new_n6121_));
  AOI21X1  g5736(.A0(new_n6121_), .A1(new_n1560_), .B0(new_n1561_), .Y(new_n6122_));
  OAI21X1  g5737(.A0(new_n6122_), .A1(new_n1559_), .B0(new_n1305_), .Y(new_n6123_));
  AOI21X1  g5738(.A0(new_n6123_), .A1(new_n1557_), .B0(new_n1558_), .Y(new_n6124_));
  OAI21X1  g5739(.A0(new_n6124_), .A1(new_n1556_), .B0(new_n1320_), .Y(new_n6125_));
  AOI21X1  g5740(.A0(new_n6125_), .A1(new_n1554_), .B0(new_n1555_), .Y(new_n6126_));
  OAI21X1  g5741(.A0(new_n6126_), .A1(new_n1553_), .B0(new_n1656_), .Y(new_n6127_));
  AOI21X1  g5742(.A0(new_n6127_), .A1(new_n1552_), .B0(new_n1893_), .Y(new_n6128_));
  OAI21X1  g5743(.A0(new_n6128_), .A1(new_n1395_), .B0(new_n403_), .Y(new_n6129_));
  AOI21X1  g5744(.A0(new_n6129_), .A1(new_n1393_), .B0(new_n1394_), .Y(new_n6130_));
  OAI21X1  g5745(.A0(new_n6130_), .A1(new_n1392_), .B0(new_n418_), .Y(new_n6131_));
  AOI21X1  g5746(.A0(new_n6131_), .A1(new_n1390_), .B0(new_n1391_), .Y(new_n6132_));
  OAI21X1  g5747(.A0(new_n6132_), .A1(new_n1389_), .B0(new_n433_), .Y(new_n6133_));
  AOI21X1  g5748(.A0(new_n6133_), .A1(new_n1387_), .B0(new_n1388_), .Y(new_n6134_));
  OAI21X1  g5749(.A0(new_n6134_), .A1(new_n1386_), .B0(new_n448_), .Y(new_n6135_));
  AOI21X1  g5750(.A0(new_n6135_), .A1(new_n1384_), .B0(new_n1385_), .Y(new_n6136_));
  OAI21X1  g5751(.A0(new_n6136_), .A1(new_n1383_), .B0(new_n463_), .Y(new_n6137_));
  AOI21X1  g5752(.A0(new_n6137_), .A1(new_n1381_), .B0(new_n1382_), .Y(new_n6138_));
  OAI21X1  g5753(.A0(new_n6138_), .A1(new_n1380_), .B0(new_n478_), .Y(new_n6139_));
  AOI21X1  g5754(.A0(new_n6139_), .A1(new_n1378_), .B0(new_n1379_), .Y(new_n6140_));
  OAI21X1  g5755(.A0(new_n6140_), .A1(new_n1377_), .B0(new_n493_), .Y(new_n6141_));
  AOI21X1  g5756(.A0(new_n6141_), .A1(new_n1375_), .B0(new_n1376_), .Y(new_n6142_));
  OAI21X1  g5757(.A0(new_n6142_), .A1(new_n1374_), .B0(new_n508_), .Y(new_n6143_));
  AOI21X1  g5758(.A0(new_n6143_), .A1(new_n1372_), .B0(new_n1373_), .Y(new_n6144_));
  OAI21X1  g5759(.A0(new_n6144_), .A1(new_n1371_), .B0(new_n523_), .Y(new_n6145_));
  AOI21X1  g5760(.A0(new_n6145_), .A1(new_n1369_), .B0(new_n1370_), .Y(new_n6146_));
  OAI21X1  g5761(.A0(new_n6146_), .A1(new_n1368_), .B0(new_n538_), .Y(new_n6147_));
  AOI21X1  g5762(.A0(new_n6147_), .A1(new_n1366_), .B0(new_n1367_), .Y(new_n6148_));
  OAI21X1  g5763(.A0(new_n6148_), .A1(new_n1365_), .B0(new_n553_), .Y(new_n6149_));
  AOI21X1  g5764(.A0(new_n6149_), .A1(new_n1363_), .B0(new_n1364_), .Y(new_n6150_));
  OAI21X1  g5765(.A0(new_n6150_), .A1(new_n1362_), .B0(new_n568_), .Y(new_n6151_));
  AOI21X1  g5766(.A0(new_n6151_), .A1(new_n1360_), .B0(new_n1361_), .Y(new_n6152_));
  OAI21X1  g5767(.A0(new_n6152_), .A1(new_n1359_), .B0(new_n583_), .Y(new_n6153_));
  AOI21X1  g5768(.A0(new_n6153_), .A1(new_n1357_), .B0(new_n1358_), .Y(new_n6154_));
  OAI21X1  g5769(.A0(new_n6154_), .A1(new_n1356_), .B0(new_n598_), .Y(new_n6155_));
  AOI21X1  g5770(.A0(new_n6155_), .A1(new_n1354_), .B0(new_n1355_), .Y(new_n6156_));
  OAI21X1  g5771(.A0(new_n6156_), .A1(new_n1353_), .B0(new_n613_), .Y(new_n6157_));
  AOI21X1  g5772(.A0(new_n6157_), .A1(new_n1351_), .B0(new_n1352_), .Y(new_n6158_));
  OAI21X1  g5773(.A0(new_n6158_), .A1(new_n1350_), .B0(new_n628_), .Y(new_n6159_));
  AOI21X1  g5774(.A0(new_n6159_), .A1(new_n1348_), .B0(new_n1349_), .Y(new_n6160_));
  OAI21X1  g5775(.A0(new_n6160_), .A1(new_n1347_), .B0(new_n643_), .Y(new_n6161_));
  OAI21X1  g5776(.A0(new_n965_), .A1(\priority[107] ), .B0(\req[107] ), .Y(new_n6162_));
  AOI21X1  g5777(.A0(new_n6161_), .A1(new_n1345_), .B0(new_n6162_), .Y(\grant[107] ));
  NOR2X1   g5778(.A(new_n973_), .B(new_n657_), .Y(new_n6164_));
  OAI21X1  g5779(.A0(new_n6164_), .A1(new_n664_), .B0(new_n666_), .Y(new_n6165_));
  AOI21X1  g5780(.A0(new_n6165_), .A1(new_n671_), .B0(new_n674_), .Y(new_n6166_));
  OAI21X1  g5781(.A0(new_n6166_), .A1(new_n679_), .B0(new_n681_), .Y(new_n6167_));
  AOI21X1  g5782(.A0(new_n6167_), .A1(new_n686_), .B0(new_n689_), .Y(new_n6168_));
  OAI21X1  g5783(.A0(new_n6168_), .A1(new_n694_), .B0(new_n696_), .Y(new_n6169_));
  AOI21X1  g5784(.A0(new_n6169_), .A1(new_n701_), .B0(new_n1662_), .Y(new_n6170_));
  OAI21X1  g5785(.A0(new_n6170_), .A1(new_n1661_), .B0(new_n1705_), .Y(new_n6171_));
  AOI21X1  g5786(.A0(new_n6171_), .A1(new_n1660_), .B0(new_n1938_), .Y(new_n6172_));
  OAI21X1  g5787(.A0(new_n6172_), .A1(new_n1504_), .B0(new_n721_), .Y(new_n6173_));
  AOI21X1  g5788(.A0(new_n6173_), .A1(new_n1502_), .B0(new_n1503_), .Y(new_n6174_));
  OAI21X1  g5789(.A0(new_n6174_), .A1(new_n1501_), .B0(new_n736_), .Y(new_n6175_));
  AOI21X1  g5790(.A0(new_n6175_), .A1(new_n1499_), .B0(new_n1500_), .Y(new_n6176_));
  OAI21X1  g5791(.A0(new_n6176_), .A1(new_n1498_), .B0(new_n751_), .Y(new_n6177_));
  AOI21X1  g5792(.A0(new_n6177_), .A1(new_n1496_), .B0(new_n1497_), .Y(new_n6178_));
  OAI21X1  g5793(.A0(new_n6178_), .A1(new_n1495_), .B0(new_n766_), .Y(new_n6179_));
  AOI21X1  g5794(.A0(new_n6179_), .A1(new_n1493_), .B0(new_n1494_), .Y(new_n6180_));
  OAI21X1  g5795(.A0(new_n6180_), .A1(new_n1492_), .B0(new_n781_), .Y(new_n6181_));
  AOI21X1  g5796(.A0(new_n6181_), .A1(new_n1490_), .B0(new_n1491_), .Y(new_n6182_));
  OAI21X1  g5797(.A0(new_n6182_), .A1(new_n1489_), .B0(new_n796_), .Y(new_n6183_));
  AOI21X1  g5798(.A0(new_n6183_), .A1(new_n1487_), .B0(new_n1488_), .Y(new_n6184_));
  OAI21X1  g5799(.A0(new_n6184_), .A1(new_n1486_), .B0(new_n811_), .Y(new_n6185_));
  AOI21X1  g5800(.A0(new_n6185_), .A1(new_n1484_), .B0(new_n1485_), .Y(new_n6186_));
  OAI21X1  g5801(.A0(new_n6186_), .A1(new_n1483_), .B0(new_n826_), .Y(new_n6187_));
  AOI21X1  g5802(.A0(new_n6187_), .A1(new_n1481_), .B0(new_n1482_), .Y(new_n6188_));
  OAI21X1  g5803(.A0(new_n6188_), .A1(new_n1480_), .B0(new_n841_), .Y(new_n6189_));
  AOI21X1  g5804(.A0(new_n6189_), .A1(new_n1478_), .B0(new_n1479_), .Y(new_n6190_));
  OAI21X1  g5805(.A0(new_n6190_), .A1(new_n1477_), .B0(new_n856_), .Y(new_n6191_));
  AOI21X1  g5806(.A0(new_n6191_), .A1(new_n1475_), .B0(new_n1476_), .Y(new_n6192_));
  OAI21X1  g5807(.A0(new_n6192_), .A1(new_n1474_), .B0(new_n871_), .Y(new_n6193_));
  AOI21X1  g5808(.A0(new_n6193_), .A1(new_n1472_), .B0(new_n1473_), .Y(new_n6194_));
  OAI21X1  g5809(.A0(new_n6194_), .A1(new_n1471_), .B0(new_n886_), .Y(new_n6195_));
  AOI21X1  g5810(.A0(new_n6195_), .A1(new_n1469_), .B0(new_n1470_), .Y(new_n6196_));
  OAI21X1  g5811(.A0(new_n6196_), .A1(new_n1468_), .B0(new_n901_), .Y(new_n6197_));
  AOI21X1  g5812(.A0(new_n6197_), .A1(new_n1466_), .B0(new_n1467_), .Y(new_n6198_));
  OAI21X1  g5813(.A0(new_n6198_), .A1(new_n1465_), .B0(new_n916_), .Y(new_n6199_));
  AOI21X1  g5814(.A0(new_n6199_), .A1(new_n1463_), .B0(new_n1464_), .Y(new_n6200_));
  OAI21X1  g5815(.A0(new_n6200_), .A1(new_n1462_), .B0(new_n931_), .Y(new_n6201_));
  AOI21X1  g5816(.A0(new_n6201_), .A1(new_n1460_), .B0(new_n1461_), .Y(new_n6202_));
  OAI21X1  g5817(.A0(new_n6202_), .A1(new_n1459_), .B0(new_n946_), .Y(new_n6203_));
  AOI21X1  g5818(.A0(new_n6203_), .A1(new_n1457_), .B0(new_n1458_), .Y(new_n6204_));
  OAI21X1  g5819(.A0(new_n6204_), .A1(new_n1456_), .B0(new_n961_), .Y(new_n6205_));
  OAI21X1  g5820(.A0(new_n1279_), .A1(\priority[108] ), .B0(\req[108] ), .Y(new_n6206_));
  AOI21X1  g5821(.A0(new_n6205_), .A1(new_n1454_), .B0(new_n6206_), .Y(\grant[108] ));
  NOR2X1   g5822(.A(new_n1287_), .B(new_n975_), .Y(new_n6208_));
  OAI21X1  g5823(.A0(new_n6208_), .A1(new_n982_), .B0(new_n984_), .Y(new_n6209_));
  AOI21X1  g5824(.A0(new_n6209_), .A1(new_n989_), .B0(new_n992_), .Y(new_n6210_));
  OAI21X1  g5825(.A0(new_n6210_), .A1(new_n997_), .B0(new_n999_), .Y(new_n6211_));
  AOI21X1  g5826(.A0(new_n6211_), .A1(new_n1004_), .B0(new_n1007_), .Y(new_n6212_));
  OAI21X1  g5827(.A0(new_n6212_), .A1(new_n1012_), .B0(new_n1014_), .Y(new_n6213_));
  AOI21X1  g5828(.A0(new_n6213_), .A1(new_n1017_), .B0(new_n1711_), .Y(new_n6214_));
  OAI21X1  g5829(.A0(new_n6214_), .A1(new_n1710_), .B0(new_n1754_), .Y(new_n6215_));
  AOI21X1  g5830(.A0(new_n6215_), .A1(new_n1709_), .B0(new_n1983_), .Y(new_n6216_));
  OAI21X1  g5831(.A0(new_n6216_), .A1(new_n1613_), .B0(new_n1035_), .Y(new_n6217_));
  AOI21X1  g5832(.A0(new_n6217_), .A1(new_n1611_), .B0(new_n1612_), .Y(new_n6218_));
  OAI21X1  g5833(.A0(new_n6218_), .A1(new_n1610_), .B0(new_n1050_), .Y(new_n6219_));
  AOI21X1  g5834(.A0(new_n6219_), .A1(new_n1608_), .B0(new_n1609_), .Y(new_n6220_));
  OAI21X1  g5835(.A0(new_n6220_), .A1(new_n1607_), .B0(new_n1065_), .Y(new_n6221_));
  AOI21X1  g5836(.A0(new_n6221_), .A1(new_n1605_), .B0(new_n1606_), .Y(new_n6222_));
  OAI21X1  g5837(.A0(new_n6222_), .A1(new_n1604_), .B0(new_n1080_), .Y(new_n6223_));
  AOI21X1  g5838(.A0(new_n6223_), .A1(new_n1602_), .B0(new_n1603_), .Y(new_n6224_));
  OAI21X1  g5839(.A0(new_n6224_), .A1(new_n1601_), .B0(new_n1095_), .Y(new_n6225_));
  AOI21X1  g5840(.A0(new_n6225_), .A1(new_n1599_), .B0(new_n1600_), .Y(new_n6226_));
  OAI21X1  g5841(.A0(new_n6226_), .A1(new_n1598_), .B0(new_n1110_), .Y(new_n6227_));
  AOI21X1  g5842(.A0(new_n6227_), .A1(new_n1596_), .B0(new_n1597_), .Y(new_n6228_));
  OAI21X1  g5843(.A0(new_n6228_), .A1(new_n1595_), .B0(new_n1125_), .Y(new_n6229_));
  AOI21X1  g5844(.A0(new_n6229_), .A1(new_n1593_), .B0(new_n1594_), .Y(new_n6230_));
  OAI21X1  g5845(.A0(new_n6230_), .A1(new_n1592_), .B0(new_n1140_), .Y(new_n6231_));
  AOI21X1  g5846(.A0(new_n6231_), .A1(new_n1590_), .B0(new_n1591_), .Y(new_n6232_));
  OAI21X1  g5847(.A0(new_n6232_), .A1(new_n1589_), .B0(new_n1155_), .Y(new_n6233_));
  AOI21X1  g5848(.A0(new_n6233_), .A1(new_n1587_), .B0(new_n1588_), .Y(new_n6234_));
  OAI21X1  g5849(.A0(new_n6234_), .A1(new_n1586_), .B0(new_n1170_), .Y(new_n6235_));
  AOI21X1  g5850(.A0(new_n6235_), .A1(new_n1584_), .B0(new_n1585_), .Y(new_n6236_));
  OAI21X1  g5851(.A0(new_n6236_), .A1(new_n1583_), .B0(new_n1185_), .Y(new_n6237_));
  AOI21X1  g5852(.A0(new_n6237_), .A1(new_n1581_), .B0(new_n1582_), .Y(new_n6238_));
  OAI21X1  g5853(.A0(new_n6238_), .A1(new_n1580_), .B0(new_n1200_), .Y(new_n6239_));
  AOI21X1  g5854(.A0(new_n6239_), .A1(new_n1578_), .B0(new_n1579_), .Y(new_n6240_));
  OAI21X1  g5855(.A0(new_n6240_), .A1(new_n1577_), .B0(new_n1215_), .Y(new_n6241_));
  AOI21X1  g5856(.A0(new_n6241_), .A1(new_n1575_), .B0(new_n1576_), .Y(new_n6242_));
  OAI21X1  g5857(.A0(new_n6242_), .A1(new_n1574_), .B0(new_n1230_), .Y(new_n6243_));
  AOI21X1  g5858(.A0(new_n6243_), .A1(new_n1572_), .B0(new_n1573_), .Y(new_n6244_));
  OAI21X1  g5859(.A0(new_n6244_), .A1(new_n1571_), .B0(new_n1245_), .Y(new_n6245_));
  AOI21X1  g5860(.A0(new_n6245_), .A1(new_n1569_), .B0(new_n1570_), .Y(new_n6246_));
  OAI21X1  g5861(.A0(new_n6246_), .A1(new_n1568_), .B0(new_n1260_), .Y(new_n6247_));
  AOI21X1  g5862(.A0(new_n6247_), .A1(new_n1566_), .B0(new_n1567_), .Y(new_n6248_));
  OAI21X1  g5863(.A0(new_n6248_), .A1(new_n1565_), .B0(new_n1275_), .Y(new_n6249_));
  OAI21X1  g5864(.A0(new_n654_), .A1(\priority[109] ), .B0(\req[109] ), .Y(new_n6250_));
  AOI21X1  g5865(.A0(new_n6249_), .A1(new_n1563_), .B0(new_n6250_), .Y(\grant[109] ));
  NOR2X1   g5866(.A(new_n1289_), .B(new_n663_), .Y(new_n6252_));
  OAI21X1  g5867(.A0(new_n6252_), .A1(new_n1296_), .B0(new_n1298_), .Y(new_n6253_));
  AOI21X1  g5868(.A0(new_n6253_), .A1(new_n1303_), .B0(new_n1306_), .Y(new_n6254_));
  OAI21X1  g5869(.A0(new_n6254_), .A1(new_n1311_), .B0(new_n1313_), .Y(new_n6255_));
  AOI21X1  g5870(.A0(new_n6255_), .A1(new_n1318_), .B0(new_n1321_), .Y(new_n6256_));
  OAI21X1  g5871(.A0(new_n6256_), .A1(new_n1326_), .B0(new_n1328_), .Y(new_n6257_));
  AOI21X1  g5872(.A0(new_n6257_), .A1(new_n1331_), .B0(new_n1758_), .Y(new_n6258_));
  OAI21X1  g5873(.A0(new_n6258_), .A1(new_n394_), .B0(new_n396_), .Y(new_n6259_));
  AOI21X1  g5874(.A0(new_n6259_), .A1(new_n401_), .B0(new_n404_), .Y(new_n6260_));
  OAI21X1  g5875(.A0(new_n6260_), .A1(new_n409_), .B0(new_n411_), .Y(new_n6261_));
  AOI21X1  g5876(.A0(new_n6261_), .A1(new_n416_), .B0(new_n419_), .Y(new_n6262_));
  OAI21X1  g5877(.A0(new_n6262_), .A1(new_n424_), .B0(new_n426_), .Y(new_n6263_));
  AOI21X1  g5878(.A0(new_n6263_), .A1(new_n431_), .B0(new_n434_), .Y(new_n6264_));
  OAI21X1  g5879(.A0(new_n6264_), .A1(new_n439_), .B0(new_n441_), .Y(new_n6265_));
  AOI21X1  g5880(.A0(new_n6265_), .A1(new_n446_), .B0(new_n449_), .Y(new_n6266_));
  OAI21X1  g5881(.A0(new_n6266_), .A1(new_n454_), .B0(new_n456_), .Y(new_n6267_));
  AOI21X1  g5882(.A0(new_n6267_), .A1(new_n461_), .B0(new_n464_), .Y(new_n6268_));
  OAI21X1  g5883(.A0(new_n6268_), .A1(new_n469_), .B0(new_n471_), .Y(new_n6269_));
  AOI21X1  g5884(.A0(new_n6269_), .A1(new_n476_), .B0(new_n479_), .Y(new_n6270_));
  OAI21X1  g5885(.A0(new_n6270_), .A1(new_n484_), .B0(new_n486_), .Y(new_n6271_));
  AOI21X1  g5886(.A0(new_n6271_), .A1(new_n491_), .B0(new_n494_), .Y(new_n6272_));
  OAI21X1  g5887(.A0(new_n6272_), .A1(new_n499_), .B0(new_n501_), .Y(new_n6273_));
  AOI21X1  g5888(.A0(new_n6273_), .A1(new_n506_), .B0(new_n509_), .Y(new_n6274_));
  OAI21X1  g5889(.A0(new_n6274_), .A1(new_n514_), .B0(new_n516_), .Y(new_n6275_));
  AOI21X1  g5890(.A0(new_n6275_), .A1(new_n521_), .B0(new_n524_), .Y(new_n6276_));
  OAI21X1  g5891(.A0(new_n6276_), .A1(new_n529_), .B0(new_n531_), .Y(new_n6277_));
  AOI21X1  g5892(.A0(new_n6277_), .A1(new_n536_), .B0(new_n539_), .Y(new_n6278_));
  OAI21X1  g5893(.A0(new_n6278_), .A1(new_n544_), .B0(new_n546_), .Y(new_n6279_));
  AOI21X1  g5894(.A0(new_n6279_), .A1(new_n551_), .B0(new_n554_), .Y(new_n6280_));
  OAI21X1  g5895(.A0(new_n6280_), .A1(new_n559_), .B0(new_n561_), .Y(new_n6281_));
  AOI21X1  g5896(.A0(new_n6281_), .A1(new_n566_), .B0(new_n569_), .Y(new_n6282_));
  OAI21X1  g5897(.A0(new_n6282_), .A1(new_n574_), .B0(new_n576_), .Y(new_n6283_));
  AOI21X1  g5898(.A0(new_n6283_), .A1(new_n581_), .B0(new_n584_), .Y(new_n6284_));
  OAI21X1  g5899(.A0(new_n6284_), .A1(new_n589_), .B0(new_n591_), .Y(new_n6285_));
  AOI21X1  g5900(.A0(new_n6285_), .A1(new_n596_), .B0(new_n599_), .Y(new_n6286_));
  OAI21X1  g5901(.A0(new_n6286_), .A1(new_n604_), .B0(new_n606_), .Y(new_n6287_));
  AOI21X1  g5902(.A0(new_n6287_), .A1(new_n611_), .B0(new_n614_), .Y(new_n6288_));
  OAI21X1  g5903(.A0(new_n6288_), .A1(new_n619_), .B0(new_n621_), .Y(new_n6289_));
  AOI21X1  g5904(.A0(new_n6289_), .A1(new_n626_), .B0(new_n629_), .Y(new_n6290_));
  OAI21X1  g5905(.A0(new_n6290_), .A1(new_n634_), .B0(new_n636_), .Y(new_n6291_));
  AOI21X1  g5906(.A0(new_n6291_), .A1(new_n641_), .B0(new_n644_), .Y(new_n6292_));
  OAI21X1  g5907(.A0(new_n6292_), .A1(new_n649_), .B0(new_n651_), .Y(new_n6293_));
  OAI21X1  g5908(.A0(new_n972_), .A1(\priority[110] ), .B0(\req[110] ), .Y(new_n6294_));
  AOI21X1  g5909(.A0(new_n6293_), .A1(new_n656_), .B0(new_n6294_), .Y(\grant[110] ));
  NOR2X1   g5910(.A(new_n981_), .B(new_n665_), .Y(new_n6296_));
  OAI21X1  g5911(.A0(new_n6296_), .A1(new_n1341_), .B0(new_n673_), .Y(new_n6297_));
  AOI21X1  g5912(.A0(new_n6297_), .A1(new_n1339_), .B0(new_n1340_), .Y(new_n6298_));
  OAI21X1  g5913(.A0(new_n6298_), .A1(new_n1338_), .B0(new_n688_), .Y(new_n6299_));
  AOI21X1  g5914(.A0(new_n6299_), .A1(new_n1336_), .B0(new_n1337_), .Y(new_n6300_));
  OAI21X1  g5915(.A0(new_n6300_), .A1(new_n1335_), .B0(new_n1438_), .Y(new_n6301_));
  AOI21X1  g5916(.A0(new_n6301_), .A1(new_n1440_), .B0(new_n1803_), .Y(new_n6302_));
  OAI21X1  g5917(.A0(new_n6302_), .A1(new_n712_), .B0(new_n714_), .Y(new_n6303_));
  AOI21X1  g5918(.A0(new_n6303_), .A1(new_n719_), .B0(new_n722_), .Y(new_n6304_));
  OAI21X1  g5919(.A0(new_n6304_), .A1(new_n727_), .B0(new_n729_), .Y(new_n6305_));
  AOI21X1  g5920(.A0(new_n6305_), .A1(new_n734_), .B0(new_n737_), .Y(new_n6306_));
  OAI21X1  g5921(.A0(new_n6306_), .A1(new_n742_), .B0(new_n744_), .Y(new_n6307_));
  AOI21X1  g5922(.A0(new_n6307_), .A1(new_n749_), .B0(new_n752_), .Y(new_n6308_));
  OAI21X1  g5923(.A0(new_n6308_), .A1(new_n757_), .B0(new_n759_), .Y(new_n6309_));
  AOI21X1  g5924(.A0(new_n6309_), .A1(new_n764_), .B0(new_n767_), .Y(new_n6310_));
  OAI21X1  g5925(.A0(new_n6310_), .A1(new_n772_), .B0(new_n774_), .Y(new_n6311_));
  AOI21X1  g5926(.A0(new_n6311_), .A1(new_n779_), .B0(new_n782_), .Y(new_n6312_));
  OAI21X1  g5927(.A0(new_n6312_), .A1(new_n787_), .B0(new_n789_), .Y(new_n6313_));
  AOI21X1  g5928(.A0(new_n6313_), .A1(new_n794_), .B0(new_n797_), .Y(new_n6314_));
  OAI21X1  g5929(.A0(new_n6314_), .A1(new_n802_), .B0(new_n804_), .Y(new_n6315_));
  AOI21X1  g5930(.A0(new_n6315_), .A1(new_n809_), .B0(new_n812_), .Y(new_n6316_));
  OAI21X1  g5931(.A0(new_n6316_), .A1(new_n817_), .B0(new_n819_), .Y(new_n6317_));
  AOI21X1  g5932(.A0(new_n6317_), .A1(new_n824_), .B0(new_n827_), .Y(new_n6318_));
  OAI21X1  g5933(.A0(new_n6318_), .A1(new_n832_), .B0(new_n834_), .Y(new_n6319_));
  AOI21X1  g5934(.A0(new_n6319_), .A1(new_n839_), .B0(new_n842_), .Y(new_n6320_));
  OAI21X1  g5935(.A0(new_n6320_), .A1(new_n847_), .B0(new_n849_), .Y(new_n6321_));
  AOI21X1  g5936(.A0(new_n6321_), .A1(new_n854_), .B0(new_n857_), .Y(new_n6322_));
  OAI21X1  g5937(.A0(new_n6322_), .A1(new_n862_), .B0(new_n864_), .Y(new_n6323_));
  AOI21X1  g5938(.A0(new_n6323_), .A1(new_n869_), .B0(new_n872_), .Y(new_n6324_));
  OAI21X1  g5939(.A0(new_n6324_), .A1(new_n877_), .B0(new_n879_), .Y(new_n6325_));
  AOI21X1  g5940(.A0(new_n6325_), .A1(new_n884_), .B0(new_n887_), .Y(new_n6326_));
  OAI21X1  g5941(.A0(new_n6326_), .A1(new_n892_), .B0(new_n894_), .Y(new_n6327_));
  AOI21X1  g5942(.A0(new_n6327_), .A1(new_n899_), .B0(new_n902_), .Y(new_n6328_));
  OAI21X1  g5943(.A0(new_n6328_), .A1(new_n907_), .B0(new_n909_), .Y(new_n6329_));
  AOI21X1  g5944(.A0(new_n6329_), .A1(new_n914_), .B0(new_n917_), .Y(new_n6330_));
  OAI21X1  g5945(.A0(new_n6330_), .A1(new_n922_), .B0(new_n924_), .Y(new_n6331_));
  AOI21X1  g5946(.A0(new_n6331_), .A1(new_n929_), .B0(new_n932_), .Y(new_n6332_));
  OAI21X1  g5947(.A0(new_n6332_), .A1(new_n937_), .B0(new_n939_), .Y(new_n6333_));
  AOI21X1  g5948(.A0(new_n6333_), .A1(new_n944_), .B0(new_n947_), .Y(new_n6334_));
  OAI21X1  g5949(.A0(new_n6334_), .A1(new_n952_), .B0(new_n954_), .Y(new_n6335_));
  AOI21X1  g5950(.A0(new_n6335_), .A1(new_n959_), .B0(new_n962_), .Y(new_n6336_));
  OAI21X1  g5951(.A0(new_n6336_), .A1(new_n967_), .B0(new_n969_), .Y(new_n6337_));
  OAI21X1  g5952(.A0(new_n1286_), .A1(\priority[111] ), .B0(\req[111] ), .Y(new_n6338_));
  AOI21X1  g5953(.A0(new_n6337_), .A1(new_n974_), .B0(new_n6338_), .Y(\grant[111] ));
  NOR2X1   g5954(.A(new_n1295_), .B(new_n983_), .Y(new_n6340_));
  OAI21X1  g5955(.A0(new_n6340_), .A1(new_n1450_), .B0(new_n991_), .Y(new_n6341_));
  AOI21X1  g5956(.A0(new_n6341_), .A1(new_n1448_), .B0(new_n1449_), .Y(new_n6342_));
  OAI21X1  g5957(.A0(new_n6342_), .A1(new_n1447_), .B0(new_n1006_), .Y(new_n6343_));
  AOI21X1  g5958(.A0(new_n6343_), .A1(new_n1445_), .B0(new_n1446_), .Y(new_n6344_));
  OAI21X1  g5959(.A0(new_n6344_), .A1(new_n1444_), .B0(new_n1547_), .Y(new_n6345_));
  AOI21X1  g5960(.A0(new_n6345_), .A1(new_n1549_), .B0(new_n1848_), .Y(new_n6346_));
  OAI21X1  g5961(.A0(new_n6346_), .A1(new_n1026_), .B0(new_n1028_), .Y(new_n6347_));
  AOI21X1  g5962(.A0(new_n6347_), .A1(new_n1033_), .B0(new_n1036_), .Y(new_n6348_));
  OAI21X1  g5963(.A0(new_n6348_), .A1(new_n1041_), .B0(new_n1043_), .Y(new_n6349_));
  AOI21X1  g5964(.A0(new_n6349_), .A1(new_n1048_), .B0(new_n1051_), .Y(new_n6350_));
  OAI21X1  g5965(.A0(new_n6350_), .A1(new_n1056_), .B0(new_n1058_), .Y(new_n6351_));
  AOI21X1  g5966(.A0(new_n6351_), .A1(new_n1063_), .B0(new_n1066_), .Y(new_n6352_));
  OAI21X1  g5967(.A0(new_n6352_), .A1(new_n1071_), .B0(new_n1073_), .Y(new_n6353_));
  AOI21X1  g5968(.A0(new_n6353_), .A1(new_n1078_), .B0(new_n1081_), .Y(new_n6354_));
  OAI21X1  g5969(.A0(new_n6354_), .A1(new_n1086_), .B0(new_n1088_), .Y(new_n6355_));
  AOI21X1  g5970(.A0(new_n6355_), .A1(new_n1093_), .B0(new_n1096_), .Y(new_n6356_));
  OAI21X1  g5971(.A0(new_n6356_), .A1(new_n1101_), .B0(new_n1103_), .Y(new_n6357_));
  AOI21X1  g5972(.A0(new_n6357_), .A1(new_n1108_), .B0(new_n1111_), .Y(new_n6358_));
  OAI21X1  g5973(.A0(new_n6358_), .A1(new_n1116_), .B0(new_n1118_), .Y(new_n6359_));
  AOI21X1  g5974(.A0(new_n6359_), .A1(new_n1123_), .B0(new_n1126_), .Y(new_n6360_));
  OAI21X1  g5975(.A0(new_n6360_), .A1(new_n1131_), .B0(new_n1133_), .Y(new_n6361_));
  AOI21X1  g5976(.A0(new_n6361_), .A1(new_n1138_), .B0(new_n1141_), .Y(new_n6362_));
  OAI21X1  g5977(.A0(new_n6362_), .A1(new_n1146_), .B0(new_n1148_), .Y(new_n6363_));
  AOI21X1  g5978(.A0(new_n6363_), .A1(new_n1153_), .B0(new_n1156_), .Y(new_n6364_));
  OAI21X1  g5979(.A0(new_n6364_), .A1(new_n1161_), .B0(new_n1163_), .Y(new_n6365_));
  AOI21X1  g5980(.A0(new_n6365_), .A1(new_n1168_), .B0(new_n1171_), .Y(new_n6366_));
  OAI21X1  g5981(.A0(new_n6366_), .A1(new_n1176_), .B0(new_n1178_), .Y(new_n6367_));
  AOI21X1  g5982(.A0(new_n6367_), .A1(new_n1183_), .B0(new_n1186_), .Y(new_n6368_));
  OAI21X1  g5983(.A0(new_n6368_), .A1(new_n1191_), .B0(new_n1193_), .Y(new_n6369_));
  AOI21X1  g5984(.A0(new_n6369_), .A1(new_n1198_), .B0(new_n1201_), .Y(new_n6370_));
  OAI21X1  g5985(.A0(new_n6370_), .A1(new_n1206_), .B0(new_n1208_), .Y(new_n6371_));
  AOI21X1  g5986(.A0(new_n6371_), .A1(new_n1213_), .B0(new_n1216_), .Y(new_n6372_));
  OAI21X1  g5987(.A0(new_n6372_), .A1(new_n1221_), .B0(new_n1223_), .Y(new_n6373_));
  AOI21X1  g5988(.A0(new_n6373_), .A1(new_n1228_), .B0(new_n1231_), .Y(new_n6374_));
  OAI21X1  g5989(.A0(new_n6374_), .A1(new_n1236_), .B0(new_n1238_), .Y(new_n6375_));
  AOI21X1  g5990(.A0(new_n6375_), .A1(new_n1243_), .B0(new_n1246_), .Y(new_n6376_));
  OAI21X1  g5991(.A0(new_n6376_), .A1(new_n1251_), .B0(new_n1253_), .Y(new_n6377_));
  AOI21X1  g5992(.A0(new_n6377_), .A1(new_n1258_), .B0(new_n1261_), .Y(new_n6378_));
  OAI21X1  g5993(.A0(new_n6378_), .A1(new_n1266_), .B0(new_n1268_), .Y(new_n6379_));
  AOI21X1  g5994(.A0(new_n6379_), .A1(new_n1273_), .B0(new_n1276_), .Y(new_n6380_));
  OAI21X1  g5995(.A0(new_n6380_), .A1(new_n1281_), .B0(new_n1283_), .Y(new_n6381_));
  OAI21X1  g5996(.A0(new_n662_), .A1(\priority[112] ), .B0(\req[112] ), .Y(new_n6382_));
  AOI21X1  g5997(.A0(new_n6381_), .A1(new_n1288_), .B0(new_n6382_), .Y(\grant[112] ));
  NOR2X1   g5998(.A(new_n1297_), .B(new_n670_), .Y(new_n6384_));
  OAI21X1  g5999(.A0(new_n6384_), .A1(new_n1559_), .B0(new_n1305_), .Y(new_n6385_));
  AOI21X1  g6000(.A0(new_n6385_), .A1(new_n1557_), .B0(new_n1558_), .Y(new_n6386_));
  OAI21X1  g6001(.A0(new_n6386_), .A1(new_n1556_), .B0(new_n1320_), .Y(new_n6387_));
  AOI21X1  g6002(.A0(new_n6387_), .A1(new_n1554_), .B0(new_n1555_), .Y(new_n6388_));
  OAI21X1  g6003(.A0(new_n6388_), .A1(new_n1553_), .B0(new_n1656_), .Y(new_n6389_));
  AOI21X1  g6004(.A0(new_n6389_), .A1(new_n1552_), .B0(new_n1893_), .Y(new_n6390_));
  OAI21X1  g6005(.A0(new_n6390_), .A1(new_n1395_), .B0(new_n403_), .Y(new_n6391_));
  AOI21X1  g6006(.A0(new_n6391_), .A1(new_n1393_), .B0(new_n1394_), .Y(new_n6392_));
  OAI21X1  g6007(.A0(new_n6392_), .A1(new_n1392_), .B0(new_n418_), .Y(new_n6393_));
  AOI21X1  g6008(.A0(new_n6393_), .A1(new_n1390_), .B0(new_n1391_), .Y(new_n6394_));
  OAI21X1  g6009(.A0(new_n6394_), .A1(new_n1389_), .B0(new_n433_), .Y(new_n6395_));
  AOI21X1  g6010(.A0(new_n6395_), .A1(new_n1387_), .B0(new_n1388_), .Y(new_n6396_));
  OAI21X1  g6011(.A0(new_n6396_), .A1(new_n1386_), .B0(new_n448_), .Y(new_n6397_));
  AOI21X1  g6012(.A0(new_n6397_), .A1(new_n1384_), .B0(new_n1385_), .Y(new_n6398_));
  OAI21X1  g6013(.A0(new_n6398_), .A1(new_n1383_), .B0(new_n463_), .Y(new_n6399_));
  AOI21X1  g6014(.A0(new_n6399_), .A1(new_n1381_), .B0(new_n1382_), .Y(new_n6400_));
  OAI21X1  g6015(.A0(new_n6400_), .A1(new_n1380_), .B0(new_n478_), .Y(new_n6401_));
  AOI21X1  g6016(.A0(new_n6401_), .A1(new_n1378_), .B0(new_n1379_), .Y(new_n6402_));
  OAI21X1  g6017(.A0(new_n6402_), .A1(new_n1377_), .B0(new_n493_), .Y(new_n6403_));
  AOI21X1  g6018(.A0(new_n6403_), .A1(new_n1375_), .B0(new_n1376_), .Y(new_n6404_));
  OAI21X1  g6019(.A0(new_n6404_), .A1(new_n1374_), .B0(new_n508_), .Y(new_n6405_));
  AOI21X1  g6020(.A0(new_n6405_), .A1(new_n1372_), .B0(new_n1373_), .Y(new_n6406_));
  OAI21X1  g6021(.A0(new_n6406_), .A1(new_n1371_), .B0(new_n523_), .Y(new_n6407_));
  AOI21X1  g6022(.A0(new_n6407_), .A1(new_n1369_), .B0(new_n1370_), .Y(new_n6408_));
  OAI21X1  g6023(.A0(new_n6408_), .A1(new_n1368_), .B0(new_n538_), .Y(new_n6409_));
  AOI21X1  g6024(.A0(new_n6409_), .A1(new_n1366_), .B0(new_n1367_), .Y(new_n6410_));
  OAI21X1  g6025(.A0(new_n6410_), .A1(new_n1365_), .B0(new_n553_), .Y(new_n6411_));
  AOI21X1  g6026(.A0(new_n6411_), .A1(new_n1363_), .B0(new_n1364_), .Y(new_n6412_));
  OAI21X1  g6027(.A0(new_n6412_), .A1(new_n1362_), .B0(new_n568_), .Y(new_n6413_));
  AOI21X1  g6028(.A0(new_n6413_), .A1(new_n1360_), .B0(new_n1361_), .Y(new_n6414_));
  OAI21X1  g6029(.A0(new_n6414_), .A1(new_n1359_), .B0(new_n583_), .Y(new_n6415_));
  AOI21X1  g6030(.A0(new_n6415_), .A1(new_n1357_), .B0(new_n1358_), .Y(new_n6416_));
  OAI21X1  g6031(.A0(new_n6416_), .A1(new_n1356_), .B0(new_n598_), .Y(new_n6417_));
  AOI21X1  g6032(.A0(new_n6417_), .A1(new_n1354_), .B0(new_n1355_), .Y(new_n6418_));
  OAI21X1  g6033(.A0(new_n6418_), .A1(new_n1353_), .B0(new_n613_), .Y(new_n6419_));
  AOI21X1  g6034(.A0(new_n6419_), .A1(new_n1351_), .B0(new_n1352_), .Y(new_n6420_));
  OAI21X1  g6035(.A0(new_n6420_), .A1(new_n1350_), .B0(new_n628_), .Y(new_n6421_));
  AOI21X1  g6036(.A0(new_n6421_), .A1(new_n1348_), .B0(new_n1349_), .Y(new_n6422_));
  OAI21X1  g6037(.A0(new_n6422_), .A1(new_n1347_), .B0(new_n643_), .Y(new_n6423_));
  AOI21X1  g6038(.A0(new_n6423_), .A1(new_n1345_), .B0(new_n1346_), .Y(new_n6424_));
  OAI21X1  g6039(.A0(new_n6424_), .A1(new_n1344_), .B0(new_n658_), .Y(new_n6425_));
  OAI21X1  g6040(.A0(new_n980_), .A1(\priority[113] ), .B0(\req[113] ), .Y(new_n6426_));
  AOI21X1  g6041(.A0(new_n6425_), .A1(new_n1342_), .B0(new_n6426_), .Y(\grant[113] ));
  NOR2X1   g6042(.A(new_n988_), .B(new_n672_), .Y(new_n6428_));
  OAI21X1  g6043(.A0(new_n6428_), .A1(new_n679_), .B0(new_n681_), .Y(new_n6429_));
  AOI21X1  g6044(.A0(new_n6429_), .A1(new_n686_), .B0(new_n689_), .Y(new_n6430_));
  OAI21X1  g6045(.A0(new_n6430_), .A1(new_n694_), .B0(new_n696_), .Y(new_n6431_));
  AOI21X1  g6046(.A0(new_n6431_), .A1(new_n701_), .B0(new_n1662_), .Y(new_n6432_));
  OAI21X1  g6047(.A0(new_n6432_), .A1(new_n1661_), .B0(new_n1705_), .Y(new_n6433_));
  AOI21X1  g6048(.A0(new_n6433_), .A1(new_n1660_), .B0(new_n1938_), .Y(new_n6434_));
  OAI21X1  g6049(.A0(new_n6434_), .A1(new_n1504_), .B0(new_n721_), .Y(new_n6435_));
  AOI21X1  g6050(.A0(new_n6435_), .A1(new_n1502_), .B0(new_n1503_), .Y(new_n6436_));
  OAI21X1  g6051(.A0(new_n6436_), .A1(new_n1501_), .B0(new_n736_), .Y(new_n6437_));
  AOI21X1  g6052(.A0(new_n6437_), .A1(new_n1499_), .B0(new_n1500_), .Y(new_n6438_));
  OAI21X1  g6053(.A0(new_n6438_), .A1(new_n1498_), .B0(new_n751_), .Y(new_n6439_));
  AOI21X1  g6054(.A0(new_n6439_), .A1(new_n1496_), .B0(new_n1497_), .Y(new_n6440_));
  OAI21X1  g6055(.A0(new_n6440_), .A1(new_n1495_), .B0(new_n766_), .Y(new_n6441_));
  AOI21X1  g6056(.A0(new_n6441_), .A1(new_n1493_), .B0(new_n1494_), .Y(new_n6442_));
  OAI21X1  g6057(.A0(new_n6442_), .A1(new_n1492_), .B0(new_n781_), .Y(new_n6443_));
  AOI21X1  g6058(.A0(new_n6443_), .A1(new_n1490_), .B0(new_n1491_), .Y(new_n6444_));
  OAI21X1  g6059(.A0(new_n6444_), .A1(new_n1489_), .B0(new_n796_), .Y(new_n6445_));
  AOI21X1  g6060(.A0(new_n6445_), .A1(new_n1487_), .B0(new_n1488_), .Y(new_n6446_));
  OAI21X1  g6061(.A0(new_n6446_), .A1(new_n1486_), .B0(new_n811_), .Y(new_n6447_));
  AOI21X1  g6062(.A0(new_n6447_), .A1(new_n1484_), .B0(new_n1485_), .Y(new_n6448_));
  OAI21X1  g6063(.A0(new_n6448_), .A1(new_n1483_), .B0(new_n826_), .Y(new_n6449_));
  AOI21X1  g6064(.A0(new_n6449_), .A1(new_n1481_), .B0(new_n1482_), .Y(new_n6450_));
  OAI21X1  g6065(.A0(new_n6450_), .A1(new_n1480_), .B0(new_n841_), .Y(new_n6451_));
  AOI21X1  g6066(.A0(new_n6451_), .A1(new_n1478_), .B0(new_n1479_), .Y(new_n6452_));
  OAI21X1  g6067(.A0(new_n6452_), .A1(new_n1477_), .B0(new_n856_), .Y(new_n6453_));
  AOI21X1  g6068(.A0(new_n6453_), .A1(new_n1475_), .B0(new_n1476_), .Y(new_n6454_));
  OAI21X1  g6069(.A0(new_n6454_), .A1(new_n1474_), .B0(new_n871_), .Y(new_n6455_));
  AOI21X1  g6070(.A0(new_n6455_), .A1(new_n1472_), .B0(new_n1473_), .Y(new_n6456_));
  OAI21X1  g6071(.A0(new_n6456_), .A1(new_n1471_), .B0(new_n886_), .Y(new_n6457_));
  AOI21X1  g6072(.A0(new_n6457_), .A1(new_n1469_), .B0(new_n1470_), .Y(new_n6458_));
  OAI21X1  g6073(.A0(new_n6458_), .A1(new_n1468_), .B0(new_n901_), .Y(new_n6459_));
  AOI21X1  g6074(.A0(new_n6459_), .A1(new_n1466_), .B0(new_n1467_), .Y(new_n6460_));
  OAI21X1  g6075(.A0(new_n6460_), .A1(new_n1465_), .B0(new_n916_), .Y(new_n6461_));
  AOI21X1  g6076(.A0(new_n6461_), .A1(new_n1463_), .B0(new_n1464_), .Y(new_n6462_));
  OAI21X1  g6077(.A0(new_n6462_), .A1(new_n1462_), .B0(new_n931_), .Y(new_n6463_));
  AOI21X1  g6078(.A0(new_n6463_), .A1(new_n1460_), .B0(new_n1461_), .Y(new_n6464_));
  OAI21X1  g6079(.A0(new_n6464_), .A1(new_n1459_), .B0(new_n946_), .Y(new_n6465_));
  AOI21X1  g6080(.A0(new_n6465_), .A1(new_n1457_), .B0(new_n1458_), .Y(new_n6466_));
  OAI21X1  g6081(.A0(new_n6466_), .A1(new_n1456_), .B0(new_n961_), .Y(new_n6467_));
  AOI21X1  g6082(.A0(new_n6467_), .A1(new_n1454_), .B0(new_n1455_), .Y(new_n6468_));
  OAI21X1  g6083(.A0(new_n6468_), .A1(new_n1453_), .B0(new_n976_), .Y(new_n6469_));
  OAI21X1  g6084(.A0(new_n1294_), .A1(\priority[114] ), .B0(\req[114] ), .Y(new_n6470_));
  AOI21X1  g6085(.A0(new_n6469_), .A1(new_n1451_), .B0(new_n6470_), .Y(\grant[114] ));
  NOR2X1   g6086(.A(new_n1302_), .B(new_n990_), .Y(new_n6472_));
  OAI21X1  g6087(.A0(new_n6472_), .A1(new_n997_), .B0(new_n999_), .Y(new_n6473_));
  AOI21X1  g6088(.A0(new_n6473_), .A1(new_n1004_), .B0(new_n1007_), .Y(new_n6474_));
  OAI21X1  g6089(.A0(new_n6474_), .A1(new_n1012_), .B0(new_n1014_), .Y(new_n6475_));
  AOI21X1  g6090(.A0(new_n6475_), .A1(new_n1017_), .B0(new_n1711_), .Y(new_n6476_));
  OAI21X1  g6091(.A0(new_n6476_), .A1(new_n1710_), .B0(new_n1754_), .Y(new_n6477_));
  AOI21X1  g6092(.A0(new_n6477_), .A1(new_n1709_), .B0(new_n1983_), .Y(new_n6478_));
  OAI21X1  g6093(.A0(new_n6478_), .A1(new_n1613_), .B0(new_n1035_), .Y(new_n6479_));
  AOI21X1  g6094(.A0(new_n6479_), .A1(new_n1611_), .B0(new_n1612_), .Y(new_n6480_));
  OAI21X1  g6095(.A0(new_n6480_), .A1(new_n1610_), .B0(new_n1050_), .Y(new_n6481_));
  AOI21X1  g6096(.A0(new_n6481_), .A1(new_n1608_), .B0(new_n1609_), .Y(new_n6482_));
  OAI21X1  g6097(.A0(new_n6482_), .A1(new_n1607_), .B0(new_n1065_), .Y(new_n6483_));
  AOI21X1  g6098(.A0(new_n6483_), .A1(new_n1605_), .B0(new_n1606_), .Y(new_n6484_));
  OAI21X1  g6099(.A0(new_n6484_), .A1(new_n1604_), .B0(new_n1080_), .Y(new_n6485_));
  AOI21X1  g6100(.A0(new_n6485_), .A1(new_n1602_), .B0(new_n1603_), .Y(new_n6486_));
  OAI21X1  g6101(.A0(new_n6486_), .A1(new_n1601_), .B0(new_n1095_), .Y(new_n6487_));
  AOI21X1  g6102(.A0(new_n6487_), .A1(new_n1599_), .B0(new_n1600_), .Y(new_n6488_));
  OAI21X1  g6103(.A0(new_n6488_), .A1(new_n1598_), .B0(new_n1110_), .Y(new_n6489_));
  AOI21X1  g6104(.A0(new_n6489_), .A1(new_n1596_), .B0(new_n1597_), .Y(new_n6490_));
  OAI21X1  g6105(.A0(new_n6490_), .A1(new_n1595_), .B0(new_n1125_), .Y(new_n6491_));
  AOI21X1  g6106(.A0(new_n6491_), .A1(new_n1593_), .B0(new_n1594_), .Y(new_n6492_));
  OAI21X1  g6107(.A0(new_n6492_), .A1(new_n1592_), .B0(new_n1140_), .Y(new_n6493_));
  AOI21X1  g6108(.A0(new_n6493_), .A1(new_n1590_), .B0(new_n1591_), .Y(new_n6494_));
  OAI21X1  g6109(.A0(new_n6494_), .A1(new_n1589_), .B0(new_n1155_), .Y(new_n6495_));
  AOI21X1  g6110(.A0(new_n6495_), .A1(new_n1587_), .B0(new_n1588_), .Y(new_n6496_));
  OAI21X1  g6111(.A0(new_n6496_), .A1(new_n1586_), .B0(new_n1170_), .Y(new_n6497_));
  AOI21X1  g6112(.A0(new_n6497_), .A1(new_n1584_), .B0(new_n1585_), .Y(new_n6498_));
  OAI21X1  g6113(.A0(new_n6498_), .A1(new_n1583_), .B0(new_n1185_), .Y(new_n6499_));
  AOI21X1  g6114(.A0(new_n6499_), .A1(new_n1581_), .B0(new_n1582_), .Y(new_n6500_));
  OAI21X1  g6115(.A0(new_n6500_), .A1(new_n1580_), .B0(new_n1200_), .Y(new_n6501_));
  AOI21X1  g6116(.A0(new_n6501_), .A1(new_n1578_), .B0(new_n1579_), .Y(new_n6502_));
  OAI21X1  g6117(.A0(new_n6502_), .A1(new_n1577_), .B0(new_n1215_), .Y(new_n6503_));
  AOI21X1  g6118(.A0(new_n6503_), .A1(new_n1575_), .B0(new_n1576_), .Y(new_n6504_));
  OAI21X1  g6119(.A0(new_n6504_), .A1(new_n1574_), .B0(new_n1230_), .Y(new_n6505_));
  AOI21X1  g6120(.A0(new_n6505_), .A1(new_n1572_), .B0(new_n1573_), .Y(new_n6506_));
  OAI21X1  g6121(.A0(new_n6506_), .A1(new_n1571_), .B0(new_n1245_), .Y(new_n6507_));
  AOI21X1  g6122(.A0(new_n6507_), .A1(new_n1569_), .B0(new_n1570_), .Y(new_n6508_));
  OAI21X1  g6123(.A0(new_n6508_), .A1(new_n1568_), .B0(new_n1260_), .Y(new_n6509_));
  AOI21X1  g6124(.A0(new_n6509_), .A1(new_n1566_), .B0(new_n1567_), .Y(new_n6510_));
  OAI21X1  g6125(.A0(new_n6510_), .A1(new_n1565_), .B0(new_n1275_), .Y(new_n6511_));
  AOI21X1  g6126(.A0(new_n6511_), .A1(new_n1563_), .B0(new_n1564_), .Y(new_n6512_));
  OAI21X1  g6127(.A0(new_n6512_), .A1(new_n1562_), .B0(new_n1290_), .Y(new_n6513_));
  OAI21X1  g6128(.A0(new_n669_), .A1(\priority[115] ), .B0(\req[115] ), .Y(new_n6514_));
  AOI21X1  g6129(.A0(new_n6513_), .A1(new_n1560_), .B0(new_n6514_), .Y(\grant[115] ));
  NOR2X1   g6130(.A(new_n1304_), .B(new_n678_), .Y(new_n6516_));
  OAI21X1  g6131(.A0(new_n6516_), .A1(new_n1311_), .B0(new_n1313_), .Y(new_n6517_));
  AOI21X1  g6132(.A0(new_n6517_), .A1(new_n1318_), .B0(new_n1321_), .Y(new_n6518_));
  OAI21X1  g6133(.A0(new_n6518_), .A1(new_n1326_), .B0(new_n1328_), .Y(new_n6519_));
  AOI21X1  g6134(.A0(new_n6519_), .A1(new_n1331_), .B0(new_n1758_), .Y(new_n6520_));
  OAI21X1  g6135(.A0(new_n6520_), .A1(new_n394_), .B0(new_n396_), .Y(new_n6521_));
  AOI21X1  g6136(.A0(new_n6521_), .A1(new_n401_), .B0(new_n404_), .Y(new_n6522_));
  OAI21X1  g6137(.A0(new_n6522_), .A1(new_n409_), .B0(new_n411_), .Y(new_n6523_));
  AOI21X1  g6138(.A0(new_n6523_), .A1(new_n416_), .B0(new_n419_), .Y(new_n6524_));
  OAI21X1  g6139(.A0(new_n6524_), .A1(new_n424_), .B0(new_n426_), .Y(new_n6525_));
  AOI21X1  g6140(.A0(new_n6525_), .A1(new_n431_), .B0(new_n434_), .Y(new_n6526_));
  OAI21X1  g6141(.A0(new_n6526_), .A1(new_n439_), .B0(new_n441_), .Y(new_n6527_));
  AOI21X1  g6142(.A0(new_n6527_), .A1(new_n446_), .B0(new_n449_), .Y(new_n6528_));
  OAI21X1  g6143(.A0(new_n6528_), .A1(new_n454_), .B0(new_n456_), .Y(new_n6529_));
  AOI21X1  g6144(.A0(new_n6529_), .A1(new_n461_), .B0(new_n464_), .Y(new_n6530_));
  OAI21X1  g6145(.A0(new_n6530_), .A1(new_n469_), .B0(new_n471_), .Y(new_n6531_));
  AOI21X1  g6146(.A0(new_n6531_), .A1(new_n476_), .B0(new_n479_), .Y(new_n6532_));
  OAI21X1  g6147(.A0(new_n6532_), .A1(new_n484_), .B0(new_n486_), .Y(new_n6533_));
  AOI21X1  g6148(.A0(new_n6533_), .A1(new_n491_), .B0(new_n494_), .Y(new_n6534_));
  OAI21X1  g6149(.A0(new_n6534_), .A1(new_n499_), .B0(new_n501_), .Y(new_n6535_));
  AOI21X1  g6150(.A0(new_n6535_), .A1(new_n506_), .B0(new_n509_), .Y(new_n6536_));
  OAI21X1  g6151(.A0(new_n6536_), .A1(new_n514_), .B0(new_n516_), .Y(new_n6537_));
  AOI21X1  g6152(.A0(new_n6537_), .A1(new_n521_), .B0(new_n524_), .Y(new_n6538_));
  OAI21X1  g6153(.A0(new_n6538_), .A1(new_n529_), .B0(new_n531_), .Y(new_n6539_));
  AOI21X1  g6154(.A0(new_n6539_), .A1(new_n536_), .B0(new_n539_), .Y(new_n6540_));
  OAI21X1  g6155(.A0(new_n6540_), .A1(new_n544_), .B0(new_n546_), .Y(new_n6541_));
  AOI21X1  g6156(.A0(new_n6541_), .A1(new_n551_), .B0(new_n554_), .Y(new_n6542_));
  OAI21X1  g6157(.A0(new_n6542_), .A1(new_n559_), .B0(new_n561_), .Y(new_n6543_));
  AOI21X1  g6158(.A0(new_n6543_), .A1(new_n566_), .B0(new_n569_), .Y(new_n6544_));
  OAI21X1  g6159(.A0(new_n6544_), .A1(new_n574_), .B0(new_n576_), .Y(new_n6545_));
  AOI21X1  g6160(.A0(new_n6545_), .A1(new_n581_), .B0(new_n584_), .Y(new_n6546_));
  OAI21X1  g6161(.A0(new_n6546_), .A1(new_n589_), .B0(new_n591_), .Y(new_n6547_));
  AOI21X1  g6162(.A0(new_n6547_), .A1(new_n596_), .B0(new_n599_), .Y(new_n6548_));
  OAI21X1  g6163(.A0(new_n6548_), .A1(new_n604_), .B0(new_n606_), .Y(new_n6549_));
  AOI21X1  g6164(.A0(new_n6549_), .A1(new_n611_), .B0(new_n614_), .Y(new_n6550_));
  OAI21X1  g6165(.A0(new_n6550_), .A1(new_n619_), .B0(new_n621_), .Y(new_n6551_));
  AOI21X1  g6166(.A0(new_n6551_), .A1(new_n626_), .B0(new_n629_), .Y(new_n6552_));
  OAI21X1  g6167(.A0(new_n6552_), .A1(new_n634_), .B0(new_n636_), .Y(new_n6553_));
  AOI21X1  g6168(.A0(new_n6553_), .A1(new_n641_), .B0(new_n644_), .Y(new_n6554_));
  OAI21X1  g6169(.A0(new_n6554_), .A1(new_n649_), .B0(new_n651_), .Y(new_n6555_));
  AOI21X1  g6170(.A0(new_n6555_), .A1(new_n656_), .B0(new_n659_), .Y(new_n6556_));
  OAI21X1  g6171(.A0(new_n6556_), .A1(new_n664_), .B0(new_n666_), .Y(new_n6557_));
  OAI21X1  g6172(.A0(new_n987_), .A1(\priority[116] ), .B0(\req[116] ), .Y(new_n6558_));
  AOI21X1  g6173(.A0(new_n6557_), .A1(new_n671_), .B0(new_n6558_), .Y(\grant[116] ));
  NOR2X1   g6174(.A(new_n996_), .B(new_n680_), .Y(new_n6560_));
  OAI21X1  g6175(.A0(new_n6560_), .A1(new_n1338_), .B0(new_n688_), .Y(new_n6561_));
  AOI21X1  g6176(.A0(new_n6561_), .A1(new_n1336_), .B0(new_n1337_), .Y(new_n6562_));
  OAI21X1  g6177(.A0(new_n6562_), .A1(new_n1335_), .B0(new_n1438_), .Y(new_n6563_));
  AOI21X1  g6178(.A0(new_n6563_), .A1(new_n1440_), .B0(new_n1803_), .Y(new_n6564_));
  OAI21X1  g6179(.A0(new_n6564_), .A1(new_n712_), .B0(new_n714_), .Y(new_n6565_));
  AOI21X1  g6180(.A0(new_n6565_), .A1(new_n719_), .B0(new_n722_), .Y(new_n6566_));
  OAI21X1  g6181(.A0(new_n6566_), .A1(new_n727_), .B0(new_n729_), .Y(new_n6567_));
  AOI21X1  g6182(.A0(new_n6567_), .A1(new_n734_), .B0(new_n737_), .Y(new_n6568_));
  OAI21X1  g6183(.A0(new_n6568_), .A1(new_n742_), .B0(new_n744_), .Y(new_n6569_));
  AOI21X1  g6184(.A0(new_n6569_), .A1(new_n749_), .B0(new_n752_), .Y(new_n6570_));
  OAI21X1  g6185(.A0(new_n6570_), .A1(new_n757_), .B0(new_n759_), .Y(new_n6571_));
  AOI21X1  g6186(.A0(new_n6571_), .A1(new_n764_), .B0(new_n767_), .Y(new_n6572_));
  OAI21X1  g6187(.A0(new_n6572_), .A1(new_n772_), .B0(new_n774_), .Y(new_n6573_));
  AOI21X1  g6188(.A0(new_n6573_), .A1(new_n779_), .B0(new_n782_), .Y(new_n6574_));
  OAI21X1  g6189(.A0(new_n6574_), .A1(new_n787_), .B0(new_n789_), .Y(new_n6575_));
  AOI21X1  g6190(.A0(new_n6575_), .A1(new_n794_), .B0(new_n797_), .Y(new_n6576_));
  OAI21X1  g6191(.A0(new_n6576_), .A1(new_n802_), .B0(new_n804_), .Y(new_n6577_));
  AOI21X1  g6192(.A0(new_n6577_), .A1(new_n809_), .B0(new_n812_), .Y(new_n6578_));
  OAI21X1  g6193(.A0(new_n6578_), .A1(new_n817_), .B0(new_n819_), .Y(new_n6579_));
  AOI21X1  g6194(.A0(new_n6579_), .A1(new_n824_), .B0(new_n827_), .Y(new_n6580_));
  OAI21X1  g6195(.A0(new_n6580_), .A1(new_n832_), .B0(new_n834_), .Y(new_n6581_));
  AOI21X1  g6196(.A0(new_n6581_), .A1(new_n839_), .B0(new_n842_), .Y(new_n6582_));
  OAI21X1  g6197(.A0(new_n6582_), .A1(new_n847_), .B0(new_n849_), .Y(new_n6583_));
  AOI21X1  g6198(.A0(new_n6583_), .A1(new_n854_), .B0(new_n857_), .Y(new_n6584_));
  OAI21X1  g6199(.A0(new_n6584_), .A1(new_n862_), .B0(new_n864_), .Y(new_n6585_));
  AOI21X1  g6200(.A0(new_n6585_), .A1(new_n869_), .B0(new_n872_), .Y(new_n6586_));
  OAI21X1  g6201(.A0(new_n6586_), .A1(new_n877_), .B0(new_n879_), .Y(new_n6587_));
  AOI21X1  g6202(.A0(new_n6587_), .A1(new_n884_), .B0(new_n887_), .Y(new_n6588_));
  OAI21X1  g6203(.A0(new_n6588_), .A1(new_n892_), .B0(new_n894_), .Y(new_n6589_));
  AOI21X1  g6204(.A0(new_n6589_), .A1(new_n899_), .B0(new_n902_), .Y(new_n6590_));
  OAI21X1  g6205(.A0(new_n6590_), .A1(new_n907_), .B0(new_n909_), .Y(new_n6591_));
  AOI21X1  g6206(.A0(new_n6591_), .A1(new_n914_), .B0(new_n917_), .Y(new_n6592_));
  OAI21X1  g6207(.A0(new_n6592_), .A1(new_n922_), .B0(new_n924_), .Y(new_n6593_));
  AOI21X1  g6208(.A0(new_n6593_), .A1(new_n929_), .B0(new_n932_), .Y(new_n6594_));
  OAI21X1  g6209(.A0(new_n6594_), .A1(new_n937_), .B0(new_n939_), .Y(new_n6595_));
  AOI21X1  g6210(.A0(new_n6595_), .A1(new_n944_), .B0(new_n947_), .Y(new_n6596_));
  OAI21X1  g6211(.A0(new_n6596_), .A1(new_n952_), .B0(new_n954_), .Y(new_n6597_));
  AOI21X1  g6212(.A0(new_n6597_), .A1(new_n959_), .B0(new_n962_), .Y(new_n6598_));
  OAI21X1  g6213(.A0(new_n6598_), .A1(new_n967_), .B0(new_n969_), .Y(new_n6599_));
  AOI21X1  g6214(.A0(new_n6599_), .A1(new_n974_), .B0(new_n977_), .Y(new_n6600_));
  OAI21X1  g6215(.A0(new_n6600_), .A1(new_n982_), .B0(new_n984_), .Y(new_n6601_));
  OAI21X1  g6216(.A0(new_n1301_), .A1(\priority[117] ), .B0(\req[117] ), .Y(new_n6602_));
  AOI21X1  g6217(.A0(new_n6601_), .A1(new_n989_), .B0(new_n6602_), .Y(\grant[117] ));
  NOR2X1   g6218(.A(new_n1310_), .B(new_n998_), .Y(new_n6604_));
  OAI21X1  g6219(.A0(new_n6604_), .A1(new_n1447_), .B0(new_n1006_), .Y(new_n6605_));
  AOI21X1  g6220(.A0(new_n6605_), .A1(new_n1445_), .B0(new_n1446_), .Y(new_n6606_));
  OAI21X1  g6221(.A0(new_n6606_), .A1(new_n1444_), .B0(new_n1547_), .Y(new_n6607_));
  AOI21X1  g6222(.A0(new_n6607_), .A1(new_n1549_), .B0(new_n1848_), .Y(new_n6608_));
  OAI21X1  g6223(.A0(new_n6608_), .A1(new_n1026_), .B0(new_n1028_), .Y(new_n6609_));
  AOI21X1  g6224(.A0(new_n6609_), .A1(new_n1033_), .B0(new_n1036_), .Y(new_n6610_));
  OAI21X1  g6225(.A0(new_n6610_), .A1(new_n1041_), .B0(new_n1043_), .Y(new_n6611_));
  AOI21X1  g6226(.A0(new_n6611_), .A1(new_n1048_), .B0(new_n1051_), .Y(new_n6612_));
  OAI21X1  g6227(.A0(new_n6612_), .A1(new_n1056_), .B0(new_n1058_), .Y(new_n6613_));
  AOI21X1  g6228(.A0(new_n6613_), .A1(new_n1063_), .B0(new_n1066_), .Y(new_n6614_));
  OAI21X1  g6229(.A0(new_n6614_), .A1(new_n1071_), .B0(new_n1073_), .Y(new_n6615_));
  AOI21X1  g6230(.A0(new_n6615_), .A1(new_n1078_), .B0(new_n1081_), .Y(new_n6616_));
  OAI21X1  g6231(.A0(new_n6616_), .A1(new_n1086_), .B0(new_n1088_), .Y(new_n6617_));
  AOI21X1  g6232(.A0(new_n6617_), .A1(new_n1093_), .B0(new_n1096_), .Y(new_n6618_));
  OAI21X1  g6233(.A0(new_n6618_), .A1(new_n1101_), .B0(new_n1103_), .Y(new_n6619_));
  AOI21X1  g6234(.A0(new_n6619_), .A1(new_n1108_), .B0(new_n1111_), .Y(new_n6620_));
  OAI21X1  g6235(.A0(new_n6620_), .A1(new_n1116_), .B0(new_n1118_), .Y(new_n6621_));
  AOI21X1  g6236(.A0(new_n6621_), .A1(new_n1123_), .B0(new_n1126_), .Y(new_n6622_));
  OAI21X1  g6237(.A0(new_n6622_), .A1(new_n1131_), .B0(new_n1133_), .Y(new_n6623_));
  AOI21X1  g6238(.A0(new_n6623_), .A1(new_n1138_), .B0(new_n1141_), .Y(new_n6624_));
  OAI21X1  g6239(.A0(new_n6624_), .A1(new_n1146_), .B0(new_n1148_), .Y(new_n6625_));
  AOI21X1  g6240(.A0(new_n6625_), .A1(new_n1153_), .B0(new_n1156_), .Y(new_n6626_));
  OAI21X1  g6241(.A0(new_n6626_), .A1(new_n1161_), .B0(new_n1163_), .Y(new_n6627_));
  AOI21X1  g6242(.A0(new_n6627_), .A1(new_n1168_), .B0(new_n1171_), .Y(new_n6628_));
  OAI21X1  g6243(.A0(new_n6628_), .A1(new_n1176_), .B0(new_n1178_), .Y(new_n6629_));
  AOI21X1  g6244(.A0(new_n6629_), .A1(new_n1183_), .B0(new_n1186_), .Y(new_n6630_));
  OAI21X1  g6245(.A0(new_n6630_), .A1(new_n1191_), .B0(new_n1193_), .Y(new_n6631_));
  AOI21X1  g6246(.A0(new_n6631_), .A1(new_n1198_), .B0(new_n1201_), .Y(new_n6632_));
  OAI21X1  g6247(.A0(new_n6632_), .A1(new_n1206_), .B0(new_n1208_), .Y(new_n6633_));
  AOI21X1  g6248(.A0(new_n6633_), .A1(new_n1213_), .B0(new_n1216_), .Y(new_n6634_));
  OAI21X1  g6249(.A0(new_n6634_), .A1(new_n1221_), .B0(new_n1223_), .Y(new_n6635_));
  AOI21X1  g6250(.A0(new_n6635_), .A1(new_n1228_), .B0(new_n1231_), .Y(new_n6636_));
  OAI21X1  g6251(.A0(new_n6636_), .A1(new_n1236_), .B0(new_n1238_), .Y(new_n6637_));
  AOI21X1  g6252(.A0(new_n6637_), .A1(new_n1243_), .B0(new_n1246_), .Y(new_n6638_));
  OAI21X1  g6253(.A0(new_n6638_), .A1(new_n1251_), .B0(new_n1253_), .Y(new_n6639_));
  AOI21X1  g6254(.A0(new_n6639_), .A1(new_n1258_), .B0(new_n1261_), .Y(new_n6640_));
  OAI21X1  g6255(.A0(new_n6640_), .A1(new_n1266_), .B0(new_n1268_), .Y(new_n6641_));
  AOI21X1  g6256(.A0(new_n6641_), .A1(new_n1273_), .B0(new_n1276_), .Y(new_n6642_));
  OAI21X1  g6257(.A0(new_n6642_), .A1(new_n1281_), .B0(new_n1283_), .Y(new_n6643_));
  AOI21X1  g6258(.A0(new_n6643_), .A1(new_n1288_), .B0(new_n1291_), .Y(new_n6644_));
  OAI21X1  g6259(.A0(new_n6644_), .A1(new_n1296_), .B0(new_n1298_), .Y(new_n6645_));
  OAI21X1  g6260(.A0(new_n677_), .A1(\priority[118] ), .B0(\req[118] ), .Y(new_n6646_));
  AOI21X1  g6261(.A0(new_n6645_), .A1(new_n1303_), .B0(new_n6646_), .Y(\grant[118] ));
  NOR2X1   g6262(.A(new_n1312_), .B(new_n685_), .Y(new_n6648_));
  OAI21X1  g6263(.A0(new_n6648_), .A1(new_n1556_), .B0(new_n1320_), .Y(new_n6649_));
  AOI21X1  g6264(.A0(new_n6649_), .A1(new_n1554_), .B0(new_n1555_), .Y(new_n6650_));
  OAI21X1  g6265(.A0(new_n6650_), .A1(new_n1553_), .B0(new_n1656_), .Y(new_n6651_));
  AOI21X1  g6266(.A0(new_n6651_), .A1(new_n1552_), .B0(new_n1893_), .Y(new_n6652_));
  OAI21X1  g6267(.A0(new_n6652_), .A1(new_n1395_), .B0(new_n403_), .Y(new_n6653_));
  AOI21X1  g6268(.A0(new_n6653_), .A1(new_n1393_), .B0(new_n1394_), .Y(new_n6654_));
  OAI21X1  g6269(.A0(new_n6654_), .A1(new_n1392_), .B0(new_n418_), .Y(new_n6655_));
  AOI21X1  g6270(.A0(new_n6655_), .A1(new_n1390_), .B0(new_n1391_), .Y(new_n6656_));
  OAI21X1  g6271(.A0(new_n6656_), .A1(new_n1389_), .B0(new_n433_), .Y(new_n6657_));
  AOI21X1  g6272(.A0(new_n6657_), .A1(new_n1387_), .B0(new_n1388_), .Y(new_n6658_));
  OAI21X1  g6273(.A0(new_n6658_), .A1(new_n1386_), .B0(new_n448_), .Y(new_n6659_));
  AOI21X1  g6274(.A0(new_n6659_), .A1(new_n1384_), .B0(new_n1385_), .Y(new_n6660_));
  OAI21X1  g6275(.A0(new_n6660_), .A1(new_n1383_), .B0(new_n463_), .Y(new_n6661_));
  AOI21X1  g6276(.A0(new_n6661_), .A1(new_n1381_), .B0(new_n1382_), .Y(new_n6662_));
  OAI21X1  g6277(.A0(new_n6662_), .A1(new_n1380_), .B0(new_n478_), .Y(new_n6663_));
  AOI21X1  g6278(.A0(new_n6663_), .A1(new_n1378_), .B0(new_n1379_), .Y(new_n6664_));
  OAI21X1  g6279(.A0(new_n6664_), .A1(new_n1377_), .B0(new_n493_), .Y(new_n6665_));
  AOI21X1  g6280(.A0(new_n6665_), .A1(new_n1375_), .B0(new_n1376_), .Y(new_n6666_));
  OAI21X1  g6281(.A0(new_n6666_), .A1(new_n1374_), .B0(new_n508_), .Y(new_n6667_));
  AOI21X1  g6282(.A0(new_n6667_), .A1(new_n1372_), .B0(new_n1373_), .Y(new_n6668_));
  OAI21X1  g6283(.A0(new_n6668_), .A1(new_n1371_), .B0(new_n523_), .Y(new_n6669_));
  AOI21X1  g6284(.A0(new_n6669_), .A1(new_n1369_), .B0(new_n1370_), .Y(new_n6670_));
  OAI21X1  g6285(.A0(new_n6670_), .A1(new_n1368_), .B0(new_n538_), .Y(new_n6671_));
  AOI21X1  g6286(.A0(new_n6671_), .A1(new_n1366_), .B0(new_n1367_), .Y(new_n6672_));
  OAI21X1  g6287(.A0(new_n6672_), .A1(new_n1365_), .B0(new_n553_), .Y(new_n6673_));
  AOI21X1  g6288(.A0(new_n6673_), .A1(new_n1363_), .B0(new_n1364_), .Y(new_n6674_));
  OAI21X1  g6289(.A0(new_n6674_), .A1(new_n1362_), .B0(new_n568_), .Y(new_n6675_));
  AOI21X1  g6290(.A0(new_n6675_), .A1(new_n1360_), .B0(new_n1361_), .Y(new_n6676_));
  OAI21X1  g6291(.A0(new_n6676_), .A1(new_n1359_), .B0(new_n583_), .Y(new_n6677_));
  AOI21X1  g6292(.A0(new_n6677_), .A1(new_n1357_), .B0(new_n1358_), .Y(new_n6678_));
  OAI21X1  g6293(.A0(new_n6678_), .A1(new_n1356_), .B0(new_n598_), .Y(new_n6679_));
  AOI21X1  g6294(.A0(new_n6679_), .A1(new_n1354_), .B0(new_n1355_), .Y(new_n6680_));
  OAI21X1  g6295(.A0(new_n6680_), .A1(new_n1353_), .B0(new_n613_), .Y(new_n6681_));
  AOI21X1  g6296(.A0(new_n6681_), .A1(new_n1351_), .B0(new_n1352_), .Y(new_n6682_));
  OAI21X1  g6297(.A0(new_n6682_), .A1(new_n1350_), .B0(new_n628_), .Y(new_n6683_));
  AOI21X1  g6298(.A0(new_n6683_), .A1(new_n1348_), .B0(new_n1349_), .Y(new_n6684_));
  OAI21X1  g6299(.A0(new_n6684_), .A1(new_n1347_), .B0(new_n643_), .Y(new_n6685_));
  AOI21X1  g6300(.A0(new_n6685_), .A1(new_n1345_), .B0(new_n1346_), .Y(new_n6686_));
  OAI21X1  g6301(.A0(new_n6686_), .A1(new_n1344_), .B0(new_n658_), .Y(new_n6687_));
  AOI21X1  g6302(.A0(new_n6687_), .A1(new_n1342_), .B0(new_n1343_), .Y(new_n6688_));
  OAI21X1  g6303(.A0(new_n6688_), .A1(new_n1341_), .B0(new_n673_), .Y(new_n6689_));
  OAI21X1  g6304(.A0(new_n995_), .A1(\priority[119] ), .B0(\req[119] ), .Y(new_n6690_));
  AOI21X1  g6305(.A0(new_n6689_), .A1(new_n1339_), .B0(new_n6690_), .Y(\grant[119] ));
  NOR2X1   g6306(.A(new_n1003_), .B(new_n687_), .Y(new_n6692_));
  OAI21X1  g6307(.A0(new_n6692_), .A1(new_n694_), .B0(new_n696_), .Y(new_n6693_));
  AOI21X1  g6308(.A0(new_n6693_), .A1(new_n701_), .B0(new_n1662_), .Y(new_n6694_));
  OAI21X1  g6309(.A0(new_n6694_), .A1(new_n1661_), .B0(new_n1705_), .Y(new_n6695_));
  AOI21X1  g6310(.A0(new_n6695_), .A1(new_n1660_), .B0(new_n1938_), .Y(new_n6696_));
  OAI21X1  g6311(.A0(new_n6696_), .A1(new_n1504_), .B0(new_n721_), .Y(new_n6697_));
  AOI21X1  g6312(.A0(new_n6697_), .A1(new_n1502_), .B0(new_n1503_), .Y(new_n6698_));
  OAI21X1  g6313(.A0(new_n6698_), .A1(new_n1501_), .B0(new_n736_), .Y(new_n6699_));
  AOI21X1  g6314(.A0(new_n6699_), .A1(new_n1499_), .B0(new_n1500_), .Y(new_n6700_));
  OAI21X1  g6315(.A0(new_n6700_), .A1(new_n1498_), .B0(new_n751_), .Y(new_n6701_));
  AOI21X1  g6316(.A0(new_n6701_), .A1(new_n1496_), .B0(new_n1497_), .Y(new_n6702_));
  OAI21X1  g6317(.A0(new_n6702_), .A1(new_n1495_), .B0(new_n766_), .Y(new_n6703_));
  AOI21X1  g6318(.A0(new_n6703_), .A1(new_n1493_), .B0(new_n1494_), .Y(new_n6704_));
  OAI21X1  g6319(.A0(new_n6704_), .A1(new_n1492_), .B0(new_n781_), .Y(new_n6705_));
  AOI21X1  g6320(.A0(new_n6705_), .A1(new_n1490_), .B0(new_n1491_), .Y(new_n6706_));
  OAI21X1  g6321(.A0(new_n6706_), .A1(new_n1489_), .B0(new_n796_), .Y(new_n6707_));
  AOI21X1  g6322(.A0(new_n6707_), .A1(new_n1487_), .B0(new_n1488_), .Y(new_n6708_));
  OAI21X1  g6323(.A0(new_n6708_), .A1(new_n1486_), .B0(new_n811_), .Y(new_n6709_));
  AOI21X1  g6324(.A0(new_n6709_), .A1(new_n1484_), .B0(new_n1485_), .Y(new_n6710_));
  OAI21X1  g6325(.A0(new_n6710_), .A1(new_n1483_), .B0(new_n826_), .Y(new_n6711_));
  AOI21X1  g6326(.A0(new_n6711_), .A1(new_n1481_), .B0(new_n1482_), .Y(new_n6712_));
  OAI21X1  g6327(.A0(new_n6712_), .A1(new_n1480_), .B0(new_n841_), .Y(new_n6713_));
  AOI21X1  g6328(.A0(new_n6713_), .A1(new_n1478_), .B0(new_n1479_), .Y(new_n6714_));
  OAI21X1  g6329(.A0(new_n6714_), .A1(new_n1477_), .B0(new_n856_), .Y(new_n6715_));
  AOI21X1  g6330(.A0(new_n6715_), .A1(new_n1475_), .B0(new_n1476_), .Y(new_n6716_));
  OAI21X1  g6331(.A0(new_n6716_), .A1(new_n1474_), .B0(new_n871_), .Y(new_n6717_));
  AOI21X1  g6332(.A0(new_n6717_), .A1(new_n1472_), .B0(new_n1473_), .Y(new_n6718_));
  OAI21X1  g6333(.A0(new_n6718_), .A1(new_n1471_), .B0(new_n886_), .Y(new_n6719_));
  AOI21X1  g6334(.A0(new_n6719_), .A1(new_n1469_), .B0(new_n1470_), .Y(new_n6720_));
  OAI21X1  g6335(.A0(new_n6720_), .A1(new_n1468_), .B0(new_n901_), .Y(new_n6721_));
  AOI21X1  g6336(.A0(new_n6721_), .A1(new_n1466_), .B0(new_n1467_), .Y(new_n6722_));
  OAI21X1  g6337(.A0(new_n6722_), .A1(new_n1465_), .B0(new_n916_), .Y(new_n6723_));
  AOI21X1  g6338(.A0(new_n6723_), .A1(new_n1463_), .B0(new_n1464_), .Y(new_n6724_));
  OAI21X1  g6339(.A0(new_n6724_), .A1(new_n1462_), .B0(new_n931_), .Y(new_n6725_));
  AOI21X1  g6340(.A0(new_n6725_), .A1(new_n1460_), .B0(new_n1461_), .Y(new_n6726_));
  OAI21X1  g6341(.A0(new_n6726_), .A1(new_n1459_), .B0(new_n946_), .Y(new_n6727_));
  AOI21X1  g6342(.A0(new_n6727_), .A1(new_n1457_), .B0(new_n1458_), .Y(new_n6728_));
  OAI21X1  g6343(.A0(new_n6728_), .A1(new_n1456_), .B0(new_n961_), .Y(new_n6729_));
  AOI21X1  g6344(.A0(new_n6729_), .A1(new_n1454_), .B0(new_n1455_), .Y(new_n6730_));
  OAI21X1  g6345(.A0(new_n6730_), .A1(new_n1453_), .B0(new_n976_), .Y(new_n6731_));
  AOI21X1  g6346(.A0(new_n6731_), .A1(new_n1451_), .B0(new_n1452_), .Y(new_n6732_));
  OAI21X1  g6347(.A0(new_n6732_), .A1(new_n1450_), .B0(new_n991_), .Y(new_n6733_));
  OAI21X1  g6348(.A0(new_n1309_), .A1(\priority[120] ), .B0(\req[120] ), .Y(new_n6734_));
  AOI21X1  g6349(.A0(new_n6733_), .A1(new_n1448_), .B0(new_n6734_), .Y(\grant[120] ));
  NOR2X1   g6350(.A(new_n1317_), .B(new_n1005_), .Y(new_n6736_));
  OAI21X1  g6351(.A0(new_n6736_), .A1(new_n1012_), .B0(new_n1014_), .Y(new_n6737_));
  AOI21X1  g6352(.A0(new_n6737_), .A1(new_n1017_), .B0(new_n1711_), .Y(new_n6738_));
  OAI21X1  g6353(.A0(new_n6738_), .A1(new_n1710_), .B0(new_n1754_), .Y(new_n6739_));
  AOI21X1  g6354(.A0(new_n6739_), .A1(new_n1709_), .B0(new_n1983_), .Y(new_n6740_));
  OAI21X1  g6355(.A0(new_n6740_), .A1(new_n1613_), .B0(new_n1035_), .Y(new_n6741_));
  AOI21X1  g6356(.A0(new_n6741_), .A1(new_n1611_), .B0(new_n1612_), .Y(new_n6742_));
  OAI21X1  g6357(.A0(new_n6742_), .A1(new_n1610_), .B0(new_n1050_), .Y(new_n6743_));
  AOI21X1  g6358(.A0(new_n6743_), .A1(new_n1608_), .B0(new_n1609_), .Y(new_n6744_));
  OAI21X1  g6359(.A0(new_n6744_), .A1(new_n1607_), .B0(new_n1065_), .Y(new_n6745_));
  AOI21X1  g6360(.A0(new_n6745_), .A1(new_n1605_), .B0(new_n1606_), .Y(new_n6746_));
  OAI21X1  g6361(.A0(new_n6746_), .A1(new_n1604_), .B0(new_n1080_), .Y(new_n6747_));
  AOI21X1  g6362(.A0(new_n6747_), .A1(new_n1602_), .B0(new_n1603_), .Y(new_n6748_));
  OAI21X1  g6363(.A0(new_n6748_), .A1(new_n1601_), .B0(new_n1095_), .Y(new_n6749_));
  AOI21X1  g6364(.A0(new_n6749_), .A1(new_n1599_), .B0(new_n1600_), .Y(new_n6750_));
  OAI21X1  g6365(.A0(new_n6750_), .A1(new_n1598_), .B0(new_n1110_), .Y(new_n6751_));
  AOI21X1  g6366(.A0(new_n6751_), .A1(new_n1596_), .B0(new_n1597_), .Y(new_n6752_));
  OAI21X1  g6367(.A0(new_n6752_), .A1(new_n1595_), .B0(new_n1125_), .Y(new_n6753_));
  AOI21X1  g6368(.A0(new_n6753_), .A1(new_n1593_), .B0(new_n1594_), .Y(new_n6754_));
  OAI21X1  g6369(.A0(new_n6754_), .A1(new_n1592_), .B0(new_n1140_), .Y(new_n6755_));
  AOI21X1  g6370(.A0(new_n6755_), .A1(new_n1590_), .B0(new_n1591_), .Y(new_n6756_));
  OAI21X1  g6371(.A0(new_n6756_), .A1(new_n1589_), .B0(new_n1155_), .Y(new_n6757_));
  AOI21X1  g6372(.A0(new_n6757_), .A1(new_n1587_), .B0(new_n1588_), .Y(new_n6758_));
  OAI21X1  g6373(.A0(new_n6758_), .A1(new_n1586_), .B0(new_n1170_), .Y(new_n6759_));
  AOI21X1  g6374(.A0(new_n6759_), .A1(new_n1584_), .B0(new_n1585_), .Y(new_n6760_));
  OAI21X1  g6375(.A0(new_n6760_), .A1(new_n1583_), .B0(new_n1185_), .Y(new_n6761_));
  AOI21X1  g6376(.A0(new_n6761_), .A1(new_n1581_), .B0(new_n1582_), .Y(new_n6762_));
  OAI21X1  g6377(.A0(new_n6762_), .A1(new_n1580_), .B0(new_n1200_), .Y(new_n6763_));
  AOI21X1  g6378(.A0(new_n6763_), .A1(new_n1578_), .B0(new_n1579_), .Y(new_n6764_));
  OAI21X1  g6379(.A0(new_n6764_), .A1(new_n1577_), .B0(new_n1215_), .Y(new_n6765_));
  AOI21X1  g6380(.A0(new_n6765_), .A1(new_n1575_), .B0(new_n1576_), .Y(new_n6766_));
  OAI21X1  g6381(.A0(new_n6766_), .A1(new_n1574_), .B0(new_n1230_), .Y(new_n6767_));
  AOI21X1  g6382(.A0(new_n6767_), .A1(new_n1572_), .B0(new_n1573_), .Y(new_n6768_));
  OAI21X1  g6383(.A0(new_n6768_), .A1(new_n1571_), .B0(new_n1245_), .Y(new_n6769_));
  AOI21X1  g6384(.A0(new_n6769_), .A1(new_n1569_), .B0(new_n1570_), .Y(new_n6770_));
  OAI21X1  g6385(.A0(new_n6770_), .A1(new_n1568_), .B0(new_n1260_), .Y(new_n6771_));
  AOI21X1  g6386(.A0(new_n6771_), .A1(new_n1566_), .B0(new_n1567_), .Y(new_n6772_));
  OAI21X1  g6387(.A0(new_n6772_), .A1(new_n1565_), .B0(new_n1275_), .Y(new_n6773_));
  AOI21X1  g6388(.A0(new_n6773_), .A1(new_n1563_), .B0(new_n1564_), .Y(new_n6774_));
  OAI21X1  g6389(.A0(new_n6774_), .A1(new_n1562_), .B0(new_n1290_), .Y(new_n6775_));
  AOI21X1  g6390(.A0(new_n6775_), .A1(new_n1560_), .B0(new_n1561_), .Y(new_n6776_));
  OAI21X1  g6391(.A0(new_n6776_), .A1(new_n1559_), .B0(new_n1305_), .Y(new_n6777_));
  OAI21X1  g6392(.A0(new_n684_), .A1(\priority[121] ), .B0(\req[121] ), .Y(new_n6778_));
  AOI21X1  g6393(.A0(new_n6777_), .A1(new_n1557_), .B0(new_n6778_), .Y(\grant[121] ));
  NOR2X1   g6394(.A(new_n1319_), .B(new_n693_), .Y(new_n6780_));
  OAI21X1  g6395(.A0(new_n6780_), .A1(new_n1326_), .B0(new_n1328_), .Y(new_n6781_));
  AOI21X1  g6396(.A0(new_n6781_), .A1(new_n1331_), .B0(new_n1758_), .Y(new_n6782_));
  OAI21X1  g6397(.A0(new_n6782_), .A1(new_n394_), .B0(new_n396_), .Y(new_n6783_));
  AOI21X1  g6398(.A0(new_n6783_), .A1(new_n401_), .B0(new_n404_), .Y(new_n6784_));
  OAI21X1  g6399(.A0(new_n6784_), .A1(new_n409_), .B0(new_n411_), .Y(new_n6785_));
  AOI21X1  g6400(.A0(new_n6785_), .A1(new_n416_), .B0(new_n419_), .Y(new_n6786_));
  OAI21X1  g6401(.A0(new_n6786_), .A1(new_n424_), .B0(new_n426_), .Y(new_n6787_));
  AOI21X1  g6402(.A0(new_n6787_), .A1(new_n431_), .B0(new_n434_), .Y(new_n6788_));
  OAI21X1  g6403(.A0(new_n6788_), .A1(new_n439_), .B0(new_n441_), .Y(new_n6789_));
  AOI21X1  g6404(.A0(new_n6789_), .A1(new_n446_), .B0(new_n449_), .Y(new_n6790_));
  OAI21X1  g6405(.A0(new_n6790_), .A1(new_n454_), .B0(new_n456_), .Y(new_n6791_));
  AOI21X1  g6406(.A0(new_n6791_), .A1(new_n461_), .B0(new_n464_), .Y(new_n6792_));
  OAI21X1  g6407(.A0(new_n6792_), .A1(new_n469_), .B0(new_n471_), .Y(new_n6793_));
  AOI21X1  g6408(.A0(new_n6793_), .A1(new_n476_), .B0(new_n479_), .Y(new_n6794_));
  OAI21X1  g6409(.A0(new_n6794_), .A1(new_n484_), .B0(new_n486_), .Y(new_n6795_));
  AOI21X1  g6410(.A0(new_n6795_), .A1(new_n491_), .B0(new_n494_), .Y(new_n6796_));
  OAI21X1  g6411(.A0(new_n6796_), .A1(new_n499_), .B0(new_n501_), .Y(new_n6797_));
  AOI21X1  g6412(.A0(new_n6797_), .A1(new_n506_), .B0(new_n509_), .Y(new_n6798_));
  OAI21X1  g6413(.A0(new_n6798_), .A1(new_n514_), .B0(new_n516_), .Y(new_n6799_));
  AOI21X1  g6414(.A0(new_n6799_), .A1(new_n521_), .B0(new_n524_), .Y(new_n6800_));
  OAI21X1  g6415(.A0(new_n6800_), .A1(new_n529_), .B0(new_n531_), .Y(new_n6801_));
  AOI21X1  g6416(.A0(new_n6801_), .A1(new_n536_), .B0(new_n539_), .Y(new_n6802_));
  OAI21X1  g6417(.A0(new_n6802_), .A1(new_n544_), .B0(new_n546_), .Y(new_n6803_));
  AOI21X1  g6418(.A0(new_n6803_), .A1(new_n551_), .B0(new_n554_), .Y(new_n6804_));
  OAI21X1  g6419(.A0(new_n6804_), .A1(new_n559_), .B0(new_n561_), .Y(new_n6805_));
  AOI21X1  g6420(.A0(new_n6805_), .A1(new_n566_), .B0(new_n569_), .Y(new_n6806_));
  OAI21X1  g6421(.A0(new_n6806_), .A1(new_n574_), .B0(new_n576_), .Y(new_n6807_));
  AOI21X1  g6422(.A0(new_n6807_), .A1(new_n581_), .B0(new_n584_), .Y(new_n6808_));
  OAI21X1  g6423(.A0(new_n6808_), .A1(new_n589_), .B0(new_n591_), .Y(new_n6809_));
  AOI21X1  g6424(.A0(new_n6809_), .A1(new_n596_), .B0(new_n599_), .Y(new_n6810_));
  OAI21X1  g6425(.A0(new_n6810_), .A1(new_n604_), .B0(new_n606_), .Y(new_n6811_));
  AOI21X1  g6426(.A0(new_n6811_), .A1(new_n611_), .B0(new_n614_), .Y(new_n6812_));
  OAI21X1  g6427(.A0(new_n6812_), .A1(new_n619_), .B0(new_n621_), .Y(new_n6813_));
  AOI21X1  g6428(.A0(new_n6813_), .A1(new_n626_), .B0(new_n629_), .Y(new_n6814_));
  OAI21X1  g6429(.A0(new_n6814_), .A1(new_n634_), .B0(new_n636_), .Y(new_n6815_));
  AOI21X1  g6430(.A0(new_n6815_), .A1(new_n641_), .B0(new_n644_), .Y(new_n6816_));
  OAI21X1  g6431(.A0(new_n6816_), .A1(new_n649_), .B0(new_n651_), .Y(new_n6817_));
  AOI21X1  g6432(.A0(new_n6817_), .A1(new_n656_), .B0(new_n659_), .Y(new_n6818_));
  OAI21X1  g6433(.A0(new_n6818_), .A1(new_n664_), .B0(new_n666_), .Y(new_n6819_));
  AOI21X1  g6434(.A0(new_n6819_), .A1(new_n671_), .B0(new_n674_), .Y(new_n6820_));
  OAI21X1  g6435(.A0(new_n6820_), .A1(new_n679_), .B0(new_n681_), .Y(new_n6821_));
  OAI21X1  g6436(.A0(new_n1002_), .A1(\priority[122] ), .B0(\req[122] ), .Y(new_n6822_));
  AOI21X1  g6437(.A0(new_n6821_), .A1(new_n686_), .B0(new_n6822_), .Y(\grant[122] ));
  NOR2X1   g6438(.A(new_n1011_), .B(new_n695_), .Y(new_n6824_));
  OAI21X1  g6439(.A0(new_n6824_), .A1(new_n1335_), .B0(new_n1438_), .Y(new_n6825_));
  AOI21X1  g6440(.A0(new_n6825_), .A1(new_n1440_), .B0(new_n1803_), .Y(new_n6826_));
  OAI21X1  g6441(.A0(new_n6826_), .A1(new_n712_), .B0(new_n714_), .Y(new_n6827_));
  AOI21X1  g6442(.A0(new_n6827_), .A1(new_n719_), .B0(new_n722_), .Y(new_n6828_));
  OAI21X1  g6443(.A0(new_n6828_), .A1(new_n727_), .B0(new_n729_), .Y(new_n6829_));
  AOI21X1  g6444(.A0(new_n6829_), .A1(new_n734_), .B0(new_n737_), .Y(new_n6830_));
  OAI21X1  g6445(.A0(new_n6830_), .A1(new_n742_), .B0(new_n744_), .Y(new_n6831_));
  AOI21X1  g6446(.A0(new_n6831_), .A1(new_n749_), .B0(new_n752_), .Y(new_n6832_));
  OAI21X1  g6447(.A0(new_n6832_), .A1(new_n757_), .B0(new_n759_), .Y(new_n6833_));
  AOI21X1  g6448(.A0(new_n6833_), .A1(new_n764_), .B0(new_n767_), .Y(new_n6834_));
  OAI21X1  g6449(.A0(new_n6834_), .A1(new_n772_), .B0(new_n774_), .Y(new_n6835_));
  AOI21X1  g6450(.A0(new_n6835_), .A1(new_n779_), .B0(new_n782_), .Y(new_n6836_));
  OAI21X1  g6451(.A0(new_n6836_), .A1(new_n787_), .B0(new_n789_), .Y(new_n6837_));
  AOI21X1  g6452(.A0(new_n6837_), .A1(new_n794_), .B0(new_n797_), .Y(new_n6838_));
  OAI21X1  g6453(.A0(new_n6838_), .A1(new_n802_), .B0(new_n804_), .Y(new_n6839_));
  AOI21X1  g6454(.A0(new_n6839_), .A1(new_n809_), .B0(new_n812_), .Y(new_n6840_));
  OAI21X1  g6455(.A0(new_n6840_), .A1(new_n817_), .B0(new_n819_), .Y(new_n6841_));
  AOI21X1  g6456(.A0(new_n6841_), .A1(new_n824_), .B0(new_n827_), .Y(new_n6842_));
  OAI21X1  g6457(.A0(new_n6842_), .A1(new_n832_), .B0(new_n834_), .Y(new_n6843_));
  AOI21X1  g6458(.A0(new_n6843_), .A1(new_n839_), .B0(new_n842_), .Y(new_n6844_));
  OAI21X1  g6459(.A0(new_n6844_), .A1(new_n847_), .B0(new_n849_), .Y(new_n6845_));
  AOI21X1  g6460(.A0(new_n6845_), .A1(new_n854_), .B0(new_n857_), .Y(new_n6846_));
  OAI21X1  g6461(.A0(new_n6846_), .A1(new_n862_), .B0(new_n864_), .Y(new_n6847_));
  AOI21X1  g6462(.A0(new_n6847_), .A1(new_n869_), .B0(new_n872_), .Y(new_n6848_));
  OAI21X1  g6463(.A0(new_n6848_), .A1(new_n877_), .B0(new_n879_), .Y(new_n6849_));
  AOI21X1  g6464(.A0(new_n6849_), .A1(new_n884_), .B0(new_n887_), .Y(new_n6850_));
  OAI21X1  g6465(.A0(new_n6850_), .A1(new_n892_), .B0(new_n894_), .Y(new_n6851_));
  AOI21X1  g6466(.A0(new_n6851_), .A1(new_n899_), .B0(new_n902_), .Y(new_n6852_));
  OAI21X1  g6467(.A0(new_n6852_), .A1(new_n907_), .B0(new_n909_), .Y(new_n6853_));
  AOI21X1  g6468(.A0(new_n6853_), .A1(new_n914_), .B0(new_n917_), .Y(new_n6854_));
  OAI21X1  g6469(.A0(new_n6854_), .A1(new_n922_), .B0(new_n924_), .Y(new_n6855_));
  AOI21X1  g6470(.A0(new_n6855_), .A1(new_n929_), .B0(new_n932_), .Y(new_n6856_));
  OAI21X1  g6471(.A0(new_n6856_), .A1(new_n937_), .B0(new_n939_), .Y(new_n6857_));
  AOI21X1  g6472(.A0(new_n6857_), .A1(new_n944_), .B0(new_n947_), .Y(new_n6858_));
  OAI21X1  g6473(.A0(new_n6858_), .A1(new_n952_), .B0(new_n954_), .Y(new_n6859_));
  AOI21X1  g6474(.A0(new_n6859_), .A1(new_n959_), .B0(new_n962_), .Y(new_n6860_));
  OAI21X1  g6475(.A0(new_n6860_), .A1(new_n967_), .B0(new_n969_), .Y(new_n6861_));
  AOI21X1  g6476(.A0(new_n6861_), .A1(new_n974_), .B0(new_n977_), .Y(new_n6862_));
  OAI21X1  g6477(.A0(new_n6862_), .A1(new_n982_), .B0(new_n984_), .Y(new_n6863_));
  AOI21X1  g6478(.A0(new_n6863_), .A1(new_n989_), .B0(new_n992_), .Y(new_n6864_));
  OAI21X1  g6479(.A0(new_n6864_), .A1(new_n997_), .B0(new_n999_), .Y(new_n6865_));
  OAI21X1  g6480(.A0(new_n1316_), .A1(\priority[123] ), .B0(\req[123] ), .Y(new_n6866_));
  AOI21X1  g6481(.A0(new_n6865_), .A1(new_n1004_), .B0(new_n6866_), .Y(\grant[123] ));
  NOR2X1   g6482(.A(new_n1325_), .B(new_n1013_), .Y(new_n6868_));
  OAI21X1  g6483(.A0(new_n6868_), .A1(new_n1444_), .B0(new_n1547_), .Y(new_n6869_));
  AOI21X1  g6484(.A0(new_n6869_), .A1(new_n1549_), .B0(new_n1848_), .Y(new_n6870_));
  OAI21X1  g6485(.A0(new_n6870_), .A1(new_n1026_), .B0(new_n1028_), .Y(new_n6871_));
  AOI21X1  g6486(.A0(new_n6871_), .A1(new_n1033_), .B0(new_n1036_), .Y(new_n6872_));
  OAI21X1  g6487(.A0(new_n6872_), .A1(new_n1041_), .B0(new_n1043_), .Y(new_n6873_));
  AOI21X1  g6488(.A0(new_n6873_), .A1(new_n1048_), .B0(new_n1051_), .Y(new_n6874_));
  OAI21X1  g6489(.A0(new_n6874_), .A1(new_n1056_), .B0(new_n1058_), .Y(new_n6875_));
  AOI21X1  g6490(.A0(new_n6875_), .A1(new_n1063_), .B0(new_n1066_), .Y(new_n6876_));
  OAI21X1  g6491(.A0(new_n6876_), .A1(new_n1071_), .B0(new_n1073_), .Y(new_n6877_));
  AOI21X1  g6492(.A0(new_n6877_), .A1(new_n1078_), .B0(new_n1081_), .Y(new_n6878_));
  OAI21X1  g6493(.A0(new_n6878_), .A1(new_n1086_), .B0(new_n1088_), .Y(new_n6879_));
  AOI21X1  g6494(.A0(new_n6879_), .A1(new_n1093_), .B0(new_n1096_), .Y(new_n6880_));
  OAI21X1  g6495(.A0(new_n6880_), .A1(new_n1101_), .B0(new_n1103_), .Y(new_n6881_));
  AOI21X1  g6496(.A0(new_n6881_), .A1(new_n1108_), .B0(new_n1111_), .Y(new_n6882_));
  OAI21X1  g6497(.A0(new_n6882_), .A1(new_n1116_), .B0(new_n1118_), .Y(new_n6883_));
  AOI21X1  g6498(.A0(new_n6883_), .A1(new_n1123_), .B0(new_n1126_), .Y(new_n6884_));
  OAI21X1  g6499(.A0(new_n6884_), .A1(new_n1131_), .B0(new_n1133_), .Y(new_n6885_));
  AOI21X1  g6500(.A0(new_n6885_), .A1(new_n1138_), .B0(new_n1141_), .Y(new_n6886_));
  OAI21X1  g6501(.A0(new_n6886_), .A1(new_n1146_), .B0(new_n1148_), .Y(new_n6887_));
  AOI21X1  g6502(.A0(new_n6887_), .A1(new_n1153_), .B0(new_n1156_), .Y(new_n6888_));
  OAI21X1  g6503(.A0(new_n6888_), .A1(new_n1161_), .B0(new_n1163_), .Y(new_n6889_));
  AOI21X1  g6504(.A0(new_n6889_), .A1(new_n1168_), .B0(new_n1171_), .Y(new_n6890_));
  OAI21X1  g6505(.A0(new_n6890_), .A1(new_n1176_), .B0(new_n1178_), .Y(new_n6891_));
  AOI21X1  g6506(.A0(new_n6891_), .A1(new_n1183_), .B0(new_n1186_), .Y(new_n6892_));
  OAI21X1  g6507(.A0(new_n6892_), .A1(new_n1191_), .B0(new_n1193_), .Y(new_n6893_));
  AOI21X1  g6508(.A0(new_n6893_), .A1(new_n1198_), .B0(new_n1201_), .Y(new_n6894_));
  OAI21X1  g6509(.A0(new_n6894_), .A1(new_n1206_), .B0(new_n1208_), .Y(new_n6895_));
  AOI21X1  g6510(.A0(new_n6895_), .A1(new_n1213_), .B0(new_n1216_), .Y(new_n6896_));
  OAI21X1  g6511(.A0(new_n6896_), .A1(new_n1221_), .B0(new_n1223_), .Y(new_n6897_));
  AOI21X1  g6512(.A0(new_n6897_), .A1(new_n1228_), .B0(new_n1231_), .Y(new_n6898_));
  OAI21X1  g6513(.A0(new_n6898_), .A1(new_n1236_), .B0(new_n1238_), .Y(new_n6899_));
  AOI21X1  g6514(.A0(new_n6899_), .A1(new_n1243_), .B0(new_n1246_), .Y(new_n6900_));
  OAI21X1  g6515(.A0(new_n6900_), .A1(new_n1251_), .B0(new_n1253_), .Y(new_n6901_));
  AOI21X1  g6516(.A0(new_n6901_), .A1(new_n1258_), .B0(new_n1261_), .Y(new_n6902_));
  OAI21X1  g6517(.A0(new_n6902_), .A1(new_n1266_), .B0(new_n1268_), .Y(new_n6903_));
  AOI21X1  g6518(.A0(new_n6903_), .A1(new_n1273_), .B0(new_n1276_), .Y(new_n6904_));
  OAI21X1  g6519(.A0(new_n6904_), .A1(new_n1281_), .B0(new_n1283_), .Y(new_n6905_));
  AOI21X1  g6520(.A0(new_n6905_), .A1(new_n1288_), .B0(new_n1291_), .Y(new_n6906_));
  OAI21X1  g6521(.A0(new_n6906_), .A1(new_n1296_), .B0(new_n1298_), .Y(new_n6907_));
  AOI21X1  g6522(.A0(new_n6907_), .A1(new_n1303_), .B0(new_n1306_), .Y(new_n6908_));
  OAI21X1  g6523(.A0(new_n6908_), .A1(new_n1311_), .B0(new_n1313_), .Y(new_n6909_));
  OAI21X1  g6524(.A0(new_n692_), .A1(\priority[124] ), .B0(\req[124] ), .Y(new_n6910_));
  AOI21X1  g6525(.A0(new_n6909_), .A1(new_n1318_), .B0(new_n6910_), .Y(\grant[124] ));
  NOR2X1   g6526(.A(new_n1327_), .B(new_n700_), .Y(new_n6912_));
  OAI21X1  g6527(.A0(new_n6912_), .A1(new_n1553_), .B0(new_n1656_), .Y(new_n6913_));
  AOI21X1  g6528(.A0(new_n6913_), .A1(new_n1552_), .B0(new_n1893_), .Y(new_n6914_));
  OAI21X1  g6529(.A0(new_n6914_), .A1(new_n1395_), .B0(new_n403_), .Y(new_n6915_));
  AOI21X1  g6530(.A0(new_n6915_), .A1(new_n1393_), .B0(new_n1394_), .Y(new_n6916_));
  OAI21X1  g6531(.A0(new_n6916_), .A1(new_n1392_), .B0(new_n418_), .Y(new_n6917_));
  AOI21X1  g6532(.A0(new_n6917_), .A1(new_n1390_), .B0(new_n1391_), .Y(new_n6918_));
  OAI21X1  g6533(.A0(new_n6918_), .A1(new_n1389_), .B0(new_n433_), .Y(new_n6919_));
  AOI21X1  g6534(.A0(new_n6919_), .A1(new_n1387_), .B0(new_n1388_), .Y(new_n6920_));
  OAI21X1  g6535(.A0(new_n6920_), .A1(new_n1386_), .B0(new_n448_), .Y(new_n6921_));
  AOI21X1  g6536(.A0(new_n6921_), .A1(new_n1384_), .B0(new_n1385_), .Y(new_n6922_));
  OAI21X1  g6537(.A0(new_n6922_), .A1(new_n1383_), .B0(new_n463_), .Y(new_n6923_));
  AOI21X1  g6538(.A0(new_n6923_), .A1(new_n1381_), .B0(new_n1382_), .Y(new_n6924_));
  OAI21X1  g6539(.A0(new_n6924_), .A1(new_n1380_), .B0(new_n478_), .Y(new_n6925_));
  AOI21X1  g6540(.A0(new_n6925_), .A1(new_n1378_), .B0(new_n1379_), .Y(new_n6926_));
  OAI21X1  g6541(.A0(new_n6926_), .A1(new_n1377_), .B0(new_n493_), .Y(new_n6927_));
  AOI21X1  g6542(.A0(new_n6927_), .A1(new_n1375_), .B0(new_n1376_), .Y(new_n6928_));
  OAI21X1  g6543(.A0(new_n6928_), .A1(new_n1374_), .B0(new_n508_), .Y(new_n6929_));
  AOI21X1  g6544(.A0(new_n6929_), .A1(new_n1372_), .B0(new_n1373_), .Y(new_n6930_));
  OAI21X1  g6545(.A0(new_n6930_), .A1(new_n1371_), .B0(new_n523_), .Y(new_n6931_));
  AOI21X1  g6546(.A0(new_n6931_), .A1(new_n1369_), .B0(new_n1370_), .Y(new_n6932_));
  OAI21X1  g6547(.A0(new_n6932_), .A1(new_n1368_), .B0(new_n538_), .Y(new_n6933_));
  AOI21X1  g6548(.A0(new_n6933_), .A1(new_n1366_), .B0(new_n1367_), .Y(new_n6934_));
  OAI21X1  g6549(.A0(new_n6934_), .A1(new_n1365_), .B0(new_n553_), .Y(new_n6935_));
  AOI21X1  g6550(.A0(new_n6935_), .A1(new_n1363_), .B0(new_n1364_), .Y(new_n6936_));
  OAI21X1  g6551(.A0(new_n6936_), .A1(new_n1362_), .B0(new_n568_), .Y(new_n6937_));
  AOI21X1  g6552(.A0(new_n6937_), .A1(new_n1360_), .B0(new_n1361_), .Y(new_n6938_));
  OAI21X1  g6553(.A0(new_n6938_), .A1(new_n1359_), .B0(new_n583_), .Y(new_n6939_));
  AOI21X1  g6554(.A0(new_n6939_), .A1(new_n1357_), .B0(new_n1358_), .Y(new_n6940_));
  OAI21X1  g6555(.A0(new_n6940_), .A1(new_n1356_), .B0(new_n598_), .Y(new_n6941_));
  AOI21X1  g6556(.A0(new_n6941_), .A1(new_n1354_), .B0(new_n1355_), .Y(new_n6942_));
  OAI21X1  g6557(.A0(new_n6942_), .A1(new_n1353_), .B0(new_n613_), .Y(new_n6943_));
  AOI21X1  g6558(.A0(new_n6943_), .A1(new_n1351_), .B0(new_n1352_), .Y(new_n6944_));
  OAI21X1  g6559(.A0(new_n6944_), .A1(new_n1350_), .B0(new_n628_), .Y(new_n6945_));
  AOI21X1  g6560(.A0(new_n6945_), .A1(new_n1348_), .B0(new_n1349_), .Y(new_n6946_));
  OAI21X1  g6561(.A0(new_n6946_), .A1(new_n1347_), .B0(new_n643_), .Y(new_n6947_));
  AOI21X1  g6562(.A0(new_n6947_), .A1(new_n1345_), .B0(new_n1346_), .Y(new_n6948_));
  OAI21X1  g6563(.A0(new_n6948_), .A1(new_n1344_), .B0(new_n658_), .Y(new_n6949_));
  AOI21X1  g6564(.A0(new_n6949_), .A1(new_n1342_), .B0(new_n1343_), .Y(new_n6950_));
  OAI21X1  g6565(.A0(new_n6950_), .A1(new_n1341_), .B0(new_n673_), .Y(new_n6951_));
  AOI21X1  g6566(.A0(new_n6951_), .A1(new_n1339_), .B0(new_n1340_), .Y(new_n6952_));
  OAI21X1  g6567(.A0(new_n6952_), .A1(new_n1338_), .B0(new_n688_), .Y(new_n6953_));
  OAI21X1  g6568(.A0(new_n1010_), .A1(\priority[125] ), .B0(\req[125] ), .Y(new_n6954_));
  AOI21X1  g6569(.A0(new_n6953_), .A1(new_n1336_), .B0(new_n6954_), .Y(\grant[125] ));
  NOR2X1   g6570(.A(new_n1437_), .B(new_n1016_), .Y(new_n6956_));
  OAI21X1  g6571(.A0(new_n6956_), .A1(new_n1661_), .B0(new_n1705_), .Y(new_n6957_));
  AOI21X1  g6572(.A0(new_n6957_), .A1(new_n1660_), .B0(new_n1938_), .Y(new_n6958_));
  OAI21X1  g6573(.A0(new_n6958_), .A1(new_n1504_), .B0(new_n721_), .Y(new_n6959_));
  AOI21X1  g6574(.A0(new_n6959_), .A1(new_n1502_), .B0(new_n1503_), .Y(new_n6960_));
  OAI21X1  g6575(.A0(new_n6960_), .A1(new_n1501_), .B0(new_n736_), .Y(new_n6961_));
  AOI21X1  g6576(.A0(new_n6961_), .A1(new_n1499_), .B0(new_n1500_), .Y(new_n6962_));
  OAI21X1  g6577(.A0(new_n6962_), .A1(new_n1498_), .B0(new_n751_), .Y(new_n6963_));
  AOI21X1  g6578(.A0(new_n6963_), .A1(new_n1496_), .B0(new_n1497_), .Y(new_n6964_));
  OAI21X1  g6579(.A0(new_n6964_), .A1(new_n1495_), .B0(new_n766_), .Y(new_n6965_));
  AOI21X1  g6580(.A0(new_n6965_), .A1(new_n1493_), .B0(new_n1494_), .Y(new_n6966_));
  OAI21X1  g6581(.A0(new_n6966_), .A1(new_n1492_), .B0(new_n781_), .Y(new_n6967_));
  AOI21X1  g6582(.A0(new_n6967_), .A1(new_n1490_), .B0(new_n1491_), .Y(new_n6968_));
  OAI21X1  g6583(.A0(new_n6968_), .A1(new_n1489_), .B0(new_n796_), .Y(new_n6969_));
  AOI21X1  g6584(.A0(new_n6969_), .A1(new_n1487_), .B0(new_n1488_), .Y(new_n6970_));
  OAI21X1  g6585(.A0(new_n6970_), .A1(new_n1486_), .B0(new_n811_), .Y(new_n6971_));
  AOI21X1  g6586(.A0(new_n6971_), .A1(new_n1484_), .B0(new_n1485_), .Y(new_n6972_));
  OAI21X1  g6587(.A0(new_n6972_), .A1(new_n1483_), .B0(new_n826_), .Y(new_n6973_));
  AOI21X1  g6588(.A0(new_n6973_), .A1(new_n1481_), .B0(new_n1482_), .Y(new_n6974_));
  OAI21X1  g6589(.A0(new_n6974_), .A1(new_n1480_), .B0(new_n841_), .Y(new_n6975_));
  AOI21X1  g6590(.A0(new_n6975_), .A1(new_n1478_), .B0(new_n1479_), .Y(new_n6976_));
  OAI21X1  g6591(.A0(new_n6976_), .A1(new_n1477_), .B0(new_n856_), .Y(new_n6977_));
  AOI21X1  g6592(.A0(new_n6977_), .A1(new_n1475_), .B0(new_n1476_), .Y(new_n6978_));
  OAI21X1  g6593(.A0(new_n6978_), .A1(new_n1474_), .B0(new_n871_), .Y(new_n6979_));
  AOI21X1  g6594(.A0(new_n6979_), .A1(new_n1472_), .B0(new_n1473_), .Y(new_n6980_));
  OAI21X1  g6595(.A0(new_n6980_), .A1(new_n1471_), .B0(new_n886_), .Y(new_n6981_));
  AOI21X1  g6596(.A0(new_n6981_), .A1(new_n1469_), .B0(new_n1470_), .Y(new_n6982_));
  OAI21X1  g6597(.A0(new_n6982_), .A1(new_n1468_), .B0(new_n901_), .Y(new_n6983_));
  AOI21X1  g6598(.A0(new_n6983_), .A1(new_n1466_), .B0(new_n1467_), .Y(new_n6984_));
  OAI21X1  g6599(.A0(new_n6984_), .A1(new_n1465_), .B0(new_n916_), .Y(new_n6985_));
  AOI21X1  g6600(.A0(new_n6985_), .A1(new_n1463_), .B0(new_n1464_), .Y(new_n6986_));
  OAI21X1  g6601(.A0(new_n6986_), .A1(new_n1462_), .B0(new_n931_), .Y(new_n6987_));
  AOI21X1  g6602(.A0(new_n6987_), .A1(new_n1460_), .B0(new_n1461_), .Y(new_n6988_));
  OAI21X1  g6603(.A0(new_n6988_), .A1(new_n1459_), .B0(new_n946_), .Y(new_n6989_));
  AOI21X1  g6604(.A0(new_n6989_), .A1(new_n1457_), .B0(new_n1458_), .Y(new_n6990_));
  OAI21X1  g6605(.A0(new_n6990_), .A1(new_n1456_), .B0(new_n961_), .Y(new_n6991_));
  AOI21X1  g6606(.A0(new_n6991_), .A1(new_n1454_), .B0(new_n1455_), .Y(new_n6992_));
  OAI21X1  g6607(.A0(new_n6992_), .A1(new_n1453_), .B0(new_n976_), .Y(new_n6993_));
  AOI21X1  g6608(.A0(new_n6993_), .A1(new_n1451_), .B0(new_n1452_), .Y(new_n6994_));
  OAI21X1  g6609(.A0(new_n6994_), .A1(new_n1450_), .B0(new_n991_), .Y(new_n6995_));
  AOI21X1  g6610(.A0(new_n6995_), .A1(new_n1448_), .B0(new_n1449_), .Y(new_n6996_));
  OAI21X1  g6611(.A0(new_n6996_), .A1(new_n1447_), .B0(new_n1006_), .Y(new_n6997_));
  OAI21X1  g6612(.A0(new_n1324_), .A1(\priority[126] ), .B0(\req[126] ), .Y(new_n6998_));
  AOI21X1  g6613(.A0(new_n6997_), .A1(new_n1445_), .B0(new_n6998_), .Y(\grant[126] ));
  NOR2X1   g6614(.A(new_n1546_), .B(new_n1330_), .Y(new_n7000_));
  OAI21X1  g6615(.A0(new_n7000_), .A1(new_n1710_), .B0(new_n1754_), .Y(new_n7001_));
  AOI21X1  g6616(.A0(new_n7001_), .A1(new_n1709_), .B0(new_n1983_), .Y(new_n7002_));
  OAI21X1  g6617(.A0(new_n7002_), .A1(new_n1613_), .B0(new_n1035_), .Y(new_n7003_));
  AOI21X1  g6618(.A0(new_n7003_), .A1(new_n1611_), .B0(new_n1612_), .Y(new_n7004_));
  OAI21X1  g6619(.A0(new_n7004_), .A1(new_n1610_), .B0(new_n1050_), .Y(new_n7005_));
  AOI21X1  g6620(.A0(new_n7005_), .A1(new_n1608_), .B0(new_n1609_), .Y(new_n7006_));
  OAI21X1  g6621(.A0(new_n7006_), .A1(new_n1607_), .B0(new_n1065_), .Y(new_n7007_));
  AOI21X1  g6622(.A0(new_n7007_), .A1(new_n1605_), .B0(new_n1606_), .Y(new_n7008_));
  OAI21X1  g6623(.A0(new_n7008_), .A1(new_n1604_), .B0(new_n1080_), .Y(new_n7009_));
  AOI21X1  g6624(.A0(new_n7009_), .A1(new_n1602_), .B0(new_n1603_), .Y(new_n7010_));
  OAI21X1  g6625(.A0(new_n7010_), .A1(new_n1601_), .B0(new_n1095_), .Y(new_n7011_));
  AOI21X1  g6626(.A0(new_n7011_), .A1(new_n1599_), .B0(new_n1600_), .Y(new_n7012_));
  OAI21X1  g6627(.A0(new_n7012_), .A1(new_n1598_), .B0(new_n1110_), .Y(new_n7013_));
  AOI21X1  g6628(.A0(new_n7013_), .A1(new_n1596_), .B0(new_n1597_), .Y(new_n7014_));
  OAI21X1  g6629(.A0(new_n7014_), .A1(new_n1595_), .B0(new_n1125_), .Y(new_n7015_));
  AOI21X1  g6630(.A0(new_n7015_), .A1(new_n1593_), .B0(new_n1594_), .Y(new_n7016_));
  OAI21X1  g6631(.A0(new_n7016_), .A1(new_n1592_), .B0(new_n1140_), .Y(new_n7017_));
  AOI21X1  g6632(.A0(new_n7017_), .A1(new_n1590_), .B0(new_n1591_), .Y(new_n7018_));
  OAI21X1  g6633(.A0(new_n7018_), .A1(new_n1589_), .B0(new_n1155_), .Y(new_n7019_));
  AOI21X1  g6634(.A0(new_n7019_), .A1(new_n1587_), .B0(new_n1588_), .Y(new_n7020_));
  OAI21X1  g6635(.A0(new_n7020_), .A1(new_n1586_), .B0(new_n1170_), .Y(new_n7021_));
  AOI21X1  g6636(.A0(new_n7021_), .A1(new_n1584_), .B0(new_n1585_), .Y(new_n7022_));
  OAI21X1  g6637(.A0(new_n7022_), .A1(new_n1583_), .B0(new_n1185_), .Y(new_n7023_));
  AOI21X1  g6638(.A0(new_n7023_), .A1(new_n1581_), .B0(new_n1582_), .Y(new_n7024_));
  OAI21X1  g6639(.A0(new_n7024_), .A1(new_n1580_), .B0(new_n1200_), .Y(new_n7025_));
  AOI21X1  g6640(.A0(new_n7025_), .A1(new_n1578_), .B0(new_n1579_), .Y(new_n7026_));
  OAI21X1  g6641(.A0(new_n7026_), .A1(new_n1577_), .B0(new_n1215_), .Y(new_n7027_));
  AOI21X1  g6642(.A0(new_n7027_), .A1(new_n1575_), .B0(new_n1576_), .Y(new_n7028_));
  OAI21X1  g6643(.A0(new_n7028_), .A1(new_n1574_), .B0(new_n1230_), .Y(new_n7029_));
  AOI21X1  g6644(.A0(new_n7029_), .A1(new_n1572_), .B0(new_n1573_), .Y(new_n7030_));
  OAI21X1  g6645(.A0(new_n7030_), .A1(new_n1571_), .B0(new_n1245_), .Y(new_n7031_));
  AOI21X1  g6646(.A0(new_n7031_), .A1(new_n1569_), .B0(new_n1570_), .Y(new_n7032_));
  OAI21X1  g6647(.A0(new_n7032_), .A1(new_n1568_), .B0(new_n1260_), .Y(new_n7033_));
  AOI21X1  g6648(.A0(new_n7033_), .A1(new_n1566_), .B0(new_n1567_), .Y(new_n7034_));
  OAI21X1  g6649(.A0(new_n7034_), .A1(new_n1565_), .B0(new_n1275_), .Y(new_n7035_));
  AOI21X1  g6650(.A0(new_n7035_), .A1(new_n1563_), .B0(new_n1564_), .Y(new_n7036_));
  OAI21X1  g6651(.A0(new_n7036_), .A1(new_n1562_), .B0(new_n1290_), .Y(new_n7037_));
  AOI21X1  g6652(.A0(new_n7037_), .A1(new_n1560_), .B0(new_n1561_), .Y(new_n7038_));
  OAI21X1  g6653(.A0(new_n7038_), .A1(new_n1559_), .B0(new_n1305_), .Y(new_n7039_));
  AOI21X1  g6654(.A0(new_n7039_), .A1(new_n1557_), .B0(new_n1558_), .Y(new_n7040_));
  OAI21X1  g6655(.A0(new_n7040_), .A1(new_n1556_), .B0(new_n1320_), .Y(new_n7041_));
  OAI21X1  g6656(.A0(new_n699_), .A1(\priority[127] ), .B0(\req[127] ), .Y(new_n7042_));
  AOI21X1  g6657(.A0(new_n7041_), .A1(new_n1554_), .B0(new_n7042_), .Y(\grant[127] ));
  OR4X1    g6658(.A(\req[123] ), .B(\req[122] ), .C(\req[7] ), .D(\req[6] ), .Y(new_n7044_));
  OR4X1    g6659(.A(\req[19] ), .B(\req[18] ), .C(\req[13] ), .D(\req[12] ), .Y(new_n7045_));
  OR4X1    g6660(.A(\req[105] ), .B(\req[104] ), .C(\req[99] ), .D(\req[98] ), .Y(new_n7046_));
  OR4X1    g6661(.A(\req[117] ), .B(\req[116] ), .C(\req[111] ), .D(\req[110] ), .Y(new_n7047_));
  OR4X1    g6662(.A(new_n7047_), .B(new_n7046_), .C(new_n7045_), .D(new_n7044_), .Y(new_n7048_));
  OR4X1    g6663(.A(\req[55] ), .B(\req[54] ), .C(\req[49] ), .D(\req[48] ), .Y(new_n7049_));
  OR4X1    g6664(.A(\req[67] ), .B(\req[66] ), .C(\req[61] ), .D(\req[60] ), .Y(new_n7050_));
  OR4X1    g6665(.A(\req[31] ), .B(\req[30] ), .C(\req[25] ), .D(\req[24] ), .Y(new_n7051_));
  OR4X1    g6666(.A(\req[43] ), .B(\req[42] ), .C(\req[37] ), .D(\req[36] ), .Y(new_n7052_));
  OR4X1    g6667(.A(new_n7052_), .B(new_n7051_), .C(new_n7050_), .D(new_n7049_), .Y(new_n7053_));
  OR4X1    g6668(.A(\req[33] ), .B(\req[32] ), .C(\req[27] ), .D(\req[26] ), .Y(new_n7054_));
  OR4X1    g6669(.A(\req[45] ), .B(\req[44] ), .C(\req[39] ), .D(\req[38] ), .Y(new_n7055_));
  OR4X1    g6670(.A(\req[9] ), .B(\req[8] ), .C(\req[3] ), .D(\req[2] ), .Y(new_n7056_));
  OR4X1    g6671(.A(\req[21] ), .B(\req[20] ), .C(\req[15] ), .D(\req[14] ), .Y(new_n7057_));
  OR4X1    g6672(.A(new_n7057_), .B(new_n7056_), .C(new_n7055_), .D(new_n7054_), .Y(new_n7058_));
  OR4X1    g6673(.A(\req[81] ), .B(\req[80] ), .C(\req[75] ), .D(\req[74] ), .Y(new_n7059_));
  OR4X1    g6674(.A(\req[93] ), .B(\req[92] ), .C(\req[87] ), .D(\req[86] ), .Y(new_n7060_));
  OR4X1    g6675(.A(\req[57] ), .B(\req[56] ), .C(\req[51] ), .D(\req[50] ), .Y(new_n7061_));
  OR4X1    g6676(.A(\req[69] ), .B(\req[68] ), .C(\req[63] ), .D(\req[62] ), .Y(new_n7062_));
  OR4X1    g6677(.A(new_n7062_), .B(new_n7061_), .C(new_n7060_), .D(new_n7059_), .Y(new_n7063_));
  OR4X1    g6678(.A(new_n7063_), .B(new_n7058_), .C(new_n7053_), .D(new_n7048_), .Y(new_n7064_));
  OR4X1    g6679(.A(\req[71] ), .B(\req[70] ), .C(\req[65] ), .D(\req[64] ), .Y(new_n7065_));
  OR4X1    g6680(.A(\req[83] ), .B(\req[82] ), .C(\req[77] ), .D(\req[76] ), .Y(new_n7066_));
  OR4X1    g6681(.A(\req[47] ), .B(\req[46] ), .C(\req[41] ), .D(\req[40] ), .Y(new_n7067_));
  OR4X1    g6682(.A(\req[59] ), .B(\req[58] ), .C(\req[53] ), .D(\req[52] ), .Y(new_n7068_));
  OR4X1    g6683(.A(new_n7068_), .B(new_n7067_), .C(new_n7066_), .D(new_n7065_), .Y(new_n7069_));
  OR4X1    g6684(.A(\req[119] ), .B(\req[118] ), .C(\req[113] ), .D(\req[112] ), .Y(new_n7070_));
  OR4X1    g6685(.A(\req[125] ), .B(\req[124] ), .C(\req[1] ), .D(\req[0] ), .Y(new_n7071_));
  OR4X1    g6686(.A(\req[95] ), .B(\req[94] ), .C(\req[89] ), .D(\req[88] ), .Y(new_n7072_));
  OR4X1    g6687(.A(\req[107] ), .B(\req[106] ), .C(\req[101] ), .D(\req[100] ), .Y(new_n7073_));
  OR4X1    g6688(.A(new_n7073_), .B(new_n7072_), .C(new_n7071_), .D(new_n7070_), .Y(new_n7074_));
  OR4X1    g6689(.A(\req[103] ), .B(\req[102] ), .C(\req[97] ), .D(\req[96] ), .Y(new_n7075_));
  OR4X1    g6690(.A(\req[115] ), .B(\req[114] ), .C(\req[109] ), .D(\req[108] ), .Y(new_n7076_));
  OR4X1    g6691(.A(\req[79] ), .B(\req[78] ), .C(\req[73] ), .D(\req[72] ), .Y(new_n7077_));
  OR4X1    g6692(.A(\req[91] ), .B(\req[90] ), .C(\req[85] ), .D(\req[84] ), .Y(new_n7078_));
  OR4X1    g6693(.A(new_n7078_), .B(new_n7077_), .C(new_n7076_), .D(new_n7075_), .Y(new_n7079_));
  OR4X1    g6694(.A(\req[23] ), .B(\req[22] ), .C(\req[17] ), .D(\req[16] ), .Y(new_n7080_));
  OR4X1    g6695(.A(\req[35] ), .B(\req[34] ), .C(\req[29] ), .D(\req[28] ), .Y(new_n7081_));
  OR4X1    g6696(.A(new_n1034_), .B(new_n1021_), .C(new_n1013_), .D(new_n998_), .Y(new_n7082_));
  OR4X1    g6697(.A(new_n7082_), .B(new_n7081_), .C(new_n7080_), .D(new_n7079_), .Y(new_n7083_));
  OR4X1    g6698(.A(new_n7083_), .B(new_n7074_), .C(new_n7069_), .D(new_n7064_), .Y(anyGrant));
endmodule


