//Converted to Combinational (Partial output: n78) , Module name: s510_n78
module s510_n78 ( cnt44, st_4, st_0, st_5, st_3, cnt261, st_1, cnt45, st_2, cnt509, cnt10, cnt283, cnt21, cnt511, cnt567, john, cnt272, cnt591, cnt284, pcnt6, n78 );
input cnt44, st_4, st_0, st_5, st_3, cnt261, st_1, cnt45, st_2, cnt509, cnt10, cnt283, cnt21, cnt511, cnt567, john, cnt272, cnt591, cnt284, pcnt6;
output n78;
wire n187, n168, n173, n181, n186, n79, n183, n161, n167, n88, n169, n172, n180, n175, n176, n179, n185, n80, n121, n184, n182, n151, n143, n160, n53_1, n166, n163, n164, n165, n141, n171, n155, n157, n84, n64, n174, n148, n177, n178, n48, n66, n51, n98, n162, n44, n170, n69;
NAND4X1  g144(.A(n181), .B(n173), .C(n168), .D(n187), .Y(n78));
AOI22X1  g143(.A0(n183), .A1(cnt44), .B0(n79), .B1(n186), .Y(n187));
OAI21X1  g124(.A0(n167), .A1(n161), .B0(st_4), .Y(n168));
OAI21X1  g129(.A0(n172), .A1(n169), .B0(n88), .Y(n173));
NOR4X1   g137(.A(n179), .B(n176), .C(n175), .D(n180), .Y(n181));
OAI22X1  g142(.A0(n184), .A1(n121), .B0(n80), .B1(n185), .Y(n186));
INVX1    g035(.A(st_0), .Y(n79));
OAI21X1  g139(.A0(n151), .A1(st_4), .B0(n182), .Y(n183));
NOR4X1   g117(.A(st_0), .B(n53_1), .C(n160), .D(n143), .Y(n161));
NAND4X1  g123(.A(n165), .B(n164), .C(n163), .D(n166), .Y(n167));
NOR2X1   g044(.A(st_4), .B(st_5), .Y(n88));
NOR4X1   g125(.A(st_0), .B(n53_1), .C(n141), .D(n143), .Y(n169));
OAI21X1  g128(.A0(n157), .A1(n155), .B0(n171), .Y(n172));
NOR4X1   g136(.A(n64), .B(n79), .C(st_4), .D(n84), .Y(n180));
NOR4X1   g131(.A(n143), .B(st_0), .C(st_3), .D(n174), .Y(n175));
NOR4X1   g132(.A(n79), .B(st_1), .C(cnt261), .D(n148), .Y(n176));
AND2X1   g135(.A(n178), .B(n177), .Y(n179));
NAND3X1  g141(.A(n66), .B(n48), .C(cnt45), .Y(n185));
AOI21X1  g036(.A0(st_3), .A1(st_4), .B0(st_5), .Y(n80));
NAND3X1  g077(.A(n66), .B(st_2), .C(st_3), .Y(n121));
NAND2X1  g140(.A(st_5), .B(cnt509), .Y(n184));
NAND4X1  g138(.A(st_1), .B(n48), .C(st_5), .D(n79), .Y(n182));
NAND4X1  g107(.A(st_1), .B(n48), .C(n53_1), .D(n79), .Y(n151));
NAND2X1  g099(.A(st_1), .B(st_2), .Y(n143));
INVX1    g116(.A(cnt10), .Y(n160));
INVX1    g009(.A(st_3), .Y(n53_1));
NAND3X1  g122(.A(n98), .B(n51), .C(cnt283), .Y(n166));
NAND4X1  g119(.A(n66), .B(st_2), .C(st_3), .D(n162), .Y(n163));
NAND3X1  g120(.A(n98), .B(n53_1), .C(cnt21), .Y(n164));
NAND4X1  g121(.A(st_2), .B(n53_1), .C(cnt45), .D(n44), .Y(n165));
INVX1    g097(.A(cnt511), .Y(n141));
OR4X1    g127(.A(n69), .B(n48), .C(st_3), .D(n170), .Y(n171));
INVX1    g111(.A(cnt567), .Y(n155));
NAND2X1  g113(.A(n98), .B(n51), .Y(n157));
XOR2X1   g040(.A(st_1), .B(st_2), .Y(n84));
OR2X1    g020(.A(st_3), .B(st_5), .Y(n64));
AOI22X1  g130(.A0(st_5), .A1(cnt10), .B0(john), .B1(st_4), .Y(n174));
NAND3X1  g104(.A(st_2), .B(n53_1), .C(st_5), .Y(n148));
MX2X1    g133(.A(cnt591), .B(cnt272), .S0(st_2), .Y(n177));
NOR4X1   g134(.A(n53_1), .B(st_4), .C(st_5), .D(n69), .Y(n178));
INVX1    g004(.A(st_2), .Y(n48));
INVX1    g022(.A(st_1), .Y(n66));
AND2X1   g007(.A(st_1), .B(st_3), .Y(n51));
NOR2X1   g054(.A(st_0), .B(st_2), .Y(n98));
OR2X1    g118(.A(st_0), .B(cnt21), .Y(n162));
NOR2X1   g000(.A(st_0), .B(st_1), .Y(n44));
NAND2X1  g126(.A(pcnt6), .B(cnt284), .Y(n170));
OR2X1    g025(.A(st_0), .B(st_1), .Y(n69));

endmodule
