//Converted to Combinational , Module name: s5378 , Timestamp: 2018-12-03T15:51:02.717824 
module s5378 ( n3065gat, n3066gat, n3067gat, n3068gat, n3069gat, n3070gat, n3071gat, n3072gat, n3073gat, n3074gat, n3075gat, n3076gat, n3077gat, n3078gat, n3079gat, n3080gat, n3081gat, n3082gat, n3083gat, n3084gat, n3085gat, n3086gat, n3087gat, n3088gat, n3089gat, n3090gat, n3091gat, n3092gat, n3093gat, n3094gat, n3095gat, n3097gat, n3098gat, n3099gat, n3100gat, n673gat, n398gat, n402gat, n919gat, n846gat, n394gat, n703gat, n722gat, n726gat, n2510gat, n271gat, n160gat, n337gat, n842gat, n341gat, n2522gat, n2472gat, n2319gat, n1821gat, n1825gat, n2029gat, n1829gat, n283gat, n165gat, n279gat, n1026gat, n275gat, n2476gat, n1068gat, n957gat, n861gat, n1294gat, n1241gat, n1298gat, n865gat, n1080gat, n1148gat, n2468gat, n618gat, n491gat, n622gat, n626gat, n834gat, n707gat, n838gat, n830gat, n614gat, n2526gat, n680gat, n816gat, n580gat, n824gat, n820gat, n883gat, n584gat, n684gat, n699gat, n2464gat, n2399gat, n2343gat, n2203gat, n2562gat, n2207gat, n2626gat, n2490gat, n2622gat, n2630gat, n2543gat, n2102gat, n1880gat, n1763gat, n2155gat, n1035gat, n1121gat, n1072gat, n1282gat, n1226gat, n931gat, n1135gat, n1045gat, n1197gat, n2518gat, n667gat, n659gat, n553gat, n777gat, n561gat, n366gat, n322gat, n318gat, n314gat, n2599gat, n2588gat, n2640gat, n2658gat, n2495gat, n2390gat, n2270gat, n2339gat, n2502gat, n2634gat, n2506gat, n1834gat, n1767gat, n2084gat, n2143gat, n2061gat, n2139gat, n1899gat, n1850gat, n2403gat, n2394gat, n2440gat, n2407gat, n2347gat, n1389gat, n2021gat, n1394gat, n1496gat, n2091gat, n1332gat, n1740gat, n2179gat, n2190gat, n2135gat, n2262gat, n2182gat, n1433gat, n1316gat, n1363gat, n1312gat, n1775gat, n1871gat, n2592gat, n1508gat, n1678gat, n2309gat, n2450gat, n2446gat, n2095gat, n2176gat, n2169gat, n2454gat, n2040gat, n2044gat, n2037gat, n2025gat, n2099gat, n2266gat, n2033gat, n2110gat, n2125gat, n2121gat, n2117gat, n1975gat, n2644gat, n156gat, n152gat, n331gat, n388gat, n463gat, n327gat, n384gat, n256gat, n470gat, n148gat, n2458gat, n2514gat, n1771gat, n1336gat, n1748gat, n1675gat, n1807gat, n1340gat, n1456gat, n1525gat, n1462gat, n1596gat, n1588gat, n3104gat, n3105gat, n3106gat, n3107gat, n3108gat, n3109gat, n3110gat, n3111gat, n3112gat, n3113gat, n3114gat, n3115gat, n3116gat, n3117gat, n3118gat, n3119gat, n3120gat, n3121gat, n3122gat, n3123gat, n3124gat, n3125gat, n3126gat, n3127gat, n3128gat, n3129gat, n3130gat, n3131gat, n3132gat, n3133gat, n3134gat, n3135gat, n3136gat, n3137gat, n3138gat, n3139gat, n3140gat, n3141gat, n3142gat, n3143gat, n3144gat, n3145gat, n3146gat, n3147gat, n3148gat, n3149gat, n3150gat, n3151gat, n3152gat, n169, n174, n179, n184, n189, n193, n197, n201, n205, n210, n215, n220, n225, n230, n235, n240, n245, n250, n255, n259, n264, n269, n273, n277, n281, n285, n289, n294, n299, n304, n309, n319, n323, n328, n333, n338, n343, n347, n351, n355, n359, n364, n369, n374, n379, n384, n389, n394, n399, n404, n409, n414, n419, n424, n429, n434, n439, n444, n449, n454, n459, n464, n469, n474, n479, n484, n489, n494, n499, n504, n509, n514, n519, n524, n529, n534, n539, n544, n549, n554, n559, n564, n569, n574, n579, n584, n589, n594, n599, n604, n609, n614, n619, n624, n629, n634, n639, n644, n649, n654, n659, n664, n669, n674, n679, n684, n689, n694, n699, n704, n709, n714, n719, n724, n729, n734, n739, n744, n749, n754, n759, n764, n769, n774, n779, n784, n789, n794, n799, n804, n809, n814, n819, n824, n829, n834, n839, n844, n849, n854, n859, n864, n869, n874, n879, n884, n889, n894, n899, n904, n909, n914, n919, n924, n929, n934, n939, n944, n949, n954, n959, n964, n969, n974, n979, n984, n989, n994, n999, n1004, n1009, n1014, n1019, n1024, n1029, n1034, n1039, n1044 );
input n3065gat, n3066gat, n3067gat, n3068gat, n3069gat, n3070gat, n3071gat, n3072gat, n3073gat, n3074gat, n3075gat, n3076gat, n3077gat, n3078gat, n3079gat, n3080gat, n3081gat, n3082gat, n3083gat, n3084gat, n3085gat, n3086gat, n3087gat, n3088gat, n3089gat, n3090gat, n3091gat, n3092gat, n3093gat, n3094gat, n3095gat, n3097gat, n3098gat, n3099gat, n3100gat, n673gat, n398gat, n402gat, n919gat, n846gat, n394gat, n703gat, n722gat, n726gat, n2510gat, n271gat, n160gat, n337gat, n842gat, n341gat, n2522gat, n2472gat, n2319gat, n1821gat, n1825gat, n2029gat, n1829gat, n283gat, n165gat, n279gat, n1026gat, n275gat, n2476gat, n1068gat, n957gat, n861gat, n1294gat, n1241gat, n1298gat, n865gat, n1080gat, n1148gat, n2468gat, n618gat, n491gat, n622gat, n626gat, n834gat, n707gat, n838gat, n830gat, n614gat, n2526gat, n680gat, n816gat, n580gat, n824gat, n820gat, n883gat, n584gat, n684gat, n699gat, n2464gat, n2399gat, n2343gat, n2203gat, n2562gat, n2207gat, n2626gat, n2490gat, n2622gat, n2630gat, n2543gat, n2102gat, n1880gat, n1763gat, n2155gat, n1035gat, n1121gat, n1072gat, n1282gat, n1226gat, n931gat, n1135gat, n1045gat, n1197gat, n2518gat, n667gat, n659gat, n553gat, n777gat, n561gat, n366gat, n322gat, n318gat, n314gat, n2599gat, n2588gat, n2640gat, n2658gat, n2495gat, n2390gat, n2270gat, n2339gat, n2502gat, n2634gat, n2506gat, n1834gat, n1767gat, n2084gat, n2143gat, n2061gat, n2139gat, n1899gat, n1850gat, n2403gat, n2394gat, n2440gat, n2407gat, n2347gat, n1389gat, n2021gat, n1394gat, n1496gat, n2091gat, n1332gat, n1740gat, n2179gat, n2190gat, n2135gat, n2262gat, n2182gat, n1433gat, n1316gat, n1363gat, n1312gat, n1775gat, n1871gat, n2592gat, n1508gat, n1678gat, n2309gat, n2450gat, n2446gat, n2095gat, n2176gat, n2169gat, n2454gat, n2040gat, n2044gat, n2037gat, n2025gat, n2099gat, n2266gat, n2033gat, n2110gat, n2125gat, n2121gat, n2117gat, n1975gat, n2644gat, n156gat, n152gat, n331gat, n388gat, n463gat, n327gat, n384gat, n256gat, n470gat, n148gat, n2458gat, n2514gat, n1771gat, n1336gat, n1748gat, n1675gat, n1807gat, n1340gat, n1456gat, n1525gat, n1462gat, n1596gat, n1588gat;
output n3104gat, n3105gat, n3106gat, n3107gat, n3108gat, n3109gat, n3110gat, n3111gat, n3112gat, n3113gat, n3114gat, n3115gat, n3116gat, n3117gat, n3118gat, n3119gat, n3120gat, n3121gat, n3122gat, n3123gat, n3124gat, n3125gat, n3126gat, n3127gat, n3128gat, n3129gat, n3130gat, n3131gat, n3132gat, n3133gat, n3134gat, n3135gat, n3136gat, n3137gat, n3138gat, n3139gat, n3140gat, n3141gat, n3142gat, n3143gat, n3144gat, n3145gat, n3146gat, n3147gat, n3148gat, n3149gat, n3150gat, n3151gat, n3152gat, n169, n174, n179, n184, n189, n193, n197, n201, n205, n210, n215, n220, n225, n230, n235, n240, n245, n250, n255, n259, n264, n269, n273, n277, n281, n285, n289, n294, n299, n304, n309, n319, n323, n328, n333, n338, n343, n347, n351, n355, n359, n364, n369, n374, n379, n384, n389, n394, n399, n404, n409, n414, n419, n424, n429, n434, n439, n444, n449, n454, n459, n464, n469, n474, n479, n484, n489, n494, n499, n504, n509, n514, n519, n524, n529, n534, n539, n544, n549, n554, n559, n564, n569, n574, n579, n584, n589, n594, n599, n604, n609, n614, n619, n624, n629, n634, n639, n644, n649, n654, n659, n664, n669, n674, n679, n684, n689, n694, n699, n704, n709, n714, n719, n724, n729, n734, n739, n744, n749, n754, n759, n764, n769, n774, n779, n784, n789, n794, n799, n804, n809, n814, n819, n824, n829, n834, n839, n844, n849, n854, n859, n864, n869, n874, n879, n884, n889, n894, n899, n904, n909, n914, n919, n924, n929, n934, n939, n944, n949, n954, n959, n964, n969, n974, n979, n984, n989, n994, n999, n1004, n1009, n1014, n1019, n1024, n1029, n1034, n1039, n1044;
wire n314, n621, n622, n624_1, n625, n626, n627, n628, n629_1, n630, n631, n632, n633, n634_1, n635, n636, n637, n638, n639_1, n641, n642, n643, n644_1, n645, n646, n647, n648, n649_1, n650, n651, n652, n653, n655, n657, n658, n660, n661, n662, n663, n664_1, n665, n667, n671, n672, n676, n677, n678, n679_1, n680, n681, n682, n683, n684_1, n685, n686, n687, n688, n689_1, n690, n691, n692, n693, n694_1, n695, n696, n697, n698, n699_1, n701, n702, n703, n704_1, n705, n706, n707, n708, n709_1, n710, n711, n712, n713, n714_1, n715, n716, n717, n718, n719_1, n720, n721, n722, n723, n724_1, n725, n726, n727, n728, n729_1, n730, n731, n732, n733, n734_1, n735, n736, n737, n738, n741, n742, n743, n744_1, n745, n746, n747, n748, n749_1, n750, n751, n752, n753, n754_1, n755, n756, n757, n758, n759_1, n760, n761, n762, n763, n764_1, n765, n766, n767, n768, n769_1, n770, n771, n772, n773, n774_1, n775, n776, n779_1, n780, n781, n782, n783, n784_1, n785, n786, n787, n788, n789_1, n790, n791, n792, n793, n794_1, n795, n796, n797, n798, n799_1, n800, n801, n802, n803, n804_1, n805, n806, n807, n808, n809_1, n810, n811, n812, n815, n816, n817, n818, n819_1, n820, n821, n822, n823, n824_1, n825, n826, n827, n828, n829_1, n830, n831, n832, n833, n834_1, n835, n836, n837, n838, n839_1, n840, n841, n842, n843, n844_1, n845, n846, n847, n848, n849_1, n850, n854_1, n855, n856, n857, n858, n859_1, n860, n861, n862, n864_1, n865, n866, n867, n868, n869_1, n872, n874_1, n875, n876, n877, n878, n879_1, n880, n881, n882, n883, n886, n887, n888, n889_1, n892, n894_1, n895, n896, n897, n898, n900, n901, n902, n903, n904_1, n905, n906, n907, n909_1, n910, n911, n912, n913, n914_1, n915, n916, n917, n918, n919_1, n920, n923, n924_1, n925, n926, n927, n928, n929_1, n930, n931, n932, n933, n934_1, n935, n936, n937, n938, n939_1, n940, n941, n942, n943, n944_1, n945, n948, n949_1, n950, n951, n952, n953, n954_1, n955, n956, n959_1, n960, n961, n962, n963, n964_1, n965, n966, n968, n973, n974_1, n975, n976, n977, n978, n979_1, n980, n981, n982, n983, n984_1, n985, n987, n988, n990, n991, n993, n994_1, n996, n997, n999_1, n1000, n1002, n1003, n1005, n1006, n1008, n1009_1, n1011, n1012, n1013, n1014_1, n1015, n1016, n1017, n1019_1, n1020, n1022, n1023, n1026, n1027, n1028, n1029_1, n1030, n1031, n1032, n1033, n1034_1, n1036, n1037, n1040, n1041, n1042, n1043, n1044_1, n1045, n1046, n1047, n1049, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1077, n1078, n1079, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1089, n1090, n1091, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1151, n1153, n1154, n1155, n1156, n1159, n1161, n1162, n1163, n1164, n1167, n1168, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1182, n1185, n1186, n1190, n1192, n1193, n1196, n1197, n1201, n1204, n1205, n1207, n1208, n1210, n1211, n1213, n1214, n1216, n1217, n1219, n1220, n1222, n1223, n1225, n1226, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1245, n1246, n1247, n1248, n1249, n1251, n1253, n1254, n1256, n1258, n1259, n1260, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1273, n1274, n1275, n1276, n1277, n1279, n1280, n1283, n1284, n1285, n1287, n1288, n1289, n1290, n1291, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1305, n1306, n1307, n1308, n1309, n1310, n1312, n1314, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1335, n1341, n1342, n1344, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1365, n1366, n1367, n1369, n1370, n1372, n1374, n1376, n1378, n1380, n1382, n1384, n1386, n1387, n1388, n1390, n1391, n1392, n1394, n1395, n1396, n1400, n1401, n1402, n1406, n1407, n1408, n1409, n1411, n1412, n1414, n1415, n1416, n1419, n1424, n1425, n1426, n1427, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1472, n1473, n1475, n1476, n1493, n1496;
INVX1    g000(.A(n3087gat), .Y(n621));
INVX1    g001(.A(n3095gat), .Y(n622));
INVX1    g002(.A(n1871gat), .Y(n3106gat));
OR2X1    g003(.A(n3085gat), .B(n3083gat), .Y(n624_1));
NOR4X1   g004(.A(n3106gat), .B(n622), .C(n3084gat), .D(n624_1), .Y(n625));
INVX1    g005(.A(n625), .Y(n626));
NOR4X1   g006(.A(n3088gat), .B(n621), .C(n3086gat), .D(n626), .Y(n627));
NAND2X1  g007(.A(n627), .B(n3094gat), .Y(n628));
NOR4X1   g008(.A(n2139gat), .B(n2061gat), .C(n2143gat), .D(n1899gat), .Y(n629_1));
XOR2X1   g009(.A(n629_1), .B(n1850gat), .Y(n630));
INVX1    g010(.A(n3086gat), .Y(n631));
INVX1    g011(.A(n3093gat), .Y(n632));
NOR4X1   g012(.A(n632), .B(n3084gat), .C(n3083gat), .D(n3106gat), .Y(n633));
INVX1    g013(.A(n633), .Y(n634_1));
NAND2X1  g014(.A(n3088gat), .B(n621), .Y(n635));
NOR4X1   g015(.A(n634_1), .B(n631), .C(n3085gat), .D(n635), .Y(n636));
NOR2X1   g016(.A(n3092gat), .B(n3091gat), .Y(n637));
INVX1    g017(.A(n637), .Y(n638));
NAND2X1  g018(.A(n638), .B(n636), .Y(n639_1));
NAND3X1  g019(.A(n639_1), .B(n630), .C(n628), .Y(n3104gat));
INVX1    g020(.A(n3094gat), .Y(n641));
INVX1    g021(.A(n3088gat), .Y(n642));
NAND4X1  g022(.A(n642), .B(n621), .C(n3086gat), .D(n625), .Y(n643));
INVX1    g023(.A(n2143gat), .Y(n644_1));
NOR4X1   g024(.A(n2139gat), .B(n2061gat), .C(n644_1), .D(n1899gat), .Y(n645));
INVX1    g025(.A(n2061gat), .Y(n646));
NOR2X1   g026(.A(n1899gat), .B(n2139gat), .Y(n647));
AOI21X1  g027(.A0(n647), .A1(n646), .B0(n2143gat), .Y(n648));
NOR2X1   g028(.A(n648), .B(n645), .Y(n649_1));
INVX1    g029(.A(n3085gat), .Y(n650));
NOR4X1   g030(.A(n3087gat), .B(n3086gat), .C(n650), .D(n642), .Y(n651));
NAND3X1  g031(.A(n651), .B(n638), .C(n633), .Y(n652));
AND2X1   g032(.A(n652), .B(n649_1), .Y(n653));
OAI21X1  g033(.A0(n643), .A1(n641), .B0(n653), .Y(n3105gat));
AND2X1   g034(.A(n1771gat), .B(n1775gat), .Y(n655));
NOR2X1   g035(.A(n655), .B(n3106gat), .Y(n3107gat));
NOR4X1   g036(.A(n2440gat), .B(n2394gat), .C(n2403gat), .D(n2347gat), .Y(n657));
XOR2X1   g037(.A(n657), .B(n2407gat), .Y(n658));
NAND2X1  g038(.A(n658), .B(n1035gat), .Y(n3108gat));
INVX1    g039(.A(n2347gat), .Y(n660));
NOR4X1   g040(.A(n2440gat), .B(n2394gat), .C(n2403gat), .D(n660), .Y(n661));
INVX1    g041(.A(n2403gat), .Y(n662));
NOR2X1   g042(.A(n2440gat), .B(n2394gat), .Y(n663));
AOI21X1  g043(.A0(n663), .A1(n662), .B0(n2347gat), .Y(n664_1));
NOR2X1   g044(.A(n664_1), .B(n661), .Y(n665));
NAND2X1  g045(.A(n665), .B(n1072gat), .Y(n3109gat));
XOR2X1   g046(.A(n663), .B(n2403gat), .Y(n667));
NAND2X1  g047(.A(n667), .B(n1121gat), .Y(n3110gat));
NAND3X1  g048(.A(n2440gat), .B(n2394gat), .C(n931gat), .Y(n3111gat));
ONE      g049(.Y(n3112gat));
NOR2X1   g050(.A(n2262gat), .B(n2190gat), .Y(n671));
XOR2X1   g051(.A(n671), .B(n2135gat), .Y(n672));
NAND2X1  g052(.A(n672), .B(n1135gat), .Y(n3113gat));
NAND3X1  g053(.A(n2262gat), .B(n2190gat), .C(n1282gat), .Y(n3114gat));
ONE      g054(.Y(n3115gat));
INVX1    g055(.A(n1035gat), .Y(n676));
INVX1    g056(.A(n1121gat), .Y(n677));
NOR3X1   g057(.A(n1072gat), .B(n677), .C(n676), .Y(n678));
INVX1    g058(.A(n1072gat), .Y(n679_1));
NOR3X1   g059(.A(n679_1), .B(n677), .C(n1035gat), .Y(n680));
NOR3X1   g060(.A(n679_1), .B(n1121gat), .C(n676), .Y(n681));
NOR3X1   g061(.A(n1072gat), .B(n1121gat), .C(n1035gat), .Y(n682));
NOR4X1   g062(.A(n681), .B(n680), .C(n678), .D(n682), .Y(n683));
INVX1    g063(.A(n683), .Y(n684_1));
INVX1    g064(.A(n931gat), .Y(n685));
INVX1    g065(.A(n1135gat), .Y(n686));
NOR3X1   g066(.A(n1045gat), .B(n686), .C(n685), .Y(n687));
INVX1    g067(.A(n1045gat), .Y(n688));
NOR3X1   g068(.A(n688), .B(n686), .C(n931gat), .Y(n689_1));
NOR3X1   g069(.A(n688), .B(n1135gat), .C(n685), .Y(n690));
NOR3X1   g070(.A(n1045gat), .B(n1135gat), .C(n931gat), .Y(n691));
NOR4X1   g071(.A(n690), .B(n689_1), .C(n687), .D(n691), .Y(n692));
XOR2X1   g072(.A(n1226gat), .B(n1282gat), .Y(n693));
INVX1    g073(.A(n693), .Y(n694_1));
NOR3X1   g074(.A(n694_1), .B(n692), .C(n684_1), .Y(n695));
INVX1    g075(.A(n692), .Y(n696));
NOR3X1   g076(.A(n694_1), .B(n696), .C(n683), .Y(n697));
NOR3X1   g077(.A(n693), .B(n696), .C(n684_1), .Y(n698));
NOR3X1   g078(.A(n693), .B(n692), .C(n683), .Y(n699_1));
OR4X1    g079(.A(n698), .B(n697), .C(n695), .D(n699_1), .Y(n3116gat));
INVX1    g080(.A(n1068gat), .Y(n701));
INVX1    g081(.A(n680gat), .Y(n702));
AOI22X1  g082(.A0(n3093gat), .A1(n3087gat), .B0(n3088gat), .B1(n3095gat), .Y(n703));
AOI22X1  g083(.A0(n3093gat), .A1(n3086gat), .B0(n3087gat), .B1(n3095gat), .Y(n704_1));
INVX1    g084(.A(n704_1), .Y(n705));
AOI22X1  g085(.A0(n3093gat), .A1(n3085gat), .B0(n3086gat), .B1(n3095gat), .Y(n706));
NOR3X1   g086(.A(n706), .B(n705), .C(n703), .Y(n707));
INVX1    g087(.A(n706), .Y(n708));
NOR3X1   g088(.A(n708), .B(n704_1), .C(n703), .Y(n709_1));
AOI22X1  g089(.A0(n707), .A1(n702), .B0(n701), .B1(n709_1), .Y(n710));
INVX1    g090(.A(n271gat), .Y(n711));
INVX1    g091(.A(n659gat), .Y(n712));
INVX1    g092(.A(n703), .Y(n713));
NOR3X1   g093(.A(n706), .B(n704_1), .C(n713), .Y(n714_1));
NOR3X1   g094(.A(n706), .B(n704_1), .C(n703), .Y(n715));
AOI22X1  g095(.A0(n714_1), .A1(n712), .B0(n711), .B1(n715), .Y(n716));
AND2X1   g096(.A(n716), .B(n710), .Y(n717));
OAI21X1  g097(.A0(n3084gat), .A1(n3083gat), .B0(n3095gat), .Y(n718));
OAI21X1  g098(.A0(n622), .A1(n650), .B0(n718), .Y(n719_1));
OAI21X1  g099(.A0(n3087gat), .A1(n3086gat), .B0(n3095gat), .Y(n720));
NOR2X1   g100(.A(n720), .B(n719_1), .Y(n721));
INVX1    g101(.A(n721), .Y(n722));
INVX1    g102(.A(n3084gat), .Y(n723));
OR2X1    g103(.A(n624_1), .B(n723), .Y(n724_1));
NAND3X1  g104(.A(n650), .B(n723), .C(n3083gat), .Y(n725));
INVX1    g105(.A(n3083gat), .Y(n726));
NAND3X1  g106(.A(n3085gat), .B(n723), .C(n726), .Y(n727));
NAND3X1  g107(.A(n3085gat), .B(n3084gat), .C(n3083gat), .Y(n728));
NAND4X1  g108(.A(n727), .B(n725), .C(n724_1), .D(n728), .Y(n729_1));
XOR2X1   g109(.A(n3087gat), .B(n3086gat), .Y(n730));
XOR2X1   g110(.A(n3089gat), .B(n3088gat), .Y(n731));
AND2X1   g111(.A(n731), .B(n730), .Y(n732));
INVX1    g112(.A(n730), .Y(n733));
AND2X1   g113(.A(n731), .B(n733), .Y(n734_1));
MX2X1    g114(.A(n732), .B(n734_1), .S0(n729_1), .Y(n735));
NOR2X1   g115(.A(n731), .B(n730), .Y(n736));
NOR2X1   g116(.A(n731), .B(n733), .Y(n737));
MX2X1    g117(.A(n736), .B(n737), .S0(n729_1), .Y(n738));
OR2X1    g118(.A(n738), .B(n735), .Y(n210));
OAI21X1  g119(.A0(n722), .A1(n717), .B0(n210), .Y(n3117gat));
INVX1    g120(.A(n861gat), .Y(n741));
INVX1    g121(.A(n580gat), .Y(n742));
AOI22X1  g122(.A0(n707), .A1(n742), .B0(n741), .B1(n709_1), .Y(n743));
INVX1    g123(.A(n337gat), .Y(n744_1));
INVX1    g124(.A(n777gat), .Y(n745));
AOI22X1  g125(.A0(n714_1), .A1(n745), .B0(n744_1), .B1(n715), .Y(n746));
AND2X1   g126(.A(n746), .B(n743), .Y(n747));
INVX1    g127(.A(n160gat), .Y(n748));
NOR3X1   g128(.A(n337gat), .B(n748), .C(n711), .Y(n749_1));
NOR3X1   g129(.A(n744_1), .B(n748), .C(n271gat), .Y(n750));
NOR3X1   g130(.A(n744_1), .B(n160gat), .C(n711), .Y(n751));
NOR3X1   g131(.A(n337gat), .B(n160gat), .C(n271gat), .Y(n752));
NOR4X1   g132(.A(n751), .B(n750), .C(n749_1), .D(n752), .Y(n753));
INVX1    g133(.A(n703gat), .Y(n754_1));
INVX1    g134(.A(n341gat), .Y(n755));
NOR3X1   g135(.A(n755), .B(n754_1), .C(n394gat), .Y(n756));
INVX1    g136(.A(n394gat), .Y(n757));
NOR3X1   g137(.A(n341gat), .B(n754_1), .C(n757), .Y(n758));
NOR3X1   g138(.A(n755), .B(n703gat), .C(n757), .Y(n759_1));
NOR3X1   g139(.A(n341gat), .B(n703gat), .C(n394gat), .Y(n760));
NOR4X1   g140(.A(n759_1), .B(n758), .C(n756), .D(n760), .Y(n761));
INVX1    g141(.A(n761), .Y(n762));
INVX1    g142(.A(n726gat), .Y(n763));
INVX1    g143(.A(n842gat), .Y(n764_1));
NOR3X1   g144(.A(n764_1), .B(n763), .C(n722gat), .Y(n765));
INVX1    g145(.A(n722gat), .Y(n766));
NOR3X1   g146(.A(n764_1), .B(n726gat), .C(n766), .Y(n767));
NOR3X1   g147(.A(n842gat), .B(n763), .C(n766), .Y(n768));
NOR3X1   g148(.A(n842gat), .B(n726gat), .C(n722gat), .Y(n769_1));
NOR4X1   g149(.A(n768), .B(n767), .C(n765), .D(n769_1), .Y(n770));
INVX1    g150(.A(n770), .Y(n771));
NAND3X1  g151(.A(n771), .B(n762), .C(n753), .Y(n772));
INVX1    g152(.A(n753), .Y(n773));
NAND3X1  g153(.A(n771), .B(n761), .C(n773), .Y(n774_1));
NAND3X1  g154(.A(n770), .B(n761), .C(n753), .Y(n775));
NAND3X1  g155(.A(n770), .B(n762), .C(n773), .Y(n776));
NAND4X1  g156(.A(n775), .B(n774_1), .C(n772), .D(n776), .Y(n240));
OAI21X1  g157(.A0(n747), .A1(n722), .B0(n240), .Y(n3118gat));
INVX1    g158(.A(n553gat), .Y(n779_1));
AOI22X1  g159(.A0(n714_1), .A1(n779_1), .B0(n748), .B1(n715), .Y(n780));
INVX1    g160(.A(n957gat), .Y(n781));
INVX1    g161(.A(n816gat), .Y(n782));
AOI22X1  g162(.A0(n707), .A1(n782), .B0(n781), .B1(n709_1), .Y(n783));
AND2X1   g163(.A(n783), .B(n780), .Y(n784_1));
NOR3X1   g164(.A(n861gat), .B(n781), .C(n701), .Y(n785));
NOR3X1   g165(.A(n741), .B(n781), .C(n1068gat), .Y(n786));
NOR3X1   g166(.A(n741), .B(n957gat), .C(n701), .Y(n787));
NOR3X1   g167(.A(n861gat), .B(n957gat), .C(n1068gat), .Y(n788));
NOR4X1   g168(.A(n787), .B(n786), .C(n785), .D(n788), .Y(n789_1));
INVX1    g169(.A(n865gat), .Y(n790));
INVX1    g170(.A(n1080gat), .Y(n791));
NOR3X1   g171(.A(n1148gat), .B(n791), .C(n790), .Y(n792));
INVX1    g172(.A(n1148gat), .Y(n793));
NOR3X1   g173(.A(n793), .B(n791), .C(n865gat), .Y(n794_1));
NOR3X1   g174(.A(n793), .B(n1080gat), .C(n790), .Y(n795));
NOR3X1   g175(.A(n1148gat), .B(n1080gat), .C(n865gat), .Y(n796));
NOR4X1   g176(.A(n795), .B(n794_1), .C(n792), .D(n796), .Y(n797));
INVX1    g177(.A(n797), .Y(n798));
INVX1    g178(.A(n1294gat), .Y(n799_1));
INVX1    g179(.A(n1241gat), .Y(n800));
NOR3X1   g180(.A(n1298gat), .B(n800), .C(n799_1), .Y(n801));
INVX1    g181(.A(n1298gat), .Y(n802));
NOR3X1   g182(.A(n802), .B(n800), .C(n1294gat), .Y(n803));
NOR3X1   g183(.A(n802), .B(n1241gat), .C(n799_1), .Y(n804_1));
NOR3X1   g184(.A(n1298gat), .B(n1241gat), .C(n1294gat), .Y(n805));
NOR4X1   g185(.A(n804_1), .B(n803), .C(n801), .D(n805), .Y(n806));
INVX1    g186(.A(n806), .Y(n807));
NAND3X1  g187(.A(n807), .B(n798), .C(n789_1), .Y(n808));
INVX1    g188(.A(n789_1), .Y(n809_1));
NAND3X1  g189(.A(n807), .B(n797), .C(n809_1), .Y(n810));
NAND3X1  g190(.A(n806), .B(n797), .C(n789_1), .Y(n811));
NAND3X1  g191(.A(n806), .B(n798), .C(n809_1), .Y(n812));
NAND4X1  g192(.A(n811), .B(n810), .C(n808), .D(n812), .Y(n343));
OAI21X1  g193(.A0(n784_1), .A1(n722), .B0(n343), .Y(n3119gat));
INVX1    g194(.A(n322gat), .Y(n815));
AOI22X1  g195(.A0(n709_1), .A1(n790), .B0(n815), .B1(n714_1), .Y(n816));
INVX1    g196(.A(n584gat), .Y(n817));
AOI22X1  g197(.A0(n707), .A1(n817), .B0(n755), .B1(n715), .Y(n818));
AND2X1   g198(.A(n818), .B(n816), .Y(n819_1));
INVX1    g199(.A(n283gat), .Y(n820));
INVX1    g200(.A(n165gat), .Y(n821));
NOR3X1   g201(.A(n279gat), .B(n821), .C(n820), .Y(n822));
INVX1    g202(.A(n279gat), .Y(n823));
NOR3X1   g203(.A(n823), .B(n821), .C(n283gat), .Y(n824_1));
NOR3X1   g204(.A(n823), .B(n165gat), .C(n820), .Y(n825));
NOR3X1   g205(.A(n279gat), .B(n165gat), .C(n283gat), .Y(n826));
NOR4X1   g206(.A(n825), .B(n824_1), .C(n822), .D(n826), .Y(n827));
INVX1    g207(.A(n402gat), .Y(n828));
INVX1    g208(.A(n275gat), .Y(n829_1));
NOR3X1   g209(.A(n829_1), .B(n828), .C(n398gat), .Y(n830));
INVX1    g210(.A(n398gat), .Y(n831));
NOR3X1   g211(.A(n275gat), .B(n828), .C(n831), .Y(n832));
NOR3X1   g212(.A(n829_1), .B(n402gat), .C(n831), .Y(n833));
NOR3X1   g213(.A(n275gat), .B(n402gat), .C(n398gat), .Y(n834_1));
NOR4X1   g214(.A(n833), .B(n832), .C(n830), .D(n834_1), .Y(n835));
INVX1    g215(.A(n835), .Y(n836));
INVX1    g216(.A(n846gat), .Y(n837));
INVX1    g217(.A(n1026gat), .Y(n838));
NOR3X1   g218(.A(n838), .B(n837), .C(n919gat), .Y(n839_1));
INVX1    g219(.A(n919gat), .Y(n840));
NOR3X1   g220(.A(n838), .B(n846gat), .C(n840), .Y(n841));
NOR3X1   g221(.A(n1026gat), .B(n837), .C(n840), .Y(n842));
NOR3X1   g222(.A(n1026gat), .B(n846gat), .C(n919gat), .Y(n843));
NOR4X1   g223(.A(n842), .B(n841), .C(n839_1), .D(n843), .Y(n844_1));
INVX1    g224(.A(n844_1), .Y(n845));
NAND3X1  g225(.A(n845), .B(n836), .C(n827), .Y(n846));
INVX1    g226(.A(n827), .Y(n847));
NAND3X1  g227(.A(n845), .B(n835), .C(n847), .Y(n848));
NAND3X1  g228(.A(n844_1), .B(n835), .C(n827), .Y(n849_1));
NAND3X1  g229(.A(n844_1), .B(n836), .C(n847), .Y(n850));
NAND4X1  g230(.A(n849_1), .B(n848), .C(n846), .D(n850), .Y(n294));
OAI21X1  g231(.A0(n819_1), .A1(n722), .B0(n294), .Y(n3120gat));
INVX1    g232(.A(n699gat), .Y(n964));
AOI22X1  g233(.A0(n707), .A1(n964), .B0(n793), .B1(n709_1), .Y(n854_1));
INVX1    g234(.A(n314gat), .Y(n855));
AOI22X1  g235(.A0(n714_1), .A1(n855), .B0(n757), .B1(n715), .Y(n856));
AND2X1   g236(.A(n856), .B(n854_1), .Y(n857));
NOR3X1   g237(.A(n580gat), .B(n782), .C(n702), .Y(n858));
NOR3X1   g238(.A(n742), .B(n782), .C(n680gat), .Y(n859_1));
NOR3X1   g239(.A(n742), .B(n816gat), .C(n702), .Y(n860));
NOR3X1   g240(.A(n580gat), .B(n816gat), .C(n680gat), .Y(n861));
NOR4X1   g241(.A(n860), .B(n859_1), .C(n858), .D(n861), .Y(n862));
INVX1    g242(.A(n684gat), .Y(n959));
NOR3X1   g243(.A(n699gat), .B(n959), .C(n817), .Y(n864_1));
NOR3X1   g244(.A(n964), .B(n959), .C(n584gat), .Y(n865));
NOR3X1   g245(.A(n964), .B(n684gat), .C(n817), .Y(n866));
NOR3X1   g246(.A(n699gat), .B(n684gat), .C(n584gat), .Y(n867));
NOR4X1   g247(.A(n866), .B(n865), .C(n864_1), .D(n867), .Y(n868));
INVX1    g248(.A(n868), .Y(n869_1));
INVX1    g249(.A(n824gat), .Y(n944));
INVX1    g250(.A(n820gat), .Y(n954));
NOR3X1   g251(.A(n883gat), .B(n954), .C(n944), .Y(n872));
INVX1    g252(.A(n883gat), .Y(n949));
NOR3X1   g253(.A(n949), .B(n954), .C(n824gat), .Y(n874_1));
NOR3X1   g254(.A(n949), .B(n820gat), .C(n944), .Y(n875));
NOR3X1   g255(.A(n883gat), .B(n820gat), .C(n824gat), .Y(n876));
NOR4X1   g256(.A(n875), .B(n874_1), .C(n872), .D(n876), .Y(n877));
INVX1    g257(.A(n877), .Y(n878));
NAND3X1  g258(.A(n878), .B(n869_1), .C(n862), .Y(n879_1));
INVX1    g259(.A(n862), .Y(n880));
NAND3X1  g260(.A(n878), .B(n868), .C(n880), .Y(n881));
NAND3X1  g261(.A(n877), .B(n868), .C(n862), .Y(n882));
NAND3X1  g262(.A(n877), .B(n869_1), .C(n880), .Y(n883));
NAND4X1  g263(.A(n882), .B(n881), .C(n879_1), .D(n883), .Y(n439));
OAI21X1  g264(.A0(n857), .A1(n722), .B0(n439), .Y(n3121gat));
AOI22X1  g265(.A0(n707), .A1(n959), .B0(n754_1), .B1(n715), .Y(n886));
INVX1    g266(.A(n318gat), .Y(n887));
AOI22X1  g267(.A0(n709_1), .A1(n791), .B0(n887), .B1(n714_1), .Y(n888));
AND2X1   g268(.A(n888), .B(n886), .Y(n889_1));
INVX1    g269(.A(n834gat), .Y(n979));
INVX1    g270(.A(n707gat), .Y(n939));
NOR3X1   g271(.A(n838gat), .B(n939), .C(n979), .Y(n892));
INVX1    g272(.A(n838gat), .Y(n969));
NOR3X1   g273(.A(n969), .B(n939), .C(n834gat), .Y(n894_1));
NOR3X1   g274(.A(n969), .B(n707gat), .C(n979), .Y(n895));
NOR3X1   g275(.A(n838gat), .B(n707gat), .C(n834gat), .Y(n896));
NOR4X1   g276(.A(n895), .B(n894_1), .C(n892), .D(n896), .Y(n897));
INVX1    g277(.A(n618gat), .Y(n898));
INVX1    g278(.A(n614gat), .Y(n934));
NOR3X1   g279(.A(n934), .B(n491gat), .C(n898), .Y(n900));
INVX1    g280(.A(n491gat), .Y(n901));
NOR3X1   g281(.A(n614gat), .B(n901), .C(n898), .Y(n902));
NOR3X1   g282(.A(n934), .B(n901), .C(n618gat), .Y(n903));
NOR3X1   g283(.A(n614gat), .B(n491gat), .C(n618gat), .Y(n904_1));
NOR4X1   g284(.A(n903), .B(n902), .C(n900), .D(n904_1), .Y(n905));
INVX1    g285(.A(n905), .Y(n906));
INVX1    g286(.A(n622gat), .Y(n907));
INVX1    g287(.A(n830gat), .Y(n974));
NOR3X1   g288(.A(n974), .B(n626gat), .C(n907), .Y(n909_1));
INVX1    g289(.A(n626gat), .Y(n910));
NOR3X1   g290(.A(n974), .B(n910), .C(n622gat), .Y(n911));
NOR3X1   g291(.A(n830gat), .B(n910), .C(n907), .Y(n912));
NOR3X1   g292(.A(n830gat), .B(n626gat), .C(n622gat), .Y(n913));
NOR4X1   g293(.A(n912), .B(n911), .C(n909_1), .D(n913), .Y(n914_1));
INVX1    g294(.A(n914_1), .Y(n915));
NAND3X1  g295(.A(n915), .B(n906), .C(n897), .Y(n916));
INVX1    g296(.A(n897), .Y(n917));
NAND3X1  g297(.A(n915), .B(n905), .C(n917), .Y(n918));
NAND3X1  g298(.A(n914_1), .B(n905), .C(n897), .Y(n919_1));
NAND3X1  g299(.A(n914_1), .B(n906), .C(n917), .Y(n920));
NAND4X1  g300(.A(n919_1), .B(n918), .C(n916), .D(n920), .Y(n389));
OAI21X1  g301(.A0(n889_1), .A1(n722), .B0(n389), .Y(n3122gat));
INVX1    g302(.A(n561gat), .Y(n923));
AOI22X1  g303(.A0(n714_1), .A1(n923), .B0(n763), .B1(n715), .Y(n924_1));
AOI22X1  g304(.A0(n707), .A1(n944), .B0(n799_1), .B1(n709_1), .Y(n925));
AND2X1   g305(.A(n925), .B(n924_1), .Y(n926));
NOR3X1   g306(.A(n777gat), .B(n779_1), .C(n712), .Y(n927));
NOR3X1   g307(.A(n745), .B(n779_1), .C(n659gat), .Y(n928));
NOR3X1   g308(.A(n745), .B(n553gat), .C(n712), .Y(n929_1));
NOR3X1   g309(.A(n777gat), .B(n553gat), .C(n659gat), .Y(n930));
OR4X1    g310(.A(n929_1), .B(n928), .C(n927), .D(n930), .Y(n931));
NOR3X1   g311(.A(n314gat), .B(n887), .C(n815), .Y(n932));
NOR3X1   g312(.A(n855), .B(n887), .C(n322gat), .Y(n933));
NOR3X1   g313(.A(n855), .B(n318gat), .C(n815), .Y(n934_1));
NOR3X1   g314(.A(n314gat), .B(n318gat), .C(n322gat), .Y(n935));
NOR4X1   g315(.A(n934_1), .B(n933), .C(n932), .D(n935), .Y(n936));
XOR2X1   g316(.A(n366gat), .B(n561gat), .Y(n937));
INVX1    g317(.A(n937), .Y(n938));
NOR3X1   g318(.A(n938), .B(n936), .C(n931), .Y(n939_1));
NOR4X1   g319(.A(n929_1), .B(n928), .C(n927), .D(n930), .Y(n940));
OR4X1    g320(.A(n934_1), .B(n933), .C(n932), .D(n935), .Y(n941));
NOR3X1   g321(.A(n938), .B(n941), .C(n940), .Y(n942));
NOR3X1   g322(.A(n937), .B(n941), .C(n931), .Y(n943));
NOR3X1   g323(.A(n937), .B(n936), .C(n940), .Y(n944_1));
NOR4X1   g324(.A(n943), .B(n942), .C(n939_1), .D(n944_1), .Y(n945));
XOR2X1   g325(.A(n945), .B(n667gat), .Y(n609));
OAI21X1  g326(.A0(n926), .A1(n722), .B0(n609), .Y(n3123gat));
INVX1    g327(.A(n714_1), .Y(n948));
OR4X1    g328(.A(n704_1), .B(n713), .C(n673gat), .D(n708), .Y(n949_1));
OAI21X1  g329(.A0(n948), .A1(n366gat), .B0(n949_1), .Y(n950));
NOR4X1   g330(.A(n704_1), .B(n703), .C(n722gat), .D(n706), .Y(n951));
INVX1    g331(.A(n707), .Y(n952));
INVX1    g332(.A(n709_1), .Y(n953));
OAI22X1  g333(.A0(n952), .A1(n883gat), .B0(n1298gat), .B1(n953), .Y(n954_1));
NOR3X1   g334(.A(n954_1), .B(n951), .C(n950), .Y(n955));
NOR4X1   g335(.A(n698), .B(n697), .C(n695), .D(n699_1), .Y(n956));
XOR2X1   g336(.A(n956), .B(n1197gat), .Y(n559));
OAI21X1  g337(.A0(n955), .A1(n722), .B0(n559), .Y(n3124gat));
NOR2X1   g338(.A(n945), .B(n948), .Y(n959_1));
NAND4X1  g339(.A(n705), .B(n703), .C(n673gat), .D(n706), .Y(n960));
NAND3X1  g340(.A(n708), .B(n704_1), .C(n703), .Y(n961));
NAND4X1  g341(.A(n705), .B(n713), .C(n800), .D(n706), .Y(n962));
AOI22X1  g342(.A0(n707), .A1(n954), .B0(n764_1), .B1(n715), .Y(n963));
NAND4X1  g343(.A(n962), .B(n961), .C(n960), .D(n963), .Y(n964_1));
NOR2X1   g344(.A(n964_1), .B(n959_1), .Y(n965));
XOR2X1   g345(.A(n2390gat), .B(n2495gat), .Y(n966));
INVX1    g346(.A(n2270gat), .Y(n3127gat));
XOR2X1   g347(.A(n2339gat), .B(n3127gat), .Y(n968));
XOR2X1   g348(.A(n968), .B(n966), .Y(n649));
OAI21X1  g349(.A0(n965), .A1(n722), .B0(n649), .Y(n3125gat));
INVX1    g350(.A(n2339gat), .Y(n3126gat));
INVX1    g351(.A(n2390gat), .Y(n3128gat));
INVX1    g352(.A(n719_1), .Y(n973));
AND2X1   g353(.A(n3093gat), .B(n3088gat), .Y(n974_1));
NAND3X1  g354(.A(n3093gat), .B(n3088gat), .C(n3087gat), .Y(n975));
NOR4X1   g355(.A(n632), .B(n631), .C(n650), .D(n975), .Y(n976));
OAI21X1  g356(.A0(n3086gat), .A1(n3085gat), .B0(n3093gat), .Y(n977));
AOI21X1  g357(.A0(n723), .A1(n726), .B0(n632), .Y(n978));
NOR4X1   g358(.A(n977), .B(n976), .C(n974_1), .D(n978), .Y(n979_1));
NOR4X1   g359(.A(n642), .B(n621), .C(n631), .D(n622), .Y(n980));
AOI21X1  g360(.A0(n980), .A1(n973), .B0(n979_1), .Y(n981));
NOR3X1   g361(.A(n978), .B(n977), .C(n976), .Y(n982));
AOI21X1  g362(.A0(n982), .A1(n974_1), .B0(n721), .Y(n983));
OAI22X1  g363(.A0(n952), .A1(n830gat), .B0(n1026gat), .B1(n953), .Y(n984_1));
AOI21X1  g364(.A0(n714_1), .A1(n3116gat), .B0(n984_1), .Y(n985));
OAI22X1  g365(.A0(n983), .A1(n985), .B0(n981), .B1(n965), .Y(n3129gat));
OAI22X1  g366(.A0(n952), .A1(n834gat), .B0(n1035gat), .B1(n948), .Y(n987));
AOI21X1  g367(.A0(n709_1), .A1(n820), .B0(n987), .Y(n988));
OAI22X1  g368(.A0(n983), .A1(n988), .B0(n981), .B1(n717), .Y(n3130gat));
OAI22X1  g369(.A0(n952), .A1(n838gat), .B0(n1072gat), .B1(n948), .Y(n990));
AOI21X1  g370(.A0(n709_1), .A1(n823), .B0(n990), .Y(n991));
OAI22X1  g371(.A0(n983), .A1(n991), .B0(n981), .B1(n747), .Y(n3131gat));
OAI22X1  g372(.A0(n952), .A1(n707gat), .B0(n1121gat), .B1(n948), .Y(n993));
AOI21X1  g373(.A0(n709_1), .A1(n821), .B0(n993), .Y(n994_1));
OAI22X1  g374(.A0(n983), .A1(n994_1), .B0(n981), .B1(n784_1), .Y(n3132gat));
OAI22X1  g375(.A0(n952), .A1(n614gat), .B0(n931gat), .B1(n948), .Y(n996));
AOI21X1  g376(.A0(n709_1), .A1(n829_1), .B0(n996), .Y(n997));
OAI22X1  g377(.A0(n983), .A1(n997), .B0(n981), .B1(n819_1), .Y(n3133gat));
OAI22X1  g378(.A0(n952), .A1(n491gat), .B0(n1045gat), .B1(n948), .Y(n999_1));
AOI21X1  g379(.A0(n709_1), .A1(n831), .B0(n999_1), .Y(n1000));
OAI22X1  g380(.A0(n983), .A1(n1000), .B0(n981), .B1(n857), .Y(n3134gat));
OAI22X1  g381(.A0(n952), .A1(n618gat), .B0(n1135gat), .B1(n948), .Y(n1002));
AOI21X1  g382(.A0(n709_1), .A1(n828), .B0(n1002), .Y(n1003));
OAI22X1  g383(.A0(n983), .A1(n1003), .B0(n981), .B1(n889_1), .Y(n3135gat));
OAI22X1  g384(.A0(n952), .A1(n622gat), .B0(n1282gat), .B1(n948), .Y(n1005));
AOI21X1  g385(.A0(n709_1), .A1(n837), .B0(n1005), .Y(n1006));
OAI22X1  g386(.A0(n983), .A1(n1006), .B0(n981), .B1(n926), .Y(n3136gat));
OAI22X1  g387(.A0(n952), .A1(n626gat), .B0(n1226gat), .B1(n948), .Y(n1008));
AOI21X1  g388(.A0(n709_1), .A1(n840), .B0(n1008), .Y(n1009_1));
OAI22X1  g389(.A0(n983), .A1(n1009_1), .B0(n981), .B1(n955), .Y(n3137gat));
NAND2X1  g390(.A(n754_1), .B(n394gat), .Y(n1011));
AND2X1   g391(.A(n726gat), .B(n722gat), .Y(n1012));
INVX1    g392(.A(n1012), .Y(n1013));
NOR3X1   g393(.A(n1013), .B(n1011), .C(n2454gat), .Y(n1014_1));
NAND2X1  g394(.A(n726gat), .B(n766), .Y(n1015));
NOR3X1   g395(.A(n1015), .B(n1011), .C(n2454gat), .Y(n1016));
NOR2X1   g396(.A(n1016), .B(n1014_1), .Y(n1017));
INVX1    g397(.A(n2562gat), .Y(n714));
NOR2X1   g398(.A(n2207gat), .B(n2203gat), .Y(n1019_1));
NAND4X1  g399(.A(n714), .B(n2343gat), .C(n2399gat), .D(n1019_1), .Y(n1020));
INVX1    g400(.A(n2626gat), .Y(n694));
AND2X1   g401(.A(n2543gat), .B(n2630gat), .Y(n1022));
NAND4X1  g402(.A(n2622gat), .B(n2490gat), .C(n694), .D(n1022), .Y(n1023));
NOR3X1   g403(.A(n1023), .B(n1020), .C(n1017), .Y(n3138gat));
INVX1    g404(.A(n2343gat), .Y(n709));
NAND4X1  g405(.A(n2562gat), .B(n709), .C(n2399gat), .D(n1019_1), .Y(n1026));
OR2X1    g406(.A(n726gat), .B(n722gat), .Y(n1027));
INVX1    g407(.A(n2454gat), .Y(n1028));
NAND3X1  g408(.A(n1028), .B(n703gat), .C(n394gat), .Y(n1029_1));
NAND2X1  g409(.A(n763), .B(n722gat), .Y(n1030));
AOI21X1  g410(.A0(n1030), .A1(n1027), .B0(n1029_1), .Y(n1031));
NAND4X1  g411(.A(n1028), .B(n703gat), .C(n757), .D(n1012), .Y(n1032));
OAI21X1  g412(.A0(n1029_1), .A1(n1015), .B0(n1032), .Y(n1033));
NOR4X1   g413(.A(n1031), .B(n1016), .C(n1014_1), .D(n1033), .Y(n1034_1));
OAI21X1  g414(.A0(n1763gat), .A1(n1880gat), .B0(n2102gat), .Y(n509));
INVX1    g415(.A(n509), .Y(n1036));
NOR3X1   g416(.A(n1036), .B(n1034_1), .C(n1340gat), .Y(n1037));
INVX1    g417(.A(n1394gat), .Y(n744));
NAND3X1  g418(.A(n1767gat), .B(n1834gat), .C(n1880gat), .Y(n3149gat));
INVX1    g419(.A(n3149gat), .Y(n1040));
NOR4X1   g420(.A(n1036), .B(n1462gat), .C(n744), .D(n1040), .Y(n1041));
AOI21X1  g421(.A0(n1037), .A1(n1026), .B0(n1041), .Y(n1042));
OR2X1    g422(.A(n1042), .B(n1508gat), .Y(n1043));
NAND2X1  g423(.A(n509), .B(n1462gat), .Y(n1044_1));
INVX1    g424(.A(n1596gat), .Y(n1045));
NAND3X1  g425(.A(n1036), .B(n1031), .C(n1045), .Y(n1046));
AOI21X1  g426(.A0(n1046), .A1(n1044_1), .B0(n1678gat), .Y(n1047));
INVX1    g427(.A(n1775gat), .Y(n819));
NAND4X1  g428(.A(n2021gat), .B(n1880gat), .C(n3097gat), .D(n819), .Y(n1049));
NAND2X1  g429(.A(n1825gat), .B(n1821gat), .Y(n264));
NOR2X1   g430(.A(n264), .B(n1829gat), .Y(n1051));
OR4X1    g431(.A(n3106gat), .B(n1775gat), .C(n3098gat), .D(n1051), .Y(n1052));
AOI21X1  g432(.A0(n1049), .A1(n1825gat), .B0(n1052), .Y(n1053));
NOR3X1   g433(.A(n1033), .B(n1016), .C(n1014_1), .Y(n1054));
NOR4X1   g434(.A(n1054), .B(n1525gat), .C(n1394gat), .D(n509), .Y(n1055));
NOR3X1   g435(.A(n1055), .B(n1053), .C(n1047), .Y(n1056));
NOR4X1   g436(.A(n2454gat), .B(n754_1), .C(n757), .D(n1027), .Y(n1057));
NOR2X1   g437(.A(n1030), .B(n1029_1), .Y(n1058));
NOR2X1   g438(.A(n1058), .B(n1057), .Y(n1059));
NOR4X1   g439(.A(n1596gat), .B(n1678gat), .C(n744), .D(n509), .Y(n1060));
NOR3X1   g440(.A(n509), .B(n1588gat), .C(n1045), .Y(n1061));
AOI21X1  g441(.A0(n1060), .A1(n1059), .B0(n1061), .Y(n1062));
NAND3X1  g442(.A(n1062), .B(n1056), .C(n1043), .Y(n3139gat));
INVX1    g443(.A(n1456gat), .Y(n1064));
AND2X1   g444(.A(n3149gat), .B(n509), .Y(n1065));
OAI21X1  g445(.A0(n1065), .A1(n1037), .B0(n1064), .Y(n1066));
INVX1    g446(.A(n1748gat), .Y(n1067));
OR2X1    g447(.A(n1763gat), .B(n1880gat), .Y(n1068));
NAND3X1  g448(.A(n1068), .B(n1336gat), .C(n2102gat), .Y(n1069));
OAI21X1  g449(.A0(n3149gat), .A1(n1031), .B0(n1036), .Y(n1070));
OAI21X1  g450(.A0(n1069), .A1(n1054), .B0(n1070), .Y(n1071));
NAND2X1  g451(.A(n1071), .B(n1067), .Y(n1072));
INVX1    g452(.A(n1807gat), .Y(n1073));
NAND3X1  g453(.A(n509), .B(n1340gat), .C(n1073), .Y(n1074));
OR4X1    g454(.A(n1054), .B(n1675gat), .C(n1394gat), .D(n509), .Y(n1075));
NAND4X1  g455(.A(n1074), .B(n1072), .C(n1066), .D(n1075), .Y(n3141gat));
XOR2X1   g456(.A(n1057), .B(n945), .Y(n1077));
NAND4X1  g457(.A(n2562gat), .B(n2343gat), .C(n2399gat), .D(n1019_1), .Y(n1078));
NAND3X1  g458(.A(n2562gat), .B(n709), .C(n2399gat), .Y(n1079));
INVX1    g459(.A(n2207gat), .Y(n719));
NAND3X1  g460(.A(n779_1), .B(n719), .C(n2203gat), .Y(n1081));
NOR2X1   g461(.A(n2562gat), .B(n2343gat), .Y(n1082));
NAND2X1  g462(.A(n1082), .B(n2399gat), .Y(n1083));
NAND3X1  g463(.A(n815), .B(n719), .C(n2203gat), .Y(n1084));
OAI22X1  g464(.A0(n1083), .A1(n1084), .B0(n1081), .B1(n1079), .Y(n1085));
NAND3X1  g465(.A(n714), .B(n2343gat), .C(n2399gat), .Y(n1086));
NAND3X1  g466(.A(n745), .B(n719), .C(n2203gat), .Y(n1087));
INVX1    g467(.A(n2203gat), .Y(n724));
NAND3X1  g468(.A(n2562gat), .B(n2343gat), .C(n2399gat), .Y(n1089));
OR4X1    g469(.A(n659gat), .B(n2207gat), .C(n724), .D(n1089), .Y(n1090));
OAI21X1  g470(.A0(n1087), .A1(n1086), .B0(n1090), .Y(n1091));
INVX1    g471(.A(n2399gat), .Y(n704));
NOR3X1   g472(.A(n366gat), .B(n2207gat), .C(n724), .Y(n1093));
NAND3X1  g473(.A(n1093), .B(n1082), .C(n704), .Y(n1094));
NAND3X1  g474(.A(n2562gat), .B(n2343gat), .C(n704), .Y(n1095));
NAND3X1  g475(.A(n855), .B(n719), .C(n2203gat), .Y(n1096));
OAI21X1  g476(.A0(n1096), .A1(n1095), .B0(n1094), .Y(n1097));
NAND3X1  g477(.A(n2562gat), .B(n709), .C(n704), .Y(n1098));
NAND3X1  g478(.A(n923), .B(n719), .C(n2203gat), .Y(n1099));
NAND3X1  g479(.A(n714), .B(n2343gat), .C(n704), .Y(n1100));
NAND3X1  g480(.A(n887), .B(n719), .C(n2203gat), .Y(n1101));
OAI22X1  g481(.A0(n1100), .A1(n1101), .B0(n1099), .B1(n1098), .Y(n1102));
NOR4X1   g482(.A(n1097), .B(n1091), .C(n1085), .D(n1102), .Y(n1103));
OAI21X1  g483(.A0(n1078), .A1(n1077), .B0(n1103), .Y(n1104));
INVX1    g484(.A(n1389gat), .Y(n1105));
MX2X1    g485(.A(n707gat), .B(n165gat), .S0(n3149gat), .Y(n1106));
OR4X1    g486(.A(n1095), .B(n719), .C(n2203gat), .D(n1106), .Y(n1107));
MX2X1    g487(.A(n838gat), .B(n279gat), .S0(n3149gat), .Y(n1108));
OR4X1    g488(.A(n1083), .B(n719), .C(n2203gat), .D(n1108), .Y(n1109));
MX2X1    g489(.A(n834gat), .B(n283gat), .S0(n3149gat), .Y(n1110));
OR4X1    g490(.A(n1079), .B(n719), .C(n2203gat), .D(n1110), .Y(n1111));
MX2X1    g491(.A(n614gat), .B(n275gat), .S0(n3149gat), .Y(n1112));
OR4X1    g492(.A(n1100), .B(n719), .C(n2203gat), .D(n1112), .Y(n1113));
NAND4X1  g493(.A(n1111), .B(n1109), .C(n1107), .D(n1113), .Y(n1114));
AND2X1   g494(.A(n2207gat), .B(n2203gat), .Y(n1115));
NAND4X1  g495(.A(n714), .B(n2343gat), .C(n2399gat), .D(n1115), .Y(n1116));
AOI21X1  g496(.A0(n1032), .A1(n1059), .B0(n1116), .Y(n1117));
NAND2X1  g497(.A(n2207gat), .B(n2203gat), .Y(n1118));
MX2X1    g498(.A(n699gat), .B(n1148gat), .S0(n3149gat), .Y(n1119));
NOR3X1   g499(.A(n1119), .B(n1118), .C(n1098), .Y(n1120));
OR2X1    g500(.A(n1118), .B(n1089), .Y(n1121));
AOI21X1  g501(.A0(n1032), .A1(n2084gat), .B0(n1121), .Y(n1122));
OR2X1    g502(.A(n1122), .B(n1120), .Y(n1123));
MX2X1    g503(.A(n959), .B(n791), .S0(n3149gat), .Y(n1124));
NAND4X1  g504(.A(n1115), .B(n1082), .C(n704), .D(n1124), .Y(n1125));
MX2X1    g505(.A(n949), .B(n802), .S0(n3149gat), .Y(n1126));
NOR3X1   g506(.A(n1086), .B(n719), .C(n2203gat), .Y(n1127));
MX2X1    g507(.A(n944), .B(n799_1), .S0(n3149gat), .Y(n1128));
NOR3X1   g508(.A(n1089), .B(n719), .C(n2203gat), .Y(n1129));
AOI22X1  g509(.A0(n1128), .A1(n1129), .B0(n1127), .B1(n1126), .Y(n1130));
MX2X1    g510(.A(n782), .B(n781), .S0(n3149gat), .Y(n1131));
NOR4X1   g511(.A(n714), .B(n709), .C(n2399gat), .D(n1118), .Y(n1132));
MX2X1    g512(.A(n702), .B(n701), .S0(n3149gat), .Y(n1133));
NOR4X1   g513(.A(n714), .B(n2343gat), .C(n704), .D(n1118), .Y(n1134));
AOI22X1  g514(.A0(n1133), .A1(n1134), .B0(n1132), .B1(n1131), .Y(n1135));
MX2X1    g515(.A(n742), .B(n741), .S0(n3149gat), .Y(n1136));
NOR4X1   g516(.A(n2562gat), .B(n2343gat), .C(n704), .D(n1118), .Y(n1137));
MX2X1    g517(.A(n817), .B(n790), .S0(n3149gat), .Y(n1138));
NOR4X1   g518(.A(n2562gat), .B(n709), .C(n2399gat), .D(n1118), .Y(n1139));
AOI22X1  g519(.A0(n1138), .A1(n1139), .B0(n1137), .B1(n1136), .Y(n1140));
NAND4X1  g520(.A(n1135), .B(n1130), .C(n1125), .D(n1140), .Y(n1141));
NOR4X1   g521(.A(n1123), .B(n1117), .C(n1114), .D(n1141), .Y(n1142));
NOR4X1   g522(.A(n1036), .B(n1508gat), .C(n1394gat), .D(n1040), .Y(n1143));
NAND3X1  g523(.A(n3149gat), .B(n1068), .C(n2102gat), .Y(n1144));
NOR3X1   g524(.A(n1144), .B(n1678gat), .C(n1394gat), .Y(n1145));
NOR3X1   g525(.A(n2592gat), .B(n3106gat), .C(n673gat), .Y(n1146));
NOR3X1   g526(.A(n1146), .B(n1145), .C(n1143), .Y(n1147));
OAI21X1  g527(.A0(n1142), .A1(n1105), .B0(n1147), .Y(n1148));
AOI21X1  g528(.A0(n1104), .A1(n1031), .B0(n1148), .Y(n1149));
INVX1    g529(.A(n2622gat), .Y(n684));
NOR3X1   g530(.A(n684), .B(n2490gat), .C(n2626gat), .Y(n1151));
INVX1    g531(.A(n2490gat), .Y(n689));
NOR3X1   g532(.A(n2622gat), .B(n689), .C(n2626gat), .Y(n1153));
NOR3X1   g533(.A(n684), .B(n689), .C(n694), .Y(n1154));
NOR3X1   g534(.A(n2622gat), .B(n2490gat), .C(n694), .Y(n1155));
NOR4X1   g535(.A(n1154), .B(n1153), .C(n1151), .D(n1155), .Y(n1156));
INVX1    g536(.A(n2630gat), .Y(n699));
INVX1    g537(.A(n2634gat), .Y(n924));
NOR3X1   g538(.A(n924), .B(n2543gat), .C(n699), .Y(n1159));
INVX1    g539(.A(n2543gat), .Y(n679));
NOR3X1   g540(.A(n924), .B(n679), .C(n2630gat), .Y(n1161));
AND2X1   g541(.A(n1022), .B(n924), .Y(n1162));
NOR3X1   g542(.A(n2634gat), .B(n2543gat), .C(n2630gat), .Y(n1163));
NOR4X1   g543(.A(n1162), .B(n1161), .C(n1159), .D(n1163), .Y(n1164));
XOR2X1   g544(.A(n1164), .B(n1156), .Y(n659));
NAND2X1  g545(.A(n659), .B(n1149), .Y(n3143gat));
NOR3X1   g546(.A(n2640gat), .B(n2562gat), .C(n709), .Y(n1167));
NOR3X1   g547(.A(n2640gat), .B(n714), .C(n2343gat), .Y(n1168));
INVX1    g548(.A(n2640gat), .Y(n929));
NOR3X1   g549(.A(n929), .B(n714), .C(n709), .Y(n1170));
AND2X1   g550(.A(n1082), .B(n2640gat), .Y(n1171));
NOR4X1   g551(.A(n1170), .B(n1168), .C(n1167), .D(n1171), .Y(n1172));
NOR3X1   g552(.A(n719), .B(n2203gat), .C(n704), .Y(n1173));
NOR3X1   g553(.A(n2207gat), .B(n724), .C(n704), .Y(n1174));
NOR2X1   g554(.A(n1118), .B(n2399gat), .Y(n1175));
NOR3X1   g555(.A(n2207gat), .B(n2203gat), .C(n2399gat), .Y(n1176));
NOR4X1   g556(.A(n1175), .B(n1174), .C(n1173), .D(n1176), .Y(n1177));
XOR2X1   g557(.A(n1177), .B(n1172), .Y(n624));
NAND2X1  g558(.A(n624), .B(n1149), .Y(n3144gat));
INVX1    g559(.A(n1034_1), .Y(n869));
AOI21X1  g560(.A0(n655), .A1(n2514gat), .B0(n869), .Y(n3145gat));
NAND4X1  g561(.A(n2514gat), .B(n1871gat), .C(n1775gat), .D(n1771gat), .Y(n1182));
INVX1    g562(.A(n2176gat), .Y(n859));
INVX1    g563(.A(n2110gat), .Y(n909));
NAND4X1  g564(.A(n2037gat), .B(n2169gat), .C(n2095gat), .D(n2033gat), .Y(n1185));
NOR3X1   g565(.A(n1185), .B(n909), .C(n859), .Y(n1186));
AND2X1   g566(.A(n1186), .B(n1182), .Y(n3146gat));
NAND2X1  g567(.A(n2446gat), .B(n2450gat), .Y(n3147gat));
INVX1    g568(.A(n2450gat), .Y(n3148gat));
XOR2X1   g569(.A(n647), .B(n2061gat), .Y(n1190));
OAI21X1  g570(.A0(n2454gat), .A1(n337gat), .B0(n1190), .Y(n3150gat));
INVX1    g571(.A(n2139gat), .Y(n1192));
INVX1    g572(.A(n1899gat), .Y(n1193));
OR4X1    g573(.A(n627), .B(n1193), .C(n1192), .D(n636), .Y(n3151gat));
ONE      g574(.Y(n3152gat));
INVX1    g575(.A(n3072gat), .Y(n1196));
INVX1    g576(.A(n3081gat), .Y(n1197));
OAI22X1  g577(.A0(n632), .A1(n1196), .B0(n1197), .B1(n622), .Y(n169));
NOR4X1   g578(.A(n766), .B(n754_1), .C(n757), .D(n763), .Y(n245));
INVX1    g579(.A(n2472gat), .Y(n250));
INVX1    g580(.A(n2319gat), .Y(n1201));
NOR2X1   g581(.A(n1201), .B(n3099gat), .Y(n255));
INVX1    g582(.A(n2029gat), .Y(n269));
INVX1    g583(.A(n3065gat), .Y(n1204));
INVX1    g584(.A(n3074gat), .Y(n1205));
OAI22X1  g585(.A0(n632), .A1(n1204), .B0(n1205), .B1(n622), .Y(n299));
INVX1    g586(.A(n3067gat), .Y(n1207));
INVX1    g587(.A(n3076gat), .Y(n1208));
OAI22X1  g588(.A0(n632), .A1(n1207), .B0(n1208), .B1(n622), .Y(n304));
INVX1    g589(.A(n3066gat), .Y(n1210));
INVX1    g590(.A(n3075gat), .Y(n1211));
OAI22X1  g591(.A0(n632), .A1(n1210), .B0(n1211), .B1(n622), .Y(n309));
INVX1    g592(.A(n3071gat), .Y(n1213));
NAND2X1  g593(.A(n3095gat), .B(n3080gat), .Y(n1214));
OAI21X1  g594(.A0(n632), .A1(n1213), .B0(n1214), .Y(n314));
INVX1    g595(.A(n3073gat), .Y(n1216));
INVX1    g596(.A(n3082gat), .Y(n1217));
OAI22X1  g597(.A0(n632), .A1(n1216), .B0(n1217), .B1(n622), .Y(n319));
INVX1    g598(.A(n3068gat), .Y(n1219));
INVX1    g599(.A(n3077gat), .Y(n1220));
OAI22X1  g600(.A0(n632), .A1(n1219), .B0(n1220), .B1(n622), .Y(n328));
INVX1    g601(.A(n3070gat), .Y(n1222));
INVX1    g602(.A(n3079gat), .Y(n1223));
OAI22X1  g603(.A0(n632), .A1(n1222), .B0(n1223), .B1(n622), .Y(n333));
INVX1    g604(.A(n3069gat), .Y(n1225));
INVX1    g605(.A(n3078gat), .Y(n1226));
OAI22X1  g606(.A0(n632), .A1(n1225), .B0(n1226), .B1(n622), .Y(n338));
AND2X1   g607(.A(n625), .B(n3086gat), .Y(n1228));
INVX1    g608(.A(n1228), .Y(n1229));
AND2X1   g609(.A(n625), .B(n3087gat), .Y(n1230));
NAND2X1  g610(.A(n625), .B(n3088gat), .Y(n1231));
NOR4X1   g611(.A(n1230), .B(n1229), .C(n641), .D(n1231), .Y(n1232));
NAND3X1  g612(.A(n638), .B(n3088gat), .C(n3087gat), .Y(n1233));
NOR4X1   g613(.A(n634_1), .B(n3086gat), .C(n650), .D(n1233), .Y(n1234));
NOR2X1   g614(.A(n1234), .B(n1232), .Y(n1235));
INVX1    g615(.A(n156gat), .Y(n1236));
INVX1    g616(.A(n256gat), .Y(n1237));
NOR4X1   g617(.A(n1011), .B(n152gat), .C(n2454gat), .D(n1015), .Y(n1238));
NAND4X1  g618(.A(n148gat), .B(n1237), .C(n1236), .D(n1238), .Y(n1239));
AND2X1   g619(.A(n1238), .B(n1236), .Y(n1240));
OR2X1    g620(.A(n1240), .B(n148gat), .Y(n1241));
OR2X1    g621(.A(n148gat), .B(n1237), .Y(n1242));
NAND3X1  g622(.A(n1242), .B(n1241), .C(n1239), .Y(n1243));
MX2X1    g623(.A(n3065gat), .B(n1243), .S0(n1235), .Y(n364));
NAND3X1  g624(.A(n1016), .B(n152gat), .C(n1236), .Y(n1245));
INVX1    g625(.A(n152gat), .Y(n1246));
NAND2X1  g626(.A(n1246), .B(n156gat), .Y(n1247));
OR2X1    g627(.A(n1016), .B(n152gat), .Y(n1248));
NAND3X1  g628(.A(n1248), .B(n1247), .C(n1245), .Y(n1249));
MX2X1    g629(.A(n3067gat), .B(n1249), .S0(n1235), .Y(n369));
XOR2X1   g630(.A(n1240), .B(n1237), .Y(n1251));
MX2X1    g631(.A(n3066gat), .B(n1251), .S0(n1235), .Y(n374));
AOI22X1  g632(.A0(n1016), .A1(n156gat), .B0(n256gat), .B1(n1238), .Y(n1253));
XOR2X1   g633(.A(n1253), .B(n470gat), .Y(n1254));
MX2X1    g634(.A(n3073gat), .B(n1254), .S0(n1235), .Y(n379));
XOR2X1   g635(.A(n1016), .B(n1236), .Y(n1256));
MX2X1    g636(.A(n3068gat), .B(n1256), .S0(n1235), .Y(n384));
INVX1    g637(.A(n1232), .Y(n1258));
NOR3X1   g638(.A(n637), .B(n3088gat), .C(n621), .Y(n1259));
NAND4X1  g639(.A(n633), .B(n631), .C(n3085gat), .D(n1259), .Y(n1260));
OAI22X1  g640(.A0(n1258), .A1(n1205), .B0(n1204), .B1(n1260), .Y(n394));
OAI22X1  g641(.A0(n1258), .A1(n1208), .B0(n1207), .B1(n1260), .Y(n399));
OAI22X1  g642(.A0(n1258), .A1(n1211), .B0(n1210), .B1(n1260), .Y(n404));
INVX1    g643(.A(n1260), .Y(n1264));
OR2X1    g644(.A(n1264), .B(n1232), .Y(n1265));
INVX1    g645(.A(n331gat), .Y(n1266));
NOR2X1   g646(.A(n388gat), .B(n1266), .Y(n1267));
INVX1    g647(.A(n388gat), .Y(n1268));
AOI21X1  g648(.A0(n1014_1), .A1(n1268), .B0(n331gat), .Y(n1269));
AOI21X1  g649(.A0(n1267), .A1(n1014_1), .B0(n1269), .Y(n1270));
AOI22X1  g650(.A0(n1232), .A1(n3080gat), .B0(n3071gat), .B1(n1264), .Y(n1271));
OAI21X1  g651(.A0(n1270), .A1(n1265), .B0(n1271), .Y(n409));
INVX1    g652(.A(n1014_1), .Y(n1273));
NAND2X1  g653(.A(n327gat), .B(n1266), .Y(n1274));
AOI21X1  g654(.A0(n1274), .A1(n1268), .B0(n1273), .Y(n1275));
XOR2X1   g655(.A(n1275), .B(n463gat), .Y(n1276));
AOI22X1  g656(.A0(n1232), .A1(n3082gat), .B0(n3073gat), .B1(n1264), .Y(n1277));
OAI21X1  g657(.A0(n1276), .A1(n1265), .B0(n1277), .Y(n414));
XOR2X1   g658(.A(n1014_1), .B(n388gat), .Y(n1279));
AOI22X1  g659(.A0(n1232), .A1(n3081gat), .B0(n3072gat), .B1(n1264), .Y(n1280));
OAI21X1  g660(.A0(n1279), .A1(n1265), .B0(n1280), .Y(n419));
OAI22X1  g661(.A0(n1258), .A1(n1220), .B0(n1219), .B1(n1260), .Y(n424));
NOR3X1   g662(.A(n1273), .B(n388gat), .C(n331gat), .Y(n1283));
XOR2X1   g663(.A(n1283), .B(n327gat), .Y(n1284));
AOI22X1  g664(.A0(n1232), .A1(n3079gat), .B0(n3070gat), .B1(n1264), .Y(n1285));
OAI21X1  g665(.A0(n1284), .A1(n1265), .B0(n1285), .Y(n429));
INVX1    g666(.A(n327gat), .Y(n1287));
AND2X1   g667(.A(n384gat), .B(n1287), .Y(n1288));
AOI21X1  g668(.A0(n1283), .A1(n1287), .B0(n384gat), .Y(n1289));
AOI21X1  g669(.A0(n1288), .A1(n1283), .B0(n1289), .Y(n1290));
AOI22X1  g670(.A0(n1232), .A1(n3078gat), .B0(n3069gat), .B1(n1264), .Y(n1291));
OAI21X1  g671(.A0(n1290), .A1(n1265), .B0(n1291), .Y(n434));
INVX1    g672(.A(n2394gat), .Y(n1293));
NAND2X1  g673(.A(n2440gat), .B(n1293), .Y(n1294));
INVX1    g674(.A(n2407gat), .Y(n1295));
NAND3X1  g675(.A(n660), .B(n1295), .C(n2403gat), .Y(n1296));
NOR2X1   g676(.A(n1296), .B(n1294), .Y(n1297));
INVX1    g677(.A(n2440gat), .Y(n1298));
NAND2X1  g678(.A(n1298), .B(n2394gat), .Y(n1299));
NOR2X1   g679(.A(n1296), .B(n1299), .Y(n1300));
MX2X1    g680(.A(n1297), .B(n1300), .S0(n1036), .Y(n1301));
INVX1    g681(.A(n2095gat), .Y(n854));
INVX1    g682(.A(n2037gat), .Y(n899));
INVX1    g683(.A(n2309gat), .Y(n839));
NAND2X1  g684(.A(n2658gat), .B(n2588gat), .Y(n1305));
NAND3X1  g685(.A(n2506gat), .B(n2502gat), .C(n2510gat), .Y(n1306));
NOR3X1   g686(.A(n1306), .B(n1305), .C(n839), .Y(n1307));
NOR2X1   g687(.A(n1307), .B(n3100gat), .Y(n1308));
NAND2X1  g688(.A(n2021gat), .B(n1880gat), .Y(n1309));
AND2X1   g689(.A(n1309), .B(n2099gat), .Y(n1310));
NOR4X1   g690(.A(n1308), .B(n899), .C(n854), .D(n1310), .Y(n634));
INVX1    g691(.A(n634), .Y(n1312));
NOR3X1   g692(.A(n1312), .B(n1301), .C(n667), .Y(n444));
AND2X1   g693(.A(n2440gat), .B(n2394gat), .Y(n1314));
NOR3X1   g694(.A(n1312), .B(n1301), .C(n1314), .Y(n449));
NOR3X1   g695(.A(n1312), .B(n1301), .C(n665), .Y(n454));
NOR2X1   g696(.A(n1312), .B(n1301), .Y(n459));
NOR3X1   g697(.A(n1312), .B(n1301), .C(n658), .Y(n464));
INVX1    g698(.A(n1740gat), .Y(n1319));
AND2X1   g699(.A(n509), .B(n1319), .Y(n1320));
NAND4X1  g700(.A(n1850gat), .B(n646), .C(n2143gat), .D(n647), .Y(n1321));
NOR3X1   g701(.A(n509), .B(n2091gat), .C(n1496gat), .Y(n1322));
AND2X1   g702(.A(n509), .B(n1740gat), .Y(n1323));
NOR4X1   g703(.A(n1322), .B(n1321), .C(n1320), .D(n1323), .Y(n1324));
NAND2X1  g704(.A(n2061gat), .B(n2143gat), .Y(n1325));
NOR4X1   g705(.A(n1850gat), .B(n1899gat), .C(n1192), .D(n1325), .Y(n1326));
AND2X1   g706(.A(n1326), .B(n1320), .Y(n1327));
NAND2X1  g707(.A(n1850gat), .B(n2139gat), .Y(n1328));
OR4X1    g708(.A(n1899gat), .B(n2061gat), .C(n644_1), .D(n1328), .Y(n1329));
NOR4X1   g709(.A(n509), .B(n2091gat), .C(n1496gat), .D(n1329), .Y(n1330));
NAND4X1  g710(.A(n1850gat), .B(n646), .C(n644_1), .D(n647), .Y(n1331));
NOR3X1   g711(.A(n1331), .B(n1036), .C(n1319), .Y(n1332));
NOR4X1   g712(.A(n1330), .B(n1327), .C(n1324), .D(n1332), .Y(n1333));
AND2X1   g713(.A(n1333), .B(n634), .Y(n469));
INVX1    g714(.A(n469), .Y(n1335));
AOI21X1  g715(.A0(n1899gat), .A1(n2139gat), .B0(n1335), .Y(n474));
NOR2X1   g716(.A(n1335), .B(n1190), .Y(n479));
NOR2X1   g717(.A(n1335), .B(n630), .Y(n484));
NOR2X1   g718(.A(n1335), .B(n649_1), .Y(n489));
NOR2X1   g719(.A(n2454gat), .B(n271gat), .Y(n494));
INVX1    g720(.A(n2117gat), .Y(n1341));
AOI21X1  g721(.A0(n2446gat), .A1(n2450gat), .B0(n3100gat), .Y(n1342));
NOR3X1   g722(.A(n1342), .B(n1341), .C(n2125gat), .Y(n499));
INVX1    g723(.A(n494), .Y(n1344));
NOR4X1   g724(.A(n1344), .B(n1051), .C(n250), .D(n1342), .Y(n504));
NOR3X1   g725(.A(n626), .B(n3088gat), .C(n621), .Y(n1346));
NOR3X1   g726(.A(n626), .B(n641), .C(n631), .Y(n1347));
NOR4X1   g727(.A(n635), .B(n631), .C(n650), .D(n637), .Y(n1348));
AOI22X1  g728(.A0(n1347), .A1(n1346), .B0(n633), .B1(n1348), .Y(n1349));
OR2X1    g729(.A(n2155gat), .B(n2490gat), .Y(n1350));
NAND4X1  g730(.A(n2630gat), .B(n684), .C(n2626gat), .D(n679), .Y(n1351));
NAND2X1  g731(.A(n2155gat), .B(n2490gat), .Y(n1352));
NAND3X1  g732(.A(n1022), .B(n684), .C(n694), .Y(n1353));
OAI22X1  g733(.A0(n1352), .A1(n1353), .B0(n1351), .B1(n1350), .Y(n1354));
NAND4X1  g734(.A(n1026), .B(n1020), .C(n719), .D(n1354), .Y(n1355));
OAI22X1  g735(.A0(n1349), .A1(n1204), .B0(n1054), .B1(n1355), .Y(n514));
OAI22X1  g736(.A0(n1349), .A1(n1207), .B0(n1054), .B1(n1355), .Y(n519));
OAI22X1  g737(.A0(n1349), .A1(n1210), .B0(n1054), .B1(n1355), .Y(n524));
OAI22X1  g738(.A0(n1349), .A1(n1213), .B0(n1054), .B1(n1355), .Y(n529));
OAI22X1  g739(.A0(n1349), .A1(n1196), .B0(n1054), .B1(n1355), .Y(n534));
OAI22X1  g740(.A0(n1349), .A1(n1219), .B0(n1054), .B1(n1355), .Y(n539));
OAI22X1  g741(.A0(n1349), .A1(n1222), .B0(n1054), .B1(n1355), .Y(n544));
OAI22X1  g742(.A0(n1349), .A1(n1225), .B0(n1054), .B1(n1355), .Y(n549));
OAI22X1  g743(.A0(n1349), .A1(n1216), .B0(n1054), .B1(n1355), .Y(n554));
OAI21X1  g744(.A0(n1355), .A1(n1054), .B0(n3095gat), .Y(n1365));
NOR2X1   g745(.A(n1355), .B(n1054), .Y(n1366));
AOI21X1  g746(.A0(n3093gat), .A1(n3073gat), .B0(n1366), .Y(n1367));
OAI21X1  g747(.A0(n1365), .A1(n1217), .B0(n1367), .Y(n564));
OAI21X1  g748(.A0(n1355), .A1(n1054), .B0(n3093gat), .Y(n1369));
AOI21X1  g749(.A0(n3095gat), .A1(n3074gat), .B0(n1366), .Y(n1370));
OAI21X1  g750(.A0(n1369), .A1(n1204), .B0(n1370), .Y(n569));
AOI21X1  g751(.A0(n3095gat), .A1(n3076gat), .B0(n1366), .Y(n1372));
OAI21X1  g752(.A0(n1369), .A1(n1207), .B0(n1372), .Y(n574));
AOI21X1  g753(.A0(n3093gat), .A1(n3066gat), .B0(n1366), .Y(n1374));
OAI21X1  g754(.A0(n1365), .A1(n1211), .B0(n1374), .Y(n579));
AOI21X1  g755(.A0(n3095gat), .A1(n3080gat), .B0(n1366), .Y(n1376));
OAI21X1  g756(.A0(n1369), .A1(n1213), .B0(n1376), .Y(n584));
AOI21X1  g757(.A0(n3093gat), .A1(n3072gat), .B0(n1366), .Y(n1378));
OAI21X1  g758(.A0(n1365), .A1(n1197), .B0(n1378), .Y(n589));
AOI21X1  g759(.A0(n3095gat), .A1(n3077gat), .B0(n1366), .Y(n1380));
OAI21X1  g760(.A0(n1369), .A1(n1219), .B0(n1380), .Y(n594));
AOI21X1  g761(.A0(n3093gat), .A1(n3070gat), .B0(n1366), .Y(n1382));
OAI21X1  g762(.A0(n1365), .A1(n1223), .B0(n1382), .Y(n599));
AOI21X1  g763(.A0(n3093gat), .A1(n3069gat), .B0(n1366), .Y(n1384));
OAI21X1  g764(.A0(n1365), .A1(n1226), .B0(n1384), .Y(n604));
INVX1    g765(.A(n2518gat), .Y(n1386));
NAND4X1  g766(.A(n2526gat), .B(n2468gat), .C(n2476gat), .D(n2464gat), .Y(n1387));
NAND2X1  g767(.A(n2599gat), .B(n2522gat), .Y(n1388));
OR4X1    g768(.A(n1387), .B(n1386), .C(n3090gat), .D(n1388), .Y(n614));
OAI21X1  g769(.A0(n2394gat), .A1(n662), .B0(n1298), .Y(n1390));
OR2X1    g770(.A(n1390), .B(n657), .Y(n1391));
XOR2X1   g771(.A(n1391), .B(n2644gat), .Y(n1392));
NAND2X1  g772(.A(n1392), .B(n459), .Y(n619));
INVX1    g773(.A(n2190gat), .Y(n1394));
OR2X1    g774(.A(n2262gat), .B(n1394), .Y(n1395));
XOR2X1   g775(.A(n1395), .B(n2266gat), .Y(n1396));
NAND2X1  g776(.A(n1396), .B(n634), .Y(n629));
AOI21X1  g777(.A0(n2262gat), .A1(n2190gat), .B0(n1312), .Y(n639));
NOR2X1   g778(.A(n1312), .B(n672), .Y(n644));
OAI21X1  g779(.A0(n2139gat), .A1(n646), .B0(n1193), .Y(n1400));
NOR2X1   g780(.A(n1400), .B(n629_1), .Y(n1401));
XOR2X1   g781(.A(n1401), .B(n1975gat), .Y(n1402));
OR2X1    g782(.A(n1402), .B(n1335), .Y(n654));
NOR4X1   g783(.A(n2454gat), .B(n703gat), .C(n757), .D(n1027), .Y(n664));
NOR3X1   g784(.A(n1030), .B(n1011), .C(n2454gat), .Y(n669));
NAND2X1  g785(.A(n1326), .B(n509), .Y(n1406));
OR2X1    g786(.A(n1321), .B(n509), .Y(n1407));
OR2X1    g787(.A(n2347gat), .B(n2403gat), .Y(n1408));
OR4X1    g788(.A(n1295), .B(n1298), .C(n2394gat), .D(n1408), .Y(n1409));
AOI21X1  g789(.A0(n1407), .A1(n1406), .B0(n1409), .Y(n729));
INVX1    g790(.A(n664), .Y(n1411));
INVX1    g791(.A(n669), .Y(n1412));
NAND3X1  g792(.A(n1412), .B(n1411), .C(n1034_1), .Y(n734));
NAND3X1  g793(.A(n1850gat), .B(n1193), .C(n2139gat), .Y(n1414));
AND2X1   g794(.A(n2347gat), .B(n2394gat), .Y(n1415));
NAND4X1  g795(.A(n1295), .B(n2440gat), .C(n2403gat), .D(n1415), .Y(n1416));
NOR3X1   g796(.A(n1416), .B(n1414), .C(n1325), .Y(n739));
INVX1    g797(.A(n1054), .Y(n749));
NAND4X1  g798(.A(n1850gat), .B(n2061gat), .C(n2143gat), .D(n647), .Y(n1419));
NOR2X1   g799(.A(n1419), .B(n1409), .Y(n754));
INVX1    g800(.A(n1332gat), .Y(n759));
INVX1    g801(.A(n1017), .Y(n764));
OR2X1    g802(.A(n1033), .B(n1031), .Y(n784));
NOR4X1   g803(.A(n2135gat), .B(n2190gat), .C(n2179gat), .D(n2262gat), .Y(n1424));
NAND2X1  g804(.A(n1424), .B(n1301), .Y(n1425));
INVX1    g805(.A(n2182gat), .Y(n1426));
NAND2X1  g806(.A(n1301), .B(n1426), .Y(n1427));
AOI21X1  g807(.A0(n1427), .A1(n1425), .B0(n1333), .Y(n789));
INVX1    g808(.A(n1433gat), .Y(n794));
INVX1    g809(.A(n1316gat), .Y(n799));
INVX1    g810(.A(n1363gat), .Y(n804));
NOR4X1   g811(.A(n1342), .B(n1051), .C(n250), .D(n1412), .Y(n809));
OAI22X1  g812(.A0(n1321), .A1(n1144), .B0(n1040), .B1(n1406), .Y(n1433));
INVX1    g813(.A(n1433), .Y(n1434));
NOR3X1   g814(.A(n919gat), .B(n402gat), .C(n831), .Y(n1435));
NOR2X1   g815(.A(n846gat), .B(n831), .Y(n1436));
NAND4X1  g816(.A(n1435), .B(n661), .C(n1295), .D(n1436), .Y(n1437));
NAND2X1  g817(.A(n2440gat), .B(n2394gat), .Y(n1438));
NOR4X1   g818(.A(n2347gat), .B(n2407gat), .C(n662), .D(n1438), .Y(n1439));
NAND2X1  g819(.A(n2347gat), .B(n662), .Y(n1440));
NAND3X1  g820(.A(n837), .B(n919gat), .C(n398gat), .Y(n1441));
NAND3X1  g821(.A(n1295), .B(n828), .C(n398gat), .Y(n1442));
NOR4X1   g822(.A(n1441), .B(n1294), .C(n1440), .D(n1442), .Y(n1443));
OAI21X1  g823(.A0(n1443), .A1(n1439), .B0(n1433), .Y(n1444));
OAI21X1  g824(.A0(n1437), .A1(n1434), .B0(n1444), .Y(n1445));
NAND3X1  g825(.A(n1295), .B(n840), .C(n398gat), .Y(n1446));
NAND3X1  g826(.A(n663), .B(n2347gat), .C(n2403gat), .Y(n1447));
NAND3X1  g827(.A(n837), .B(n402gat), .C(n398gat), .Y(n1448));
NOR3X1   g828(.A(n1448), .B(n1447), .C(n1446), .Y(n1449));
NAND3X1  g829(.A(n2347gat), .B(n1295), .C(n662), .Y(n1450));
NOR3X1   g830(.A(n1450), .B(n1436), .C(n1299), .Y(n1451));
AND2X1   g831(.A(n1451), .B(n1435), .Y(n1452));
OAI21X1  g832(.A0(n1452), .A1(n1449), .B0(n1433), .Y(n1453));
NOR2X1   g833(.A(n402gat), .B(n831), .Y(n1454));
NAND4X1  g834(.A(n2440gat), .B(n1293), .C(n2403gat), .D(n2347gat), .Y(n1455));
NOR4X1   g835(.A(n1441), .B(n1454), .C(n2407gat), .D(n1455), .Y(n1456));
AOI21X1  g836(.A0(n846gat), .A1(n919gat), .B0(n831), .Y(n1457));
NOR4X1   g837(.A(n1442), .B(n1438), .C(n1440), .D(n1457), .Y(n1458));
OAI21X1  g838(.A0(n1458), .A1(n1456), .B0(n1433), .Y(n1459));
NAND4X1  g839(.A(n1295), .B(n2403gat), .C(n398gat), .D(n2347gat), .Y(n1460));
NOR4X1   g840(.A(n1457), .B(n1438), .C(n1454), .D(n1460), .Y(n1461));
NAND4X1  g841(.A(n1298), .B(n2394gat), .C(n2403gat), .D(n2347gat), .Y(n1462));
NOR4X1   g842(.A(n1446), .B(n1436), .C(n1454), .D(n1462), .Y(n1463));
OAI21X1  g843(.A0(n1463), .A1(n1461), .B0(n1433), .Y(n1464));
NAND3X1  g844(.A(n1464), .B(n1459), .C(n1453), .Y(n1465));
OAI21X1  g845(.A0(n819), .A1(n1312gat), .B0(n1309), .Y(n1466));
NOR4X1   g846(.A(n1465), .B(n1445), .C(n1308), .D(n1466), .Y(n814));
NOR4X1   g847(.A(n1036), .B(n646), .C(n2143gat), .D(n1414), .Y(n824));
NOR4X1   g848(.A(n1193), .B(n2061gat), .C(n644_1), .D(n1328), .Y(n829));
ONE      g849(.Y(n834));
OR2X1    g850(.A(n1306), .B(n1305), .Y(n844));
NAND4X1  g851(.A(n633), .B(n3086gat), .C(n3085gat), .D(n1259), .Y(n1472));
NAND4X1  g852(.A(n625), .B(n3088gat), .C(n3087gat), .D(n1347), .Y(n1473));
NAND2X1  g853(.A(n1473), .B(n1472), .Y(n849));
INVX1    g854(.A(n1312gat), .Y(n1475));
OR2X1    g855(.A(n1465), .B(n1445), .Y(n1476));
NOR4X1   g856(.A(n1308), .B(n2169gat), .C(n1475), .D(n1476), .Y(n864));
NOR3X1   g857(.A(n2040gat), .B(n1775gat), .C(n1316gat), .Y(n874));
INVX1    g858(.A(n2044gat), .Y(n879));
AOI21X1  g859(.A0(n2021gat), .A1(n1880gat), .B0(n1476), .Y(n884));
INVX1    g860(.A(n2025gat), .Y(n889));
INVX1    g861(.A(n2495gat), .Y(n894));
INVX1    g862(.A(n2033gat), .Y(n904));
INVX1    g863(.A(n2125gat), .Y(n914));
INVX1    g864(.A(n2121gat), .Y(n919));
INVX1    g865(.A(n2592gat), .Y(n984));
INVX1    g866(.A(n2458gat), .Y(n989));
NOR4X1   g867(.A(n1342), .B(n1051), .C(n250), .D(n1411), .Y(n994));
NOR4X1   g868(.A(n1023), .B(n2207gat), .C(n724), .D(n1089), .Y(n999));
NOR3X1   g869(.A(n1465), .B(n1445), .C(n1321), .Y(n1004));
INVX1    g870(.A(n1329), .Y(n1009));
INVX1    g871(.A(n1331), .Y(n1014));
NOR4X1   g872(.A(n1295), .B(n1298), .C(n2394gat), .D(n1408), .Y(n1493));
AND2X1   g873(.A(n829), .B(n1493), .Y(n1019));
NOR4X1   g874(.A(n1445), .B(n1406), .C(n1297), .D(n1465), .Y(n1024));
NAND3X1  g875(.A(n1850gat), .B(n2061gat), .C(n2143gat), .Y(n1496));
NOR3X1   g876(.A(n1496), .B(n1193), .C(n2139gat), .Y(n1029));
NOR4X1   g877(.A(n1299), .B(n1408), .C(n1295), .D(n1331), .Y(n1034));
NOR4X1   g878(.A(n1299), .B(n1408), .C(n1295), .D(n1321), .Y(n1039));
NOR3X1   g879(.A(n1414), .B(n1325), .C(n1475), .Y(n1044));
NAND3X1  g880(.A(n1062), .B(n1056), .C(n1043), .Y(n3140gat));
NAND4X1  g881(.A(n1074), .B(n1072), .C(n1066), .D(n1075), .Y(n3142gat));
BUFX1    g882(.A(n3069gat), .Y(n174));
BUFX1    g883(.A(n3070gat), .Y(n179));
BUFX1    g884(.A(n3072gat), .Y(n184));
BUFX1    g885(.A(n3071gat), .Y(n189));
BUFX1    g886(.A(n3069gat), .Y(n193));
BUFX1    g887(.A(n3070gat), .Y(n197));
BUFX1    g888(.A(n3072gat), .Y(n201));
BUFX1    g889(.A(n3071gat), .Y(n205));
BUFX1    g890(.A(n3065gat), .Y(n215));
BUFX1    g891(.A(n3067gat), .Y(n220));
BUFX1    g892(.A(n3066gat), .Y(n225));
BUFX1    g893(.A(n3073gat), .Y(n230));
BUFX1    g894(.A(n3068gat), .Y(n235));
NOR2X1   g895(.A(n1201), .B(n3099gat), .Y(n259));
BUFX1    g896(.A(n3065gat), .Y(n273));
BUFX1    g897(.A(n3067gat), .Y(n277));
BUFX1    g898(.A(n3066gat), .Y(n281));
BUFX1    g899(.A(n3073gat), .Y(n285));
BUFX1    g900(.A(n3068gat), .Y(n289));
OAI22X1  g901(.A0(n632), .A1(n1196), .B0(n1197), .B1(n622), .Y(n323));
BUFX1    g902(.A(n3070gat), .Y(n347));
BUFX1    g903(.A(n3069gat), .Y(n351));
BUFX1    g904(.A(n3071gat), .Y(n355));
BUFX1    g905(.A(n3072gat), .Y(n359));
NAND3X1  g906(.A(n1767gat), .B(n1834gat), .C(n1880gat), .Y(n674));
INVX1    g907(.A(n2270gat), .Y(n769));
INVX1    g908(.A(n2339gat), .Y(n774));
INVX1    g909(.A(n2390gat), .Y(n779));
endmodule
