//Converted to Combinational (Partial output: n510) , Module name: s15850_n510 , Timestamp: 2018-12-03T15:51:04.849239 
module s15850_n510 ( g599, g591, g605, g611, g695, g731, g617, g722, g700, g627, g639, g677, g686, g668, g658, g654, g646, g650, g643, g713, g704, n510 );
input g599, g591, g605, g611, g695, g731, g617, g722, g700, g627, g639, g677, g686, g668, g658, g654, g646, g650, g643, g713, g704;
output n510;
wire n2478, n2473, n2516, n2477, n2474, n2462, n2475_1, n2472, n2446, n2515_1, n2448, n2476, n2437, n2442, n2465_1, n2471, n2445_1, n2514, n2441, n2434, n2438, n2464, n2452, n2453, n2470_1, n2466, n2467, n2454, n2444, n2513, n2511, n2439, n2440_1, n2433, n2435, n2436_1, n2463, n2469, n2443, n2512, n2468, n2431_1, n2432, n2450_1, n2430, n2449;
OAI21X1  g0677(.A0(n2516), .A1(n2473), .B0(n2478), .Y(n510));
OR4X1    g0638(.A(n2475_1), .B(n2462), .C(n2474), .D(n2477), .Y(n2478));
OR2X1    g0633(.A(n2472), .B(n2462), .Y(n2473));
MX2X1    g0676(.A(n2448), .B(n2515_1), .S0(n2446), .Y(n2516));
INVX1    g0637(.A(n2476), .Y(n2477));
NOR3X1   g0634(.A(n2437), .B(g591), .C(g599), .Y(n2474));
NOR4X1   g0622(.A(g591), .B(g599), .C(g611), .D(g605), .Y(n2462));
INVX1    g0635(.A(n2472), .Y(n2475_1));
AOI21X1  g0632(.A0(n2471), .A1(n2465_1), .B0(n2442), .Y(n2472));
NAND2X1  g0606(.A(n2445_1), .B(n2442), .Y(n2446));
XOR2X1   g0675(.A(n2514), .B(g695), .Y(n2515_1));
INVX1    g0608(.A(g695), .Y(n2448));
AOI21X1  g0636(.A0(n2437), .A1(g599), .B0(n2441), .Y(n2476));
INVX1    g0597(.A(g605), .Y(n2437));
OAI21X1  g0602(.A0(n2441), .A1(n2438), .B0(n2434), .Y(n2442));
OR4X1    g0625(.A(n2453), .B(n2452), .C(g731), .D(n2464), .Y(n2465_1));
OR4X1    g0631(.A(n2454), .B(n2467), .C(n2466), .D(n2470_1), .Y(n2471));
OAI21X1  g0605(.A0(n2444), .A1(g617), .B0(n2434), .Y(n2445_1));
MX2X1    g0674(.A(n2511), .B(n2513), .S0(n2445_1), .Y(n2514));
NOR3X1   g0601(.A(n2440_1), .B(g617), .C(n2439), .Y(n2441));
INVX1    g0594(.A(n2433), .Y(n2434));
AOI21X1  g0598(.A0(n2437), .A1(n2436_1), .B0(n2435), .Y(n2438));
OR2X1    g0624(.A(n2463), .B(g722), .Y(n2464));
NOR3X1   g0612(.A(g605), .B(g591), .C(n2436_1), .Y(n2452));
AOI21X1  g0613(.A0(n2437), .A1(n2440_1), .B0(g599), .Y(n2453));
INVX1    g0630(.A(n2469), .Y(n2470_1));
INVX1    g0626(.A(g722), .Y(n2466));
INVX1    g0627(.A(g731), .Y(n2467));
NOR2X1   g0614(.A(n2453), .B(n2452), .Y(n2454));
NOR4X1   g0604(.A(n2440_1), .B(g599), .C(g617), .D(n2443), .Y(n2444));
MX2X1    g0673(.A(n2468), .B(n2512), .S0(n2454), .Y(n2513));
INVX1    g0671(.A(g700), .Y(n2511));
INVX1    g0599(.A(g611), .Y(n2439));
INVX1    g0600(.A(g591), .Y(n2440_1));
NAND3X1  g0593(.A(n2432), .B(n2431_1), .C(g627), .Y(n2433));
INVX1    g0595(.A(g639), .Y(n2435));
INVX1    g0596(.A(g599), .Y(n2436_1));
NAND4X1  g0623(.A(n2449), .B(n2448), .C(n2430), .D(n2450_1), .Y(n2463));
NOR4X1   g0629(.A(n2449), .B(n2448), .C(n2430), .D(n2468), .Y(n2469));
OR2X1    g0603(.A(g605), .B(g611), .Y(n2443));
INVX1    g0672(.A(n2450_1), .Y(n2512));
NAND4X1  g0628(.A(g658), .B(g668), .C(g686), .D(g677), .Y(n2468));
INVX1    g0591(.A(g654), .Y(n2431_1));
NOR3X1   g0592(.A(g643), .B(g650), .C(g646), .Y(n2432));
NOR4X1   g0610(.A(g658), .B(g668), .C(g686), .D(g677), .Y(n2450_1));
INVX1    g0590(.A(g713), .Y(n2430));
INVX1    g0609(.A(g704), .Y(n2449));

endmodule
