//Converted to Combinational , Module name: s1423 , Timestamp: 2018-12-03T15:51:02.400016 
module s1423 ( G0, G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G40, G41, G42, G43, G44, G45, G46, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G58, G59, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G70, G71, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G83, G84, G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G726, G729, G702, G727, G701BF, n45, n50, n55, n60, n65, n70, n75, n80, n85, n90, n95, n100, n105, n110, n115, n120, n125, n130, n135, n140, n145, n150, n155, n160, n165, n170, n175, n180, n185, n190, n195, n200, n205, n210, n215, n220, n225, n230, n235, n240, n245, n250, n255, n260, n265, n270, n275, n280, n285, n290, n295, n300, n305, n310, n315, n320, n325, n330, n335, n340, n345, n350, n355, n360, n365, n370, n375, n380, n385, n390, n395, n400, n405, n410 );
input G0, G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G40, G41, G42, G43, G44, G45, G46, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G58, G59, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G70, G71, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G83, G84, G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95;
output G726, G729, G702, G727, G701BF, n45, n50, n55, n60, n65, n70, n75, n80, n85, n90, n95, n100, n105, n110, n115, n120, n125, n130, n135, n140, n145, n150, n155, n160, n165, n170, n175, n180, n185, n190, n195, n200, n205, n210, n215, n220, n225, n230, n235, n240, n245, n250, n255, n260, n265, n270, n275, n280, n285, n290, n295, n300, n305, n310, n315, n320, n325, n330, n335, n340, n345, n350, n355, n360, n365, n370, n375, n380, n385, n390, n395, n400, n405, n410;
wire n244, n245_1, n246, n247, n248, n249, n250_1, n251, n252, n253, n254, n255_1, n256, n257, n258, n259, n260_1, n261, n262, n263, n264, n265_1, n266, n267, n268, n269, n270_1, n271, n272, n273, n274, n275_1, n276, n277, n278, n279, n280_1, n281, n282, n283, n284, n285_1, n286, n287, n288, n289, n290_1, n291, n292, n293, n294, n295_1, n296, n297, n298, n299, n300_1, n301, n302, n303, n304, n305_1, n306, n307, n308, n309, n310_1, n311, n312, n313, n314, n315_1, n316, n317, n318, n319, n320_1, n321, n322, n323, n324, n325_1, n326, n327, n328, n329, n331, n332, n333, n334, n335_1, n336, n337, n338, n339, n342, n343, n344, n345_1, n346, n347, n348, n349, n350_1, n351, n353, n354, n355_1, n357, n359, n360_1, n361, n363, n365_1, n367, n368, n370_1, n371, n373, n374, n376, n377, n379, n381, n382, n384, n385_1, n388, n390_1, n391, n393, n395_1, n397, n398, n399, n401, n403, n404, n405_1, n406, n407, n409, n410_1, n412, n413, n415, n416, n418, n419, n421, n422, n423, n424, n426, n428, n430, n432, n433, n434, n435, n437, n438, n439, n441, n442, n444, n445, n446, n448, n449, n450, n452, n453, n455, n456, n458, n459, n460, n462, n463, n465, n466, n467, n469, n470, n471, n473, n475, n476, n477, n479, n480, n481, n483, n485, n486, n488, n489, n490, n491, n492, n494, n495, n497, n498, n499, n501, n503, n504, n506, n508, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n522, n523, n525, n526, n527, n529, n531, n532, n534, n539, n540, n545, n546, n548, n549, n551, n552, n554, n555, n557, n558, n559, n561, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n582, n584;
INVX1    g000(.A(G53), .Y(n244));
INVX1    g001(.A(G92), .Y(n245_1));
INVX1    g002(.A(G33), .Y(n246));
INVX1    g003(.A(G27), .Y(n247));
INVX1    g004(.A(G25), .Y(n248));
INVX1    g005(.A(G26), .Y(n249));
INVX1    g006(.A(G78), .Y(n250_1));
INVX1    g007(.A(G90), .Y(n251));
NAND2X1  g008(.A(G90), .B(G64), .Y(n252));
OR2X1    g009(.A(G90), .B(G8), .Y(n253));
AOI21X1  g010(.A0(n253), .A1(n252), .B0(G85), .Y(n254));
AND2X1   g011(.A(G90), .B(G64), .Y(n255_1));
NOR2X1   g012(.A(G90), .B(G8), .Y(n256));
NOR3X1   g013(.A(n256), .B(n255_1), .C(G84), .Y(n257));
OR4X1    g014(.A(n254), .B(n251), .C(n250_1), .D(n257), .Y(n258));
OR2X1    g015(.A(G90), .B(G4), .Y(n259));
AOI21X1  g016(.A0(n259), .A1(n258), .B0(G46), .Y(n260_1));
AND2X1   g017(.A(n259), .B(n258), .Y(n261));
XOR2X1   g018(.A(n261), .B(G46), .Y(n262));
INVX1    g019(.A(G77), .Y(n263));
OR4X1    g020(.A(n254), .B(n251), .C(n263), .D(n257), .Y(n264));
OR2X1    g021(.A(G90), .B(G3), .Y(n265_1));
AND2X1   g022(.A(n265_1), .B(n264), .Y(n266));
OR2X1    g023(.A(n266), .B(G45), .Y(n267));
INVX1    g024(.A(G45), .Y(n268));
XOR2X1   g025(.A(n266), .B(n268), .Y(n269));
INVX1    g026(.A(G76), .Y(n270_1));
OR4X1    g027(.A(n254), .B(n251), .C(n270_1), .D(n257), .Y(n271));
OR2X1    g028(.A(G90), .B(G2), .Y(n272));
AOI21X1  g029(.A0(n272), .A1(n271), .B0(G44), .Y(n273));
AND2X1   g030(.A(n272), .B(n271), .Y(n274));
XOR2X1   g031(.A(n274), .B(G44), .Y(n275_1));
INVX1    g032(.A(G43), .Y(n276));
NAND2X1  g033(.A(G90), .B(G75), .Y(n277));
NOR3X1   g034(.A(n277), .B(n257), .C(n254), .Y(n278));
NOR2X1   g035(.A(G90), .B(G1), .Y(n279));
OAI21X1  g036(.A0(n279), .A1(n278), .B0(n276), .Y(n280_1));
NOR3X1   g037(.A(n279), .B(n278), .C(n276), .Y(n281));
INVX1    g038(.A(G42), .Y(n282));
NAND2X1  g039(.A(G90), .B(G74), .Y(n283));
NOR3X1   g040(.A(n283), .B(n257), .C(n254), .Y(n284));
NOR2X1   g041(.A(G90), .B(G0), .Y(n285_1));
NOR3X1   g042(.A(n285_1), .B(n284), .C(n282), .Y(n286));
OAI21X1  g043(.A0(n286), .A1(n281), .B0(n280_1), .Y(n287));
AOI21X1  g044(.A0(n287), .A1(n275_1), .B0(n273), .Y(n288));
OAI21X1  g045(.A0(n288), .A1(n269), .B0(n267), .Y(n289));
AOI21X1  g046(.A0(n289), .A1(n262), .B0(n260_1), .Y(n290_1));
NOR4X1   g047(.A(n249), .B(n248), .C(G24), .D(n290_1), .Y(n291));
NAND3X1  g048(.A(n291), .B(G28), .C(n247), .Y(n292));
AOI21X1  g049(.A0(n292), .A1(G92), .B0(G29), .Y(n293));
NAND4X1  g050(.A(G32), .B(G31), .C(G30), .D(n293), .Y(n294));
NOR3X1   g051(.A(n294), .B(G34), .C(n246), .Y(n295_1));
NOR2X1   g052(.A(n295_1), .B(n245_1), .Y(n296));
INVX1    g053(.A(n296), .Y(n297));
INVX1    g054(.A(G37), .Y(n298));
INVX1    g055(.A(G38), .Y(n299));
INVX1    g056(.A(G36), .Y(n300_1));
INVX1    g057(.A(G91), .Y(n301));
INVX1    g058(.A(G41), .Y(n302));
NOR4X1   g059(.A(n302), .B(G40), .C(G39), .D(n296), .Y(n303));
OAI21X1  g060(.A0(n303), .A1(n301), .B0(n300_1), .Y(n304));
NOR3X1   g061(.A(n304), .B(n299), .C(n298), .Y(n305_1));
INVX1    g062(.A(G16), .Y(n306));
INVX1    g063(.A(G83), .Y(n307));
NOR4X1   g064(.A(G81), .B(G80), .C(G79), .D(G82), .Y(n308));
XOR2X1   g065(.A(n308), .B(G78), .Y(n309));
XOR2X1   g066(.A(G81), .B(G76), .Y(n310_1));
XOR2X1   g067(.A(G79), .B(G74), .Y(n311));
XOR2X1   g068(.A(G80), .B(G75), .Y(n312));
XOR2X1   g069(.A(G82), .B(G77), .Y(n313));
NOR4X1   g070(.A(n312), .B(n311), .C(n310_1), .D(n313), .Y(n314));
INVX1    g071(.A(n314), .Y(n315_1));
NOR2X1   g072(.A(n315_1), .B(n309), .Y(n316));
NAND2X1  g073(.A(n316), .B(n307), .Y(n317));
NOR3X1   g074(.A(n317), .B(G66), .C(n306), .Y(n318));
NOR2X1   g075(.A(n318), .B(n251), .Y(n319));
MX2X1    g076(.A(n297), .B(n305_1), .S0(n319), .Y(n320_1));
NAND3X1  g077(.A(n320_1), .B(G59), .C(G58), .Y(n321));
AOI21X1  g078(.A0(n321), .A1(G91), .B0(n244), .Y(n322));
NAND3X1  g079(.A(n322), .B(G62), .C(G61), .Y(n323));
INVX1    g080(.A(n323), .Y(n324));
INVX1    g081(.A(G88), .Y(n325_1));
INVX1    g082(.A(n303), .Y(n326));
OAI21X1  g083(.A0(n292), .A1(G94), .B0(n251), .Y(n327));
AOI21X1  g084(.A0(n295_1), .A1(G87), .B0(n327), .Y(n328));
OAI21X1  g085(.A0(n326), .A1(n325_1), .B0(n328), .Y(n329));
AOI21X1  g086(.A0(n324), .A1(G89), .B0(n329), .Y(G702));
INVX1    g087(.A(G14), .Y(n331));
INVX1    g088(.A(G70), .Y(n332));
NOR3X1   g089(.A(G73), .B(G72), .C(G71), .Y(n333));
XOR2X1   g090(.A(n333), .B(n332), .Y(n334));
XOR2X1   g091(.A(G71), .B(G67), .Y(n335_1));
XOR2X1   g092(.A(G73), .B(G69), .Y(n336));
XOR2X1   g093(.A(G72), .B(G68), .Y(n337));
NOR3X1   g094(.A(n337), .B(n336), .C(n335_1), .Y(n338));
AOI21X1  g095(.A0(n338), .A1(n334), .B0(n331), .Y(n339));
NOR2X1   g096(.A(n339), .B(G90), .Y(G727));
INVX1    g097(.A(G15), .Y(G701BF));
INVX1    g098(.A(G22), .Y(n342));
INVX1    g099(.A(G47), .Y(n343));
INVX1    g100(.A(G48), .Y(n344));
INVX1    g101(.A(G49), .Y(n345_1));
INVX1    g102(.A(G50), .Y(n346));
NOR4X1   g103(.A(n345_1), .B(n344), .C(n343), .D(n346), .Y(n347));
INVX1    g104(.A(n347), .Y(n348));
NOR2X1   g105(.A(G50), .B(G15), .Y(n349));
NOR3X1   g106(.A(G49), .B(G48), .C(G47), .Y(n350_1));
AND2X1   g107(.A(n350_1), .B(n349), .Y(n351));
OAI22X1  g108(.A0(n348), .A1(G15), .B0(n342), .B1(n351), .Y(n45));
INVX1    g109(.A(G23), .Y(n353));
NOR2X1   g110(.A(G22), .B(G701BF), .Y(n354));
NAND2X1  g111(.A(G22), .B(G15), .Y(n355_1));
AOI21X1  g112(.A0(n355_1), .A1(n353), .B0(n354), .Y(n50));
XOR2X1   g113(.A(n290_1), .B(G24), .Y(n357));
NOR2X1   g114(.A(n357), .B(n331), .Y(n55));
NOR3X1   g115(.A(n290_1), .B(n248), .C(G24), .Y(n359));
NOR2X1   g116(.A(n290_1), .B(G24), .Y(n360_1));
OAI21X1  g117(.A0(n360_1), .A1(G25), .B0(G14), .Y(n361));
NOR2X1   g118(.A(n361), .B(n359), .Y(n60));
OAI21X1  g119(.A0(n359), .A1(G26), .B0(G14), .Y(n363));
NOR2X1   g120(.A(n363), .B(n291), .Y(n65));
XOR2X1   g121(.A(n291), .B(n247), .Y(n365_1));
NOR2X1   g122(.A(n365_1), .B(n331), .Y(n70));
AOI21X1  g123(.A0(n291), .A1(n247), .B0(G28), .Y(n367));
NOR2X1   g124(.A(n367), .B(n331), .Y(n368));
AND2X1   g125(.A(n368), .B(n292), .Y(n75));
AND2X1   g126(.A(n292), .B(G92), .Y(n370_1));
XOR2X1   g127(.A(n370_1), .B(G29), .Y(n371));
NOR2X1   g128(.A(n371), .B(n331), .Y(n80));
AND2X1   g129(.A(n293), .B(G30), .Y(n373));
OAI21X1  g130(.A0(n293), .A1(G30), .B0(G14), .Y(n374));
NOR2X1   g131(.A(n374), .B(n373), .Y(n85));
AND2X1   g132(.A(n373), .B(G31), .Y(n376));
AOI21X1  g133(.A0(n293), .A1(G30), .B0(G31), .Y(n377));
NOR3X1   g134(.A(n377), .B(n376), .C(n331), .Y(n90));
OAI21X1  g135(.A0(n376), .A1(G32), .B0(G14), .Y(n379));
AOI21X1  g136(.A0(n376), .A1(G32), .B0(n379), .Y(n95));
NOR2X1   g137(.A(n294), .B(n246), .Y(n381));
AND2X1   g138(.A(n294), .B(n246), .Y(n382));
NOR3X1   g139(.A(n382), .B(n381), .C(n331), .Y(n100));
INVX1    g140(.A(G34), .Y(n384));
XOR2X1   g141(.A(n381), .B(n384), .Y(n385_1));
NOR2X1   g142(.A(n385_1), .B(n331), .Y(n105));
NOR2X1   g143(.A(G35), .B(n331), .Y(n110));
NAND3X1  g144(.A(n326), .B(G91), .C(G36), .Y(n388));
AOI21X1  g145(.A0(n388), .A1(n304), .B0(n331), .Y(n115));
INVX1    g146(.A(n304), .Y(n390_1));
OAI21X1  g147(.A0(n390_1), .A1(G37), .B0(G14), .Y(n391));
AOI21X1  g148(.A0(n390_1), .A1(G37), .B0(n391), .Y(n120));
AOI21X1  g149(.A0(n390_1), .A1(G37), .B0(G38), .Y(n393));
NOR3X1   g150(.A(n393), .B(n305_1), .C(n331), .Y(n125));
XOR2X1   g151(.A(n296), .B(G39), .Y(n395_1));
NOR2X1   g152(.A(n395_1), .B(n331), .Y(n130));
INVX1    g153(.A(G40), .Y(n397));
NOR2X1   g154(.A(n296), .B(G39), .Y(n398));
XOR2X1   g155(.A(n398), .B(n397), .Y(n399));
NOR2X1   g156(.A(n399), .B(n331), .Y(n135));
AOI21X1  g157(.A0(n398), .A1(n397), .B0(G41), .Y(n401));
NOR3X1   g158(.A(n401), .B(n303), .C(n331), .Y(n140));
NOR3X1   g159(.A(n50), .B(n348), .C(n282), .Y(n403));
NOR2X1   g160(.A(n50), .B(n348), .Y(n404));
NOR2X1   g161(.A(n404), .B(G42), .Y(n405_1));
INVX1    g162(.A(n339), .Y(n406));
MX2X1    g163(.A(G7), .B(n406), .S0(G90), .Y(n407));
NOR3X1   g164(.A(n407), .B(n405_1), .C(n403), .Y(n145));
NOR2X1   g165(.A(n403), .B(G43), .Y(n409));
NOR4X1   g166(.A(n348), .B(n276), .C(n282), .D(n50), .Y(n410_1));
NOR3X1   g167(.A(n410_1), .B(n409), .C(n407), .Y(n150));
NOR2X1   g168(.A(n410_1), .B(G44), .Y(n412));
AND2X1   g169(.A(n410_1), .B(G44), .Y(n413));
NOR3X1   g170(.A(n413), .B(n412), .C(n407), .Y(n155));
AOI21X1  g171(.A0(n410_1), .A1(G44), .B0(G45), .Y(n415));
AND2X1   g172(.A(n413), .B(G45), .Y(n416));
NOR3X1   g173(.A(n416), .B(n415), .C(n407), .Y(n160));
OR2X1    g174(.A(n416), .B(G46), .Y(n418));
AOI21X1  g175(.A0(n416), .A1(G46), .B0(n407), .Y(n419));
AND2X1   g176(.A(n419), .B(n418), .Y(n165));
INVX1    g177(.A(G54), .Y(n421));
NOR2X1   g178(.A(n296), .B(n421), .Y(n422));
AOI21X1  g179(.A0(n422), .A1(G56), .B0(n301), .Y(n423));
OAI21X1  g180(.A0(n423), .A1(G12), .B0(G14), .Y(n424));
AOI21X1  g181(.A0(n423), .A1(n343), .B0(n424), .Y(n170));
OAI21X1  g182(.A0(n423), .A1(G47), .B0(G14), .Y(n426));
AOI21X1  g183(.A0(n423), .A1(n344), .B0(n426), .Y(n175));
OAI21X1  g184(.A0(n423), .A1(G48), .B0(G14), .Y(n428));
AOI21X1  g185(.A0(n423), .A1(n345_1), .B0(n428), .Y(n180));
OAI21X1  g186(.A0(n423), .A1(G49), .B0(G14), .Y(n430));
AOI21X1  g187(.A0(n423), .A1(n346), .B0(n430), .Y(n185));
NOR2X1   g188(.A(n322), .B(n331), .Y(n432));
INVX1    g189(.A(G51), .Y(n433));
AND2X1   g190(.A(n321), .B(G91), .Y(n434));
XOR2X1   g191(.A(n434), .B(n433), .Y(n435));
AND2X1   g192(.A(n435), .B(n432), .Y(n190));
AOI21X1  g193(.A0(n321), .A1(G91), .B0(n433), .Y(n437));
NOR2X1   g194(.A(n437), .B(G52), .Y(n438));
AND2X1   g195(.A(n437), .B(G52), .Y(n439));
NOR4X1   g196(.A(n438), .B(n322), .C(n331), .D(n439), .Y(n195));
AOI21X1  g197(.A0(n437), .A1(G52), .B0(G53), .Y(n441));
AND2X1   g198(.A(n439), .B(G53), .Y(n442));
NOR4X1   g199(.A(n441), .B(n322), .C(n331), .D(n442), .Y(n200));
INVX1    g200(.A(G56), .Y(n444));
NOR3X1   g201(.A(n296), .B(n444), .C(n421), .Y(n445));
XOR2X1   g202(.A(n296), .B(G54), .Y(n446));
NOR3X1   g203(.A(n446), .B(n445), .C(n331), .Y(n205));
OR2X1    g204(.A(n445), .B(n331), .Y(n448));
INVX1    g205(.A(G55), .Y(n449));
XOR2X1   g206(.A(n422), .B(n449), .Y(n450));
NOR2X1   g207(.A(n450), .B(n448), .Y(n210));
AOI21X1  g208(.A0(n422), .A1(G55), .B0(G56), .Y(n452));
NOR4X1   g209(.A(n444), .B(n449), .C(n421), .D(n296), .Y(n453));
NOR3X1   g210(.A(n453), .B(n452), .C(n448), .Y(n215));
AOI21X1  g211(.A0(n320_1), .A1(G58), .B0(n331), .Y(n455));
XOR2X1   g212(.A(n320_1), .B(G57), .Y(n456));
AND2X1   g213(.A(n456), .B(n455), .Y(n220));
AOI21X1  g214(.A0(n320_1), .A1(G57), .B0(G58), .Y(n458));
NAND3X1  g215(.A(n320_1), .B(G58), .C(G57), .Y(n459));
NAND2X1  g216(.A(n459), .B(n455), .Y(n460));
NOR2X1   g217(.A(n460), .B(n458), .Y(n225));
INVX1    g218(.A(n321), .Y(n462));
AOI21X1  g219(.A0(n320_1), .A1(G58), .B0(G59), .Y(n463));
NOR3X1   g220(.A(n463), .B(n462), .C(n331), .Y(n230));
AND2X1   g221(.A(n322), .B(G61), .Y(n465));
INVX1    g222(.A(G60), .Y(n466));
XOR2X1   g223(.A(n322), .B(n466), .Y(n467));
NOR3X1   g224(.A(n467), .B(n465), .C(n331), .Y(n235));
AOI21X1  g225(.A0(n322), .A1(G60), .B0(G61), .Y(n469));
INVX1    g226(.A(G61), .Y(n470));
NOR4X1   g227(.A(n470), .B(n466), .C(n244), .D(n434), .Y(n471));
NOR4X1   g228(.A(n469), .B(n465), .C(n331), .D(n471), .Y(n240));
AOI21X1  g229(.A0(n322), .A1(G61), .B0(G62), .Y(n473));
NOR3X1   g230(.A(n473), .B(n324), .C(n331), .Y(n245));
MX2X1    g231(.A(n384), .B(G35), .S0(n245_1), .Y(n475));
MX2X1    g232(.A(n475), .B(G38), .S0(n319), .Y(n476));
NOR2X1   g233(.A(n476), .B(G63), .Y(n477));
NOR2X1   g234(.A(n477), .B(n331), .Y(n250));
INVX1    g235(.A(G63), .Y(n479));
AND2X1   g236(.A(n338), .B(n334), .Y(n480));
OAI21X1  g237(.A0(n480), .A1(G64), .B0(G14), .Y(n481));
AOI21X1  g238(.A0(n480), .A1(n479), .B0(n481), .Y(n255));
AOI21X1  g239(.A0(n338), .A1(n334), .B0(G65), .Y(n483));
NOR2X1   g240(.A(n483), .B(n331), .Y(n260));
INVX1    g241(.A(G65), .Y(n485));
OAI21X1  g242(.A0(n480), .A1(G66), .B0(G14), .Y(n486));
AOI21X1  g243(.A0(n480), .A1(n485), .B0(n486), .Y(n265));
MX2X1    g244(.A(n321), .B(n323), .S0(G91), .Y(n488));
NAND2X1  g245(.A(n488), .B(G90), .Y(n489));
NOR2X1   g246(.A(n489), .B(G67), .Y(n490));
INVX1    g247(.A(G67), .Y(n491));
AOI21X1  g248(.A0(n488), .A1(G90), .B0(n491), .Y(n492));
NOR3X1   g249(.A(n492), .B(n490), .C(n406), .Y(n270));
OR2X1    g250(.A(n492), .B(G68), .Y(n494));
AOI21X1  g251(.A0(n492), .A1(G68), .B0(n406), .Y(n495));
AND2X1   g252(.A(n495), .B(n494), .Y(n275));
AOI21X1  g253(.A0(n492), .A1(G68), .B0(G69), .Y(n497));
NAND3X1  g254(.A(n492), .B(G69), .C(G68), .Y(n498));
NAND2X1  g255(.A(n498), .B(n339), .Y(n499));
NOR2X1   g256(.A(n499), .B(n497), .Y(n280));
OAI21X1  g257(.A0(n498), .A1(n332), .B0(n339), .Y(n501));
AOI21X1  g258(.A0(n498), .A1(n332), .B0(n501), .Y(n285));
OAI21X1  g259(.A0(n339), .A1(n251), .B0(G14), .Y(n503));
MX2X1    g260(.A(G0), .B(G3), .S0(G63), .Y(n504));
MX2X1    g261(.A(G71), .B(n504), .S0(n503), .Y(n290));
MX2X1    g262(.A(G1), .B(G4), .S0(G63), .Y(n506));
MX2X1    g263(.A(G72), .B(n506), .S0(n503), .Y(n295));
MX2X1    g264(.A(G2), .B(G5), .S0(G63), .Y(n508));
MX2X1    g265(.A(G73), .B(n508), .S0(n503), .Y(n300));
NAND3X1  g266(.A(n390_1), .B(n299), .C(G37), .Y(n510));
INVX1    g267(.A(n316), .Y(n511));
NOR3X1   g268(.A(n294), .B(n384), .C(n246), .Y(n512));
NOR2X1   g269(.A(n319), .B(n245_1), .Y(n513));
INVX1    g270(.A(n513), .Y(n514));
OAI21X1  g271(.A0(n514), .A1(n512), .B0(n511), .Y(n515));
AOI21X1  g272(.A0(n510), .A1(n319), .B0(n515), .Y(n516));
AND2X1   g273(.A(n516), .B(G74), .Y(n517));
MX2X1    g274(.A(G9), .B(n406), .S0(G90), .Y(n518));
INVX1    g275(.A(n518), .Y(n519));
OAI21X1  g276(.A0(n516), .A1(G74), .B0(n519), .Y(n520));
NOR2X1   g277(.A(n520), .B(n517), .Y(n305));
OR2X1    g278(.A(n517), .B(G75), .Y(n522));
AOI21X1  g279(.A0(n517), .A1(G75), .B0(n518), .Y(n523));
AND2X1   g280(.A(n523), .B(n522), .Y(n310));
AOI21X1  g281(.A0(n517), .A1(G75), .B0(G76), .Y(n525));
NAND4X1  g282(.A(G76), .B(G75), .C(G74), .D(n516), .Y(n526));
NAND2X1  g283(.A(n526), .B(n519), .Y(n527));
NOR2X1   g284(.A(n527), .B(n525), .Y(n315));
OAI21X1  g285(.A0(n526), .A1(n263), .B0(n519), .Y(n529));
AOI21X1  g286(.A0(n526), .A1(n263), .B0(n529), .Y(n320));
OR2X1    g287(.A(n526), .B(n263), .Y(n531));
OAI21X1  g288(.A0(n531), .A1(n250_1), .B0(n519), .Y(n532));
AOI21X1  g289(.A0(n531), .A1(n250_1), .B0(n532), .Y(n325));
OAI21X1  g290(.A0(n339), .A1(n301), .B0(G14), .Y(n534));
MX2X1    g291(.A(G79), .B(G6), .S0(n534), .Y(n330));
MX2X1    g292(.A(G80), .B(G7), .S0(n534), .Y(n335));
MX2X1    g293(.A(G81), .B(G8), .S0(n534), .Y(n340));
MX2X1    g294(.A(G82), .B(G9), .S0(n534), .Y(n345));
INVX1    g295(.A(n516), .Y(n539));
OAI21X1  g296(.A0(n476), .A1(n511), .B0(G83), .Y(n540));
AOI21X1  g297(.A0(n540), .A1(n539), .B0(n518), .Y(n350));
MX2X1    g298(.A(G84), .B(G10), .S0(n534), .Y(n355));
MX2X1    g299(.A(G85), .B(G11), .S0(n534), .Y(n360));
AND2X1   g300(.A(G14), .B(G13), .Y(n365));
NOR2X1   g301(.A(G87), .B(G11), .Y(n545));
AND2X1   g302(.A(G94), .B(G11), .Y(n546));
NOR3X1   g303(.A(n546), .B(n545), .C(n331), .Y(n370));
INVX1    g304(.A(G11), .Y(n548));
OAI21X1  g305(.A0(G87), .A1(n548), .B0(G14), .Y(n549));
AOI21X1  g306(.A0(n325_1), .A1(n548), .B0(n549), .Y(n375));
NOR2X1   g307(.A(G89), .B(G11), .Y(n551));
OAI21X1  g308(.A0(G88), .A1(n548), .B0(G14), .Y(n552));
NOR2X1   g309(.A(n552), .B(n551), .Y(n380));
INVX1    g310(.A(G13), .Y(n554));
OAI22X1  g311(.A0(G86), .A1(n554), .B0(G10), .B1(G90), .Y(n555));
NAND2X1  g312(.A(n555), .B(n365), .Y(n385));
NOR2X1   g313(.A(G86), .B(n554), .Y(n557));
INVX1    g314(.A(G10), .Y(n558));
MX2X1    g315(.A(n251), .B(n301), .S0(n558), .Y(n559));
OAI21X1  g316(.A0(n559), .A1(n557), .B0(n365), .Y(n390));
MX2X1    g317(.A(n301), .B(n245_1), .S0(n558), .Y(n561));
OAI21X1  g318(.A0(n561), .A1(n557), .B0(n365), .Y(n395));
MX2X1    g319(.A(G6), .B(n318), .S0(G90), .Y(n563));
MX2X1    g320(.A(G59), .B(G62), .S0(G91), .Y(n564));
MX2X1    g321(.A(G35), .B(n564), .S0(G90), .Y(n565));
NAND2X1  g322(.A(n565), .B(n563), .Y(n566));
NOR2X1   g323(.A(n285_1), .B(n284), .Y(n567));
XOR2X1   g324(.A(n567), .B(G42), .Y(n568));
NAND2X1  g325(.A(n568), .B(n275_1), .Y(n569));
NAND3X1  g326(.A(n265_1), .B(n264), .C(G45), .Y(n570));
NOR2X1   g327(.A(n279), .B(n278), .Y(n571));
XOR2X1   g328(.A(n571), .B(G43), .Y(n572));
NAND4X1  g329(.A(n570), .B(n267), .C(n262), .D(n572), .Y(n573));
NOR2X1   g330(.A(n573), .B(n569), .Y(n574));
NOR2X1   g331(.A(n574), .B(n290_1), .Y(n575));
NAND2X1  g332(.A(n574), .B(n476), .Y(n576));
MX2X1    g333(.A(G5), .B(n317), .S0(G90), .Y(n577));
AND2X1   g334(.A(n577), .B(n476), .Y(n578));
NOR3X1   g335(.A(n578), .B(n563), .C(n290_1), .Y(n579));
OAI21X1  g336(.A0(n576), .A1(n575), .B0(n579), .Y(n580));
AOI21X1  g337(.A0(n580), .A1(n566), .B0(n331), .Y(n400));
OAI21X1  g338(.A0(G94), .A1(G11), .B0(G14), .Y(n582));
AOI21X1  g339(.A0(G89), .A1(G11), .B0(n582), .Y(n405));
NOR4X1   g340(.A(n254), .B(n307), .C(n331), .D(n257), .Y(n584));
AND2X1   g341(.A(n584), .B(n476), .Y(n410));
BUFX1    g342(.A(G93), .Y(G726));
BUFX1    g343(.A(G95), .Y(G729));
endmodule
