// Benchmark "mem_ctrl" written by ABC on Mon Sep 21 04:04:28 2020

module mem_ctrl ( 
    pi0000, pi0001, pi0002, pi0003, pi0004, pi0005, pi0006, pi0007, pi0008,
    pi0009, pi0010, pi0011, pi0012, pi0013, pi0014, pi0015, pi0016, pi0017,
    pi0018, pi0019, pi0020, pi0021, pi0022, pi0023, pi0024, pi0025, pi0026,
    pi0027, pi0028, pi0029, pi0030, pi0031, pi0032, pi0033, pi0034, pi0035,
    pi0036, pi0037, pi0038, pi0039, pi0040, pi0041, pi0042, pi0043, pi0044,
    pi0045, pi0046, pi0047, pi0048, pi0049, pi0050, pi0051, pi0052, pi0053,
    pi0054, pi0055, pi0056, pi0057, pi0058, pi0059, pi0060, pi0061, pi0062,
    pi0063, pi0064, pi0065, pi0066, pi0067, pi0068, pi0069, pi0070, pi0071,
    pi0072, pi0073, pi0074, pi0075, pi0076, pi0077, pi0078, pi0079, pi0080,
    pi0081, pi0082, pi0083, pi0084, pi0085, pi0086, pi0087, pi0088, pi0089,
    pi0090, pi0091, pi0092, pi0093, pi0094, pi0095, pi0096, pi0097, pi0098,
    pi0099, pi0100, pi0101, pi0102, pi0103, pi0104, pi0105, pi0106, pi0107,
    pi0108, pi0109, pi0110, pi0111, pi0112, pi0113, pi0114, pi0115, pi0116,
    pi0117, pi0118, pi0119, pi0120, pi0121, pi0122, pi0123, pi0124, pi0125,
    pi0126, pi0127, pi0128, pi0129, pi0130, pi0131, pi0132, pi0133, pi0134,
    pi0135, pi0136, pi0137, pi0138, pi0139, pi0140, pi0141, pi0142, pi0143,
    pi0144, pi0145, pi0146, pi0147, pi0148, pi0149, pi0150, pi0151, pi0152,
    pi0153, pi0154, pi0155, pi0156, pi0157, pi0158, pi0159, pi0160, pi0161,
    pi0162, pi0163, pi0164, pi0165, pi0166, pi0167, pi0168, pi0169, pi0170,
    pi0171, pi0172, pi0173, pi0174, pi0175, pi0176, pi0177, pi0178, pi0179,
    pi0180, pi0181, pi0182, pi0183, pi0184, pi0185, pi0186, pi0187, pi0188,
    pi0189, pi0190, pi0191, pi0192, pi0193, pi0194, pi0195, pi0196, pi0197,
    pi0198, pi0199, pi0200, pi0201, pi0202, pi0203, pi0204, pi0205, pi0206,
    pi0207, pi0208, pi0209, pi0210, pi0211, pi0212, pi0213, pi0214, pi0215,
    pi0216, pi0217, pi0218, pi0219, pi0220, pi0221, pi0222, pi0223, pi0224,
    pi0225, pi0226, pi0227, pi0228, pi0229, pi0230, pi0231, pi0232, pi0233,
    pi0234, pi0235, pi0236, pi0237, pi0238, pi0239, pi0240, pi0241, pi0242,
    pi0243, pi0244, pi0245, pi0246, pi0247, pi0248, pi0249, pi0250, pi0251,
    pi0252, pi0253, pi0254, pi0255, pi0256, pi0257, pi0258, pi0259, pi0260,
    pi0261, pi0262, pi0263, pi0264, pi0265, pi0266, pi0267, pi0268, pi0269,
    pi0270, pi0271, pi0272, pi0273, pi0274, pi0275, pi0276, pi0277, pi0278,
    pi0279, pi0280, pi0281, pi0282, pi0283, pi0284, pi0285, pi0286, pi0287,
    pi0288, pi0289, pi0290, pi0291, pi0292, pi0293, pi0294, pi0295, pi0296,
    pi0297, pi0298, pi0299, pi0300, pi0301, pi0302, pi0303, pi0304, pi0305,
    pi0306, pi0307, pi0308, pi0309, pi0310, pi0311, pi0312, pi0313, pi0314,
    pi0315, pi0316, pi0317, pi0318, pi0319, pi0320, pi0321, pi0322, pi0323,
    pi0324, pi0325, pi0326, pi0327, pi0328, pi0329, pi0330, pi0331, pi0332,
    pi0333, pi0334, pi0335, pi0336, pi0337, pi0338, pi0339, pi0340, pi0341,
    pi0342, pi0343, pi0344, pi0345, pi0346, pi0347, pi0348, pi0349, pi0350,
    pi0351, pi0352, pi0353, pi0354, pi0355, pi0356, pi0357, pi0358, pi0359,
    pi0360, pi0361, pi0362, pi0363, pi0364, pi0365, pi0366, pi0367, pi0368,
    pi0369, pi0370, pi0371, pi0372, pi0373, pi0374, pi0375, pi0376, pi0377,
    pi0378, pi0379, pi0380, pi0381, pi0382, pi0383, pi0384, pi0385, pi0386,
    pi0387, pi0388, pi0389, pi0390, pi0391, pi0392, pi0393, pi0394, pi0395,
    pi0396, pi0397, pi0398, pi0399, pi0400, pi0401, pi0402, pi0403, pi0404,
    pi0405, pi0406, pi0407, pi0408, pi0409, pi0410, pi0411, pi0412, pi0413,
    pi0414, pi0415, pi0416, pi0417, pi0418, pi0419, pi0420, pi0421, pi0422,
    pi0423, pi0424, pi0425, pi0426, pi0427, pi0428, pi0429, pi0430, pi0431,
    pi0432, pi0433, pi0434, pi0435, pi0436, pi0437, pi0438, pi0439, pi0440,
    pi0441, pi0442, pi0443, pi0444, pi0445, pi0446, pi0447, pi0448, pi0449,
    pi0450, pi0451, pi0452, pi0453, pi0454, pi0455, pi0456, pi0457, pi0458,
    pi0459, pi0460, pi0461, pi0462, pi0463, pi0464, pi0465, pi0466, pi0467,
    pi0468, pi0469, pi0470, pi0471, pi0472, pi0473, pi0474, pi0475, pi0476,
    pi0477, pi0478, pi0479, pi0480, pi0481, pi0482, pi0483, pi0484, pi0485,
    pi0486, pi0487, pi0488, pi0489, pi0490, pi0491, pi0492, pi0493, pi0494,
    pi0495, pi0496, pi0497, pi0498, pi0499, pi0500, pi0501, pi0502, pi0503,
    pi0504, pi0505, pi0506, pi0507, pi0508, pi0509, pi0510, pi0511, pi0512,
    pi0513, pi0514, pi0515, pi0516, pi0517, pi0518, pi0519, pi0520, pi0521,
    pi0522, pi0523, pi0524, pi0525, pi0526, pi0527, pi0528, pi0529, pi0530,
    pi0531, pi0532, pi0533, pi0534, pi0535, pi0536, pi0537, pi0538, pi0539,
    pi0540, pi0541, pi0542, pi0543, pi0544, pi0545, pi0546, pi0547, pi0548,
    pi0549, pi0550, pi0551, pi0552, pi0553, pi0554, pi0555, pi0556, pi0557,
    pi0558, pi0559, pi0560, pi0561, pi0562, pi0563, pi0564, pi0565, pi0566,
    pi0567, pi0568, pi0569, pi0570, pi0571, pi0572, pi0573, pi0574, pi0575,
    pi0576, pi0577, pi0578, pi0579, pi0580, pi0581, pi0582, pi0583, pi0584,
    pi0585, pi0586, pi0587, pi0588, pi0589, pi0590, pi0591, pi0592, pi0593,
    pi0594, pi0595, pi0596, pi0597, pi0598, pi0599, pi0600, pi0601, pi0602,
    pi0603, pi0604, pi0605, pi0606, pi0607, pi0608, pi0609, pi0610, pi0611,
    pi0612, pi0613, pi0614, pi0615, pi0616, pi0617, pi0618, pi0619, pi0620,
    pi0621, pi0622, pi0623, pi0624, pi0625, pi0626, pi0627, pi0628, pi0629,
    pi0630, pi0631, pi0632, pi0633, pi0634, pi0635, pi0636, pi0637, pi0638,
    pi0639, pi0640, pi0641, pi0642, pi0643, pi0644, pi0645, pi0646, pi0647,
    pi0648, pi0649, pi0650, pi0651, pi0652, pi0653, pi0654, pi0655, pi0656,
    pi0657, pi0658, pi0659, pi0660, pi0661, pi0662, pi0663, pi0664, pi0665,
    pi0666, pi0667, pi0668, pi0669, pi0670, pi0671, pi0672, pi0673, pi0674,
    pi0675, pi0676, pi0677, pi0678, pi0679, pi0680, pi0681, pi0682, pi0683,
    pi0684, pi0685, pi0686, pi0687, pi0688, pi0689, pi0690, pi0691, pi0692,
    pi0693, pi0694, pi0695, pi0696, pi0697, pi0698, pi0699, pi0700, pi0701,
    pi0702, pi0703, pi0704, pi0705, pi0706, pi0707, pi0708, pi0709, pi0710,
    pi0711, pi0712, pi0713, pi0714, pi0715, pi0716, pi0717, pi0718, pi0719,
    pi0720, pi0721, pi0722, pi0723, pi0724, pi0725, pi0726, pi0727, pi0728,
    pi0729, pi0730, pi0731, pi0732, pi0733, pi0734, pi0735, pi0736, pi0737,
    pi0738, pi0739, pi0740, pi0741, pi0742, pi0743, pi0744, pi0745, pi0746,
    pi0747, pi0748, pi0749, pi0750, pi0751, pi0752, pi0753, pi0754, pi0755,
    pi0756, pi0757, pi0758, pi0759, pi0760, pi0761, pi0762, pi0763, pi0764,
    pi0765, pi0766, pi0767, pi0768, pi0769, pi0770, pi0771, pi0772, pi0773,
    pi0774, pi0775, pi0776, pi0777, pi0778, pi0779, pi0780, pi0781, pi0782,
    pi0783, pi0784, pi0785, pi0786, pi0787, pi0788, pi0789, pi0790, pi0791,
    pi0792, pi0793, pi0794, pi0795, pi0796, pi0797, pi0798, pi0799, pi0800,
    pi0801, pi0802, pi0803, pi0804, pi0805, pi0806, pi0807, pi0808, pi0809,
    pi0810, pi0811, pi0812, pi0813, pi0814, pi0815, pi0816, pi0817, pi0818,
    pi0819, pi0820, pi0821, pi0822, pi0823, pi0824, pi0825, pi0826, pi0827,
    pi0828, pi0829, pi0830, pi0831, pi0832, pi0833, pi0834, pi0835, pi0836,
    pi0837, pi0838, pi0839, pi0840, pi0841, pi0842, pi0843, pi0844, pi0845,
    pi0846, pi0847, pi0848, pi0849, pi0850, pi0851, pi0852, pi0853, pi0854,
    pi0855, pi0856, pi0857, pi0858, pi0859, pi0860, pi0861, pi0862, pi0863,
    pi0864, pi0865, pi0866, pi0867, pi0868, pi0869, pi0870, pi0871, pi0872,
    pi0873, pi0874, pi0875, pi0876, pi0877, pi0878, pi0879, pi0880, pi0881,
    pi0882, pi0883, pi0884, pi0885, pi0886, pi0887, pi0888, pi0889, pi0890,
    pi0891, pi0892, pi0893, pi0894, pi0895, pi0896, pi0897, pi0898, pi0899,
    pi0900, pi0901, pi0902, pi0903, pi0904, pi0905, pi0906, pi0907, pi0908,
    pi0909, pi0910, pi0911, pi0912, pi0913, pi0914, pi0915, pi0916, pi0917,
    pi0918, pi0919, pi0920, pi0921, pi0922, pi0923, pi0924, pi0925, pi0926,
    pi0927, pi0928, pi0929, pi0930, pi0931, pi0932, pi0933, pi0934, pi0935,
    pi0936, pi0937, pi0938, pi0939, pi0940, pi0941, pi0942, pi0943, pi0944,
    pi0945, pi0946, pi0947, pi0948, pi0949, pi0950, pi0951, pi0952, pi0953,
    pi0954, pi0955, pi0956, pi0957, pi0958, pi0959, pi0960, pi0961, pi0962,
    pi0963, pi0964, pi0965, pi0966, pi0967, pi0968, pi0969, pi0970, pi0971,
    pi0972, pi0973, pi0974, pi0975, pi0976, pi0977, pi0978, pi0979, pi0980,
    pi0981, pi0982, pi0983, pi0984, pi0985, pi0986, pi0987, pi0988, pi0989,
    pi0990, pi0991, pi0992, pi0993, pi0994, pi0995, pi0996, pi0997, pi0998,
    pi0999, pi1000, pi1001, pi1002, pi1003, pi1004, pi1005, pi1006, pi1007,
    pi1008, pi1009, pi1010, pi1011, pi1012, pi1013, pi1014, pi1015, pi1016,
    pi1017, pi1018, pi1019, pi1020, pi1021, pi1022, pi1023, pi1024, pi1025,
    pi1026, pi1027, pi1028, pi1029, pi1030, pi1031, pi1032, pi1033, pi1034,
    pi1035, pi1036, pi1037, pi1038, pi1039, pi1040, pi1041, pi1042, pi1043,
    pi1044, pi1045, pi1046, pi1047, pi1048, pi1049, pi1050, pi1051, pi1052,
    pi1053, pi1054, pi1055, pi1056, pi1057, pi1058, pi1059, pi1060, pi1061,
    pi1062, pi1063, pi1064, pi1065, pi1066, pi1067, pi1068, pi1069, pi1070,
    pi1071, pi1072, pi1073, pi1074, pi1075, pi1076, pi1077, pi1078, pi1079,
    pi1080, pi1081, pi1082, pi1083, pi1084, pi1085, pi1086, pi1087, pi1088,
    pi1089, pi1090, pi1091, pi1092, pi1093, pi1094, pi1095, pi1096, pi1097,
    pi1098, pi1099, pi1100, pi1101, pi1102, pi1103, pi1104, pi1105, pi1106,
    pi1107, pi1108, pi1109, pi1110, pi1111, pi1112, pi1113, pi1114, pi1115,
    pi1116, pi1117, pi1118, pi1119, pi1120, pi1121, pi1122, pi1123, pi1124,
    pi1125, pi1126, pi1127, pi1128, pi1129, pi1130, pi1131, pi1132, pi1133,
    pi1134, pi1135, pi1136, pi1137, pi1138, pi1139, pi1140, pi1141, pi1142,
    pi1143, pi1144, pi1145, pi1146, pi1147, pi1148, pi1149, pi1150, pi1151,
    pi1152, pi1153, pi1154, pi1155, pi1156, pi1157, pi1158, pi1159, pi1160,
    pi1161, pi1162, pi1163, pi1164, pi1165, pi1166, pi1167, pi1168, pi1169,
    pi1170, pi1171, pi1172, pi1173, pi1174, pi1175, pi1176, pi1177, pi1178,
    pi1179, pi1180, pi1181, pi1182, pi1183, pi1184, pi1185, pi1186, pi1187,
    pi1188, pi1189, pi1190, pi1191, pi1192, pi1193, pi1194, pi1195, pi1196,
    pi1197, pi1198, pi1199, pi1200, pi1201, pi1202, pi1203,
    po0000, po0001, po0002, po0003, po0004, po0005, po0006, po0007, po0008,
    po0009, po0010, po0011, po0012, po0013, po0014, po0015, po0016, po0017,
    po0018, po0019, po0020, po0021, po0022, po0023, po0024, po0025, po0026,
    po0027, po0028, po0029, po0030, po0031, po0032, po0033, po0034, po0035,
    po0036, po0037, po0038, po0039, po0040, po0041, po0042, po0043, po0044,
    po0045, po0046, po0047, po0048, po0049, po0050, po0051, po0052, po0053,
    po0054, po0055, po0056, po0057, po0058, po0059, po0060, po0061, po0062,
    po0063, po0064, po0065, po0066, po0067, po0068, po0069, po0070, po0071,
    po0072, po0073, po0074, po0075, po0076, po0077, po0078, po0079, po0080,
    po0081, po0082, po0083, po0084, po0085, po0086, po0087, po0088, po0089,
    po0090, po0091, po0092, po0093, po0094, po0095, po0096, po0097, po0098,
    po0099, po0100, po0101, po0102, po0103, po0104, po0105, po0106, po0107,
    po0108, po0109, po0110, po0111, po0112, po0113, po0114, po0115, po0116,
    po0117, po0118, po0119, po0120, po0121, po0122, po0123, po0124, po0125,
    po0126, po0127, po0128, po0129, po0130, po0131, po0132, po0133, po0134,
    po0135, po0136, po0137, po0138, po0139, po0140, po0141, po0142, po0143,
    po0144, po0145, po0146, po0147, po0148, po0149, po0150, po0151, po0152,
    po0153, po0154, po0155, po0156, po0157, po0158, po0159, po0160, po0161,
    po0162, po0163, po0164, po0165, po0166, po0167, po0168, po0169, po0170,
    po0171, po0172, po0173, po0174, po0175, po0176, po0177, po0178, po0179,
    po0180, po0181, po0182, po0183, po0184, po0185, po0186, po0187, po0188,
    po0189, po0190, po0191, po0192, po0193, po0194, po0195, po0196, po0197,
    po0198, po0199, po0200, po0201, po0202, po0203, po0204, po0205, po0206,
    po0207, po0208, po0209, po0210, po0211, po0212, po0213, po0214, po0215,
    po0216, po0217, po0218, po0219, po0220, po0221, po0222, po0223, po0224,
    po0225, po0226, po0227, po0228, po0229, po0230, po0231, po0232, po0233,
    po0234, po0235, po0236, po0237, po0238, po0239, po0240, po0241, po0242,
    po0243, po0244, po0245, po0246, po0247, po0248, po0249, po0250, po0251,
    po0252, po0253, po0254, po0255, po0256, po0257, po0258, po0259, po0260,
    po0261, po0262, po0263, po0264, po0265, po0266, po0267, po0268, po0269,
    po0270, po0271, po0272, po0273, po0274, po0275, po0276, po0277, po0278,
    po0279, po0280, po0281, po0282, po0283, po0284, po0285, po0286, po0287,
    po0288, po0289, po0290, po0291, po0292, po0293, po0294, po0295, po0296,
    po0297, po0298, po0299, po0300, po0301, po0302, po0303, po0304, po0305,
    po0306, po0307, po0308, po0309, po0310, po0311, po0312, po0313, po0314,
    po0315, po0316, po0317, po0318, po0319, po0320, po0321, po0322, po0323,
    po0324, po0325, po0326, po0327, po0328, po0329, po0330, po0331, po0332,
    po0333, po0334, po0335, po0336, po0337, po0338, po0339, po0340, po0341,
    po0342, po0343, po0344, po0345, po0346, po0347, po0348, po0349, po0350,
    po0351, po0352, po0353, po0354, po0355, po0356, po0357, po0358, po0359,
    po0360, po0361, po0362, po0363, po0364, po0365, po0366, po0367, po0368,
    po0369, po0370, po0371, po0372, po0373, po0374, po0375, po0376, po0377,
    po0378, po0379, po0380, po0381, po0382, po0383, po0384, po0385, po0386,
    po0387, po0388, po0389, po0390, po0391, po0392, po0393, po0394, po0395,
    po0396, po0397, po0398, po0399, po0400, po0401, po0402, po0403, po0404,
    po0405, po0406, po0407, po0408, po0409, po0410, po0411, po0412, po0413,
    po0414, po0415, po0416, po0417, po0418, po0419, po0420, po0421, po0422,
    po0423, po0424, po0425, po0426, po0427, po0428, po0429, po0430, po0431,
    po0432, po0433, po0434, po0435, po0436, po0437, po0438, po0439, po0440,
    po0441, po0442, po0443, po0444, po0445, po0446, po0447, po0448, po0449,
    po0450, po0451, po0452, po0453, po0454, po0455, po0456, po0457, po0458,
    po0459, po0460, po0461, po0462, po0463, po0464, po0465, po0466, po0467,
    po0468, po0469, po0470, po0471, po0472, po0473, po0474, po0475, po0476,
    po0477, po0478, po0479, po0480, po0481, po0482, po0483, po0484, po0485,
    po0486, po0487, po0488, po0489, po0490, po0491, po0492, po0493, po0494,
    po0495, po0496, po0497, po0498, po0499, po0500, po0501, po0502, po0503,
    po0504, po0505, po0506, po0507, po0508, po0509, po0510, po0511, po0512,
    po0513, po0514, po0515, po0516, po0517, po0518, po0519, po0520, po0521,
    po0522, po0523, po0524, po0525, po0526, po0527, po0528, po0529, po0530,
    po0531, po0532, po0533, po0534, po0535, po0536, po0537, po0538, po0539,
    po0540, po0541, po0542, po0543, po0544, po0545, po0546, po0547, po0548,
    po0549, po0550, po0551, po0552, po0553, po0554, po0555, po0556, po0557,
    po0558, po0559, po0560, po0561, po0562, po0563, po0564, po0565, po0566,
    po0567, po0568, po0569, po0570, po0571, po0572, po0573, po0574, po0575,
    po0576, po0577, po0578, po0579, po0580, po0581, po0582, po0583, po0584,
    po0585, po0586, po0587, po0588, po0589, po0590, po0591, po0592, po0593,
    po0594, po0595, po0596, po0597, po0598, po0599, po0600, po0601, po0602,
    po0603, po0604, po0605, po0606, po0607, po0608, po0609, po0610, po0611,
    po0612, po0613, po0614, po0615, po0616, po0617, po0618, po0619, po0620,
    po0621, po0622, po0623, po0624, po0625, po0626, po0627, po0628, po0629,
    po0630, po0631, po0632, po0633, po0634, po0635, po0636, po0637, po0638,
    po0639, po0640, po0641, po0642, po0643, po0644, po0645, po0646, po0647,
    po0648, po0649, po0650, po0651, po0652, po0653, po0654, po0655, po0656,
    po0657, po0658, po0659, po0660, po0661, po0662, po0663, po0664, po0665,
    po0666, po0667, po0668, po0669, po0670, po0671, po0672, po0673, po0674,
    po0675, po0676, po0677, po0678, po0679, po0680, po0681, po0682, po0683,
    po0684, po0685, po0686, po0687, po0688, po0689, po0690, po0691, po0692,
    po0693, po0694, po0695, po0696, po0697, po0698, po0699, po0700, po0701,
    po0702, po0703, po0704, po0705, po0706, po0707, po0708, po0709, po0710,
    po0711, po0712, po0713, po0714, po0715, po0716, po0717, po0718, po0719,
    po0720, po0721, po0722, po0723, po0724, po0725, po0726, po0727, po0728,
    po0729, po0730, po0731, po0732, po0733, po0734, po0735, po0736, po0737,
    po0738, po0739, po0740, po0741, po0742, po0743, po0744, po0745, po0746,
    po0747, po0748, po0749, po0750, po0751, po0752, po0753, po0754, po0755,
    po0756, po0757, po0758, po0759, po0760, po0761, po0762, po0763, po0764,
    po0765, po0766, po0767, po0768, po0769, po0770, po0771, po0772, po0773,
    po0774, po0775, po0776, po0777, po0778, po0779, po0780, po0781, po0782,
    po0783, po0784, po0785, po0786, po0787, po0788, po0789, po0790, po0791,
    po0792, po0793, po0794, po0795, po0796, po0797, po0798, po0799, po0800,
    po0801, po0802, po0803, po0804, po0805, po0806, po0807, po0808, po0809,
    po0810, po0811, po0812, po0813, po0814, po0815, po0816, po0817, po0818,
    po0819, po0820, po0821, po0822, po0823, po0824, po0825, po0826, po0827,
    po0828, po0829, po0830, po0831, po0832, po0833, po0834, po0835, po0836,
    po0837, po0838, po0839, po0840, po0841, po0842, po0843, po0844, po0845,
    po0846, po0847, po0848, po0849, po0850, po0851, po0852, po0853, po0854,
    po0855, po0856, po0857, po0858, po0859, po0860, po0861, po0862, po0863,
    po0864, po0865, po0866, po0867, po0868, po0869, po0870, po0871, po0872,
    po0873, po0874, po0875, po0876, po0877, po0878, po0879, po0880, po0881,
    po0882, po0883, po0884, po0885, po0886, po0887, po0888, po0889, po0890,
    po0891, po0892, po0893, po0894, po0895, po0896, po0897, po0898, po0899,
    po0900, po0901, po0902, po0903, po0904, po0905, po0906, po0907, po0908,
    po0909, po0910, po0911, po0912, po0913, po0914, po0915, po0916, po0917,
    po0918, po0919, po0920, po0921, po0922, po0923, po0924, po0925, po0926,
    po0927, po0928, po0929, po0930, po0931, po0932, po0933, po0934, po0935,
    po0936, po0937, po0938, po0939, po0940, po0941, po0942, po0943, po0944,
    po0945, po0946, po0947, po0948, po0949, po0950, po0951, po0952, po0953,
    po0954, po0955, po0956, po0957, po0958, po0959, po0960, po0961, po0962,
    po0963, po0964, po0965, po0966, po0967, po0968, po0969, po0970, po0971,
    po0972, po0973, po0974, po0975, po0976, po0977, po0978, po0979, po0980,
    po0981, po0982, po0983, po0984, po0985, po0986, po0987, po0988, po0989,
    po0990, po0991, po0992, po0993, po0994, po0995, po0996, po0997, po0998,
    po0999, po1000, po1001, po1002, po1003, po1004, po1005, po1006, po1007,
    po1008, po1009, po1010, po1011, po1012, po1013, po1014, po1015, po1016,
    po1017, po1018, po1019, po1020, po1021, po1022, po1023, po1024, po1025,
    po1026, po1027, po1028, po1029, po1030, po1031, po1032, po1033, po1034,
    po1035, po1036, po1037, po1038, po1039, po1040, po1041, po1042, po1043,
    po1044, po1045, po1046, po1047, po1048, po1049, po1050, po1051, po1052,
    po1053, po1054, po1055, po1056, po1057, po1058, po1059, po1060, po1061,
    po1062, po1063, po1064, po1065, po1066, po1067, po1068, po1069, po1070,
    po1071, po1072, po1073, po1074, po1075, po1076, po1077, po1078, po1079,
    po1080, po1081, po1082, po1083, po1084, po1085, po1086, po1087, po1088,
    po1089, po1090, po1091, po1092, po1093, po1094, po1095, po1096, po1097,
    po1098, po1099, po1100, po1101, po1102, po1103, po1104, po1105, po1106,
    po1107, po1108, po1109, po1110, po1111, po1112, po1113, po1114, po1115,
    po1116, po1117, po1118, po1119, po1120, po1121, po1122, po1123, po1124,
    po1125, po1126, po1127, po1128, po1129, po1130, po1131, po1132, po1133,
    po1134, po1135, po1136, po1137, po1138, po1139, po1140, po1141, po1142,
    po1143, po1144, po1145, po1146, po1147, po1148, po1149, po1150, po1151,
    po1152, po1153, po1154, po1155, po1156, po1157, po1158, po1159, po1160,
    po1161, po1162, po1163, po1164, po1165, po1166, po1167, po1168, po1169,
    po1170, po1171, po1172, po1173, po1174, po1175, po1176, po1177, po1178,
    po1179, po1180, po1181, po1182, po1183, po1184, po1185, po1186, po1187,
    po1188, po1189, po1190, po1191, po1192, po1193, po1194, po1195, po1196,
    po1197, po1198, po1199, po1200, po1201, po1202, po1203, po1204, po1205,
    po1206, po1207, po1208, po1209, po1210, po1211, po1212, po1213, po1214,
    po1215, po1216, po1217, po1218, po1219, po1220, po1221, po1222, po1223,
    po1224, po1225, po1226, po1227, po1228, po1229, po1230  );
  input  pi0000, pi0001, pi0002, pi0003, pi0004, pi0005, pi0006, pi0007,
    pi0008, pi0009, pi0010, pi0011, pi0012, pi0013, pi0014, pi0015, pi0016,
    pi0017, pi0018, pi0019, pi0020, pi0021, pi0022, pi0023, pi0024, pi0025,
    pi0026, pi0027, pi0028, pi0029, pi0030, pi0031, pi0032, pi0033, pi0034,
    pi0035, pi0036, pi0037, pi0038, pi0039, pi0040, pi0041, pi0042, pi0043,
    pi0044, pi0045, pi0046, pi0047, pi0048, pi0049, pi0050, pi0051, pi0052,
    pi0053, pi0054, pi0055, pi0056, pi0057, pi0058, pi0059, pi0060, pi0061,
    pi0062, pi0063, pi0064, pi0065, pi0066, pi0067, pi0068, pi0069, pi0070,
    pi0071, pi0072, pi0073, pi0074, pi0075, pi0076, pi0077, pi0078, pi0079,
    pi0080, pi0081, pi0082, pi0083, pi0084, pi0085, pi0086, pi0087, pi0088,
    pi0089, pi0090, pi0091, pi0092, pi0093, pi0094, pi0095, pi0096, pi0097,
    pi0098, pi0099, pi0100, pi0101, pi0102, pi0103, pi0104, pi0105, pi0106,
    pi0107, pi0108, pi0109, pi0110, pi0111, pi0112, pi0113, pi0114, pi0115,
    pi0116, pi0117, pi0118, pi0119, pi0120, pi0121, pi0122, pi0123, pi0124,
    pi0125, pi0126, pi0127, pi0128, pi0129, pi0130, pi0131, pi0132, pi0133,
    pi0134, pi0135, pi0136, pi0137, pi0138, pi0139, pi0140, pi0141, pi0142,
    pi0143, pi0144, pi0145, pi0146, pi0147, pi0148, pi0149, pi0150, pi0151,
    pi0152, pi0153, pi0154, pi0155, pi0156, pi0157, pi0158, pi0159, pi0160,
    pi0161, pi0162, pi0163, pi0164, pi0165, pi0166, pi0167, pi0168, pi0169,
    pi0170, pi0171, pi0172, pi0173, pi0174, pi0175, pi0176, pi0177, pi0178,
    pi0179, pi0180, pi0181, pi0182, pi0183, pi0184, pi0185, pi0186, pi0187,
    pi0188, pi0189, pi0190, pi0191, pi0192, pi0193, pi0194, pi0195, pi0196,
    pi0197, pi0198, pi0199, pi0200, pi0201, pi0202, pi0203, pi0204, pi0205,
    pi0206, pi0207, pi0208, pi0209, pi0210, pi0211, pi0212, pi0213, pi0214,
    pi0215, pi0216, pi0217, pi0218, pi0219, pi0220, pi0221, pi0222, pi0223,
    pi0224, pi0225, pi0226, pi0227, pi0228, pi0229, pi0230, pi0231, pi0232,
    pi0233, pi0234, pi0235, pi0236, pi0237, pi0238, pi0239, pi0240, pi0241,
    pi0242, pi0243, pi0244, pi0245, pi0246, pi0247, pi0248, pi0249, pi0250,
    pi0251, pi0252, pi0253, pi0254, pi0255, pi0256, pi0257, pi0258, pi0259,
    pi0260, pi0261, pi0262, pi0263, pi0264, pi0265, pi0266, pi0267, pi0268,
    pi0269, pi0270, pi0271, pi0272, pi0273, pi0274, pi0275, pi0276, pi0277,
    pi0278, pi0279, pi0280, pi0281, pi0282, pi0283, pi0284, pi0285, pi0286,
    pi0287, pi0288, pi0289, pi0290, pi0291, pi0292, pi0293, pi0294, pi0295,
    pi0296, pi0297, pi0298, pi0299, pi0300, pi0301, pi0302, pi0303, pi0304,
    pi0305, pi0306, pi0307, pi0308, pi0309, pi0310, pi0311, pi0312, pi0313,
    pi0314, pi0315, pi0316, pi0317, pi0318, pi0319, pi0320, pi0321, pi0322,
    pi0323, pi0324, pi0325, pi0326, pi0327, pi0328, pi0329, pi0330, pi0331,
    pi0332, pi0333, pi0334, pi0335, pi0336, pi0337, pi0338, pi0339, pi0340,
    pi0341, pi0342, pi0343, pi0344, pi0345, pi0346, pi0347, pi0348, pi0349,
    pi0350, pi0351, pi0352, pi0353, pi0354, pi0355, pi0356, pi0357, pi0358,
    pi0359, pi0360, pi0361, pi0362, pi0363, pi0364, pi0365, pi0366, pi0367,
    pi0368, pi0369, pi0370, pi0371, pi0372, pi0373, pi0374, pi0375, pi0376,
    pi0377, pi0378, pi0379, pi0380, pi0381, pi0382, pi0383, pi0384, pi0385,
    pi0386, pi0387, pi0388, pi0389, pi0390, pi0391, pi0392, pi0393, pi0394,
    pi0395, pi0396, pi0397, pi0398, pi0399, pi0400, pi0401, pi0402, pi0403,
    pi0404, pi0405, pi0406, pi0407, pi0408, pi0409, pi0410, pi0411, pi0412,
    pi0413, pi0414, pi0415, pi0416, pi0417, pi0418, pi0419, pi0420, pi0421,
    pi0422, pi0423, pi0424, pi0425, pi0426, pi0427, pi0428, pi0429, pi0430,
    pi0431, pi0432, pi0433, pi0434, pi0435, pi0436, pi0437, pi0438, pi0439,
    pi0440, pi0441, pi0442, pi0443, pi0444, pi0445, pi0446, pi0447, pi0448,
    pi0449, pi0450, pi0451, pi0452, pi0453, pi0454, pi0455, pi0456, pi0457,
    pi0458, pi0459, pi0460, pi0461, pi0462, pi0463, pi0464, pi0465, pi0466,
    pi0467, pi0468, pi0469, pi0470, pi0471, pi0472, pi0473, pi0474, pi0475,
    pi0476, pi0477, pi0478, pi0479, pi0480, pi0481, pi0482, pi0483, pi0484,
    pi0485, pi0486, pi0487, pi0488, pi0489, pi0490, pi0491, pi0492, pi0493,
    pi0494, pi0495, pi0496, pi0497, pi0498, pi0499, pi0500, pi0501, pi0502,
    pi0503, pi0504, pi0505, pi0506, pi0507, pi0508, pi0509, pi0510, pi0511,
    pi0512, pi0513, pi0514, pi0515, pi0516, pi0517, pi0518, pi0519, pi0520,
    pi0521, pi0522, pi0523, pi0524, pi0525, pi0526, pi0527, pi0528, pi0529,
    pi0530, pi0531, pi0532, pi0533, pi0534, pi0535, pi0536, pi0537, pi0538,
    pi0539, pi0540, pi0541, pi0542, pi0543, pi0544, pi0545, pi0546, pi0547,
    pi0548, pi0549, pi0550, pi0551, pi0552, pi0553, pi0554, pi0555, pi0556,
    pi0557, pi0558, pi0559, pi0560, pi0561, pi0562, pi0563, pi0564, pi0565,
    pi0566, pi0567, pi0568, pi0569, pi0570, pi0571, pi0572, pi0573, pi0574,
    pi0575, pi0576, pi0577, pi0578, pi0579, pi0580, pi0581, pi0582, pi0583,
    pi0584, pi0585, pi0586, pi0587, pi0588, pi0589, pi0590, pi0591, pi0592,
    pi0593, pi0594, pi0595, pi0596, pi0597, pi0598, pi0599, pi0600, pi0601,
    pi0602, pi0603, pi0604, pi0605, pi0606, pi0607, pi0608, pi0609, pi0610,
    pi0611, pi0612, pi0613, pi0614, pi0615, pi0616, pi0617, pi0618, pi0619,
    pi0620, pi0621, pi0622, pi0623, pi0624, pi0625, pi0626, pi0627, pi0628,
    pi0629, pi0630, pi0631, pi0632, pi0633, pi0634, pi0635, pi0636, pi0637,
    pi0638, pi0639, pi0640, pi0641, pi0642, pi0643, pi0644, pi0645, pi0646,
    pi0647, pi0648, pi0649, pi0650, pi0651, pi0652, pi0653, pi0654, pi0655,
    pi0656, pi0657, pi0658, pi0659, pi0660, pi0661, pi0662, pi0663, pi0664,
    pi0665, pi0666, pi0667, pi0668, pi0669, pi0670, pi0671, pi0672, pi0673,
    pi0674, pi0675, pi0676, pi0677, pi0678, pi0679, pi0680, pi0681, pi0682,
    pi0683, pi0684, pi0685, pi0686, pi0687, pi0688, pi0689, pi0690, pi0691,
    pi0692, pi0693, pi0694, pi0695, pi0696, pi0697, pi0698, pi0699, pi0700,
    pi0701, pi0702, pi0703, pi0704, pi0705, pi0706, pi0707, pi0708, pi0709,
    pi0710, pi0711, pi0712, pi0713, pi0714, pi0715, pi0716, pi0717, pi0718,
    pi0719, pi0720, pi0721, pi0722, pi0723, pi0724, pi0725, pi0726, pi0727,
    pi0728, pi0729, pi0730, pi0731, pi0732, pi0733, pi0734, pi0735, pi0736,
    pi0737, pi0738, pi0739, pi0740, pi0741, pi0742, pi0743, pi0744, pi0745,
    pi0746, pi0747, pi0748, pi0749, pi0750, pi0751, pi0752, pi0753, pi0754,
    pi0755, pi0756, pi0757, pi0758, pi0759, pi0760, pi0761, pi0762, pi0763,
    pi0764, pi0765, pi0766, pi0767, pi0768, pi0769, pi0770, pi0771, pi0772,
    pi0773, pi0774, pi0775, pi0776, pi0777, pi0778, pi0779, pi0780, pi0781,
    pi0782, pi0783, pi0784, pi0785, pi0786, pi0787, pi0788, pi0789, pi0790,
    pi0791, pi0792, pi0793, pi0794, pi0795, pi0796, pi0797, pi0798, pi0799,
    pi0800, pi0801, pi0802, pi0803, pi0804, pi0805, pi0806, pi0807, pi0808,
    pi0809, pi0810, pi0811, pi0812, pi0813, pi0814, pi0815, pi0816, pi0817,
    pi0818, pi0819, pi0820, pi0821, pi0822, pi0823, pi0824, pi0825, pi0826,
    pi0827, pi0828, pi0829, pi0830, pi0831, pi0832, pi0833, pi0834, pi0835,
    pi0836, pi0837, pi0838, pi0839, pi0840, pi0841, pi0842, pi0843, pi0844,
    pi0845, pi0846, pi0847, pi0848, pi0849, pi0850, pi0851, pi0852, pi0853,
    pi0854, pi0855, pi0856, pi0857, pi0858, pi0859, pi0860, pi0861, pi0862,
    pi0863, pi0864, pi0865, pi0866, pi0867, pi0868, pi0869, pi0870, pi0871,
    pi0872, pi0873, pi0874, pi0875, pi0876, pi0877, pi0878, pi0879, pi0880,
    pi0881, pi0882, pi0883, pi0884, pi0885, pi0886, pi0887, pi0888, pi0889,
    pi0890, pi0891, pi0892, pi0893, pi0894, pi0895, pi0896, pi0897, pi0898,
    pi0899, pi0900, pi0901, pi0902, pi0903, pi0904, pi0905, pi0906, pi0907,
    pi0908, pi0909, pi0910, pi0911, pi0912, pi0913, pi0914, pi0915, pi0916,
    pi0917, pi0918, pi0919, pi0920, pi0921, pi0922, pi0923, pi0924, pi0925,
    pi0926, pi0927, pi0928, pi0929, pi0930, pi0931, pi0932, pi0933, pi0934,
    pi0935, pi0936, pi0937, pi0938, pi0939, pi0940, pi0941, pi0942, pi0943,
    pi0944, pi0945, pi0946, pi0947, pi0948, pi0949, pi0950, pi0951, pi0952,
    pi0953, pi0954, pi0955, pi0956, pi0957, pi0958, pi0959, pi0960, pi0961,
    pi0962, pi0963, pi0964, pi0965, pi0966, pi0967, pi0968, pi0969, pi0970,
    pi0971, pi0972, pi0973, pi0974, pi0975, pi0976, pi0977, pi0978, pi0979,
    pi0980, pi0981, pi0982, pi0983, pi0984, pi0985, pi0986, pi0987, pi0988,
    pi0989, pi0990, pi0991, pi0992, pi0993, pi0994, pi0995, pi0996, pi0997,
    pi0998, pi0999, pi1000, pi1001, pi1002, pi1003, pi1004, pi1005, pi1006,
    pi1007, pi1008, pi1009, pi1010, pi1011, pi1012, pi1013, pi1014, pi1015,
    pi1016, pi1017, pi1018, pi1019, pi1020, pi1021, pi1022, pi1023, pi1024,
    pi1025, pi1026, pi1027, pi1028, pi1029, pi1030, pi1031, pi1032, pi1033,
    pi1034, pi1035, pi1036, pi1037, pi1038, pi1039, pi1040, pi1041, pi1042,
    pi1043, pi1044, pi1045, pi1046, pi1047, pi1048, pi1049, pi1050, pi1051,
    pi1052, pi1053, pi1054, pi1055, pi1056, pi1057, pi1058, pi1059, pi1060,
    pi1061, pi1062, pi1063, pi1064, pi1065, pi1066, pi1067, pi1068, pi1069,
    pi1070, pi1071, pi1072, pi1073, pi1074, pi1075, pi1076, pi1077, pi1078,
    pi1079, pi1080, pi1081, pi1082, pi1083, pi1084, pi1085, pi1086, pi1087,
    pi1088, pi1089, pi1090, pi1091, pi1092, pi1093, pi1094, pi1095, pi1096,
    pi1097, pi1098, pi1099, pi1100, pi1101, pi1102, pi1103, pi1104, pi1105,
    pi1106, pi1107, pi1108, pi1109, pi1110, pi1111, pi1112, pi1113, pi1114,
    pi1115, pi1116, pi1117, pi1118, pi1119, pi1120, pi1121, pi1122, pi1123,
    pi1124, pi1125, pi1126, pi1127, pi1128, pi1129, pi1130, pi1131, pi1132,
    pi1133, pi1134, pi1135, pi1136, pi1137, pi1138, pi1139, pi1140, pi1141,
    pi1142, pi1143, pi1144, pi1145, pi1146, pi1147, pi1148, pi1149, pi1150,
    pi1151, pi1152, pi1153, pi1154, pi1155, pi1156, pi1157, pi1158, pi1159,
    pi1160, pi1161, pi1162, pi1163, pi1164, pi1165, pi1166, pi1167, pi1168,
    pi1169, pi1170, pi1171, pi1172, pi1173, pi1174, pi1175, pi1176, pi1177,
    pi1178, pi1179, pi1180, pi1181, pi1182, pi1183, pi1184, pi1185, pi1186,
    pi1187, pi1188, pi1189, pi1190, pi1191, pi1192, pi1193, pi1194, pi1195,
    pi1196, pi1197, pi1198, pi1199, pi1200, pi1201, pi1202, pi1203;
  output po0000, po0001, po0002, po0003, po0004, po0005, po0006, po0007,
    po0008, po0009, po0010, po0011, po0012, po0013, po0014, po0015, po0016,
    po0017, po0018, po0019, po0020, po0021, po0022, po0023, po0024, po0025,
    po0026, po0027, po0028, po0029, po0030, po0031, po0032, po0033, po0034,
    po0035, po0036, po0037, po0038, po0039, po0040, po0041, po0042, po0043,
    po0044, po0045, po0046, po0047, po0048, po0049, po0050, po0051, po0052,
    po0053, po0054, po0055, po0056, po0057, po0058, po0059, po0060, po0061,
    po0062, po0063, po0064, po0065, po0066, po0067, po0068, po0069, po0070,
    po0071, po0072, po0073, po0074, po0075, po0076, po0077, po0078, po0079,
    po0080, po0081, po0082, po0083, po0084, po0085, po0086, po0087, po0088,
    po0089, po0090, po0091, po0092, po0093, po0094, po0095, po0096, po0097,
    po0098, po0099, po0100, po0101, po0102, po0103, po0104, po0105, po0106,
    po0107, po0108, po0109, po0110, po0111, po0112, po0113, po0114, po0115,
    po0116, po0117, po0118, po0119, po0120, po0121, po0122, po0123, po0124,
    po0125, po0126, po0127, po0128, po0129, po0130, po0131, po0132, po0133,
    po0134, po0135, po0136, po0137, po0138, po0139, po0140, po0141, po0142,
    po0143, po0144, po0145, po0146, po0147, po0148, po0149, po0150, po0151,
    po0152, po0153, po0154, po0155, po0156, po0157, po0158, po0159, po0160,
    po0161, po0162, po0163, po0164, po0165, po0166, po0167, po0168, po0169,
    po0170, po0171, po0172, po0173, po0174, po0175, po0176, po0177, po0178,
    po0179, po0180, po0181, po0182, po0183, po0184, po0185, po0186, po0187,
    po0188, po0189, po0190, po0191, po0192, po0193, po0194, po0195, po0196,
    po0197, po0198, po0199, po0200, po0201, po0202, po0203, po0204, po0205,
    po0206, po0207, po0208, po0209, po0210, po0211, po0212, po0213, po0214,
    po0215, po0216, po0217, po0218, po0219, po0220, po0221, po0222, po0223,
    po0224, po0225, po0226, po0227, po0228, po0229, po0230, po0231, po0232,
    po0233, po0234, po0235, po0236, po0237, po0238, po0239, po0240, po0241,
    po0242, po0243, po0244, po0245, po0246, po0247, po0248, po0249, po0250,
    po0251, po0252, po0253, po0254, po0255, po0256, po0257, po0258, po0259,
    po0260, po0261, po0262, po0263, po0264, po0265, po0266, po0267, po0268,
    po0269, po0270, po0271, po0272, po0273, po0274, po0275, po0276, po0277,
    po0278, po0279, po0280, po0281, po0282, po0283, po0284, po0285, po0286,
    po0287, po0288, po0289, po0290, po0291, po0292, po0293, po0294, po0295,
    po0296, po0297, po0298, po0299, po0300, po0301, po0302, po0303, po0304,
    po0305, po0306, po0307, po0308, po0309, po0310, po0311, po0312, po0313,
    po0314, po0315, po0316, po0317, po0318, po0319, po0320, po0321, po0322,
    po0323, po0324, po0325, po0326, po0327, po0328, po0329, po0330, po0331,
    po0332, po0333, po0334, po0335, po0336, po0337, po0338, po0339, po0340,
    po0341, po0342, po0343, po0344, po0345, po0346, po0347, po0348, po0349,
    po0350, po0351, po0352, po0353, po0354, po0355, po0356, po0357, po0358,
    po0359, po0360, po0361, po0362, po0363, po0364, po0365, po0366, po0367,
    po0368, po0369, po0370, po0371, po0372, po0373, po0374, po0375, po0376,
    po0377, po0378, po0379, po0380, po0381, po0382, po0383, po0384, po0385,
    po0386, po0387, po0388, po0389, po0390, po0391, po0392, po0393, po0394,
    po0395, po0396, po0397, po0398, po0399, po0400, po0401, po0402, po0403,
    po0404, po0405, po0406, po0407, po0408, po0409, po0410, po0411, po0412,
    po0413, po0414, po0415, po0416, po0417, po0418, po0419, po0420, po0421,
    po0422, po0423, po0424, po0425, po0426, po0427, po0428, po0429, po0430,
    po0431, po0432, po0433, po0434, po0435, po0436, po0437, po0438, po0439,
    po0440, po0441, po0442, po0443, po0444, po0445, po0446, po0447, po0448,
    po0449, po0450, po0451, po0452, po0453, po0454, po0455, po0456, po0457,
    po0458, po0459, po0460, po0461, po0462, po0463, po0464, po0465, po0466,
    po0467, po0468, po0469, po0470, po0471, po0472, po0473, po0474, po0475,
    po0476, po0477, po0478, po0479, po0480, po0481, po0482, po0483, po0484,
    po0485, po0486, po0487, po0488, po0489, po0490, po0491, po0492, po0493,
    po0494, po0495, po0496, po0497, po0498, po0499, po0500, po0501, po0502,
    po0503, po0504, po0505, po0506, po0507, po0508, po0509, po0510, po0511,
    po0512, po0513, po0514, po0515, po0516, po0517, po0518, po0519, po0520,
    po0521, po0522, po0523, po0524, po0525, po0526, po0527, po0528, po0529,
    po0530, po0531, po0532, po0533, po0534, po0535, po0536, po0537, po0538,
    po0539, po0540, po0541, po0542, po0543, po0544, po0545, po0546, po0547,
    po0548, po0549, po0550, po0551, po0552, po0553, po0554, po0555, po0556,
    po0557, po0558, po0559, po0560, po0561, po0562, po0563, po0564, po0565,
    po0566, po0567, po0568, po0569, po0570, po0571, po0572, po0573, po0574,
    po0575, po0576, po0577, po0578, po0579, po0580, po0581, po0582, po0583,
    po0584, po0585, po0586, po0587, po0588, po0589, po0590, po0591, po0592,
    po0593, po0594, po0595, po0596, po0597, po0598, po0599, po0600, po0601,
    po0602, po0603, po0604, po0605, po0606, po0607, po0608, po0609, po0610,
    po0611, po0612, po0613, po0614, po0615, po0616, po0617, po0618, po0619,
    po0620, po0621, po0622, po0623, po0624, po0625, po0626, po0627, po0628,
    po0629, po0630, po0631, po0632, po0633, po0634, po0635, po0636, po0637,
    po0638, po0639, po0640, po0641, po0642, po0643, po0644, po0645, po0646,
    po0647, po0648, po0649, po0650, po0651, po0652, po0653, po0654, po0655,
    po0656, po0657, po0658, po0659, po0660, po0661, po0662, po0663, po0664,
    po0665, po0666, po0667, po0668, po0669, po0670, po0671, po0672, po0673,
    po0674, po0675, po0676, po0677, po0678, po0679, po0680, po0681, po0682,
    po0683, po0684, po0685, po0686, po0687, po0688, po0689, po0690, po0691,
    po0692, po0693, po0694, po0695, po0696, po0697, po0698, po0699, po0700,
    po0701, po0702, po0703, po0704, po0705, po0706, po0707, po0708, po0709,
    po0710, po0711, po0712, po0713, po0714, po0715, po0716, po0717, po0718,
    po0719, po0720, po0721, po0722, po0723, po0724, po0725, po0726, po0727,
    po0728, po0729, po0730, po0731, po0732, po0733, po0734, po0735, po0736,
    po0737, po0738, po0739, po0740, po0741, po0742, po0743, po0744, po0745,
    po0746, po0747, po0748, po0749, po0750, po0751, po0752, po0753, po0754,
    po0755, po0756, po0757, po0758, po0759, po0760, po0761, po0762, po0763,
    po0764, po0765, po0766, po0767, po0768, po0769, po0770, po0771, po0772,
    po0773, po0774, po0775, po0776, po0777, po0778, po0779, po0780, po0781,
    po0782, po0783, po0784, po0785, po0786, po0787, po0788, po0789, po0790,
    po0791, po0792, po0793, po0794, po0795, po0796, po0797, po0798, po0799,
    po0800, po0801, po0802, po0803, po0804, po0805, po0806, po0807, po0808,
    po0809, po0810, po0811, po0812, po0813, po0814, po0815, po0816, po0817,
    po0818, po0819, po0820, po0821, po0822, po0823, po0824, po0825, po0826,
    po0827, po0828, po0829, po0830, po0831, po0832, po0833, po0834, po0835,
    po0836, po0837, po0838, po0839, po0840, po0841, po0842, po0843, po0844,
    po0845, po0846, po0847, po0848, po0849, po0850, po0851, po0852, po0853,
    po0854, po0855, po0856, po0857, po0858, po0859, po0860, po0861, po0862,
    po0863, po0864, po0865, po0866, po0867, po0868, po0869, po0870, po0871,
    po0872, po0873, po0874, po0875, po0876, po0877, po0878, po0879, po0880,
    po0881, po0882, po0883, po0884, po0885, po0886, po0887, po0888, po0889,
    po0890, po0891, po0892, po0893, po0894, po0895, po0896, po0897, po0898,
    po0899, po0900, po0901, po0902, po0903, po0904, po0905, po0906, po0907,
    po0908, po0909, po0910, po0911, po0912, po0913, po0914, po0915, po0916,
    po0917, po0918, po0919, po0920, po0921, po0922, po0923, po0924, po0925,
    po0926, po0927, po0928, po0929, po0930, po0931, po0932, po0933, po0934,
    po0935, po0936, po0937, po0938, po0939, po0940, po0941, po0942, po0943,
    po0944, po0945, po0946, po0947, po0948, po0949, po0950, po0951, po0952,
    po0953, po0954, po0955, po0956, po0957, po0958, po0959, po0960, po0961,
    po0962, po0963, po0964, po0965, po0966, po0967, po0968, po0969, po0970,
    po0971, po0972, po0973, po0974, po0975, po0976, po0977, po0978, po0979,
    po0980, po0981, po0982, po0983, po0984, po0985, po0986, po0987, po0988,
    po0989, po0990, po0991, po0992, po0993, po0994, po0995, po0996, po0997,
    po0998, po0999, po1000, po1001, po1002, po1003, po1004, po1005, po1006,
    po1007, po1008, po1009, po1010, po1011, po1012, po1013, po1014, po1015,
    po1016, po1017, po1018, po1019, po1020, po1021, po1022, po1023, po1024,
    po1025, po1026, po1027, po1028, po1029, po1030, po1031, po1032, po1033,
    po1034, po1035, po1036, po1037, po1038, po1039, po1040, po1041, po1042,
    po1043, po1044, po1045, po1046, po1047, po1048, po1049, po1050, po1051,
    po1052, po1053, po1054, po1055, po1056, po1057, po1058, po1059, po1060,
    po1061, po1062, po1063, po1064, po1065, po1066, po1067, po1068, po1069,
    po1070, po1071, po1072, po1073, po1074, po1075, po1076, po1077, po1078,
    po1079, po1080, po1081, po1082, po1083, po1084, po1085, po1086, po1087,
    po1088, po1089, po1090, po1091, po1092, po1093, po1094, po1095, po1096,
    po1097, po1098, po1099, po1100, po1101, po1102, po1103, po1104, po1105,
    po1106, po1107, po1108, po1109, po1110, po1111, po1112, po1113, po1114,
    po1115, po1116, po1117, po1118, po1119, po1120, po1121, po1122, po1123,
    po1124, po1125, po1126, po1127, po1128, po1129, po1130, po1131, po1132,
    po1133, po1134, po1135, po1136, po1137, po1138, po1139, po1140, po1141,
    po1142, po1143, po1144, po1145, po1146, po1147, po1148, po1149, po1150,
    po1151, po1152, po1153, po1154, po1155, po1156, po1157, po1158, po1159,
    po1160, po1161, po1162, po1163, po1164, po1165, po1166, po1167, po1168,
    po1169, po1170, po1171, po1172, po1173, po1174, po1175, po1176, po1177,
    po1178, po1179, po1180, po1181, po1182, po1183, po1184, po1185, po1186,
    po1187, po1188, po1189, po1190, po1191, po1192, po1193, po1194, po1195,
    po1196, po1197, po1198, po1199, po1200, po1201, po1202, po1203, po1204,
    po1205, po1206, po1207, po1208, po1209, po1210, po1211, po1212, po1213,
    po1214, po1215, po1216, po1217, po1218, po1219, po1220, po1221, po1222,
    po1223, po1224, po1225, po1226, po1227, po1228, po1229, po1230;
  wire new_n2436_, new_n2437_, new_n2438_, new_n2439_, new_n2440_,
    new_n2441_, new_n2442_, new_n2443_, new_n2444_, new_n2445_, new_n2446_,
    new_n2447_, new_n2448_, new_n2449_, new_n2450_, new_n2451_, new_n2452_,
    new_n2453_, new_n2454_, new_n2455_, new_n2456_, new_n2457_, new_n2458_,
    new_n2459_, new_n2460_, new_n2461_, new_n2462_, new_n2463_, new_n2464_,
    new_n2465_, new_n2466_, new_n2467_, new_n2468_, new_n2469_, new_n2470_,
    new_n2471_, new_n2472_, new_n2473_, new_n2474_, new_n2475_, new_n2476_,
    new_n2477_, new_n2478_, new_n2479_, new_n2480_, new_n2481_, new_n2482_,
    new_n2483_, new_n2484_, new_n2485_, new_n2486_, new_n2487_, new_n2488_,
    new_n2489_, new_n2490_, new_n2491_, new_n2492_, new_n2493_, new_n2494_,
    new_n2495_, new_n2496_, new_n2497_, new_n2498_, new_n2499_, new_n2500_,
    new_n2501_, new_n2502_, new_n2503_, new_n2504_, new_n2505_, new_n2506_,
    new_n2507_, new_n2508_, new_n2509_, new_n2510_, new_n2511_, new_n2512_,
    new_n2513_, new_n2514_, new_n2515_, new_n2516_, new_n2517_, new_n2518_,
    new_n2519_, new_n2520_, new_n2521_, new_n2522_, new_n2523_, new_n2524_,
    new_n2525_, new_n2526_, new_n2527_, new_n2528_, new_n2529_, new_n2530_,
    new_n2531_, new_n2532_, new_n2533_, new_n2534_, new_n2535_, new_n2536_,
    new_n2537_, new_n2538_, new_n2539_, new_n2540_, new_n2541_, new_n2542_,
    new_n2543_, new_n2544_, new_n2545_, new_n2546_, new_n2547_, new_n2548_,
    new_n2549_, new_n2550_, new_n2551_, new_n2552_, new_n2553_, new_n2554_,
    new_n2555_, new_n2556_, new_n2557_, new_n2558_, new_n2559_, new_n2560_,
    new_n2561_, new_n2562_, new_n2563_, new_n2564_, new_n2565_, new_n2566_,
    new_n2567_, new_n2568_, new_n2569_, new_n2570_, new_n2571_, new_n2572_,
    new_n2573_, new_n2574_, new_n2575_, new_n2576_, new_n2577_, new_n2578_,
    new_n2579_, new_n2580_, new_n2581_, new_n2582_, new_n2583_, new_n2584_,
    new_n2585_, new_n2586_, new_n2587_, new_n2588_, new_n2589_, new_n2590_,
    new_n2591_, new_n2592_, new_n2593_, new_n2594_, new_n2595_, new_n2596_,
    new_n2597_, new_n2598_, new_n2599_, new_n2600_, new_n2601_, new_n2602_,
    new_n2603_, new_n2604_, new_n2605_, new_n2606_, new_n2607_, new_n2608_,
    new_n2609_, new_n2610_, new_n2611_, new_n2612_, new_n2613_, new_n2614_,
    new_n2615_, new_n2616_, new_n2617_, new_n2618_, new_n2619_, new_n2620_,
    new_n2621_, new_n2622_, new_n2623_, new_n2624_, new_n2625_, new_n2626_,
    new_n2627_, new_n2628_, new_n2629_, new_n2630_, new_n2631_, new_n2632_,
    new_n2633_, new_n2634_, new_n2635_, new_n2636_, new_n2637_, new_n2638_,
    new_n2639_, new_n2640_, new_n2641_, new_n2642_, new_n2643_, new_n2644_,
    new_n2645_, new_n2646_, new_n2647_, new_n2648_, new_n2649_, new_n2650_,
    new_n2651_, new_n2652_, new_n2653_, new_n2654_, new_n2655_, new_n2656_,
    new_n2657_, new_n2658_, new_n2659_, new_n2660_, new_n2661_, new_n2662_,
    new_n2663_, new_n2664_, new_n2665_, new_n2666_, new_n2667_, new_n2668_,
    new_n2669_, new_n2670_, new_n2671_, new_n2672_, new_n2673_, new_n2674_,
    new_n2675_, new_n2676_, new_n2677_, new_n2678_, new_n2679_, new_n2680_,
    new_n2681_, new_n2682_, new_n2683_, new_n2684_, new_n2685_, new_n2686_,
    new_n2687_, new_n2688_, new_n2689_, new_n2690_, new_n2691_, new_n2692_,
    new_n2693_, new_n2694_, new_n2695_, new_n2696_, new_n2697_, new_n2698_,
    new_n2699_, new_n2700_, new_n2701_, new_n2702_, new_n2703_, new_n2704_,
    new_n2705_, new_n2706_, new_n2707_, new_n2708_, new_n2709_, new_n2710_,
    new_n2711_, new_n2712_, new_n2713_, new_n2714_, new_n2715_, new_n2716_,
    new_n2717_, new_n2718_, new_n2719_, new_n2720_, new_n2721_, new_n2722_,
    new_n2723_, new_n2724_, new_n2725_, new_n2726_, new_n2727_, new_n2728_,
    new_n2729_, new_n2730_, new_n2731_, new_n2732_, new_n2733_, new_n2734_,
    new_n2735_, new_n2736_, new_n2737_, new_n2738_, new_n2739_, new_n2740_,
    new_n2741_, new_n2742_, new_n2743_, new_n2744_, new_n2745_, new_n2746_,
    new_n2747_, new_n2748_, new_n2749_, new_n2750_, new_n2751_, new_n2752_,
    new_n2753_, new_n2754_, new_n2755_, new_n2756_, new_n2757_, new_n2758_,
    new_n2759_, new_n2760_, new_n2761_, new_n2762_, new_n2763_, new_n2764_,
    new_n2765_, new_n2766_, new_n2767_, new_n2768_, new_n2769_, new_n2770_,
    new_n2771_, new_n2772_, new_n2773_, new_n2774_, new_n2775_, new_n2776_,
    new_n2777_, new_n2778_, new_n2779_, new_n2780_, new_n2781_, new_n2782_,
    new_n2783_, new_n2784_, new_n2785_, new_n2786_, new_n2787_, new_n2788_,
    new_n2789_, new_n2790_, new_n2791_, new_n2792_, new_n2793_, new_n2794_,
    new_n2795_, new_n2796_, new_n2797_, new_n2798_, new_n2799_, new_n2800_,
    new_n2801_, new_n2802_, new_n2803_, new_n2804_, new_n2805_, new_n2806_,
    new_n2807_, new_n2808_, new_n2809_, new_n2810_, new_n2811_, new_n2812_,
    new_n2813_, new_n2814_, new_n2815_, new_n2816_, new_n2817_, new_n2818_,
    new_n2819_, new_n2820_, new_n2821_, new_n2822_, new_n2823_, new_n2824_,
    new_n2825_, new_n2826_, new_n2827_, new_n2828_, new_n2829_, new_n2830_,
    new_n2831_, new_n2832_, new_n2833_, new_n2834_, new_n2835_, new_n2836_,
    new_n2837_, new_n2838_, new_n2839_, new_n2840_, new_n2841_, new_n2842_,
    new_n2843_, new_n2844_, new_n2845_, new_n2846_, new_n2847_, new_n2848_,
    new_n2849_, new_n2850_, new_n2851_, new_n2852_, new_n2853_, new_n2854_,
    new_n2855_, new_n2856_, new_n2857_, new_n2858_, new_n2859_, new_n2860_,
    new_n2861_, new_n2862_, new_n2863_, new_n2864_, new_n2865_, new_n2866_,
    new_n2867_, new_n2868_, new_n2869_, new_n2870_, new_n2871_, new_n2872_,
    new_n2873_, new_n2874_, new_n2875_, new_n2876_, new_n2877_, new_n2878_,
    new_n2879_, new_n2880_, new_n2881_, new_n2882_, new_n2883_, new_n2884_,
    new_n2885_, new_n2886_, new_n2887_, new_n2888_, new_n2889_, new_n2890_,
    new_n2891_, new_n2892_, new_n2893_, new_n2894_, new_n2895_, new_n2896_,
    new_n2897_, new_n2898_, new_n2899_, new_n2900_, new_n2901_, new_n2902_,
    new_n2903_, new_n2904_, new_n2905_, new_n2906_, new_n2907_, new_n2908_,
    new_n2909_, new_n2910_, new_n2911_, new_n2912_, new_n2913_, new_n2914_,
    new_n2915_, new_n2916_, new_n2917_, new_n2918_, new_n2919_, new_n2920_,
    new_n2921_, new_n2922_, new_n2923_, new_n2924_, new_n2925_, new_n2926_,
    new_n2927_, new_n2928_, new_n2929_, new_n2930_, new_n2931_, new_n2932_,
    new_n2933_, new_n2934_, new_n2935_, new_n2936_, new_n2937_, new_n2938_,
    new_n2939_, new_n2940_, new_n2941_, new_n2942_, new_n2943_, new_n2944_,
    new_n2945_, new_n2946_, new_n2947_, new_n2948_, new_n2949_, new_n2950_,
    new_n2951_, new_n2952_, new_n2953_, new_n2954_, new_n2955_, new_n2956_,
    new_n2957_, new_n2958_, new_n2959_, new_n2960_, new_n2961_, new_n2962_,
    new_n2963_, new_n2964_, new_n2965_, new_n2966_, new_n2967_, new_n2968_,
    new_n2969_, new_n2970_, new_n2971_, new_n2972_, new_n2973_, new_n2974_,
    new_n2975_, new_n2976_, new_n2977_, new_n2978_, new_n2979_, new_n2980_,
    new_n2981_, new_n2982_, new_n2983_, new_n2984_, new_n2985_, new_n2986_,
    new_n2987_, new_n2988_, new_n2989_, new_n2990_, new_n2991_, new_n2992_,
    new_n2993_, new_n2994_, new_n2995_, new_n2996_, new_n2997_, new_n2998_,
    new_n2999_, new_n3000_, new_n3001_, new_n3002_, new_n3003_, new_n3004_,
    new_n3005_, new_n3006_, new_n3007_, new_n3008_, new_n3009_, new_n3010_,
    new_n3011_, new_n3012_, new_n3013_, new_n3014_, new_n3015_, new_n3016_,
    new_n3017_, new_n3018_, new_n3019_, new_n3020_, new_n3021_, new_n3022_,
    new_n3023_, new_n3024_, new_n3025_, new_n3026_, new_n3027_, new_n3028_,
    new_n3029_, new_n3030_, new_n3031_, new_n3032_, new_n3033_, new_n3034_,
    new_n3035_, new_n3036_, new_n3037_, new_n3038_, new_n3039_, new_n3040_,
    new_n3041_, new_n3042_, new_n3043_, new_n3044_, new_n3045_, new_n3046_,
    new_n3047_, new_n3048_, new_n3049_, new_n3050_, new_n3051_, new_n3052_,
    new_n3053_, new_n3054_, new_n3055_, new_n3056_, new_n3057_, new_n3058_,
    new_n3059_, new_n3060_, new_n3061_, new_n3062_, new_n3063_, new_n3064_,
    new_n3065_, new_n3066_, new_n3067_, new_n3068_, new_n3069_, new_n3070_,
    new_n3071_, new_n3072_, new_n3073_, new_n3074_, new_n3075_, new_n3076_,
    new_n3077_, new_n3078_, new_n3079_, new_n3080_, new_n3081_, new_n3082_,
    new_n3083_, new_n3084_, new_n3085_, new_n3086_, new_n3087_, new_n3088_,
    new_n3089_, new_n3090_, new_n3091_, new_n3092_, new_n3093_, new_n3094_,
    new_n3095_, new_n3096_, new_n3097_, new_n3098_, new_n3099_, new_n3100_,
    new_n3101_, new_n3102_, new_n3103_, new_n3104_, new_n3105_, new_n3106_,
    new_n3107_, new_n3108_, new_n3109_, new_n3110_, new_n3111_, new_n3112_,
    new_n3113_, new_n3114_, new_n3115_, new_n3116_, new_n3117_, new_n3118_,
    new_n3119_, new_n3120_, new_n3121_, new_n3122_, new_n3123_, new_n3124_,
    new_n3125_, new_n3126_, new_n3127_, new_n3128_, new_n3129_, new_n3130_,
    new_n3131_, new_n3132_, new_n3133_, new_n3134_, new_n3135_, new_n3136_,
    new_n3137_, new_n3138_, new_n3139_, new_n3140_, new_n3141_, new_n3142_,
    new_n3143_, new_n3144_, new_n3145_, new_n3146_, new_n3147_, new_n3148_,
    new_n3149_, new_n3150_, new_n3151_, new_n3152_, new_n3153_, new_n3154_,
    new_n3156_, new_n3157_, new_n3158_, new_n3159_, new_n3160_, new_n3161_,
    new_n3162_, new_n3163_, new_n3164_, new_n3165_, new_n3166_, new_n3167_,
    new_n3168_, new_n3169_, new_n3170_, new_n3171_, new_n3172_, new_n3173_,
    new_n3174_, new_n3175_, new_n3176_, new_n3177_, new_n3178_, new_n3179_,
    new_n3180_, new_n3181_, new_n3182_, new_n3183_, new_n3184_, new_n3185_,
    new_n3186_, new_n3187_, new_n3188_, new_n3189_, new_n3190_, new_n3191_,
    new_n3192_, new_n3193_, new_n3194_, new_n3195_, new_n3196_, new_n3197_,
    new_n3198_, new_n3199_, new_n3200_, new_n3201_, new_n3202_, new_n3203_,
    new_n3204_, new_n3205_, new_n3206_, new_n3207_, new_n3208_, new_n3209_,
    new_n3210_, new_n3211_, new_n3212_, new_n3213_, new_n3214_, new_n3215_,
    new_n3216_, new_n3217_, new_n3218_, new_n3219_, new_n3220_, new_n3221_,
    new_n3222_, new_n3223_, new_n3224_, new_n3225_, new_n3226_, new_n3227_,
    new_n3228_, new_n3229_, new_n3230_, new_n3231_, new_n3232_, new_n3233_,
    new_n3234_, new_n3235_, new_n3236_, new_n3237_, new_n3238_, new_n3239_,
    new_n3240_, new_n3241_, new_n3242_, new_n3243_, new_n3244_, new_n3245_,
    new_n3246_, new_n3247_, new_n3248_, new_n3249_, new_n3250_, new_n3251_,
    new_n3252_, new_n3253_, new_n3254_, new_n3255_, new_n3256_, new_n3257_,
    new_n3258_, new_n3259_, new_n3260_, new_n3261_, new_n3262_, new_n3263_,
    new_n3264_, new_n3265_, new_n3266_, new_n3267_, new_n3268_, new_n3269_,
    new_n3270_, new_n3271_, new_n3272_, new_n3273_, new_n3274_, new_n3275_,
    new_n3276_, new_n3277_, new_n3278_, new_n3279_, new_n3280_, new_n3281_,
    new_n3282_, new_n3283_, new_n3284_, new_n3285_, new_n3286_, new_n3287_,
    new_n3288_, new_n3289_, new_n3290_, new_n3291_, new_n3292_, new_n3293_,
    new_n3294_, new_n3295_, new_n3296_, new_n3297_, new_n3298_, new_n3299_,
    new_n3300_, new_n3301_, new_n3302_, new_n3303_, new_n3304_, new_n3305_,
    new_n3306_, new_n3307_, new_n3308_, new_n3309_, new_n3310_, new_n3311_,
    new_n3312_, new_n3313_, new_n3314_, new_n3315_, new_n3316_, new_n3317_,
    new_n3318_, new_n3320_, new_n3321_, new_n3322_, new_n3323_, new_n3324_,
    new_n3325_, new_n3326_, new_n3327_, new_n3328_, new_n3329_, new_n3330_,
    new_n3331_, new_n3332_, new_n3333_, new_n3334_, new_n3335_, new_n3336_,
    new_n3337_, new_n3338_, new_n3339_, new_n3340_, new_n3341_, new_n3342_,
    new_n3343_, new_n3344_, new_n3345_, new_n3346_, new_n3347_, new_n3348_,
    new_n3349_, new_n3350_, new_n3351_, new_n3352_, new_n3353_, new_n3354_,
    new_n3355_, new_n3356_, new_n3357_, new_n3358_, new_n3359_, new_n3360_,
    new_n3361_, new_n3362_, new_n3363_, new_n3364_, new_n3365_, new_n3366_,
    new_n3367_, new_n3368_, new_n3369_, new_n3370_, new_n3371_, new_n3372_,
    new_n3373_, new_n3374_, new_n3375_, new_n3376_, new_n3377_, new_n3378_,
    new_n3379_, new_n3380_, new_n3381_, new_n3382_, new_n3383_, new_n3384_,
    new_n3385_, new_n3386_, new_n3387_, new_n3388_, new_n3389_, new_n3390_,
    new_n3391_, new_n3392_, new_n3393_, new_n3394_, new_n3395_, new_n3396_,
    new_n3397_, new_n3398_, new_n3399_, new_n3400_, new_n3401_, new_n3402_,
    new_n3403_, new_n3404_, new_n3405_, new_n3406_, new_n3407_, new_n3408_,
    new_n3409_, new_n3410_, new_n3411_, new_n3412_, new_n3413_, new_n3414_,
    new_n3415_, new_n3416_, new_n3417_, new_n3418_, new_n3419_, new_n3420_,
    new_n3421_, new_n3422_, new_n3423_, new_n3424_, new_n3425_, new_n3426_,
    new_n3427_, new_n3428_, new_n3429_, new_n3430_, new_n3431_, new_n3432_,
    new_n3433_, new_n3434_, new_n3436_, new_n3437_, new_n3438_, new_n3439_,
    new_n3440_, new_n3441_, new_n3442_, new_n3443_, new_n3444_, new_n3445_,
    new_n3446_, new_n3447_, new_n3448_, new_n3449_, new_n3450_, new_n3451_,
    new_n3452_, new_n3453_, new_n3454_, new_n3455_, new_n3456_, new_n3457_,
    new_n3458_, new_n3459_, new_n3460_, new_n3461_, new_n3462_, new_n3463_,
    new_n3464_, new_n3465_, new_n3466_, new_n3467_, new_n3468_, new_n3469_,
    new_n3470_, new_n3471_, new_n3472_, new_n3473_, new_n3474_, new_n3475_,
    new_n3476_, new_n3477_, new_n3478_, new_n3479_, new_n3480_, new_n3481_,
    new_n3482_, new_n3483_, new_n3484_, new_n3485_, new_n3486_, new_n3487_,
    new_n3488_, new_n3489_, new_n3490_, new_n3491_, new_n3492_, new_n3493_,
    new_n3494_, new_n3495_, new_n3496_, new_n3497_, new_n3498_, new_n3499_,
    new_n3500_, new_n3501_, new_n3502_, new_n3503_, new_n3504_, new_n3505_,
    new_n3506_, new_n3507_, new_n3508_, new_n3509_, new_n3510_, new_n3511_,
    new_n3512_, new_n3513_, new_n3514_, new_n3515_, new_n3516_, new_n3517_,
    new_n3518_, new_n3519_, new_n3520_, new_n3521_, new_n3522_, new_n3523_,
    new_n3524_, new_n3525_, new_n3526_, new_n3527_, new_n3528_, new_n3529_,
    new_n3530_, new_n3531_, new_n3532_, new_n3533_, new_n3534_, new_n3535_,
    new_n3536_, new_n3537_, new_n3538_, new_n3539_, new_n3540_, new_n3541_,
    new_n3542_, new_n3543_, new_n3544_, new_n3545_, new_n3546_, new_n3547_,
    new_n3548_, new_n3549_, new_n3550_, new_n3551_, new_n3552_, new_n3553_,
    new_n3554_, new_n3555_, new_n3556_, new_n3557_, new_n3558_, new_n3559_,
    new_n3560_, new_n3561_, new_n3562_, new_n3563_, new_n3564_, new_n3565_,
    new_n3566_, new_n3567_, new_n3568_, new_n3569_, new_n3570_, new_n3571_,
    new_n3572_, new_n3573_, new_n3574_, new_n3575_, new_n3576_, new_n3577_,
    new_n3578_, new_n3579_, new_n3580_, new_n3581_, new_n3582_, new_n3583_,
    new_n3584_, new_n3586_, new_n3587_, new_n3588_, new_n3589_, new_n3590_,
    new_n3591_, new_n3592_, new_n3593_, new_n3594_, new_n3595_, new_n3596_,
    new_n3597_, new_n3598_, new_n3599_, new_n3600_, new_n3601_, new_n3602_,
    new_n3603_, new_n3604_, new_n3605_, new_n3606_, new_n3607_, new_n3608_,
    new_n3609_, new_n3610_, new_n3611_, new_n3612_, new_n3613_, new_n3614_,
    new_n3615_, new_n3616_, new_n3617_, new_n3618_, new_n3619_, new_n3620_,
    new_n3621_, new_n3622_, new_n3623_, new_n3624_, new_n3625_, new_n3626_,
    new_n3627_, new_n3628_, new_n3629_, new_n3630_, new_n3631_, new_n3632_,
    new_n3633_, new_n3634_, new_n3635_, new_n3636_, new_n3637_, new_n3638_,
    new_n3639_, new_n3640_, new_n3641_, new_n3642_, new_n3643_, new_n3644_,
    new_n3645_, new_n3646_, new_n3647_, new_n3648_, new_n3649_, new_n3650_,
    new_n3651_, new_n3652_, new_n3653_, new_n3654_, new_n3655_, new_n3656_,
    new_n3657_, new_n3658_, new_n3659_, new_n3660_, new_n3661_, new_n3662_,
    new_n3663_, new_n3664_, new_n3665_, new_n3666_, new_n3667_, new_n3668_,
    new_n3669_, new_n3670_, new_n3671_, new_n3672_, new_n3673_, new_n3674_,
    new_n3675_, new_n3676_, new_n3677_, new_n3678_, new_n3679_, new_n3680_,
    new_n3681_, new_n3682_, new_n3683_, new_n3684_, new_n3685_, new_n3686_,
    new_n3687_, new_n3688_, new_n3689_, new_n3690_, new_n3691_, new_n3692_,
    new_n3693_, new_n3694_, new_n3695_, new_n3696_, new_n3697_, new_n3698_,
    new_n3699_, new_n3700_, new_n3701_, new_n3702_, new_n3703_, new_n3704_,
    new_n3705_, new_n3706_, new_n3707_, new_n3708_, new_n3709_, new_n3710_,
    new_n3711_, new_n3712_, new_n3713_, new_n3714_, new_n3715_, new_n3716_,
    new_n3717_, new_n3718_, new_n3719_, new_n3720_, new_n3721_, new_n3722_,
    new_n3723_, new_n3724_, new_n3725_, new_n3726_, new_n3727_, new_n3728_,
    new_n3729_, new_n3730_, new_n3731_, new_n3732_, new_n3733_, new_n3734_,
    new_n3735_, new_n3737_, new_n3738_, new_n3739_, new_n3740_, new_n3741_,
    new_n3742_, new_n3743_, new_n3744_, new_n3745_, new_n3746_, new_n3747_,
    new_n3748_, new_n3749_, new_n3750_, new_n3751_, new_n3752_, new_n3753_,
    new_n3754_, new_n3755_, new_n3756_, new_n3757_, new_n3758_, new_n3759_,
    new_n3760_, new_n3761_, new_n3762_, new_n3763_, new_n3764_, new_n3765_,
    new_n3766_, new_n3767_, new_n3768_, new_n3769_, new_n3770_, new_n3771_,
    new_n3772_, new_n3773_, new_n3774_, new_n3775_, new_n3776_, new_n3777_,
    new_n3778_, new_n3779_, new_n3780_, new_n3781_, new_n3782_, new_n3783_,
    new_n3784_, new_n3785_, new_n3786_, new_n3787_, new_n3788_, new_n3789_,
    new_n3790_, new_n3791_, new_n3792_, new_n3793_, new_n3794_, new_n3795_,
    new_n3796_, new_n3797_, new_n3798_, new_n3799_, new_n3800_, new_n3801_,
    new_n3802_, new_n3803_, new_n3804_, new_n3805_, new_n3806_, new_n3807_,
    new_n3808_, new_n3809_, new_n3810_, new_n3811_, new_n3812_, new_n3813_,
    new_n3814_, new_n3815_, new_n3816_, new_n3817_, new_n3818_, new_n3819_,
    new_n3820_, new_n3821_, new_n3822_, new_n3823_, new_n3824_, new_n3825_,
    new_n3826_, new_n3827_, new_n3828_, new_n3829_, new_n3830_, new_n3831_,
    new_n3832_, new_n3833_, new_n3834_, new_n3835_, new_n3836_, new_n3837_,
    new_n3838_, new_n3839_, new_n3840_, new_n3841_, new_n3842_, new_n3843_,
    new_n3844_, new_n3845_, new_n3846_, new_n3847_, new_n3848_, new_n3849_,
    new_n3850_, new_n3851_, new_n3852_, new_n3853_, new_n3854_, new_n3855_,
    new_n3856_, new_n3857_, new_n3858_, new_n3859_, new_n3860_, new_n3861_,
    new_n3862_, new_n3863_, new_n3864_, new_n3865_, new_n3866_, new_n3867_,
    new_n3868_, new_n3869_, new_n3870_, new_n3871_, new_n3872_, new_n3873_,
    new_n3874_, new_n3875_, new_n3876_, new_n3877_, new_n3878_, new_n3880_,
    new_n3881_, new_n3882_, new_n3883_, new_n3884_, new_n3885_, new_n3886_,
    new_n3887_, new_n3888_, new_n3889_, new_n3890_, new_n3891_, new_n3892_,
    new_n3893_, new_n3894_, new_n3895_, new_n3896_, new_n3897_, new_n3898_,
    new_n3899_, new_n3900_, new_n3901_, new_n3902_, new_n3903_, new_n3904_,
    new_n3905_, new_n3906_, new_n3907_, new_n3908_, new_n3909_, new_n3910_,
    new_n3911_, new_n3912_, new_n3913_, new_n3914_, new_n3915_, new_n3916_,
    new_n3917_, new_n3918_, new_n3919_, new_n3920_, new_n3921_, new_n3922_,
    new_n3923_, new_n3924_, new_n3925_, new_n3926_, new_n3927_, new_n3928_,
    new_n3929_, new_n3930_, new_n3931_, new_n3932_, new_n3933_, new_n3934_,
    new_n3935_, new_n3936_, new_n3937_, new_n3938_, new_n3939_, new_n3940_,
    new_n3941_, new_n3942_, new_n3943_, new_n3944_, new_n3945_, new_n3946_,
    new_n3947_, new_n3948_, new_n3949_, new_n3950_, new_n3951_, new_n3952_,
    new_n3953_, new_n3954_, new_n3955_, new_n3956_, new_n3957_, new_n3958_,
    new_n3959_, new_n3960_, new_n3961_, new_n3962_, new_n3963_, new_n3964_,
    new_n3965_, new_n3966_, new_n3967_, new_n3968_, new_n3969_, new_n3970_,
    new_n3971_, new_n3972_, new_n3973_, new_n3974_, new_n3975_, new_n3976_,
    new_n3977_, new_n3978_, new_n3979_, new_n3980_, new_n3981_, new_n3982_,
    new_n3983_, new_n3984_, new_n3985_, new_n3986_, new_n3987_, new_n3988_,
    new_n3989_, new_n3990_, new_n3991_, new_n3992_, new_n3993_, new_n3994_,
    new_n3995_, new_n3996_, new_n3997_, new_n3998_, new_n3999_, new_n4000_,
    new_n4001_, new_n4002_, new_n4003_, new_n4004_, new_n4005_, new_n4006_,
    new_n4007_, new_n4008_, new_n4009_, new_n4010_, new_n4011_, new_n4012_,
    new_n4013_, new_n4014_, new_n4015_, new_n4016_, new_n4017_, new_n4018_,
    new_n4019_, new_n4021_, new_n4022_, new_n4023_, new_n4024_, new_n4025_,
    new_n4026_, new_n4027_, new_n4028_, new_n4029_, new_n4030_, new_n4031_,
    new_n4032_, new_n4033_, new_n4034_, new_n4035_, new_n4036_, new_n4037_,
    new_n4038_, new_n4039_, new_n4040_, new_n4041_, new_n4042_, new_n4043_,
    new_n4044_, new_n4045_, new_n4046_, new_n4047_, new_n4048_, new_n4049_,
    new_n4050_, new_n4051_, new_n4052_, new_n4053_, new_n4054_, new_n4055_,
    new_n4056_, new_n4057_, new_n4058_, new_n4059_, new_n4060_, new_n4061_,
    new_n4062_, new_n4063_, new_n4064_, new_n4065_, new_n4066_, new_n4067_,
    new_n4068_, new_n4069_, new_n4070_, new_n4071_, new_n4072_, new_n4073_,
    new_n4074_, new_n4075_, new_n4076_, new_n4077_, new_n4078_, new_n4079_,
    new_n4080_, new_n4081_, new_n4082_, new_n4083_, new_n4084_, new_n4085_,
    new_n4086_, new_n4087_, new_n4088_, new_n4089_, new_n4090_, new_n4091_,
    new_n4092_, new_n4093_, new_n4094_, new_n4095_, new_n4096_, new_n4097_,
    new_n4098_, new_n4099_, new_n4100_, new_n4101_, new_n4102_, new_n4103_,
    new_n4104_, new_n4105_, new_n4106_, new_n4107_, new_n4108_, new_n4109_,
    new_n4110_, new_n4111_, new_n4112_, new_n4113_, new_n4114_, new_n4115_,
    new_n4116_, new_n4117_, new_n4118_, new_n4119_, new_n4120_, new_n4121_,
    new_n4122_, new_n4123_, new_n4124_, new_n4125_, new_n4126_, new_n4127_,
    new_n4128_, new_n4129_, new_n4130_, new_n4131_, new_n4132_, new_n4133_,
    new_n4134_, new_n4135_, new_n4136_, new_n4137_, new_n4138_, new_n4139_,
    new_n4140_, new_n4141_, new_n4142_, new_n4143_, new_n4144_, new_n4145_,
    new_n4146_, new_n4147_, new_n4148_, new_n4149_, new_n4150_, new_n4151_,
    new_n4152_, new_n4153_, new_n4154_, new_n4155_, new_n4156_, new_n4157_,
    new_n4158_, new_n4159_, new_n4160_, new_n4161_, new_n4162_, new_n4163_,
    new_n4164_, new_n4165_, new_n4166_, new_n4167_, new_n4168_, new_n4169_,
    new_n4170_, new_n4171_, new_n4173_, new_n4174_, new_n4175_, new_n4176_,
    new_n4177_, new_n4178_, new_n4179_, new_n4180_, new_n4181_, new_n4182_,
    new_n4183_, new_n4184_, new_n4185_, new_n4186_, new_n4187_, new_n4188_,
    new_n4189_, new_n4190_, new_n4191_, new_n4192_, new_n4193_, new_n4194_,
    new_n4195_, new_n4196_, new_n4197_, new_n4198_, new_n4199_, new_n4200_,
    new_n4201_, new_n4202_, new_n4203_, new_n4204_, new_n4205_, new_n4206_,
    new_n4207_, new_n4208_, new_n4209_, new_n4210_, new_n4211_, new_n4212_,
    new_n4213_, new_n4214_, new_n4215_, new_n4216_, new_n4217_, new_n4218_,
    new_n4219_, new_n4220_, new_n4221_, new_n4222_, new_n4223_, new_n4224_,
    new_n4225_, new_n4226_, new_n4227_, new_n4228_, new_n4229_, new_n4230_,
    new_n4231_, new_n4232_, new_n4233_, new_n4234_, new_n4235_, new_n4236_,
    new_n4237_, new_n4238_, new_n4239_, new_n4240_, new_n4241_, new_n4242_,
    new_n4243_, new_n4244_, new_n4245_, new_n4246_, new_n4247_, new_n4248_,
    new_n4249_, new_n4250_, new_n4251_, new_n4252_, new_n4253_, new_n4254_,
    new_n4255_, new_n4256_, new_n4257_, new_n4258_, new_n4259_, new_n4260_,
    new_n4261_, new_n4262_, new_n4263_, new_n4264_, new_n4265_, new_n4266_,
    new_n4267_, new_n4268_, new_n4269_, new_n4270_, new_n4271_, new_n4272_,
    new_n4273_, new_n4274_, new_n4275_, new_n4276_, new_n4277_, new_n4278_,
    new_n4279_, new_n4280_, new_n4281_, new_n4282_, new_n4283_, new_n4284_,
    new_n4285_, new_n4286_, new_n4287_, new_n4288_, new_n4289_, new_n4290_,
    new_n4291_, new_n4292_, new_n4293_, new_n4294_, new_n4295_, new_n4296_,
    new_n4297_, new_n4298_, new_n4299_, new_n4300_, new_n4301_, new_n4302_,
    new_n4303_, new_n4304_, new_n4305_, new_n4306_, new_n4307_, new_n4308_,
    new_n4309_, new_n4310_, new_n4311_, new_n4312_, new_n4314_, new_n4315_,
    new_n4316_, new_n4317_, new_n4318_, new_n4319_, new_n4320_, new_n4321_,
    new_n4322_, new_n4323_, new_n4324_, new_n4325_, new_n4326_, new_n4327_,
    new_n4328_, new_n4329_, new_n4330_, new_n4331_, new_n4332_, new_n4333_,
    new_n4334_, new_n4335_, new_n4336_, new_n4337_, new_n4338_, new_n4339_,
    new_n4340_, new_n4341_, new_n4342_, new_n4343_, new_n4344_, new_n4345_,
    new_n4346_, new_n4347_, new_n4348_, new_n4349_, new_n4350_, new_n4351_,
    new_n4352_, new_n4353_, new_n4354_, new_n4355_, new_n4356_, new_n4357_,
    new_n4358_, new_n4359_, new_n4360_, new_n4361_, new_n4362_, new_n4363_,
    new_n4364_, new_n4365_, new_n4366_, new_n4367_, new_n4368_, new_n4369_,
    new_n4370_, new_n4371_, new_n4372_, new_n4373_, new_n4374_, new_n4375_,
    new_n4376_, new_n4377_, new_n4378_, new_n4379_, new_n4380_, new_n4381_,
    new_n4382_, new_n4383_, new_n4384_, new_n4385_, new_n4386_, new_n4387_,
    new_n4388_, new_n4389_, new_n4390_, new_n4391_, new_n4392_, new_n4393_,
    new_n4394_, new_n4395_, new_n4396_, new_n4397_, new_n4398_, new_n4399_,
    new_n4400_, new_n4401_, new_n4402_, new_n4403_, new_n4404_, new_n4405_,
    new_n4406_, new_n4407_, new_n4408_, new_n4409_, new_n4410_, new_n4411_,
    new_n4412_, new_n4413_, new_n4414_, new_n4415_, new_n4416_, new_n4417_,
    new_n4418_, new_n4419_, new_n4420_, new_n4421_, new_n4422_, new_n4423_,
    new_n4424_, new_n4425_, new_n4426_, new_n4427_, new_n4428_, new_n4429_,
    new_n4430_, new_n4431_, new_n4432_, new_n4433_, new_n4434_, new_n4435_,
    new_n4436_, new_n4437_, new_n4438_, new_n4439_, new_n4440_, new_n4441_,
    new_n4442_, new_n4443_, new_n4444_, new_n4445_, new_n4446_, new_n4447_,
    new_n4448_, new_n4449_, new_n4450_, new_n4451_, new_n4452_, new_n4453_,
    new_n4455_, new_n4456_, new_n4457_, new_n4458_, new_n4459_, new_n4460_,
    new_n4461_, new_n4462_, new_n4463_, new_n4464_, new_n4465_, new_n4466_,
    new_n4467_, new_n4468_, new_n4469_, new_n4470_, new_n4471_, new_n4472_,
    new_n4473_, new_n4474_, new_n4475_, new_n4476_, new_n4477_, new_n4478_,
    new_n4479_, new_n4480_, new_n4481_, new_n4482_, new_n4483_, new_n4484_,
    new_n4485_, new_n4486_, new_n4487_, new_n4488_, new_n4489_, new_n4490_,
    new_n4491_, new_n4492_, new_n4493_, new_n4494_, new_n4495_, new_n4496_,
    new_n4497_, new_n4498_, new_n4499_, new_n4500_, new_n4501_, new_n4502_,
    new_n4503_, new_n4504_, new_n4505_, new_n4506_, new_n4507_, new_n4508_,
    new_n4509_, new_n4510_, new_n4511_, new_n4512_, new_n4513_, new_n4514_,
    new_n4515_, new_n4516_, new_n4517_, new_n4518_, new_n4519_, new_n4520_,
    new_n4521_, new_n4522_, new_n4523_, new_n4524_, new_n4525_, new_n4526_,
    new_n4527_, new_n4528_, new_n4529_, new_n4530_, new_n4531_, new_n4532_,
    new_n4533_, new_n4534_, new_n4535_, new_n4536_, new_n4537_, new_n4538_,
    new_n4539_, new_n4540_, new_n4541_, new_n4542_, new_n4543_, new_n4544_,
    new_n4545_, new_n4546_, new_n4547_, new_n4548_, new_n4549_, new_n4550_,
    new_n4551_, new_n4552_, new_n4553_, new_n4554_, new_n4555_, new_n4556_,
    new_n4557_, new_n4558_, new_n4559_, new_n4560_, new_n4561_, new_n4562_,
    new_n4563_, new_n4564_, new_n4565_, new_n4566_, new_n4567_, new_n4568_,
    new_n4569_, new_n4570_, new_n4571_, new_n4572_, new_n4573_, new_n4574_,
    new_n4575_, new_n4576_, new_n4577_, new_n4578_, new_n4579_, new_n4580_,
    new_n4581_, new_n4582_, new_n4583_, new_n4584_, new_n4585_, new_n4586_,
    new_n4587_, new_n4588_, new_n4589_, new_n4590_, new_n4591_, new_n4592_,
    new_n4593_, new_n4594_, new_n4595_, new_n4596_, new_n4597_, new_n4598_,
    new_n4599_, new_n4600_, new_n4601_, new_n4602_, new_n4603_, new_n4605_,
    new_n4606_, new_n4607_, new_n4608_, new_n4609_, new_n4610_, new_n4611_,
    new_n4612_, new_n4613_, new_n4614_, new_n4615_, new_n4616_, new_n4617_,
    new_n4618_, new_n4619_, new_n4620_, new_n4621_, new_n4622_, new_n4623_,
    new_n4624_, new_n4625_, new_n4626_, new_n4627_, new_n4628_, new_n4629_,
    new_n4630_, new_n4631_, new_n4632_, new_n4633_, new_n4634_, new_n4635_,
    new_n4636_, new_n4637_, new_n4638_, new_n4639_, new_n4640_, new_n4641_,
    new_n4642_, new_n4643_, new_n4644_, new_n4645_, new_n4646_, new_n4647_,
    new_n4648_, new_n4649_, new_n4650_, new_n4651_, new_n4652_, new_n4653_,
    new_n4654_, new_n4655_, new_n4656_, new_n4657_, new_n4658_, new_n4659_,
    new_n4660_, new_n4661_, new_n4662_, new_n4663_, new_n4664_, new_n4665_,
    new_n4666_, new_n4667_, new_n4668_, new_n4669_, new_n4670_, new_n4671_,
    new_n4672_, new_n4673_, new_n4674_, new_n4675_, new_n4676_, new_n4677_,
    new_n4678_, new_n4679_, new_n4680_, new_n4681_, new_n4682_, new_n4683_,
    new_n4684_, new_n4685_, new_n4686_, new_n4687_, new_n4688_, new_n4689_,
    new_n4690_, new_n4691_, new_n4692_, new_n4693_, new_n4694_, new_n4695_,
    new_n4696_, new_n4697_, new_n4698_, new_n4699_, new_n4700_, new_n4701_,
    new_n4702_, new_n4703_, new_n4704_, new_n4705_, new_n4706_, new_n4707_,
    new_n4708_, new_n4709_, new_n4710_, new_n4711_, new_n4712_, new_n4713_,
    new_n4714_, new_n4715_, new_n4716_, new_n4717_, new_n4718_, new_n4719_,
    new_n4720_, new_n4721_, new_n4722_, new_n4723_, new_n4724_, new_n4725_,
    new_n4726_, new_n4727_, new_n4728_, new_n4729_, new_n4730_, new_n4731_,
    new_n4732_, new_n4733_, new_n4734_, new_n4735_, new_n4736_, new_n4737_,
    new_n4738_, new_n4739_, new_n4740_, new_n4741_, new_n4742_, new_n4743_,
    new_n4744_, new_n4745_, new_n4746_, new_n4747_, new_n4748_, new_n4749_,
    new_n4750_, new_n4751_, new_n4752_, new_n4753_, new_n4755_, new_n4756_,
    new_n4757_, new_n4758_, new_n4759_, new_n4760_, new_n4761_, new_n4762_,
    new_n4763_, new_n4764_, new_n4765_, new_n4766_, new_n4767_, new_n4768_,
    new_n4769_, new_n4770_, new_n4771_, new_n4772_, new_n4773_, new_n4774_,
    new_n4775_, new_n4776_, new_n4777_, new_n4778_, new_n4779_, new_n4780_,
    new_n4781_, new_n4782_, new_n4783_, new_n4784_, new_n4785_, new_n4786_,
    new_n4787_, new_n4788_, new_n4789_, new_n4790_, new_n4791_, new_n4792_,
    new_n4793_, new_n4794_, new_n4795_, new_n4796_, new_n4797_, new_n4798_,
    new_n4799_, new_n4800_, new_n4801_, new_n4802_, new_n4803_, new_n4804_,
    new_n4805_, new_n4806_, new_n4807_, new_n4808_, new_n4809_, new_n4810_,
    new_n4811_, new_n4812_, new_n4813_, new_n4814_, new_n4815_, new_n4816_,
    new_n4817_, new_n4818_, new_n4819_, new_n4820_, new_n4821_, new_n4822_,
    new_n4823_, new_n4824_, new_n4825_, new_n4826_, new_n4827_, new_n4828_,
    new_n4829_, new_n4830_, new_n4831_, new_n4832_, new_n4833_, new_n4834_,
    new_n4835_, new_n4836_, new_n4837_, new_n4838_, new_n4839_, new_n4840_,
    new_n4841_, new_n4842_, new_n4843_, new_n4844_, new_n4845_, new_n4846_,
    new_n4847_, new_n4848_, new_n4849_, new_n4850_, new_n4851_, new_n4852_,
    new_n4853_, new_n4854_, new_n4855_, new_n4856_, new_n4857_, new_n4858_,
    new_n4859_, new_n4860_, new_n4861_, new_n4862_, new_n4863_, new_n4864_,
    new_n4865_, new_n4866_, new_n4867_, new_n4868_, new_n4869_, new_n4870_,
    new_n4871_, new_n4872_, new_n4873_, new_n4874_, new_n4875_, new_n4876_,
    new_n4877_, new_n4878_, new_n4879_, new_n4880_, new_n4881_, new_n4882_,
    new_n4883_, new_n4884_, new_n4885_, new_n4886_, new_n4887_, new_n4888_,
    new_n4889_, new_n4890_, new_n4891_, new_n4892_, new_n4893_, new_n4894_,
    new_n4895_, new_n4896_, new_n4897_, new_n4898_, new_n4899_, new_n4900_,
    new_n4901_, new_n4902_, new_n4903_, new_n4904_, new_n4905_, new_n4906_,
    new_n4907_, new_n4908_, new_n4909_, new_n4910_, new_n4911_, new_n4912_,
    new_n4913_, new_n4914_, new_n4915_, new_n4916_, new_n4917_, new_n4918_,
    new_n4919_, new_n4920_, new_n4921_, new_n4922_, new_n4923_, new_n4924_,
    new_n4925_, new_n4926_, new_n4927_, new_n4928_, new_n4929_, new_n4930_,
    new_n4931_, new_n4932_, new_n4933_, new_n4934_, new_n4935_, new_n4936_,
    new_n4937_, new_n4938_, new_n4939_, new_n4940_, new_n4941_, new_n4942_,
    new_n4943_, new_n4944_, new_n4945_, new_n4946_, new_n4947_, new_n4948_,
    new_n4949_, new_n4950_, new_n4951_, new_n4952_, new_n4953_, new_n4954_,
    new_n4955_, new_n4956_, new_n4957_, new_n4958_, new_n4959_, new_n4960_,
    new_n4961_, new_n4962_, new_n4963_, new_n4964_, new_n4965_, new_n4966_,
    new_n4967_, new_n4968_, new_n4969_, new_n4970_, new_n4971_, new_n4972_,
    new_n4973_, new_n4974_, new_n4975_, new_n4976_, new_n4977_, new_n4978_,
    new_n4979_, new_n4982_, new_n4983_, new_n4984_, new_n4985_, new_n4986_,
    new_n4987_, new_n4988_, new_n4989_, new_n4990_, new_n4991_, new_n4992_,
    new_n4993_, new_n4994_, new_n4995_, new_n4996_, new_n4997_, new_n4998_,
    new_n4999_, new_n5000_, new_n5001_, new_n5002_, new_n5003_, new_n5004_,
    new_n5005_, new_n5006_, new_n5007_, new_n5008_, new_n5009_, new_n5010_,
    new_n5011_, new_n5012_, new_n5013_, new_n5014_, new_n5015_, new_n5016_,
    new_n5017_, new_n5018_, new_n5019_, new_n5020_, new_n5021_, new_n5022_,
    new_n5023_, new_n5024_, new_n5025_, new_n5026_, new_n5027_, new_n5028_,
    new_n5029_, new_n5030_, new_n5031_, new_n5033_, new_n5034_, new_n5035_,
    new_n5036_, new_n5037_, new_n5038_, new_n5039_, new_n5040_, new_n5041_,
    new_n5042_, new_n5043_, new_n5044_, new_n5045_, new_n5046_, new_n5047_,
    new_n5048_, new_n5049_, new_n5050_, new_n5051_, new_n5052_, new_n5053_,
    new_n5054_, new_n5055_, new_n5056_, new_n5057_, new_n5058_, new_n5059_,
    new_n5060_, new_n5061_, new_n5062_, new_n5063_, new_n5064_, new_n5065_,
    new_n5066_, new_n5067_, new_n5068_, new_n5069_, new_n5070_, new_n5071_,
    new_n5072_, new_n5073_, new_n5074_, new_n5075_, new_n5076_, new_n5077_,
    new_n5078_, new_n5079_, new_n5080_, new_n5081_, new_n5082_, new_n5083_,
    new_n5084_, new_n5085_, new_n5086_, new_n5087_, new_n5088_, new_n5089_,
    new_n5090_, new_n5091_, new_n5092_, new_n5093_, new_n5094_, new_n5095_,
    new_n5096_, new_n5098_, new_n5099_, new_n5100_, new_n5101_, new_n5102_,
    new_n5103_, new_n5104_, new_n5105_, new_n5106_, new_n5107_, new_n5108_,
    new_n5109_, new_n5110_, new_n5111_, new_n5112_, new_n5113_, new_n5114_,
    new_n5117_, new_n5118_, new_n5119_, new_n5120_, new_n5121_, new_n5122_,
    new_n5123_, new_n5124_, new_n5125_, new_n5126_, new_n5127_, new_n5128_,
    new_n5129_, new_n5130_, new_n5131_, new_n5132_, new_n5133_, new_n5134_,
    new_n5135_, new_n5136_, new_n5137_, new_n5138_, new_n5139_, new_n5140_,
    new_n5141_, new_n5142_, new_n5143_, new_n5144_, new_n5145_, new_n5146_,
    new_n5147_, new_n5148_, new_n5149_, new_n5150_, new_n5151_, new_n5152_,
    new_n5153_, new_n5154_, new_n5155_, new_n5156_, new_n5158_, new_n5159_,
    new_n5160_, new_n5161_, new_n5162_, new_n5163_, new_n5164_, new_n5165_,
    new_n5166_, new_n5167_, new_n5168_, new_n5169_, new_n5170_, new_n5171_,
    new_n5172_, new_n5173_, new_n5174_, new_n5175_, new_n5176_, new_n5177_,
    new_n5178_, new_n5179_, new_n5180_, new_n5181_, new_n5182_, new_n5183_,
    new_n5184_, new_n5185_, new_n5186_, new_n5187_, new_n5188_, new_n5189_,
    new_n5190_, new_n5191_, new_n5192_, new_n5193_, new_n5194_, new_n5195_,
    new_n5196_, new_n5197_, new_n5198_, new_n5199_, new_n5200_, new_n5201_,
    new_n5202_, new_n5203_, new_n5204_, new_n5205_, new_n5206_, new_n5207_,
    new_n5208_, new_n5209_, new_n5210_, new_n5211_, new_n5212_, new_n5213_,
    new_n5214_, new_n5215_, new_n5216_, new_n5217_, new_n5218_, new_n5219_,
    new_n5220_, new_n5221_, new_n5222_, new_n5223_, new_n5224_, new_n5225_,
    new_n5226_, new_n5227_, new_n5228_, new_n5229_, new_n5230_, new_n5231_,
    new_n5232_, new_n5233_, new_n5234_, new_n5235_, new_n5236_, new_n5237_,
    new_n5238_, new_n5239_, new_n5240_, new_n5241_, new_n5242_, new_n5243_,
    new_n5244_, new_n5245_, new_n5246_, new_n5247_, new_n5248_, new_n5249_,
    new_n5250_, new_n5251_, new_n5252_, new_n5253_, new_n5254_, new_n5255_,
    new_n5256_, new_n5257_, new_n5258_, new_n5259_, new_n5260_, new_n5261_,
    new_n5262_, new_n5263_, new_n5264_, new_n5265_, new_n5266_, new_n5267_,
    new_n5268_, new_n5269_, new_n5270_, new_n5271_, new_n5272_, new_n5273_,
    new_n5274_, new_n5275_, new_n5276_, new_n5277_, new_n5278_, new_n5279_,
    new_n5280_, new_n5281_, new_n5282_, new_n5283_, new_n5284_, new_n5285_,
    new_n5286_, new_n5287_, new_n5288_, new_n5289_, new_n5290_, new_n5291_,
    new_n5292_, new_n5293_, new_n5294_, new_n5295_, new_n5296_, new_n5297_,
    new_n5298_, new_n5299_, new_n5300_, new_n5301_, new_n5302_, new_n5303_,
    new_n5304_, new_n5305_, new_n5306_, new_n5307_, new_n5308_, new_n5309_,
    new_n5310_, new_n5311_, new_n5312_, new_n5313_, new_n5314_, new_n5315_,
    new_n5316_, new_n5317_, new_n5318_, new_n5319_, new_n5320_, new_n5321_,
    new_n5322_, new_n5323_, new_n5324_, new_n5325_, new_n5326_, new_n5327_,
    new_n5328_, new_n5329_, new_n5331_, new_n5332_, new_n5333_, new_n5334_,
    new_n5335_, new_n5336_, new_n5337_, new_n5338_, new_n5339_, new_n5340_,
    new_n5341_, new_n5342_, new_n5343_, new_n5344_, new_n5345_, new_n5346_,
    new_n5347_, new_n5348_, new_n5349_, new_n5350_, new_n5351_, new_n5352_,
    new_n5353_, new_n5354_, new_n5355_, new_n5356_, new_n5357_, new_n5358_,
    new_n5359_, new_n5360_, new_n5361_, new_n5362_, new_n5363_, new_n5364_,
    new_n5365_, new_n5366_, new_n5367_, new_n5368_, new_n5369_, new_n5370_,
    new_n5371_, new_n5372_, new_n5373_, new_n5374_, new_n5375_, new_n5376_,
    new_n5377_, new_n5378_, new_n5379_, new_n5380_, new_n5381_, new_n5382_,
    new_n5383_, new_n5384_, new_n5385_, new_n5386_, new_n5387_, new_n5388_,
    new_n5389_, new_n5390_, new_n5391_, new_n5392_, new_n5393_, new_n5394_,
    new_n5395_, new_n5396_, new_n5397_, new_n5398_, new_n5399_, new_n5400_,
    new_n5401_, new_n5402_, new_n5403_, new_n5404_, new_n5405_, new_n5406_,
    new_n5407_, new_n5408_, new_n5410_, new_n5411_, new_n5412_, new_n5413_,
    new_n5414_, new_n5415_, new_n5416_, new_n5417_, new_n5418_, new_n5419_,
    new_n5420_, new_n5421_, new_n5422_, new_n5423_, new_n5424_, new_n5425_,
    new_n5426_, new_n5427_, new_n5428_, new_n5429_, new_n5430_, new_n5431_,
    new_n5432_, new_n5433_, new_n5434_, new_n5435_, new_n5436_, new_n5437_,
    new_n5438_, new_n5439_, new_n5440_, new_n5441_, new_n5442_, new_n5443_,
    new_n5444_, new_n5445_, new_n5446_, new_n5447_, new_n5448_, new_n5449_,
    new_n5450_, new_n5451_, new_n5452_, new_n5453_, new_n5454_, new_n5455_,
    new_n5456_, new_n5457_, new_n5458_, new_n5459_, new_n5460_, new_n5461_,
    new_n5462_, new_n5463_, new_n5464_, new_n5465_, new_n5466_, new_n5467_,
    new_n5468_, new_n5469_, new_n5470_, new_n5471_, new_n5472_, new_n5473_,
    new_n5474_, new_n5475_, new_n5476_, new_n5477_, new_n5478_, new_n5479_,
    new_n5480_, new_n5481_, new_n5482_, new_n5483_, new_n5484_, new_n5485_,
    new_n5486_, new_n5487_, new_n5488_, new_n5489_, new_n5490_, new_n5491_,
    new_n5492_, new_n5493_, new_n5494_, new_n5496_, new_n5497_, new_n5498_,
    new_n5499_, new_n5500_, new_n5501_, new_n5502_, new_n5503_, new_n5504_,
    new_n5505_, new_n5506_, new_n5507_, new_n5508_, new_n5509_, new_n5510_,
    new_n5511_, new_n5512_, new_n5513_, new_n5514_, new_n5515_, new_n5516_,
    new_n5517_, new_n5518_, new_n5519_, new_n5520_, new_n5521_, new_n5522_,
    new_n5523_, new_n5524_, new_n5525_, new_n5526_, new_n5527_, new_n5528_,
    new_n5529_, new_n5530_, new_n5531_, new_n5532_, new_n5533_, new_n5534_,
    new_n5535_, new_n5536_, new_n5537_, new_n5538_, new_n5539_, new_n5540_,
    new_n5541_, new_n5542_, new_n5543_, new_n5544_, new_n5545_, new_n5546_,
    new_n5547_, new_n5548_, new_n5549_, new_n5550_, new_n5551_, new_n5552_,
    new_n5553_, new_n5555_, new_n5556_, new_n5557_, new_n5558_, new_n5559_,
    new_n5560_, new_n5561_, new_n5562_, new_n5563_, new_n5564_, new_n5565_,
    new_n5566_, new_n5567_, new_n5568_, new_n5569_, new_n5570_, new_n5571_,
    new_n5572_, new_n5573_, new_n5574_, new_n5575_, new_n5576_, new_n5577_,
    new_n5578_, new_n5579_, new_n5580_, new_n5581_, new_n5582_, new_n5583_,
    new_n5584_, new_n5585_, new_n5586_, new_n5587_, new_n5588_, new_n5589_,
    new_n5590_, new_n5591_, new_n5592_, new_n5593_, new_n5594_, new_n5595_,
    new_n5596_, new_n5597_, new_n5598_, new_n5599_, new_n5600_, new_n5601_,
    new_n5602_, new_n5603_, new_n5604_, new_n5605_, new_n5606_, new_n5607_,
    new_n5608_, new_n5609_, new_n5610_, new_n5611_, new_n5613_, new_n5614_,
    new_n5615_, new_n5616_, new_n5617_, new_n5618_, new_n5619_, new_n5620_,
    new_n5621_, new_n5622_, new_n5623_, new_n5624_, new_n5625_, new_n5626_,
    new_n5627_, new_n5628_, new_n5629_, new_n5630_, new_n5631_, new_n5632_,
    new_n5633_, new_n5634_, new_n5635_, new_n5636_, new_n5637_, new_n5638_,
    new_n5639_, new_n5640_, new_n5641_, new_n5642_, new_n5643_, new_n5644_,
    new_n5645_, new_n5646_, new_n5647_, new_n5648_, new_n5649_, new_n5650_,
    new_n5651_, new_n5652_, new_n5653_, new_n5654_, new_n5655_, new_n5656_,
    new_n5657_, new_n5658_, new_n5659_, new_n5660_, new_n5661_, new_n5662_,
    new_n5663_, new_n5664_, new_n5665_, new_n5666_, new_n5667_, new_n5668_,
    new_n5669_, new_n5671_, new_n5672_, new_n5673_, new_n5674_, new_n5675_,
    new_n5676_, new_n5677_, new_n5678_, new_n5679_, new_n5680_, new_n5681_,
    new_n5682_, new_n5683_, new_n5684_, new_n5685_, new_n5686_, new_n5687_,
    new_n5688_, new_n5689_, new_n5690_, new_n5691_, new_n5692_, new_n5693_,
    new_n5694_, new_n5695_, new_n5696_, new_n5697_, new_n5698_, new_n5699_,
    new_n5700_, new_n5701_, new_n5702_, new_n5703_, new_n5704_, new_n5705_,
    new_n5706_, new_n5707_, new_n5708_, new_n5709_, new_n5710_, new_n5711_,
    new_n5712_, new_n5713_, new_n5714_, new_n5715_, new_n5716_, new_n5717_,
    new_n5718_, new_n5719_, new_n5720_, new_n5721_, new_n5722_, new_n5723_,
    new_n5724_, new_n5725_, new_n5726_, new_n5727_, new_n5728_, new_n5730_,
    new_n5731_, new_n5732_, new_n5733_, new_n5734_, new_n5735_, new_n5736_,
    new_n5737_, new_n5738_, new_n5739_, new_n5740_, new_n5741_, new_n5742_,
    new_n5743_, new_n5744_, new_n5745_, new_n5746_, new_n5747_, new_n5748_,
    new_n5749_, new_n5750_, new_n5751_, new_n5752_, new_n5753_, new_n5754_,
    new_n5755_, new_n5756_, new_n5757_, new_n5758_, new_n5759_, new_n5760_,
    new_n5761_, new_n5762_, new_n5763_, new_n5764_, new_n5765_, new_n5766_,
    new_n5767_, new_n5768_, new_n5769_, new_n5770_, new_n5771_, new_n5772_,
    new_n5773_, new_n5774_, new_n5775_, new_n5776_, new_n5777_, new_n5778_,
    new_n5779_, new_n5780_, new_n5781_, new_n5782_, new_n5783_, new_n5784_,
    new_n5785_, new_n5787_, new_n5788_, new_n5789_, new_n5790_, new_n5791_,
    new_n5792_, new_n5793_, new_n5794_, new_n5795_, new_n5796_, new_n5797_,
    new_n5798_, new_n5799_, new_n5800_, new_n5801_, new_n5802_, new_n5803_,
    new_n5804_, new_n5805_, new_n5806_, new_n5807_, new_n5808_, new_n5809_,
    new_n5810_, new_n5811_, new_n5812_, new_n5813_, new_n5814_, new_n5815_,
    new_n5816_, new_n5817_, new_n5818_, new_n5819_, new_n5820_, new_n5821_,
    new_n5822_, new_n5823_, new_n5824_, new_n5827_, new_n5828_, new_n5829_,
    new_n5830_, new_n5831_, new_n5832_, new_n5833_, new_n5834_, new_n5835_,
    new_n5836_, new_n5837_, new_n5838_, new_n5839_, new_n5840_, new_n5841_,
    new_n5842_, new_n5843_, new_n5844_, new_n5845_, new_n5846_, new_n5847_,
    new_n5848_, new_n5849_, new_n5850_, new_n5851_, new_n5852_, new_n5853_,
    new_n5854_, new_n5855_, new_n5856_, new_n5857_, new_n5858_, new_n5860_,
    new_n5861_, new_n5862_, new_n5863_, new_n5865_, new_n5867_, new_n5869_,
    new_n5871_, new_n5872_, new_n5873_, new_n5874_, new_n5875_, new_n5876_,
    new_n5877_, new_n5878_, new_n5879_, new_n5880_, new_n5881_, new_n5882_,
    new_n5883_, new_n5884_, new_n5885_, new_n5886_, new_n5887_, new_n5888_,
    new_n5889_, new_n5890_, new_n5891_, new_n5892_, new_n5893_, new_n5894_,
    new_n5895_, new_n5896_, new_n5897_, new_n5898_, new_n5899_, new_n5900_,
    new_n5901_, new_n5902_, new_n5903_, new_n5904_, new_n5905_, new_n5906_,
    new_n5907_, new_n5908_, new_n5909_, new_n5910_, new_n5911_, new_n5912_,
    new_n5913_, new_n5914_, new_n5915_, new_n5916_, new_n5917_, new_n5918_,
    new_n5919_, new_n5920_, new_n5921_, new_n5922_, new_n5923_, new_n5924_,
    new_n5925_, new_n5926_, new_n5927_, new_n5928_, new_n5929_, new_n5930_,
    new_n5931_, new_n5932_, new_n5933_, new_n5934_, new_n5935_, new_n5936_,
    new_n5937_, new_n5938_, new_n5939_, new_n5940_, new_n5941_, new_n5942_,
    new_n5943_, new_n5944_, new_n5945_, new_n5946_, new_n5947_, new_n5948_,
    new_n5949_, new_n5950_, new_n5951_, new_n5952_, new_n5953_, new_n5954_,
    new_n5955_, new_n5956_, new_n5957_, new_n5958_, new_n5959_, new_n5960_,
    new_n5961_, new_n5962_, new_n5963_, new_n5964_, new_n5965_, new_n5966_,
    new_n5967_, new_n5968_, new_n5969_, new_n5970_, new_n5971_, new_n5972_,
    new_n5973_, new_n5974_, new_n5975_, new_n5976_, new_n5977_, new_n5978_,
    new_n5979_, new_n5980_, new_n5981_, new_n5982_, new_n5983_, new_n5984_,
    new_n5985_, new_n5986_, new_n5987_, new_n5988_, new_n5989_, new_n5990_,
    new_n5991_, new_n5992_, new_n5993_, new_n5994_, new_n5995_, new_n5996_,
    new_n5997_, new_n5998_, new_n5999_, new_n6000_, new_n6001_, new_n6002_,
    new_n6003_, new_n6004_, new_n6005_, new_n6006_, new_n6007_, new_n6008_,
    new_n6009_, new_n6010_, new_n6011_, new_n6012_, new_n6013_, new_n6014_,
    new_n6015_, new_n6016_, new_n6017_, new_n6018_, new_n6019_, new_n6020_,
    new_n6021_, new_n6022_, new_n6023_, new_n6024_, new_n6025_, new_n6026_,
    new_n6027_, new_n6028_, new_n6029_, new_n6030_, new_n6031_, new_n6032_,
    new_n6033_, new_n6034_, new_n6035_, new_n6036_, new_n6037_, new_n6038_,
    new_n6039_, new_n6040_, new_n6041_, new_n6042_, new_n6043_, new_n6044_,
    new_n6045_, new_n6046_, new_n6047_, new_n6048_, new_n6049_, new_n6050_,
    new_n6051_, new_n6052_, new_n6053_, new_n6054_, new_n6055_, new_n6056_,
    new_n6057_, new_n6058_, new_n6059_, new_n6060_, new_n6061_, new_n6062_,
    new_n6063_, new_n6064_, new_n6065_, new_n6066_, new_n6067_, new_n6068_,
    new_n6069_, new_n6070_, new_n6071_, new_n6072_, new_n6073_, new_n6074_,
    new_n6075_, new_n6076_, new_n6077_, new_n6078_, new_n6079_, new_n6080_,
    new_n6081_, new_n6082_, new_n6083_, new_n6084_, new_n6085_, new_n6086_,
    new_n6087_, new_n6088_, new_n6089_, new_n6090_, new_n6091_, new_n6092_,
    new_n6093_, new_n6094_, new_n6095_, new_n6096_, new_n6097_, new_n6098_,
    new_n6099_, new_n6100_, new_n6101_, new_n6102_, new_n6103_, new_n6104_,
    new_n6105_, new_n6106_, new_n6107_, new_n6108_, new_n6109_, new_n6110_,
    new_n6111_, new_n6112_, new_n6113_, new_n6114_, new_n6115_, new_n6116_,
    new_n6117_, new_n6118_, new_n6119_, new_n6120_, new_n6121_, new_n6122_,
    new_n6123_, new_n6124_, new_n6125_, new_n6126_, new_n6127_, new_n6128_,
    new_n6129_, new_n6130_, new_n6131_, new_n6132_, new_n6133_, new_n6134_,
    new_n6135_, new_n6136_, new_n6137_, new_n6138_, new_n6139_, new_n6140_,
    new_n6141_, new_n6142_, new_n6143_, new_n6144_, new_n6145_, new_n6146_,
    new_n6147_, new_n6148_, new_n6149_, new_n6150_, new_n6151_, new_n6152_,
    new_n6153_, new_n6154_, new_n6155_, new_n6156_, new_n6157_, new_n6158_,
    new_n6159_, new_n6160_, new_n6161_, new_n6162_, new_n6163_, new_n6164_,
    new_n6165_, new_n6166_, new_n6167_, new_n6168_, new_n6169_, new_n6170_,
    new_n6171_, new_n6172_, new_n6173_, new_n6174_, new_n6175_, new_n6176_,
    new_n6177_, new_n6178_, new_n6179_, new_n6180_, new_n6181_, new_n6182_,
    new_n6183_, new_n6184_, new_n6185_, new_n6186_, new_n6187_, new_n6188_,
    new_n6189_, new_n6190_, new_n6191_, new_n6192_, new_n6193_, new_n6194_,
    new_n6195_, new_n6196_, new_n6197_, new_n6198_, new_n6199_, new_n6200_,
    new_n6201_, new_n6202_, new_n6203_, new_n6204_, new_n6205_, new_n6206_,
    new_n6207_, new_n6208_, new_n6209_, new_n6210_, new_n6211_, new_n6212_,
    new_n6213_, new_n6214_, new_n6215_, new_n6216_, new_n6217_, new_n6218_,
    new_n6219_, new_n6220_, new_n6221_, new_n6222_, new_n6223_, new_n6224_,
    new_n6225_, new_n6226_, new_n6227_, new_n6228_, new_n6229_, new_n6230_,
    new_n6231_, new_n6232_, new_n6233_, new_n6234_, new_n6235_, new_n6236_,
    new_n6237_, new_n6238_, new_n6239_, new_n6240_, new_n6241_, new_n6242_,
    new_n6243_, new_n6244_, new_n6245_, new_n6246_, new_n6247_, new_n6248_,
    new_n6249_, new_n6250_, new_n6251_, new_n6252_, new_n6253_, new_n6254_,
    new_n6255_, new_n6256_, new_n6257_, new_n6258_, new_n6259_, new_n6260_,
    new_n6261_, new_n6262_, new_n6263_, new_n6264_, new_n6265_, new_n6266_,
    new_n6267_, new_n6268_, new_n6269_, new_n6270_, new_n6271_, new_n6272_,
    new_n6273_, new_n6274_, new_n6275_, new_n6276_, new_n6277_, new_n6278_,
    new_n6279_, new_n6280_, new_n6281_, new_n6282_, new_n6283_, new_n6284_,
    new_n6285_, new_n6286_, new_n6287_, new_n6288_, new_n6289_, new_n6290_,
    new_n6291_, new_n6292_, new_n6293_, new_n6294_, new_n6295_, new_n6296_,
    new_n6297_, new_n6298_, new_n6299_, new_n6300_, new_n6301_, new_n6302_,
    new_n6303_, new_n6304_, new_n6305_, new_n6306_, new_n6307_, new_n6308_,
    new_n6309_, new_n6310_, new_n6311_, new_n6312_, new_n6313_, new_n6314_,
    new_n6315_, new_n6316_, new_n6317_, new_n6318_, new_n6319_, new_n6320_,
    new_n6321_, new_n6322_, new_n6323_, new_n6324_, new_n6325_, new_n6326_,
    new_n6327_, new_n6328_, new_n6329_, new_n6330_, new_n6331_, new_n6332_,
    new_n6333_, new_n6334_, new_n6335_, new_n6336_, new_n6337_, new_n6338_,
    new_n6339_, new_n6340_, new_n6341_, new_n6342_, new_n6343_, new_n6344_,
    new_n6345_, new_n6346_, new_n6347_, new_n6348_, new_n6349_, new_n6350_,
    new_n6351_, new_n6352_, new_n6353_, new_n6354_, new_n6355_, new_n6356_,
    new_n6357_, new_n6358_, new_n6359_, new_n6360_, new_n6361_, new_n6362_,
    new_n6363_, new_n6364_, new_n6365_, new_n6366_, new_n6367_, new_n6368_,
    new_n6369_, new_n6370_, new_n6371_, new_n6372_, new_n6373_, new_n6374_,
    new_n6375_, new_n6376_, new_n6377_, new_n6378_, new_n6379_, new_n6380_,
    new_n6381_, new_n6382_, new_n6383_, new_n6384_, new_n6385_, new_n6386_,
    new_n6387_, new_n6388_, new_n6389_, new_n6390_, new_n6391_, new_n6392_,
    new_n6393_, new_n6394_, new_n6395_, new_n6396_, new_n6397_, new_n6398_,
    new_n6399_, new_n6400_, new_n6401_, new_n6402_, new_n6403_, new_n6404_,
    new_n6405_, new_n6406_, new_n6407_, new_n6408_, new_n6409_, new_n6410_,
    new_n6411_, new_n6412_, new_n6413_, new_n6414_, new_n6415_, new_n6416_,
    new_n6417_, new_n6418_, new_n6419_, new_n6420_, new_n6421_, new_n6422_,
    new_n6423_, new_n6424_, new_n6425_, new_n6426_, new_n6427_, new_n6428_,
    new_n6429_, new_n6430_, new_n6431_, new_n6432_, new_n6433_, new_n6434_,
    new_n6435_, new_n6436_, new_n6437_, new_n6438_, new_n6439_, new_n6440_,
    new_n6441_, new_n6442_, new_n6443_, new_n6444_, new_n6445_, new_n6446_,
    new_n6447_, new_n6448_, new_n6449_, new_n6450_, new_n6451_, new_n6452_,
    new_n6453_, new_n6454_, new_n6455_, new_n6456_, new_n6457_, new_n6458_,
    new_n6459_, new_n6460_, new_n6461_, new_n6462_, new_n6463_, new_n6464_,
    new_n6465_, new_n6466_, new_n6467_, new_n6468_, new_n6469_, new_n6470_,
    new_n6471_, new_n6472_, new_n6473_, new_n6474_, new_n6475_, new_n6476_,
    new_n6477_, new_n6478_, new_n6479_, new_n6480_, new_n6481_, new_n6482_,
    new_n6483_, new_n6484_, new_n6485_, new_n6486_, new_n6487_, new_n6488_,
    new_n6489_, new_n6490_, new_n6491_, new_n6492_, new_n6493_, new_n6494_,
    new_n6495_, new_n6496_, new_n6497_, new_n6498_, new_n6499_, new_n6500_,
    new_n6501_, new_n6502_, new_n6503_, new_n6504_, new_n6505_, new_n6506_,
    new_n6507_, new_n6508_, new_n6509_, new_n6510_, new_n6511_, new_n6512_,
    new_n6513_, new_n6514_, new_n6515_, new_n6516_, new_n6517_, new_n6518_,
    new_n6519_, new_n6520_, new_n6522_, new_n6523_, new_n6524_, new_n6525_,
    new_n6526_, new_n6527_, new_n6528_, new_n6529_, new_n6530_, new_n6531_,
    new_n6532_, new_n6533_, new_n6534_, new_n6535_, new_n6536_, new_n6537_,
    new_n6538_, new_n6539_, new_n6540_, new_n6541_, new_n6542_, new_n6543_,
    new_n6544_, new_n6545_, new_n6546_, new_n6547_, new_n6548_, new_n6549_,
    new_n6550_, new_n6551_, new_n6552_, new_n6553_, new_n6554_, new_n6555_,
    new_n6556_, new_n6557_, new_n6558_, new_n6559_, new_n6560_, new_n6561_,
    new_n6562_, new_n6563_, new_n6564_, new_n6565_, new_n6566_, new_n6567_,
    new_n6568_, new_n6569_, new_n6570_, new_n6571_, new_n6572_, new_n6573_,
    new_n6574_, new_n6575_, new_n6576_, new_n6577_, new_n6578_, new_n6579_,
    new_n6580_, new_n6581_, new_n6582_, new_n6583_, new_n6584_, new_n6585_,
    new_n6586_, new_n6587_, new_n6588_, new_n6589_, new_n6590_, new_n6591_,
    new_n6592_, new_n6593_, new_n6594_, new_n6595_, new_n6596_, new_n6597_,
    new_n6598_, new_n6599_, new_n6600_, new_n6601_, new_n6602_, new_n6603_,
    new_n6604_, new_n6605_, new_n6606_, new_n6607_, new_n6608_, new_n6609_,
    new_n6610_, new_n6611_, new_n6612_, new_n6613_, new_n6614_, new_n6615_,
    new_n6616_, new_n6617_, new_n6618_, new_n6619_, new_n6620_, new_n6621_,
    new_n6622_, new_n6623_, new_n6624_, new_n6625_, new_n6626_, new_n6627_,
    new_n6628_, new_n6629_, new_n6630_, new_n6631_, new_n6632_, new_n6633_,
    new_n6634_, new_n6635_, new_n6636_, new_n6637_, new_n6638_, new_n6639_,
    new_n6640_, new_n6641_, new_n6642_, new_n6643_, new_n6644_, new_n6645_,
    new_n6646_, new_n6647_, new_n6648_, new_n6649_, new_n6650_, new_n6651_,
    new_n6652_, new_n6653_, new_n6654_, new_n6655_, new_n6656_, new_n6657_,
    new_n6658_, new_n6659_, new_n6660_, new_n6661_, new_n6662_, new_n6663_,
    new_n6664_, new_n6665_, new_n6666_, new_n6667_, new_n6668_, new_n6669_,
    new_n6670_, new_n6671_, new_n6672_, new_n6673_, new_n6674_, new_n6675_,
    new_n6676_, new_n6677_, new_n6678_, new_n6679_, new_n6680_, new_n6681_,
    new_n6682_, new_n6683_, new_n6684_, new_n6685_, new_n6686_, new_n6687_,
    new_n6688_, new_n6689_, new_n6690_, new_n6691_, new_n6692_, new_n6693_,
    new_n6694_, new_n6695_, new_n6696_, new_n6697_, new_n6698_, new_n6699_,
    new_n6700_, new_n6701_, new_n6702_, new_n6703_, new_n6704_, new_n6705_,
    new_n6706_, new_n6707_, new_n6708_, new_n6709_, new_n6710_, new_n6711_,
    new_n6712_, new_n6713_, new_n6714_, new_n6715_, new_n6716_, new_n6717_,
    new_n6718_, new_n6719_, new_n6720_, new_n6721_, new_n6722_, new_n6723_,
    new_n6724_, new_n6725_, new_n6726_, new_n6727_, new_n6728_, new_n6729_,
    new_n6730_, new_n6731_, new_n6732_, new_n6733_, new_n6734_, new_n6735_,
    new_n6736_, new_n6737_, new_n6738_, new_n6739_, new_n6740_, new_n6741_,
    new_n6742_, new_n6743_, new_n6744_, new_n6745_, new_n6746_, new_n6747_,
    new_n6748_, new_n6749_, new_n6750_, new_n6751_, new_n6752_, new_n6753_,
    new_n6755_, new_n6756_, new_n6757_, new_n6759_, new_n6760_, new_n6761_,
    new_n6762_, new_n6763_, new_n6764_, new_n6765_, new_n6766_, new_n6767_,
    new_n6768_, new_n6769_, new_n6770_, new_n6771_, new_n6772_, new_n6773_,
    new_n6774_, new_n6775_, new_n6776_, new_n6777_, new_n6778_, new_n6779_,
    new_n6780_, new_n6781_, new_n6782_, new_n6783_, new_n6784_, new_n6785_,
    new_n6786_, new_n6787_, new_n6788_, new_n6789_, new_n6790_, new_n6791_,
    new_n6792_, new_n6793_, new_n6794_, new_n6795_, new_n6796_, new_n6797_,
    new_n6798_, new_n6799_, new_n6800_, new_n6801_, new_n6802_, new_n6803_,
    new_n6805_, new_n6806_, new_n6807_, new_n6808_, new_n6809_, new_n6810_,
    new_n6811_, new_n6812_, new_n6813_, new_n6814_, new_n6816_, new_n6817_,
    new_n6818_, new_n6819_, new_n6820_, new_n6821_, new_n6822_, new_n6823_,
    new_n6824_, new_n6825_, new_n6826_, new_n6827_, new_n6828_, new_n6829_,
    new_n6830_, new_n6831_, new_n6832_, new_n6833_, new_n6834_, new_n6835_,
    new_n6836_, new_n6837_, new_n6838_, new_n6839_, new_n6840_, new_n6841_,
    new_n6842_, new_n6843_, new_n6844_, new_n6845_, new_n6846_, new_n6847_,
    new_n6848_, new_n6849_, new_n6850_, new_n6851_, new_n6852_, new_n6853_,
    new_n6854_, new_n6855_, new_n6856_, new_n6857_, new_n6858_, new_n6859_,
    new_n6860_, new_n6861_, new_n6862_, new_n6863_, new_n6864_, new_n6865_,
    new_n6866_, new_n6867_, new_n6868_, new_n6869_, new_n6870_, new_n6871_,
    new_n6872_, new_n6873_, new_n6874_, new_n6875_, new_n6876_, new_n6877_,
    new_n6878_, new_n6879_, new_n6880_, new_n6881_, new_n6882_, new_n6883_,
    new_n6884_, new_n6885_, new_n6886_, new_n6887_, new_n6888_, new_n6889_,
    new_n6890_, new_n6891_, new_n6892_, new_n6893_, new_n6894_, new_n6895_,
    new_n6896_, new_n6897_, new_n6898_, new_n6899_, new_n6900_, new_n6901_,
    new_n6902_, new_n6903_, new_n6904_, new_n6905_, new_n6906_, new_n6907_,
    new_n6908_, new_n6909_, new_n6910_, new_n6911_, new_n6912_, new_n6913_,
    new_n6914_, new_n6915_, new_n6916_, new_n6917_, new_n6918_, new_n6919_,
    new_n6920_, new_n6921_, new_n6922_, new_n6923_, new_n6924_, new_n6925_,
    new_n6926_, new_n6927_, new_n6928_, new_n6929_, new_n6930_, new_n6931_,
    new_n6932_, new_n6933_, new_n6934_, new_n6935_, new_n6936_, new_n6937_,
    new_n6938_, new_n6939_, new_n6940_, new_n6941_, new_n6942_, new_n6943_,
    new_n6944_, new_n6945_, new_n6946_, new_n6947_, new_n6948_, new_n6949_,
    new_n6950_, new_n6951_, new_n6952_, new_n6953_, new_n6954_, new_n6955_,
    new_n6956_, new_n6957_, new_n6958_, new_n6959_, new_n6960_, new_n6961_,
    new_n6962_, new_n6963_, new_n6964_, new_n6965_, new_n6966_, new_n6967_,
    new_n6968_, new_n6969_, new_n6970_, new_n6971_, new_n6972_, new_n6973_,
    new_n6974_, new_n6975_, new_n6976_, new_n6977_, new_n6978_, new_n6979_,
    new_n6980_, new_n6981_, new_n6982_, new_n6983_, new_n6984_, new_n6985_,
    new_n6986_, new_n6987_, new_n6988_, new_n6989_, new_n6990_, new_n6991_,
    new_n6992_, new_n6993_, new_n6994_, new_n6995_, new_n6996_, new_n6997_,
    new_n6998_, new_n6999_, new_n7000_, new_n7001_, new_n7002_, new_n7003_,
    new_n7004_, new_n7005_, new_n7006_, new_n7007_, new_n7008_, new_n7009_,
    new_n7010_, new_n7011_, new_n7012_, new_n7013_, new_n7014_, new_n7015_,
    new_n7016_, new_n7017_, new_n7018_, new_n7019_, new_n7020_, new_n7021_,
    new_n7022_, new_n7023_, new_n7024_, new_n7025_, new_n7026_, new_n7027_,
    new_n7028_, new_n7029_, new_n7030_, new_n7031_, new_n7032_, new_n7033_,
    new_n7034_, new_n7035_, new_n7036_, new_n7037_, new_n7038_, new_n7039_,
    new_n7040_, new_n7041_, new_n7042_, new_n7043_, new_n7044_, new_n7045_,
    new_n7046_, new_n7047_, new_n7048_, new_n7049_, new_n7050_, new_n7051_,
    new_n7052_, new_n7053_, new_n7054_, new_n7055_, new_n7056_, new_n7057_,
    new_n7058_, new_n7059_, new_n7060_, new_n7061_, new_n7062_, new_n7063_,
    new_n7064_, new_n7065_, new_n7066_, new_n7067_, new_n7068_, new_n7069_,
    new_n7070_, new_n7071_, new_n7072_, new_n7073_, new_n7074_, new_n7075_,
    new_n7076_, new_n7077_, new_n7078_, new_n7079_, new_n7080_, new_n7081_,
    new_n7082_, new_n7083_, new_n7084_, new_n7085_, new_n7086_, new_n7087_,
    new_n7088_, new_n7089_, new_n7090_, new_n7091_, new_n7092_, new_n7093_,
    new_n7094_, new_n7095_, new_n7096_, new_n7097_, new_n7098_, new_n7099_,
    new_n7100_, new_n7101_, new_n7102_, new_n7103_, new_n7104_, new_n7105_,
    new_n7106_, new_n7107_, new_n7108_, new_n7109_, new_n7110_, new_n7111_,
    new_n7112_, new_n7113_, new_n7114_, new_n7115_, new_n7116_, new_n7117_,
    new_n7118_, new_n7119_, new_n7120_, new_n7121_, new_n7122_, new_n7123_,
    new_n7124_, new_n7125_, new_n7126_, new_n7127_, new_n7128_, new_n7129_,
    new_n7130_, new_n7131_, new_n7132_, new_n7133_, new_n7134_, new_n7135_,
    new_n7136_, new_n7137_, new_n7138_, new_n7139_, new_n7140_, new_n7141_,
    new_n7142_, new_n7143_, new_n7144_, new_n7145_, new_n7146_, new_n7147_,
    new_n7148_, new_n7149_, new_n7150_, new_n7151_, new_n7152_, new_n7153_,
    new_n7154_, new_n7155_, new_n7156_, new_n7157_, new_n7158_, new_n7159_,
    new_n7160_, new_n7161_, new_n7162_, new_n7163_, new_n7164_, new_n7165_,
    new_n7166_, new_n7167_, new_n7168_, new_n7169_, new_n7170_, new_n7171_,
    new_n7172_, new_n7173_, new_n7174_, new_n7175_, new_n7176_, new_n7177_,
    new_n7178_, new_n7179_, new_n7180_, new_n7181_, new_n7182_, new_n7183_,
    new_n7184_, new_n7185_, new_n7186_, new_n7187_, new_n7188_, new_n7189_,
    new_n7190_, new_n7191_, new_n7192_, new_n7193_, new_n7194_, new_n7195_,
    new_n7196_, new_n7197_, new_n7198_, new_n7199_, new_n7200_, new_n7201_,
    new_n7202_, new_n7203_, new_n7204_, new_n7205_, new_n7206_, new_n7207_,
    new_n7208_, new_n7209_, new_n7210_, new_n7211_, new_n7212_, new_n7213_,
    new_n7214_, new_n7215_, new_n7216_, new_n7217_, new_n7218_, new_n7219_,
    new_n7220_, new_n7221_, new_n7222_, new_n7223_, new_n7224_, new_n7225_,
    new_n7226_, new_n7227_, new_n7228_, new_n7229_, new_n7230_, new_n7231_,
    new_n7232_, new_n7233_, new_n7234_, new_n7235_, new_n7236_, new_n7237_,
    new_n7238_, new_n7239_, new_n7240_, new_n7241_, new_n7242_, new_n7243_,
    new_n7244_, new_n7245_, new_n7246_, new_n7247_, new_n7248_, new_n7249_,
    new_n7250_, new_n7251_, new_n7252_, new_n7253_, new_n7254_, new_n7255_,
    new_n7256_, new_n7257_, new_n7258_, new_n7259_, new_n7260_, new_n7261_,
    new_n7262_, new_n7263_, new_n7264_, new_n7265_, new_n7266_, new_n7267_,
    new_n7268_, new_n7269_, new_n7270_, new_n7271_, new_n7272_, new_n7273_,
    new_n7274_, new_n7275_, new_n7276_, new_n7277_, new_n7278_, new_n7279_,
    new_n7280_, new_n7281_, new_n7282_, new_n7283_, new_n7284_, new_n7285_,
    new_n7286_, new_n7287_, new_n7288_, new_n7289_, new_n7290_, new_n7291_,
    new_n7292_, new_n7293_, new_n7294_, new_n7295_, new_n7296_, new_n7297_,
    new_n7298_, new_n7299_, new_n7300_, new_n7301_, new_n7302_, new_n7303_,
    new_n7304_, new_n7305_, new_n7306_, new_n7307_, new_n7308_, new_n7309_,
    new_n7310_, new_n7311_, new_n7312_, new_n7313_, new_n7314_, new_n7315_,
    new_n7316_, new_n7317_, new_n7318_, new_n7319_, new_n7320_, new_n7321_,
    new_n7322_, new_n7323_, new_n7324_, new_n7325_, new_n7326_, new_n7327_,
    new_n7328_, new_n7329_, new_n7330_, new_n7331_, new_n7332_, new_n7333_,
    new_n7334_, new_n7335_, new_n7336_, new_n7337_, new_n7338_, new_n7339_,
    new_n7341_, new_n7342_, new_n7344_, new_n7345_, new_n7346_, new_n7347_,
    new_n7348_, new_n7349_, new_n7350_, new_n7351_, new_n7352_, new_n7353_,
    new_n7354_, new_n7355_, new_n7356_, new_n7357_, new_n7358_, new_n7359_,
    new_n7360_, new_n7361_, new_n7362_, new_n7363_, new_n7364_, new_n7365_,
    new_n7366_, new_n7367_, new_n7368_, new_n7369_, new_n7370_, new_n7371_,
    new_n7372_, new_n7373_, new_n7374_, new_n7375_, new_n7376_, new_n7377_,
    new_n7378_, new_n7379_, new_n7380_, new_n7381_, new_n7382_, new_n7383_,
    new_n7384_, new_n7385_, new_n7386_, new_n7387_, new_n7388_, new_n7389_,
    new_n7390_, new_n7391_, new_n7392_, new_n7393_, new_n7394_, new_n7395_,
    new_n7396_, new_n7397_, new_n7398_, new_n7399_, new_n7400_, new_n7401_,
    new_n7402_, new_n7403_, new_n7404_, new_n7405_, new_n7406_, new_n7407_,
    new_n7408_, new_n7409_, new_n7410_, new_n7411_, new_n7412_, new_n7413_,
    new_n7414_, new_n7415_, new_n7416_, new_n7417_, new_n7418_, new_n7419_,
    new_n7420_, new_n7421_, new_n7422_, new_n7423_, new_n7424_, new_n7425_,
    new_n7426_, new_n7427_, new_n7428_, new_n7429_, new_n7430_, new_n7431_,
    new_n7432_, new_n7433_, new_n7434_, new_n7435_, new_n7436_, new_n7437_,
    new_n7438_, new_n7439_, new_n7440_, new_n7441_, new_n7442_, new_n7443_,
    new_n7444_, new_n7445_, new_n7446_, new_n7447_, new_n7448_, new_n7449_,
    new_n7450_, new_n7451_, new_n7452_, new_n7453_, new_n7454_, new_n7455_,
    new_n7456_, new_n7457_, new_n7458_, new_n7459_, new_n7460_, new_n7461_,
    new_n7462_, new_n7463_, new_n7464_, new_n7465_, new_n7466_, new_n7467_,
    new_n7468_, new_n7469_, new_n7470_, new_n7471_, new_n7472_, new_n7473_,
    new_n7474_, new_n7475_, new_n7476_, new_n7477_, new_n7478_, new_n7479_,
    new_n7480_, new_n7481_, new_n7482_, new_n7483_, new_n7484_, new_n7485_,
    new_n7486_, new_n7487_, new_n7488_, new_n7489_, new_n7490_, new_n7491_,
    new_n7492_, new_n7493_, new_n7494_, new_n7495_, new_n7496_, new_n7497_,
    new_n7498_, new_n7499_, new_n7500_, new_n7501_, new_n7502_, new_n7503_,
    new_n7504_, new_n7505_, new_n7506_, new_n7507_, new_n7508_, new_n7509_,
    new_n7510_, new_n7511_, new_n7512_, new_n7513_, new_n7514_, new_n7515_,
    new_n7516_, new_n7517_, new_n7518_, new_n7519_, new_n7520_, new_n7521_,
    new_n7522_, new_n7523_, new_n7524_, new_n7525_, new_n7526_, new_n7527_,
    new_n7528_, new_n7529_, new_n7530_, new_n7531_, new_n7532_, new_n7533_,
    new_n7534_, new_n7535_, new_n7536_, new_n7537_, new_n7538_, new_n7539_,
    new_n7540_, new_n7541_, new_n7542_, new_n7543_, new_n7544_, new_n7545_,
    new_n7546_, new_n7547_, new_n7548_, new_n7549_, new_n7550_, new_n7551_,
    new_n7552_, new_n7553_, new_n7554_, new_n7555_, new_n7556_, new_n7557_,
    new_n7558_, new_n7559_, new_n7560_, new_n7561_, new_n7562_, new_n7563_,
    new_n7564_, new_n7565_, new_n7566_, new_n7567_, new_n7568_, new_n7569_,
    new_n7570_, new_n7571_, new_n7572_, new_n7573_, new_n7574_, new_n7575_,
    new_n7576_, new_n7577_, new_n7578_, new_n7579_, new_n7580_, new_n7581_,
    new_n7582_, new_n7583_, new_n7584_, new_n7585_, new_n7586_, new_n7587_,
    new_n7588_, new_n7589_, new_n7590_, new_n7591_, new_n7592_, new_n7593_,
    new_n7594_, new_n7595_, new_n7596_, new_n7597_, new_n7598_, new_n7599_,
    new_n7600_, new_n7601_, new_n7602_, new_n7604_, new_n7605_, new_n7606_,
    new_n7607_, new_n7608_, new_n7609_, new_n7610_, new_n7611_, new_n7612_,
    new_n7613_, new_n7614_, new_n7615_, new_n7616_, new_n7617_, new_n7618_,
    new_n7619_, new_n7620_, new_n7621_, new_n7622_, new_n7623_, new_n7624_,
    new_n7625_, new_n7626_, new_n7627_, new_n7628_, new_n7629_, new_n7630_,
    new_n7631_, new_n7632_, new_n7633_, new_n7634_, new_n7635_, new_n7636_,
    new_n7637_, new_n7638_, new_n7639_, new_n7640_, new_n7641_, new_n7642_,
    new_n7643_, new_n7644_, new_n7645_, new_n7646_, new_n7647_, new_n7648_,
    new_n7649_, new_n7650_, new_n7651_, new_n7652_, new_n7653_, new_n7654_,
    new_n7656_, new_n7657_, new_n7658_, new_n7659_, new_n7660_, new_n7661_,
    new_n7662_, new_n7663_, new_n7664_, new_n7665_, new_n7666_, new_n7667_,
    new_n7668_, new_n7669_, new_n7670_, new_n7672_, new_n7673_, new_n7674_,
    new_n7675_, new_n7676_, new_n7677_, new_n7678_, new_n7679_, new_n7680_,
    new_n7681_, new_n7682_, new_n7683_, new_n7684_, new_n7685_, new_n7686_,
    new_n7687_, new_n7689_, new_n7690_, new_n7691_, new_n7692_, new_n7693_,
    new_n7694_, new_n7695_, new_n7696_, new_n7697_, new_n7698_, new_n7699_,
    new_n7700_, new_n7701_, new_n7702_, new_n7703_, new_n7704_, new_n7705_,
    new_n7706_, new_n7707_, new_n7708_, new_n7709_, new_n7710_, new_n7711_,
    new_n7712_, new_n7713_, new_n7714_, new_n7715_, new_n7716_, new_n7717_,
    new_n7718_, new_n7719_, new_n7720_, new_n7721_, new_n7722_, new_n7723_,
    new_n7724_, new_n7725_, new_n7726_, new_n7727_, new_n7728_, new_n7729_,
    new_n7730_, new_n7731_, new_n7732_, new_n7733_, new_n7734_, new_n7735_,
    new_n7736_, new_n7737_, new_n7738_, new_n7739_, new_n7740_, new_n7741_,
    new_n7742_, new_n7743_, new_n7744_, new_n7745_, new_n7746_, new_n7747_,
    new_n7749_, new_n7750_, new_n7751_, new_n7752_, new_n7753_, new_n7754_,
    new_n7755_, new_n7756_, new_n7757_, new_n7759_, new_n7760_, new_n7761_,
    new_n7762_, new_n7763_, new_n7764_, new_n7765_, new_n7766_, new_n7767_,
    new_n7768_, new_n7769_, new_n7770_, new_n7771_, new_n7772_, new_n7773_,
    new_n7774_, new_n7775_, new_n7776_, new_n7777_, new_n7778_, new_n7779_,
    new_n7780_, new_n7781_, new_n7782_, new_n7783_, new_n7784_, new_n7785_,
    new_n7786_, new_n7787_, new_n7788_, new_n7789_, new_n7790_, new_n7791_,
    new_n7792_, new_n7793_, new_n7794_, new_n7795_, new_n7796_, new_n7797_,
    new_n7798_, new_n7799_, new_n7800_, new_n7801_, new_n7802_, new_n7803_,
    new_n7804_, new_n7805_, new_n7806_, new_n7807_, new_n7808_, new_n7809_,
    new_n7810_, new_n7811_, new_n7812_, new_n7813_, new_n7814_, new_n7815_,
    new_n7816_, new_n7817_, new_n7818_, new_n7819_, new_n7820_, new_n7821_,
    new_n7822_, new_n7823_, new_n7824_, new_n7825_, new_n7826_, new_n7827_,
    new_n7828_, new_n7829_, new_n7830_, new_n7831_, new_n7832_, new_n7833_,
    new_n7834_, new_n7835_, new_n7836_, new_n7837_, new_n7838_, new_n7839_,
    new_n7840_, new_n7841_, new_n7842_, new_n7843_, new_n7844_, new_n7845_,
    new_n7846_, new_n7847_, new_n7848_, new_n7849_, new_n7850_, new_n7851_,
    new_n7852_, new_n7853_, new_n7854_, new_n7855_, new_n7856_, new_n7857_,
    new_n7858_, new_n7859_, new_n7860_, new_n7861_, new_n7862_, new_n7863_,
    new_n7864_, new_n7865_, new_n7866_, new_n7867_, new_n7868_, new_n7869_,
    new_n7870_, new_n7871_, new_n7872_, new_n7873_, new_n7874_, new_n7875_,
    new_n7876_, new_n7877_, new_n7878_, new_n7879_, new_n7880_, new_n7881_,
    new_n7882_, new_n7883_, new_n7884_, new_n7885_, new_n7886_, new_n7887_,
    new_n7888_, new_n7889_, new_n7890_, new_n7891_, new_n7892_, new_n7893_,
    new_n7894_, new_n7896_, new_n7897_, new_n7898_, new_n7899_, new_n7900_,
    new_n7901_, new_n7902_, new_n7903_, new_n7904_, new_n7905_, new_n7906_,
    new_n7907_, new_n7908_, new_n7909_, new_n7910_, new_n7911_, new_n7912_,
    new_n7913_, new_n7914_, new_n7915_, new_n7916_, new_n7917_, new_n7918_,
    new_n7919_, new_n7920_, new_n7921_, new_n7922_, new_n7923_, new_n7924_,
    new_n7925_, new_n7926_, new_n7927_, new_n7928_, new_n7929_, new_n7930_,
    new_n7931_, new_n7932_, new_n7933_, new_n7934_, new_n7935_, new_n7936_,
    new_n7937_, new_n7938_, new_n7939_, new_n7940_, new_n7941_, new_n7942_,
    new_n7943_, new_n7944_, new_n7945_, new_n7946_, new_n7947_, new_n7948_,
    new_n7949_, new_n7950_, new_n7951_, new_n7952_, new_n7953_, new_n7954_,
    new_n7955_, new_n7956_, new_n7957_, new_n7958_, new_n7959_, new_n7960_,
    new_n7961_, new_n7962_, new_n7963_, new_n7964_, new_n7965_, new_n7966_,
    new_n7967_, new_n7968_, new_n7969_, new_n7970_, new_n7971_, new_n7972_,
    new_n7973_, new_n7974_, new_n7975_, new_n7976_, new_n7977_, new_n7978_,
    new_n7979_, new_n7980_, new_n7981_, new_n7982_, new_n7983_, new_n7984_,
    new_n7985_, new_n7986_, new_n7987_, new_n7988_, new_n7989_, new_n7990_,
    new_n7991_, new_n7992_, new_n7993_, new_n7994_, new_n7995_, new_n7996_,
    new_n7997_, new_n7998_, new_n7999_, new_n8000_, new_n8001_, new_n8002_,
    new_n8003_, new_n8004_, new_n8005_, new_n8006_, new_n8007_, new_n8008_,
    new_n8009_, new_n8010_, new_n8011_, new_n8012_, new_n8013_, new_n8014_,
    new_n8015_, new_n8016_, new_n8017_, new_n8018_, new_n8019_, new_n8020_,
    new_n8021_, new_n8022_, new_n8023_, new_n8024_, new_n8025_, new_n8026_,
    new_n8027_, new_n8028_, new_n8029_, new_n8030_, new_n8031_, new_n8032_,
    new_n8033_, new_n8034_, new_n8035_, new_n8036_, new_n8037_, new_n8038_,
    new_n8039_, new_n8040_, new_n8041_, new_n8042_, new_n8043_, new_n8044_,
    new_n8045_, new_n8046_, new_n8047_, new_n8048_, new_n8049_, new_n8050_,
    new_n8051_, new_n8052_, new_n8053_, new_n8054_, new_n8055_, new_n8056_,
    new_n8057_, new_n8058_, new_n8059_, new_n8060_, new_n8061_, new_n8062_,
    new_n8063_, new_n8064_, new_n8065_, new_n8066_, new_n8067_, new_n8068_,
    new_n8069_, new_n8070_, new_n8071_, new_n8072_, new_n8074_, new_n8075_,
    new_n8076_, new_n8077_, new_n8078_, new_n8079_, new_n8080_, new_n8081_,
    new_n8082_, new_n8083_, new_n8084_, new_n8085_, new_n8086_, new_n8087_,
    new_n8088_, new_n8089_, new_n8090_, new_n8091_, new_n8092_, new_n8093_,
    new_n8094_, new_n8095_, new_n8096_, new_n8097_, new_n8098_, new_n8099_,
    new_n8100_, new_n8101_, new_n8102_, new_n8103_, new_n8104_, new_n8105_,
    new_n8106_, new_n8107_, new_n8108_, new_n8109_, new_n8110_, new_n8111_,
    new_n8112_, new_n8113_, new_n8114_, new_n8115_, new_n8116_, new_n8117_,
    new_n8118_, new_n8119_, new_n8120_, new_n8121_, new_n8122_, new_n8123_,
    new_n8124_, new_n8125_, new_n8126_, new_n8127_, new_n8128_, new_n8129_,
    new_n8130_, new_n8131_, new_n8132_, new_n8133_, new_n8134_, new_n8135_,
    new_n8136_, new_n8137_, new_n8138_, new_n8139_, new_n8140_, new_n8141_,
    new_n8142_, new_n8143_, new_n8144_, new_n8145_, new_n8146_, new_n8147_,
    new_n8148_, new_n8149_, new_n8150_, new_n8151_, new_n8152_, new_n8153_,
    new_n8154_, new_n8155_, new_n8156_, new_n8157_, new_n8158_, new_n8159_,
    new_n8160_, new_n8161_, new_n8162_, new_n8163_, new_n8164_, new_n8165_,
    new_n8166_, new_n8167_, new_n8168_, new_n8169_, new_n8170_, new_n8171_,
    new_n8172_, new_n8173_, new_n8174_, new_n8175_, new_n8176_, new_n8177_,
    new_n8178_, new_n8179_, new_n8180_, new_n8181_, new_n8182_, new_n8183_,
    new_n8184_, new_n8185_, new_n8186_, new_n8187_, new_n8188_, new_n8189_,
    new_n8190_, new_n8192_, new_n8193_, new_n8194_, new_n8195_, new_n8196_,
    new_n8197_, new_n8198_, new_n8199_, new_n8200_, new_n8201_, new_n8202_,
    new_n8203_, new_n8204_, new_n8205_, new_n8206_, new_n8207_, new_n8208_,
    new_n8209_, new_n8210_, new_n8211_, new_n8212_, new_n8213_, new_n8214_,
    new_n8215_, new_n8216_, new_n8217_, new_n8218_, new_n8219_, new_n8220_,
    new_n8221_, new_n8222_, new_n8223_, new_n8224_, new_n8225_, new_n8226_,
    new_n8227_, new_n8228_, new_n8229_, new_n8230_, new_n8231_, new_n8232_,
    new_n8233_, new_n8234_, new_n8235_, new_n8236_, new_n8237_, new_n8238_,
    new_n8239_, new_n8240_, new_n8241_, new_n8242_, new_n8244_, new_n8245_,
    new_n8247_, new_n8248_, new_n8249_, new_n8250_, new_n8251_, new_n8252_,
    new_n8253_, new_n8254_, new_n8255_, new_n8256_, new_n8257_, new_n8259_,
    new_n8260_, new_n8261_, new_n8262_, new_n8263_, new_n8264_, new_n8265_,
    new_n8266_, new_n8267_, new_n8268_, new_n8269_, new_n8270_, new_n8271_,
    new_n8272_, new_n8273_, new_n8274_, new_n8275_, new_n8276_, new_n8277_,
    new_n8278_, new_n8279_, new_n8280_, new_n8281_, new_n8282_, new_n8283_,
    new_n8284_, new_n8285_, new_n8286_, new_n8287_, new_n8288_, new_n8290_,
    new_n8292_, new_n8293_, new_n8294_, new_n8295_, new_n8296_, new_n8297_,
    new_n8298_, new_n8299_, new_n8300_, new_n8301_, new_n8302_, new_n8303_,
    new_n8304_, new_n8306_, new_n8307_, new_n8308_, new_n8309_, new_n8310_,
    new_n8311_, new_n8312_, new_n8313_, new_n8314_, new_n8315_, new_n8316_,
    new_n8317_, new_n8318_, new_n8319_, new_n8320_, new_n8321_, new_n8323_,
    new_n8324_, new_n8325_, new_n8326_, new_n8328_, new_n8329_, new_n8330_,
    new_n8331_, new_n8332_, new_n8333_, new_n8334_, new_n8335_, new_n8336_,
    new_n8337_, new_n8338_, new_n8339_, new_n8340_, new_n8341_, new_n8342_,
    new_n8343_, new_n8344_, new_n8345_, new_n8346_, new_n8347_, new_n8348_,
    new_n8349_, new_n8350_, new_n8351_, new_n8352_, new_n8353_, new_n8354_,
    new_n8355_, new_n8356_, new_n8357_, new_n8358_, new_n8359_, new_n8360_,
    new_n8361_, new_n8362_, new_n8363_, new_n8364_, new_n8365_, new_n8366_,
    new_n8367_, new_n8368_, new_n8369_, new_n8370_, new_n8371_, new_n8372_,
    new_n8373_, new_n8374_, new_n8375_, new_n8376_, new_n8377_, new_n8378_,
    new_n8379_, new_n8380_, new_n8381_, new_n8382_, new_n8383_, new_n8384_,
    new_n8385_, new_n8386_, new_n8387_, new_n8388_, new_n8389_, new_n8390_,
    new_n8391_, new_n8392_, new_n8393_, new_n8394_, new_n8395_, new_n8396_,
    new_n8397_, new_n8398_, new_n8399_, new_n8400_, new_n8401_, new_n8402_,
    new_n8403_, new_n8404_, new_n8405_, new_n8406_, new_n8407_, new_n8408_,
    new_n8409_, new_n8410_, new_n8411_, new_n8412_, new_n8413_, new_n8414_,
    new_n8415_, new_n8416_, new_n8417_, new_n8418_, new_n8419_, new_n8420_,
    new_n8421_, new_n8422_, new_n8423_, new_n8424_, new_n8425_, new_n8426_,
    new_n8427_, new_n8429_, new_n8430_, new_n8431_, new_n8432_, new_n8433_,
    new_n8435_, new_n8436_, new_n8437_, new_n8438_, new_n8439_, new_n8440_,
    new_n8441_, new_n8442_, new_n8443_, new_n8444_, new_n8445_, new_n8446_,
    new_n8447_, new_n8449_, new_n8450_, new_n8451_, new_n8452_, new_n8453_,
    new_n8454_, new_n8455_, new_n8456_, new_n8458_, new_n8459_, new_n8460_,
    new_n8461_, new_n8463_, new_n8464_, new_n8465_, new_n8466_, new_n8467_,
    new_n8468_, new_n8470_, new_n8472_, new_n8473_, new_n8474_, new_n8476_,
    new_n8477_, new_n8478_, new_n8479_, new_n8481_, new_n8482_, new_n8484_,
    new_n8485_, new_n8486_, new_n8488_, new_n8489_, new_n8490_, new_n8491_,
    new_n8493_, new_n8494_, new_n8495_, new_n8496_, new_n8497_, new_n8499_,
    new_n8500_, new_n8502_, new_n8503_, new_n8504_, new_n8505_, new_n8506_,
    new_n8507_, new_n8508_, new_n8509_, new_n8510_, new_n8512_, new_n8513_,
    new_n8515_, new_n8516_, new_n8517_, new_n8518_, new_n8519_, new_n8520_,
    new_n8522_, new_n8523_, new_n8524_, new_n8525_, new_n8526_, new_n8527_,
    new_n8529_, new_n8530_, new_n8531_, new_n8532_, new_n8533_, new_n8534_,
    new_n8535_, new_n8536_, new_n8537_, new_n8538_, new_n8539_, new_n8541_,
    new_n8542_, new_n8543_, new_n8544_, new_n8545_, new_n8546_, new_n8547_,
    new_n8548_, new_n8549_, new_n8550_, new_n8551_, new_n8552_, new_n8553_,
    new_n8554_, new_n8555_, new_n8557_, new_n8558_, new_n8559_, new_n8560_,
    new_n8561_, new_n8562_, new_n8563_, new_n8564_, new_n8565_, new_n8566_,
    new_n8567_, new_n8568_, new_n8569_, new_n8571_, new_n8572_, new_n8573_,
    new_n8574_, new_n8575_, new_n8576_, new_n8577_, new_n8578_, new_n8579_,
    new_n8581_, new_n8582_, new_n8583_, new_n8584_, new_n8585_, new_n8586_,
    new_n8587_, new_n8588_, new_n8590_, new_n8591_, new_n8592_, new_n8593_,
    new_n8595_, new_n8596_, new_n8597_, new_n8598_, new_n8599_, new_n8600_,
    new_n8601_, new_n8602_, new_n8603_, new_n8604_, new_n8605_, new_n8606_,
    new_n8607_, new_n8608_, new_n8609_, new_n8610_, new_n8611_, new_n8612_,
    new_n8613_, new_n8614_, new_n8615_, new_n8616_, new_n8617_, new_n8618_,
    new_n8619_, new_n8620_, new_n8621_, new_n8622_, new_n8623_, new_n8624_,
    new_n8625_, new_n8626_, new_n8627_, new_n8628_, new_n8629_, new_n8630_,
    new_n8631_, new_n8632_, new_n8633_, new_n8634_, new_n8635_, new_n8636_,
    new_n8637_, new_n8638_, new_n8639_, new_n8640_, new_n8641_, new_n8642_,
    new_n8643_, new_n8644_, new_n8645_, new_n8646_, new_n8647_, new_n8648_,
    new_n8649_, new_n8650_, new_n8651_, new_n8652_, new_n8653_, new_n8654_,
    new_n8655_, new_n8656_, new_n8657_, new_n8658_, new_n8659_, new_n8660_,
    new_n8661_, new_n8662_, new_n8663_, new_n8664_, new_n8665_, new_n8666_,
    new_n8667_, new_n8668_, new_n8669_, new_n8670_, new_n8671_, new_n8672_,
    new_n8673_, new_n8674_, new_n8675_, new_n8676_, new_n8677_, new_n8678_,
    new_n8679_, new_n8680_, new_n8681_, new_n8682_, new_n8683_, new_n8684_,
    new_n8685_, new_n8686_, new_n8687_, new_n8688_, new_n8689_, new_n8690_,
    new_n8691_, new_n8692_, new_n8693_, new_n8694_, new_n8695_, new_n8697_,
    new_n8698_, new_n8699_, new_n8700_, new_n8701_, new_n8702_, new_n8705_,
    new_n8706_, new_n8707_, new_n8708_, new_n8709_, new_n8710_, new_n8711_,
    new_n8712_, new_n8713_, new_n8714_, new_n8715_, new_n8716_, new_n8717_,
    new_n8718_, new_n8719_, new_n8720_, new_n8721_, new_n8722_, new_n8723_,
    new_n8724_, new_n8725_, new_n8726_, new_n8727_, new_n8728_, new_n8729_,
    new_n8730_, new_n8731_, new_n8732_, new_n8733_, new_n8734_, new_n8735_,
    new_n8736_, new_n8737_, new_n8738_, new_n8739_, new_n8740_, new_n8741_,
    new_n8742_, new_n8743_, new_n8744_, new_n8745_, new_n8746_, new_n8747_,
    new_n8748_, new_n8749_, new_n8750_, new_n8751_, new_n8752_, new_n8753_,
    new_n8754_, new_n8755_, new_n8756_, new_n8757_, new_n8758_, new_n8759_,
    new_n8760_, new_n8761_, new_n8762_, new_n8763_, new_n8764_, new_n8765_,
    new_n8766_, new_n8767_, new_n8768_, new_n8769_, new_n8770_, new_n8771_,
    new_n8772_, new_n8773_, new_n8774_, new_n8775_, new_n8776_, new_n8777_,
    new_n8778_, new_n8779_, new_n8780_, new_n8781_, new_n8782_, new_n8783_,
    new_n8784_, new_n8785_, new_n8786_, new_n8787_, new_n8788_, new_n8789_,
    new_n8790_, new_n8791_, new_n8792_, new_n8793_, new_n8794_, new_n8795_,
    new_n8796_, new_n8797_, new_n8798_, new_n8799_, new_n8800_, new_n8801_,
    new_n8802_, new_n8803_, new_n8804_, new_n8805_, new_n8806_, new_n8807_,
    new_n8808_, new_n8809_, new_n8810_, new_n8811_, new_n8812_, new_n8813_,
    new_n8814_, new_n8815_, new_n8816_, new_n8817_, new_n8818_, new_n8819_,
    new_n8820_, new_n8821_, new_n8822_, new_n8823_, new_n8824_, new_n8825_,
    new_n8826_, new_n8827_, new_n8828_, new_n8829_, new_n8830_, new_n8831_,
    new_n8832_, new_n8833_, new_n8834_, new_n8835_, new_n8836_, new_n8837_,
    new_n8838_, new_n8839_, new_n8840_, new_n8841_, new_n8842_, new_n8843_,
    new_n8844_, new_n8845_, new_n8846_, new_n8847_, new_n8848_, new_n8849_,
    new_n8850_, new_n8851_, new_n8852_, new_n8853_, new_n8854_, new_n8855_,
    new_n8856_, new_n8857_, new_n8858_, new_n8859_, new_n8860_, new_n8861_,
    new_n8862_, new_n8863_, new_n8864_, new_n8865_, new_n8866_, new_n8867_,
    new_n8868_, new_n8869_, new_n8870_, new_n8871_, new_n8872_, new_n8873_,
    new_n8874_, new_n8875_, new_n8876_, new_n8877_, new_n8878_, new_n8879_,
    new_n8880_, new_n8881_, new_n8882_, new_n8883_, new_n8884_, new_n8885_,
    new_n8886_, new_n8887_, new_n8888_, new_n8889_, new_n8890_, new_n8891_,
    new_n8892_, new_n8893_, new_n8894_, new_n8895_, new_n8896_, new_n8897_,
    new_n8898_, new_n8899_, new_n8900_, new_n8901_, new_n8902_, new_n8903_,
    new_n8904_, new_n8905_, new_n8906_, new_n8907_, new_n8908_, new_n8909_,
    new_n8910_, new_n8911_, new_n8912_, new_n8913_, new_n8914_, new_n8915_,
    new_n8916_, new_n8917_, new_n8918_, new_n8919_, new_n8920_, new_n8921_,
    new_n8922_, new_n8923_, new_n8924_, new_n8925_, new_n8926_, new_n8927_,
    new_n8928_, new_n8929_, new_n8930_, new_n8931_, new_n8932_, new_n8933_,
    new_n8934_, new_n8935_, new_n8936_, new_n8937_, new_n8938_, new_n8939_,
    new_n8940_, new_n8941_, new_n8942_, new_n8943_, new_n8944_, new_n8945_,
    new_n8946_, new_n8947_, new_n8948_, new_n8949_, new_n8950_, new_n8951_,
    new_n8952_, new_n8953_, new_n8954_, new_n8955_, new_n8956_, new_n8957_,
    new_n8958_, new_n8959_, new_n8960_, new_n8961_, new_n8962_, new_n8963_,
    new_n8964_, new_n8965_, new_n8966_, new_n8967_, new_n8968_, new_n8969_,
    new_n8970_, new_n8971_, new_n8972_, new_n8973_, new_n8974_, new_n8975_,
    new_n8976_, new_n8977_, new_n8978_, new_n8979_, new_n8980_, new_n8981_,
    new_n8982_, new_n8983_, new_n8984_, new_n8985_, new_n8986_, new_n8987_,
    new_n8988_, new_n8989_, new_n8990_, new_n8991_, new_n8992_, new_n8993_,
    new_n8994_, new_n8995_, new_n8996_, new_n8997_, new_n8998_, new_n8999_,
    new_n9000_, new_n9001_, new_n9002_, new_n9003_, new_n9004_, new_n9005_,
    new_n9006_, new_n9007_, new_n9008_, new_n9009_, new_n9010_, new_n9011_,
    new_n9012_, new_n9013_, new_n9014_, new_n9015_, new_n9016_, new_n9017_,
    new_n9018_, new_n9019_, new_n9020_, new_n9021_, new_n9022_, new_n9023_,
    new_n9024_, new_n9025_, new_n9026_, new_n9028_, new_n9029_, new_n9030_,
    new_n9031_, new_n9032_, new_n9033_, new_n9034_, new_n9035_, new_n9036_,
    new_n9037_, new_n9038_, new_n9039_, new_n9040_, new_n9041_, new_n9042_,
    new_n9043_, new_n9044_, new_n9045_, new_n9046_, new_n9047_, new_n9048_,
    new_n9049_, new_n9050_, new_n9051_, new_n9052_, new_n9053_, new_n9054_,
    new_n9055_, new_n9056_, new_n9057_, new_n9058_, new_n9059_, new_n9060_,
    new_n9061_, new_n9062_, new_n9063_, new_n9064_, new_n9065_, new_n9066_,
    new_n9067_, new_n9068_, new_n9069_, new_n9070_, new_n9071_, new_n9072_,
    new_n9073_, new_n9074_, new_n9075_, new_n9076_, new_n9077_, new_n9078_,
    new_n9079_, new_n9080_, new_n9081_, new_n9082_, new_n9083_, new_n9084_,
    new_n9085_, new_n9086_, new_n9087_, new_n9088_, new_n9089_, new_n9090_,
    new_n9091_, new_n9092_, new_n9093_, new_n9094_, new_n9095_, new_n9096_,
    new_n9097_, new_n9098_, new_n9099_, new_n9100_, new_n9101_, new_n9102_,
    new_n9103_, new_n9104_, new_n9105_, new_n9106_, new_n9107_, new_n9108_,
    new_n9109_, new_n9110_, new_n9111_, new_n9112_, new_n9113_, new_n9114_,
    new_n9115_, new_n9116_, new_n9117_, new_n9118_, new_n9119_, new_n9120_,
    new_n9121_, new_n9122_, new_n9123_, new_n9124_, new_n9125_, new_n9126_,
    new_n9127_, new_n9128_, new_n9129_, new_n9130_, new_n9131_, new_n9132_,
    new_n9133_, new_n9134_, new_n9135_, new_n9136_, new_n9137_, new_n9138_,
    new_n9139_, new_n9140_, new_n9141_, new_n9142_, new_n9143_, new_n9144_,
    new_n9145_, new_n9146_, new_n9147_, new_n9148_, new_n9149_, new_n9150_,
    new_n9151_, new_n9152_, new_n9153_, new_n9154_, new_n9155_, new_n9156_,
    new_n9157_, new_n9158_, new_n9159_, new_n9160_, new_n9161_, new_n9162_,
    new_n9163_, new_n9164_, new_n9165_, new_n9166_, new_n9167_, new_n9168_,
    new_n9169_, new_n9170_, new_n9171_, new_n9172_, new_n9173_, new_n9174_,
    new_n9175_, new_n9176_, new_n9177_, new_n9178_, new_n9179_, new_n9180_,
    new_n9181_, new_n9182_, new_n9183_, new_n9184_, new_n9185_, new_n9186_,
    new_n9187_, new_n9188_, new_n9189_, new_n9190_, new_n9191_, new_n9192_,
    new_n9193_, new_n9194_, new_n9195_, new_n9196_, new_n9197_, new_n9198_,
    new_n9199_, new_n9200_, new_n9201_, new_n9202_, new_n9203_, new_n9204_,
    new_n9205_, new_n9206_, new_n9207_, new_n9208_, new_n9209_, new_n9210_,
    new_n9211_, new_n9212_, new_n9213_, new_n9214_, new_n9215_, new_n9216_,
    new_n9217_, new_n9218_, new_n9219_, new_n9220_, new_n9221_, new_n9222_,
    new_n9223_, new_n9224_, new_n9225_, new_n9226_, new_n9227_, new_n9228_,
    new_n9229_, new_n9230_, new_n9231_, new_n9232_, new_n9233_, new_n9234_,
    new_n9235_, new_n9236_, new_n9237_, new_n9238_, new_n9239_, new_n9240_,
    new_n9241_, new_n9242_, new_n9243_, new_n9244_, new_n9245_, new_n9246_,
    new_n9247_, new_n9248_, new_n9249_, new_n9250_, new_n9251_, new_n9252_,
    new_n9253_, new_n9254_, new_n9255_, new_n9256_, new_n9257_, new_n9258_,
    new_n9259_, new_n9260_, new_n9261_, new_n9262_, new_n9263_, new_n9264_,
    new_n9265_, new_n9266_, new_n9267_, new_n9268_, new_n9269_, new_n9270_,
    new_n9271_, new_n9272_, new_n9273_, new_n9274_, new_n9275_, new_n9276_,
    new_n9277_, new_n9278_, new_n9279_, new_n9280_, new_n9281_, new_n9282_,
    new_n9283_, new_n9284_, new_n9285_, new_n9286_, new_n9287_, new_n9288_,
    new_n9289_, new_n9290_, new_n9291_, new_n9292_, new_n9293_, new_n9294_,
    new_n9295_, new_n9296_, new_n9297_, new_n9298_, new_n9299_, new_n9300_,
    new_n9301_, new_n9302_, new_n9303_, new_n9304_, new_n9305_, new_n9306_,
    new_n9307_, new_n9308_, new_n9309_, new_n9310_, new_n9311_, new_n9312_,
    new_n9313_, new_n9314_, new_n9315_, new_n9316_, new_n9317_, new_n9318_,
    new_n9319_, new_n9320_, new_n9321_, new_n9322_, new_n9323_, new_n9324_,
    new_n9325_, new_n9326_, new_n9327_, new_n9328_, new_n9329_, new_n9330_,
    new_n9331_, new_n9332_, new_n9333_, new_n9334_, new_n9335_, new_n9336_,
    new_n9337_, new_n9338_, new_n9339_, new_n9340_, new_n9341_, new_n9342_,
    new_n9343_, new_n9344_, new_n9345_, new_n9346_, new_n9347_, new_n9348_,
    new_n9349_, new_n9350_, new_n9351_, new_n9352_, new_n9353_, new_n9354_,
    new_n9355_, new_n9356_, new_n9357_, new_n9358_, new_n9359_, new_n9360_,
    new_n9361_, new_n9362_, new_n9363_, new_n9364_, new_n9365_, new_n9366_,
    new_n9367_, new_n9368_, new_n9369_, new_n9370_, new_n9371_, new_n9372_,
    new_n9373_, new_n9374_, new_n9375_, new_n9376_, new_n9377_, new_n9378_,
    new_n9379_, new_n9380_, new_n9381_, new_n9382_, new_n9383_, new_n9384_,
    new_n9385_, new_n9386_, new_n9387_, new_n9388_, new_n9389_, new_n9390_,
    new_n9391_, new_n9392_, new_n9393_, new_n9394_, new_n9395_, new_n9396_,
    new_n9397_, new_n9398_, new_n9399_, new_n9400_, new_n9401_, new_n9402_,
    new_n9403_, new_n9404_, new_n9405_, new_n9406_, new_n9407_, new_n9408_,
    new_n9409_, new_n9410_, new_n9411_, new_n9412_, new_n9413_, new_n9414_,
    new_n9415_, new_n9416_, new_n9417_, new_n9418_, new_n9419_, new_n9420_,
    new_n9421_, new_n9422_, new_n9423_, new_n9424_, new_n9425_, new_n9426_,
    new_n9427_, new_n9428_, new_n9429_, new_n9430_, new_n9431_, new_n9432_,
    new_n9433_, new_n9434_, new_n9435_, new_n9436_, new_n9437_, new_n9438_,
    new_n9439_, new_n9440_, new_n9441_, new_n9442_, new_n9443_, new_n9444_,
    new_n9445_, new_n9446_, new_n9447_, new_n9448_, new_n9449_, new_n9450_,
    new_n9451_, new_n9452_, new_n9453_, new_n9454_, new_n9455_, new_n9456_,
    new_n9457_, new_n9458_, new_n9459_, new_n9460_, new_n9461_, new_n9462_,
    new_n9463_, new_n9464_, new_n9465_, new_n9466_, new_n9467_, new_n9468_,
    new_n9469_, new_n9470_, new_n9471_, new_n9472_, new_n9473_, new_n9474_,
    new_n9475_, new_n9476_, new_n9477_, new_n9478_, new_n9479_, new_n9480_,
    new_n9481_, new_n9482_, new_n9483_, new_n9484_, new_n9485_, new_n9486_,
    new_n9487_, new_n9488_, new_n9489_, new_n9490_, new_n9491_, new_n9492_,
    new_n9493_, new_n9494_, new_n9495_, new_n9496_, new_n9497_, new_n9498_,
    new_n9499_, new_n9500_, new_n9501_, new_n9502_, new_n9503_, new_n9504_,
    new_n9505_, new_n9506_, new_n9507_, new_n9508_, new_n9509_, new_n9510_,
    new_n9511_, new_n9512_, new_n9513_, new_n9514_, new_n9515_, new_n9516_,
    new_n9517_, new_n9518_, new_n9519_, new_n9521_, new_n9522_, new_n9523_,
    new_n9524_, new_n9525_, new_n9526_, new_n9528_, new_n9529_, new_n9530_,
    new_n9531_, new_n9533_, new_n9534_, new_n9535_, new_n9536_, new_n9537_,
    new_n9538_, new_n9539_, new_n9540_, new_n9541_, new_n9543_, new_n9544_,
    new_n9545_, new_n9546_, new_n9547_, new_n9549_, new_n9550_, new_n9551_,
    new_n9552_, new_n9554_, new_n9556_, new_n9557_, new_n9559_, new_n9560_,
    new_n9561_, new_n9562_, new_n9563_, new_n9564_, new_n9565_, new_n9566_,
    new_n9567_, new_n9568_, new_n9570_, new_n9571_, new_n9572_, new_n9573_,
    new_n9574_, new_n9575_, new_n9577_, new_n9578_, new_n9580_, new_n9581_,
    new_n9582_, new_n9583_, new_n9584_, new_n9585_, new_n9586_, new_n9588_,
    new_n9589_, new_n9590_, new_n9591_, new_n9592_, new_n9593_, new_n9594_,
    new_n9596_, new_n9597_, new_n9598_, new_n9599_, new_n9600_, new_n9602_,
    new_n9603_, new_n9604_, new_n9605_, new_n9606_, new_n9607_, new_n9608_,
    new_n9609_, new_n9610_, new_n9611_, new_n9613_, new_n9614_, new_n9615_,
    new_n9616_, new_n9617_, new_n9618_, new_n9619_, new_n9620_, new_n9622_,
    new_n9623_, new_n9624_, new_n9625_, new_n9626_, new_n9627_, new_n9629_,
    new_n9630_, new_n9631_, new_n9632_, new_n9634_, new_n9635_, new_n9637_,
    new_n9638_, new_n9639_, new_n9640_, new_n9641_, new_n9642_, new_n9643_,
    new_n9644_, new_n9645_, new_n9646_, new_n9647_, new_n9648_, new_n9649_,
    new_n9650_, new_n9651_, new_n9652_, new_n9653_, new_n9654_, new_n9655_,
    new_n9656_, new_n9657_, new_n9658_, new_n9659_, new_n9660_, new_n9661_,
    new_n9662_, new_n9663_, new_n9664_, new_n9665_, new_n9666_, new_n9667_,
    new_n9668_, new_n9669_, new_n9670_, new_n9671_, new_n9672_, new_n9673_,
    new_n9674_, new_n9675_, new_n9676_, new_n9677_, new_n9678_, new_n9679_,
    new_n9680_, new_n9681_, new_n9682_, new_n9683_, new_n9684_, new_n9685_,
    new_n9686_, new_n9687_, new_n9689_, new_n9690_, new_n9691_, new_n9692_,
    new_n9693_, new_n9694_, new_n9695_, new_n9696_, new_n9697_, new_n9698_,
    new_n9699_, new_n9701_, new_n9702_, new_n9703_, new_n9704_, new_n9705_,
    new_n9706_, new_n9707_, new_n9708_, new_n9709_, new_n9710_, new_n9711_,
    new_n9712_, new_n9713_, new_n9714_, new_n9715_, new_n9716_, new_n9717_,
    new_n9718_, new_n9719_, new_n9720_, new_n9721_, new_n9722_, new_n9723_,
    new_n9724_, new_n9725_, new_n9726_, new_n9727_, new_n9728_, new_n9729_,
    new_n9730_, new_n9731_, new_n9732_, new_n9733_, new_n9734_, new_n9735_,
    new_n9736_, new_n9737_, new_n9738_, new_n9739_, new_n9740_, new_n9741_,
    new_n9742_, new_n9743_, new_n9744_, new_n9745_, new_n9746_, new_n9747_,
    new_n9748_, new_n9749_, new_n9750_, new_n9751_, new_n9753_, new_n9754_,
    new_n9756_, new_n9757_, new_n9758_, new_n9759_, new_n9761_, new_n9762_,
    new_n9763_, new_n9764_, new_n9765_, new_n9766_, new_n9767_, new_n9768_,
    new_n9769_, new_n9770_, new_n9771_, new_n9772_, new_n9774_, new_n9775_,
    new_n9776_, new_n9777_, new_n9778_, new_n9779_, new_n9782_, new_n9783_,
    new_n9784_, new_n9785_, new_n9786_, new_n9787_, new_n9788_, new_n9789_,
    new_n9790_, new_n9791_, new_n9792_, new_n9793_, new_n9795_, new_n9797_,
    new_n9798_, new_n9799_, new_n9800_, new_n9801_, new_n9803_, new_n9804_,
    new_n9807_, new_n9808_, new_n9809_, new_n9810_, new_n9811_, new_n9812_,
    new_n9813_, new_n9814_, new_n9815_, new_n9816_, new_n9817_, new_n9818_,
    new_n9819_, new_n9820_, new_n9821_, new_n9822_, new_n9823_, new_n9824_,
    new_n9825_, new_n9826_, new_n9827_, new_n9828_, new_n9829_, new_n9830_,
    new_n9831_, new_n9832_, new_n9833_, new_n9834_, new_n9835_, new_n9836_,
    new_n9837_, new_n9838_, new_n9839_, new_n9840_, new_n9841_, new_n9843_,
    new_n9844_, new_n9845_, new_n9846_, new_n9847_, new_n9848_, new_n9849_,
    new_n9850_, new_n9851_, new_n9852_, new_n9853_, new_n9854_, new_n9855_,
    new_n9856_, new_n9857_, new_n9858_, new_n9859_, new_n9860_, new_n9861_,
    new_n9862_, new_n9863_, new_n9864_, new_n9865_, new_n9866_, new_n9868_,
    new_n9869_, new_n9870_, new_n9871_, new_n9872_, new_n9873_, new_n9874_,
    new_n9875_, new_n9876_, new_n9877_, new_n9878_, new_n9879_, new_n9880_,
    new_n9881_, new_n9882_, new_n9883_, new_n9884_, new_n9885_, new_n9886_,
    new_n9887_, new_n9888_, new_n9889_, new_n9890_, new_n9892_, new_n9893_,
    new_n9894_, new_n9895_, new_n9896_, new_n9897_, new_n9898_, new_n9899_,
    new_n9900_, new_n9901_, new_n9902_, new_n9903_, new_n9904_, new_n9905_,
    new_n9906_, new_n9907_, new_n9908_, new_n9909_, new_n9910_, new_n9911_,
    new_n9912_, new_n9913_, new_n9914_, new_n9915_, new_n9916_, new_n9917_,
    new_n9918_, new_n9919_, new_n9920_, new_n9921_, new_n9922_, new_n9924_,
    new_n9925_, new_n9926_, new_n9927_, new_n9928_, new_n9929_, new_n9930_,
    new_n9931_, new_n9933_, new_n9934_, new_n9935_, new_n9936_, new_n9937_,
    new_n9938_, new_n9939_, new_n9940_, new_n9941_, new_n9942_, new_n9943_,
    new_n9944_, new_n9945_, new_n9946_, new_n9947_, new_n9948_, new_n9949_,
    new_n9950_, new_n9951_, new_n9952_, new_n9953_, new_n9954_, new_n9955_,
    new_n9956_, new_n9957_, new_n9958_, new_n9959_, new_n9960_, new_n9961_,
    new_n9962_, new_n9963_, new_n9964_, new_n9965_, new_n9966_, new_n9967_,
    new_n9968_, new_n9969_, new_n9970_, new_n9971_, new_n9972_, new_n9973_,
    new_n9974_, new_n9975_, new_n9976_, new_n9977_, new_n9978_, new_n9979_,
    new_n9980_, new_n9981_, new_n9982_, new_n9983_, new_n9984_, new_n9985_,
    new_n9986_, new_n9987_, new_n9988_, new_n9989_, new_n9990_, new_n9991_,
    new_n9992_, new_n9993_, new_n9994_, new_n9995_, new_n9996_, new_n9997_,
    new_n9998_, new_n9999_, new_n10000_, new_n10001_, new_n10002_,
    new_n10003_, new_n10004_, new_n10005_, new_n10006_, new_n10007_,
    new_n10008_, new_n10009_, new_n10010_, new_n10011_, new_n10012_,
    new_n10013_, new_n10014_, new_n10015_, new_n10016_, new_n10017_,
    new_n10018_, new_n10019_, new_n10020_, new_n10021_, new_n10022_,
    new_n10023_, new_n10024_, new_n10025_, new_n10026_, new_n10027_,
    new_n10028_, new_n10029_, new_n10030_, new_n10031_, new_n10032_,
    new_n10033_, new_n10034_, new_n10035_, new_n10036_, new_n10037_,
    new_n10038_, new_n10039_, new_n10040_, new_n10041_, new_n10042_,
    new_n10043_, new_n10044_, new_n10045_, new_n10046_, new_n10047_,
    new_n10048_, new_n10049_, new_n10050_, new_n10051_, new_n10052_,
    new_n10053_, new_n10054_, new_n10055_, new_n10056_, new_n10057_,
    new_n10058_, new_n10059_, new_n10060_, new_n10061_, new_n10062_,
    new_n10063_, new_n10064_, new_n10065_, new_n10066_, new_n10067_,
    new_n10068_, new_n10069_, new_n10070_, new_n10071_, new_n10072_,
    new_n10073_, new_n10074_, new_n10075_, new_n10076_, new_n10077_,
    new_n10078_, new_n10079_, new_n10080_, new_n10081_, new_n10082_,
    new_n10083_, new_n10084_, new_n10085_, new_n10086_, new_n10087_,
    new_n10088_, new_n10089_, new_n10090_, new_n10091_, new_n10092_,
    new_n10093_, new_n10094_, new_n10095_, new_n10096_, new_n10097_,
    new_n10098_, new_n10099_, new_n10100_, new_n10101_, new_n10102_,
    new_n10103_, new_n10104_, new_n10105_, new_n10106_, new_n10107_,
    new_n10108_, new_n10109_, new_n10110_, new_n10111_, new_n10112_,
    new_n10113_, new_n10114_, new_n10115_, new_n10116_, new_n10117_,
    new_n10118_, new_n10119_, new_n10120_, new_n10121_, new_n10122_,
    new_n10123_, new_n10124_, new_n10125_, new_n10126_, new_n10127_,
    new_n10128_, new_n10129_, new_n10130_, new_n10131_, new_n10133_,
    new_n10134_, new_n10135_, new_n10136_, new_n10137_, new_n10138_,
    new_n10139_, new_n10140_, new_n10141_, new_n10142_, new_n10143_,
    new_n10144_, new_n10145_, new_n10146_, new_n10147_, new_n10148_,
    new_n10149_, new_n10150_, new_n10151_, new_n10152_, new_n10153_,
    new_n10154_, new_n10155_, new_n10156_, new_n10157_, new_n10158_,
    new_n10159_, new_n10160_, new_n10161_, new_n10162_, new_n10163_,
    new_n10165_, new_n10166_, new_n10167_, new_n10168_, new_n10169_,
    new_n10170_, new_n10171_, new_n10172_, new_n10173_, new_n10174_,
    new_n10175_, new_n10176_, new_n10177_, new_n10178_, new_n10179_,
    new_n10180_, new_n10181_, new_n10182_, new_n10183_, new_n10184_,
    new_n10185_, new_n10186_, new_n10187_, new_n10188_, new_n10189_,
    new_n10190_, new_n10191_, new_n10192_, new_n10193_, new_n10194_,
    new_n10195_, new_n10196_, new_n10197_, new_n10198_, new_n10199_,
    new_n10200_, new_n10201_, new_n10202_, new_n10203_, new_n10204_,
    new_n10205_, new_n10206_, new_n10207_, new_n10208_, new_n10209_,
    new_n10210_, new_n10211_, new_n10212_, new_n10213_, new_n10214_,
    new_n10215_, new_n10216_, new_n10217_, new_n10218_, new_n10219_,
    new_n10220_, new_n10221_, new_n10222_, new_n10223_, new_n10224_,
    new_n10225_, new_n10226_, new_n10227_, new_n10228_, new_n10229_,
    new_n10230_, new_n10231_, new_n10232_, new_n10233_, new_n10234_,
    new_n10235_, new_n10236_, new_n10237_, new_n10238_, new_n10239_,
    new_n10240_, new_n10241_, new_n10242_, new_n10243_, new_n10244_,
    new_n10245_, new_n10246_, new_n10247_, new_n10248_, new_n10249_,
    new_n10250_, new_n10251_, new_n10252_, new_n10253_, new_n10254_,
    new_n10255_, new_n10256_, new_n10257_, new_n10258_, new_n10259_,
    new_n10260_, new_n10261_, new_n10262_, new_n10263_, new_n10264_,
    new_n10265_, new_n10266_, new_n10267_, new_n10268_, new_n10269_,
    new_n10270_, new_n10271_, new_n10272_, new_n10273_, new_n10274_,
    new_n10275_, new_n10276_, new_n10277_, new_n10278_, new_n10279_,
    new_n10280_, new_n10281_, new_n10282_, new_n10283_, new_n10284_,
    new_n10285_, new_n10286_, new_n10287_, new_n10288_, new_n10289_,
    new_n10290_, new_n10291_, new_n10292_, new_n10293_, new_n10294_,
    new_n10295_, new_n10296_, new_n10297_, new_n10298_, new_n10299_,
    new_n10300_, new_n10301_, new_n10302_, new_n10303_, new_n10304_,
    new_n10305_, new_n10306_, new_n10307_, new_n10308_, new_n10309_,
    new_n10310_, new_n10311_, new_n10312_, new_n10313_, new_n10314_,
    new_n10315_, new_n10316_, new_n10317_, new_n10318_, new_n10319_,
    new_n10320_, new_n10321_, new_n10322_, new_n10323_, new_n10324_,
    new_n10325_, new_n10326_, new_n10327_, new_n10328_, new_n10329_,
    new_n10330_, new_n10331_, new_n10332_, new_n10333_, new_n10334_,
    new_n10335_, new_n10336_, new_n10337_, new_n10338_, new_n10339_,
    new_n10340_, new_n10341_, new_n10342_, new_n10343_, new_n10344_,
    new_n10345_, new_n10346_, new_n10347_, new_n10348_, new_n10349_,
    new_n10350_, new_n10351_, new_n10352_, new_n10353_, new_n10354_,
    new_n10355_, new_n10356_, new_n10357_, new_n10358_, new_n10359_,
    new_n10360_, new_n10361_, new_n10362_, new_n10363_, new_n10364_,
    new_n10365_, new_n10366_, new_n10367_, new_n10368_, new_n10369_,
    new_n10370_, new_n10371_, new_n10372_, new_n10373_, new_n10374_,
    new_n10375_, new_n10376_, new_n10377_, new_n10378_, new_n10379_,
    new_n10380_, new_n10381_, new_n10382_, new_n10383_, new_n10384_,
    new_n10385_, new_n10386_, new_n10387_, new_n10388_, new_n10389_,
    new_n10390_, new_n10391_, new_n10392_, new_n10393_, new_n10394_,
    new_n10395_, new_n10396_, new_n10397_, new_n10398_, new_n10399_,
    new_n10400_, new_n10401_, new_n10402_, new_n10403_, new_n10404_,
    new_n10405_, new_n10406_, new_n10407_, new_n10408_, new_n10409_,
    new_n10410_, new_n10411_, new_n10412_, new_n10413_, new_n10414_,
    new_n10415_, new_n10416_, new_n10417_, new_n10418_, new_n10419_,
    new_n10420_, new_n10421_, new_n10422_, new_n10423_, new_n10424_,
    new_n10425_, new_n10426_, new_n10427_, new_n10428_, new_n10429_,
    new_n10431_, new_n10432_, new_n10433_, new_n10434_, new_n10435_,
    new_n10436_, new_n10437_, new_n10438_, new_n10439_, new_n10440_,
    new_n10441_, new_n10442_, new_n10443_, new_n10444_, new_n10445_,
    new_n10446_, new_n10447_, new_n10448_, new_n10449_, new_n10450_,
    new_n10451_, new_n10452_, new_n10453_, new_n10454_, new_n10455_,
    new_n10456_, new_n10457_, new_n10458_, new_n10459_, new_n10460_,
    new_n10461_, new_n10462_, new_n10463_, new_n10464_, new_n10465_,
    new_n10466_, new_n10467_, new_n10468_, new_n10469_, new_n10470_,
    new_n10471_, new_n10472_, new_n10473_, new_n10474_, new_n10475_,
    new_n10476_, new_n10477_, new_n10478_, new_n10479_, new_n10480_,
    new_n10481_, new_n10482_, new_n10483_, new_n10484_, new_n10485_,
    new_n10486_, new_n10487_, new_n10488_, new_n10489_, new_n10490_,
    new_n10491_, new_n10492_, new_n10493_, new_n10494_, new_n10495_,
    new_n10496_, new_n10497_, new_n10498_, new_n10499_, new_n10500_,
    new_n10501_, new_n10502_, new_n10503_, new_n10504_, new_n10505_,
    new_n10506_, new_n10507_, new_n10508_, new_n10509_, new_n10510_,
    new_n10511_, new_n10512_, new_n10513_, new_n10514_, new_n10515_,
    new_n10516_, new_n10517_, new_n10518_, new_n10519_, new_n10520_,
    new_n10521_, new_n10522_, new_n10523_, new_n10524_, new_n10525_,
    new_n10526_, new_n10527_, new_n10528_, new_n10529_, new_n10530_,
    new_n10531_, new_n10532_, new_n10533_, new_n10534_, new_n10535_,
    new_n10536_, new_n10537_, new_n10538_, new_n10539_, new_n10540_,
    new_n10541_, new_n10542_, new_n10543_, new_n10544_, new_n10545_,
    new_n10546_, new_n10547_, new_n10548_, new_n10549_, new_n10550_,
    new_n10551_, new_n10552_, new_n10553_, new_n10554_, new_n10555_,
    new_n10556_, new_n10557_, new_n10558_, new_n10559_, new_n10560_,
    new_n10561_, new_n10562_, new_n10563_, new_n10564_, new_n10565_,
    new_n10566_, new_n10567_, new_n10568_, new_n10569_, new_n10570_,
    new_n10571_, new_n10572_, new_n10573_, new_n10574_, new_n10575_,
    new_n10576_, new_n10577_, new_n10578_, new_n10579_, new_n10580_,
    new_n10581_, new_n10582_, new_n10583_, new_n10584_, new_n10585_,
    new_n10586_, new_n10587_, new_n10588_, new_n10589_, new_n10590_,
    new_n10591_, new_n10592_, new_n10593_, new_n10594_, new_n10595_,
    new_n10596_, new_n10597_, new_n10598_, new_n10599_, new_n10600_,
    new_n10601_, new_n10602_, new_n10603_, new_n10604_, new_n10605_,
    new_n10606_, new_n10607_, new_n10608_, new_n10609_, new_n10610_,
    new_n10611_, new_n10612_, new_n10613_, new_n10614_, new_n10615_,
    new_n10616_, new_n10617_, new_n10618_, new_n10619_, new_n10620_,
    new_n10621_, new_n10622_, new_n10623_, new_n10624_, new_n10625_,
    new_n10626_, new_n10627_, new_n10628_, new_n10629_, new_n10630_,
    new_n10631_, new_n10632_, new_n10633_, new_n10634_, new_n10635_,
    new_n10636_, new_n10637_, new_n10638_, new_n10639_, new_n10640_,
    new_n10641_, new_n10642_, new_n10643_, new_n10644_, new_n10645_,
    new_n10646_, new_n10647_, new_n10648_, new_n10649_, new_n10650_,
    new_n10651_, new_n10652_, new_n10653_, new_n10654_, new_n10655_,
    new_n10656_, new_n10657_, new_n10658_, new_n10659_, new_n10660_,
    new_n10661_, new_n10662_, new_n10663_, new_n10664_, new_n10665_,
    new_n10666_, new_n10667_, new_n10668_, new_n10669_, new_n10670_,
    new_n10671_, new_n10672_, new_n10673_, new_n10674_, new_n10675_,
    new_n10676_, new_n10677_, new_n10678_, new_n10679_, new_n10680_,
    new_n10681_, new_n10682_, new_n10683_, new_n10684_, new_n10685_,
    new_n10686_, new_n10687_, new_n10688_, new_n10689_, new_n10690_,
    new_n10691_, new_n10692_, new_n10693_, new_n10694_, new_n10695_,
    new_n10696_, new_n10697_, new_n10698_, new_n10699_, new_n10700_,
    new_n10701_, new_n10702_, new_n10703_, new_n10704_, new_n10705_,
    new_n10706_, new_n10707_, new_n10708_, new_n10709_, new_n10710_,
    new_n10711_, new_n10712_, new_n10713_, new_n10714_, new_n10715_,
    new_n10716_, new_n10717_, new_n10718_, new_n10719_, new_n10720_,
    new_n10721_, new_n10722_, new_n10723_, new_n10724_, new_n10726_,
    new_n10727_, new_n10728_, new_n10730_, new_n10731_, new_n10732_,
    new_n10733_, new_n10734_, new_n10735_, new_n10736_, new_n10737_,
    new_n10738_, new_n10739_, new_n10740_, new_n10741_, new_n10742_,
    new_n10743_, new_n10744_, new_n10745_, new_n10746_, new_n10747_,
    new_n10748_, new_n10749_, new_n10750_, new_n10751_, new_n10752_,
    new_n10753_, new_n10754_, new_n10755_, new_n10756_, new_n10757_,
    new_n10758_, new_n10759_, new_n10760_, new_n10761_, new_n10762_,
    new_n10763_, new_n10764_, new_n10766_, new_n10767_, new_n10768_,
    new_n10769_, new_n10770_, new_n10771_, new_n10772_, new_n10773_,
    new_n10774_, new_n10775_, new_n10776_, new_n10777_, new_n10778_,
    new_n10779_, new_n10780_, new_n10781_, new_n10782_, new_n10783_,
    new_n10784_, new_n10785_, new_n10786_, new_n10787_, new_n10788_,
    new_n10789_, new_n10790_, new_n10791_, new_n10792_, new_n10793_,
    new_n10794_, new_n10795_, new_n10796_, new_n10797_, new_n10798_,
    new_n10799_, new_n10800_, new_n10801_, new_n10802_, new_n10803_,
    new_n10804_, new_n10805_, new_n10806_, new_n10807_, new_n10808_,
    new_n10809_, new_n10810_, new_n10811_, new_n10812_, new_n10813_,
    new_n10814_, new_n10815_, new_n10816_, new_n10817_, new_n10818_,
    new_n10819_, new_n10820_, new_n10821_, new_n10822_, new_n10823_,
    new_n10824_, new_n10825_, new_n10826_, new_n10827_, new_n10828_,
    new_n10829_, new_n10830_, new_n10831_, new_n10832_, new_n10833_,
    new_n10834_, new_n10835_, new_n10836_, new_n10837_, new_n10838_,
    new_n10839_, new_n10840_, new_n10841_, new_n10842_, new_n10843_,
    new_n10844_, new_n10845_, new_n10846_, new_n10847_, new_n10848_,
    new_n10849_, new_n10850_, new_n10851_, new_n10852_, new_n10853_,
    new_n10854_, new_n10855_, new_n10856_, new_n10857_, new_n10858_,
    new_n10859_, new_n10860_, new_n10861_, new_n10862_, new_n10863_,
    new_n10864_, new_n10865_, new_n10866_, new_n10867_, new_n10868_,
    new_n10869_, new_n10870_, new_n10871_, new_n10872_, new_n10873_,
    new_n10874_, new_n10875_, new_n10876_, new_n10877_, new_n10878_,
    new_n10879_, new_n10880_, new_n10881_, new_n10882_, new_n10883_,
    new_n10884_, new_n10885_, new_n10886_, new_n10887_, new_n10888_,
    new_n10889_, new_n10890_, new_n10891_, new_n10892_, new_n10893_,
    new_n10894_, new_n10895_, new_n10896_, new_n10897_, new_n10898_,
    new_n10899_, new_n10900_, new_n10901_, new_n10902_, new_n10903_,
    new_n10904_, new_n10905_, new_n10906_, new_n10907_, new_n10908_,
    new_n10909_, new_n10910_, new_n10911_, new_n10912_, new_n10913_,
    new_n10914_, new_n10915_, new_n10916_, new_n10917_, new_n10918_,
    new_n10919_, new_n10920_, new_n10921_, new_n10922_, new_n10923_,
    new_n10924_, new_n10925_, new_n10926_, new_n10927_, new_n10928_,
    new_n10929_, new_n10930_, new_n10931_, new_n10932_, new_n10933_,
    new_n10934_, new_n10935_, new_n10936_, new_n10937_, new_n10938_,
    new_n10939_, new_n10940_, new_n10941_, new_n10942_, new_n10943_,
    new_n10944_, new_n10945_, new_n10946_, new_n10947_, new_n10948_,
    new_n10949_, new_n10950_, new_n10951_, new_n10952_, new_n10953_,
    new_n10954_, new_n10955_, new_n10956_, new_n10957_, new_n10958_,
    new_n10959_, new_n10960_, new_n10961_, new_n10962_, new_n10963_,
    new_n10964_, new_n10965_, new_n10966_, new_n10967_, new_n10968_,
    new_n10969_, new_n10970_, new_n10971_, new_n10972_, new_n10973_,
    new_n10974_, new_n10975_, new_n10976_, new_n10977_, new_n10978_,
    new_n10979_, new_n10980_, new_n10981_, new_n10982_, new_n10983_,
    new_n10984_, new_n10985_, new_n10986_, new_n10987_, new_n10988_,
    new_n10989_, new_n10990_, new_n10991_, new_n10992_, new_n10993_,
    new_n10994_, new_n10995_, new_n10996_, new_n10997_, new_n10998_,
    new_n10999_, new_n11000_, new_n11001_, new_n11002_, new_n11003_,
    new_n11004_, new_n11005_, new_n11006_, new_n11007_, new_n11008_,
    new_n11009_, new_n11010_, new_n11011_, new_n11012_, new_n11013_,
    new_n11014_, new_n11015_, new_n11016_, new_n11017_, new_n11018_,
    new_n11019_, new_n11020_, new_n11021_, new_n11022_, new_n11023_,
    new_n11024_, new_n11025_, new_n11026_, new_n11027_, new_n11028_,
    new_n11029_, new_n11031_, new_n11032_, new_n11033_, new_n11034_,
    new_n11035_, new_n11036_, new_n11037_, new_n11038_, new_n11039_,
    new_n11040_, new_n11041_, new_n11042_, new_n11043_, new_n11044_,
    new_n11045_, new_n11046_, new_n11047_, new_n11048_, new_n11049_,
    new_n11050_, new_n11051_, new_n11052_, new_n11053_, new_n11054_,
    new_n11055_, new_n11056_, new_n11057_, new_n11058_, new_n11059_,
    new_n11060_, new_n11061_, new_n11062_, new_n11063_, new_n11064_,
    new_n11065_, new_n11066_, new_n11067_, new_n11068_, new_n11069_,
    new_n11070_, new_n11071_, new_n11072_, new_n11073_, new_n11074_,
    new_n11075_, new_n11076_, new_n11077_, new_n11078_, new_n11079_,
    new_n11080_, new_n11081_, new_n11082_, new_n11083_, new_n11084_,
    new_n11085_, new_n11086_, new_n11087_, new_n11088_, new_n11089_,
    new_n11090_, new_n11091_, new_n11092_, new_n11093_, new_n11094_,
    new_n11095_, new_n11096_, new_n11097_, new_n11098_, new_n11099_,
    new_n11100_, new_n11101_, new_n11102_, new_n11103_, new_n11104_,
    new_n11105_, new_n11106_, new_n11107_, new_n11108_, new_n11109_,
    new_n11110_, new_n11111_, new_n11112_, new_n11113_, new_n11114_,
    new_n11115_, new_n11116_, new_n11117_, new_n11118_, new_n11119_,
    new_n11120_, new_n11121_, new_n11122_, new_n11123_, new_n11124_,
    new_n11125_, new_n11126_, new_n11127_, new_n11128_, new_n11129_,
    new_n11130_, new_n11131_, new_n11132_, new_n11133_, new_n11134_,
    new_n11135_, new_n11136_, new_n11137_, new_n11138_, new_n11139_,
    new_n11140_, new_n11141_, new_n11142_, new_n11143_, new_n11144_,
    new_n11145_, new_n11146_, new_n11147_, new_n11148_, new_n11149_,
    new_n11150_, new_n11151_, new_n11152_, new_n11153_, new_n11154_,
    new_n11155_, new_n11156_, new_n11157_, new_n11158_, new_n11159_,
    new_n11160_, new_n11161_, new_n11162_, new_n11163_, new_n11164_,
    new_n11165_, new_n11166_, new_n11167_, new_n11168_, new_n11169_,
    new_n11170_, new_n11171_, new_n11172_, new_n11173_, new_n11174_,
    new_n11175_, new_n11176_, new_n11177_, new_n11178_, new_n11179_,
    new_n11180_, new_n11181_, new_n11182_, new_n11183_, new_n11184_,
    new_n11185_, new_n11186_, new_n11187_, new_n11188_, new_n11189_,
    new_n11190_, new_n11191_, new_n11192_, new_n11193_, new_n11194_,
    new_n11195_, new_n11196_, new_n11197_, new_n11198_, new_n11199_,
    new_n11200_, new_n11201_, new_n11202_, new_n11203_, new_n11204_,
    new_n11205_, new_n11206_, new_n11207_, new_n11208_, new_n11209_,
    new_n11210_, new_n11211_, new_n11212_, new_n11213_, new_n11214_,
    new_n11215_, new_n11216_, new_n11217_, new_n11218_, new_n11219_,
    new_n11220_, new_n11221_, new_n11222_, new_n11224_, new_n11225_,
    new_n11226_, new_n11227_, new_n11228_, new_n11229_, new_n11230_,
    new_n11231_, new_n11232_, new_n11233_, new_n11234_, new_n11235_,
    new_n11236_, new_n11237_, new_n11238_, new_n11239_, new_n11240_,
    new_n11241_, new_n11242_, new_n11243_, new_n11244_, new_n11245_,
    new_n11246_, new_n11247_, new_n11248_, new_n11249_, new_n11250_,
    new_n11251_, new_n11252_, new_n11253_, new_n11254_, new_n11255_,
    new_n11256_, new_n11257_, new_n11258_, new_n11259_, new_n11260_,
    new_n11261_, new_n11262_, new_n11263_, new_n11264_, new_n11265_,
    new_n11266_, new_n11267_, new_n11268_, new_n11269_, new_n11270_,
    new_n11271_, new_n11272_, new_n11273_, new_n11274_, new_n11275_,
    new_n11276_, new_n11277_, new_n11278_, new_n11279_, new_n11280_,
    new_n11282_, new_n11283_, new_n11284_, new_n11285_, new_n11286_,
    new_n11287_, new_n11288_, new_n11289_, new_n11290_, new_n11291_,
    new_n11292_, new_n11293_, new_n11294_, new_n11295_, new_n11296_,
    new_n11298_, new_n11299_, new_n11300_, new_n11301_, new_n11302_,
    new_n11303_, new_n11304_, new_n11305_, new_n11306_, new_n11307_,
    new_n11308_, new_n11309_, new_n11310_, new_n11311_, new_n11312_,
    new_n11313_, new_n11314_, new_n11315_, new_n11316_, new_n11317_,
    new_n11318_, new_n11319_, new_n11320_, new_n11321_, new_n11322_,
    new_n11323_, new_n11324_, new_n11325_, new_n11326_, new_n11327_,
    new_n11328_, new_n11329_, new_n11330_, new_n11331_, new_n11332_,
    new_n11333_, new_n11334_, new_n11335_, new_n11336_, new_n11337_,
    new_n11338_, new_n11339_, new_n11340_, new_n11341_, new_n11342_,
    new_n11343_, new_n11344_, new_n11345_, new_n11346_, new_n11347_,
    new_n11348_, new_n11349_, new_n11350_, new_n11351_, new_n11352_,
    new_n11353_, new_n11354_, new_n11355_, new_n11356_, new_n11357_,
    new_n11358_, new_n11359_, new_n11360_, new_n11361_, new_n11362_,
    new_n11363_, new_n11364_, new_n11365_, new_n11366_, new_n11367_,
    new_n11368_, new_n11369_, new_n11370_, new_n11371_, new_n11372_,
    new_n11373_, new_n11374_, new_n11375_, new_n11376_, new_n11377_,
    new_n11378_, new_n11379_, new_n11380_, new_n11381_, new_n11382_,
    new_n11383_, new_n11384_, new_n11385_, new_n11386_, new_n11388_,
    new_n11389_, new_n11390_, new_n11391_, new_n11393_, new_n11394_,
    new_n11395_, new_n11396_, new_n11397_, new_n11398_, new_n11399_,
    new_n11400_, new_n11401_, new_n11402_, new_n11403_, new_n11404_,
    new_n11405_, new_n11406_, new_n11407_, new_n11408_, new_n11409_,
    new_n11410_, new_n11411_, new_n11412_, new_n11413_, new_n11414_,
    new_n11415_, new_n11416_, new_n11417_, new_n11418_, new_n11419_,
    new_n11420_, new_n11421_, new_n11422_, new_n11423_, new_n11424_,
    new_n11425_, new_n11426_, new_n11427_, new_n11428_, new_n11429_,
    new_n11430_, new_n11431_, new_n11432_, new_n11433_, new_n11434_,
    new_n11435_, new_n11436_, new_n11437_, new_n11438_, new_n11439_,
    new_n11440_, new_n11441_, new_n11442_, new_n11443_, new_n11444_,
    new_n11445_, new_n11446_, new_n11447_, new_n11448_, new_n11449_,
    new_n11450_, new_n11451_, new_n11452_, new_n11453_, new_n11454_,
    new_n11455_, new_n11456_, new_n11457_, new_n11458_, new_n11459_,
    new_n11460_, new_n11461_, new_n11462_, new_n11463_, new_n11464_,
    new_n11465_, new_n11466_, new_n11467_, new_n11468_, new_n11469_,
    new_n11470_, new_n11471_, new_n11472_, new_n11473_, new_n11474_,
    new_n11475_, new_n11476_, new_n11477_, new_n11478_, new_n11479_,
    new_n11480_, new_n11481_, new_n11482_, new_n11483_, new_n11484_,
    new_n11485_, new_n11486_, new_n11487_, new_n11488_, new_n11489_,
    new_n11490_, new_n11491_, new_n11492_, new_n11493_, new_n11494_,
    new_n11495_, new_n11496_, new_n11497_, new_n11498_, new_n11499_,
    new_n11500_, new_n11501_, new_n11502_, new_n11503_, new_n11504_,
    new_n11505_, new_n11506_, new_n11507_, new_n11508_, new_n11509_,
    new_n11510_, new_n11511_, new_n11512_, new_n11513_, new_n11514_,
    new_n11515_, new_n11516_, new_n11517_, new_n11518_, new_n11519_,
    new_n11520_, new_n11521_, new_n11522_, new_n11523_, new_n11525_,
    new_n11526_, new_n11527_, new_n11528_, new_n11529_, new_n11530_,
    new_n11531_, new_n11532_, new_n11533_, new_n11534_, new_n11535_,
    new_n11536_, new_n11537_, new_n11538_, new_n11539_, new_n11540_,
    new_n11541_, new_n11542_, new_n11543_, new_n11544_, new_n11545_,
    new_n11546_, new_n11547_, new_n11548_, new_n11549_, new_n11550_,
    new_n11551_, new_n11552_, new_n11553_, new_n11554_, new_n11555_,
    new_n11556_, new_n11557_, new_n11558_, new_n11559_, new_n11560_,
    new_n11561_, new_n11563_, new_n11564_, new_n11565_, new_n11566_,
    new_n11567_, new_n11568_, new_n11569_, new_n11570_, new_n11571_,
    new_n11572_, new_n11573_, new_n11574_, new_n11575_, new_n11576_,
    new_n11577_, new_n11578_, new_n11579_, new_n11580_, new_n11581_,
    new_n11582_, new_n11583_, new_n11584_, new_n11585_, new_n11586_,
    new_n11587_, new_n11588_, new_n11589_, new_n11590_, new_n11591_,
    new_n11592_, new_n11593_, new_n11594_, new_n11595_, new_n11596_,
    new_n11597_, new_n11598_, new_n11599_, new_n11600_, new_n11601_,
    new_n11602_, new_n11603_, new_n11604_, new_n11605_, new_n11606_,
    new_n11607_, new_n11608_, new_n11609_, new_n11610_, new_n11611_,
    new_n11612_, new_n11613_, new_n11614_, new_n11615_, new_n11616_,
    new_n11617_, new_n11618_, new_n11619_, new_n11620_, new_n11621_,
    new_n11622_, new_n11623_, new_n11624_, new_n11625_, new_n11626_,
    new_n11627_, new_n11628_, new_n11629_, new_n11630_, new_n11631_,
    new_n11632_, new_n11633_, new_n11634_, new_n11635_, new_n11636_,
    new_n11637_, new_n11638_, new_n11639_, new_n11641_, new_n11642_,
    new_n11643_, new_n11644_, new_n11645_, new_n11646_, new_n11647_,
    new_n11648_, new_n11649_, new_n11650_, new_n11651_, new_n11652_,
    new_n11653_, new_n11654_, new_n11655_, new_n11656_, new_n11657_,
    new_n11658_, new_n11659_, new_n11660_, new_n11661_, new_n11662_,
    new_n11663_, new_n11664_, new_n11665_, new_n11666_, new_n11667_,
    new_n11668_, new_n11669_, new_n11670_, new_n11671_, new_n11672_,
    new_n11673_, new_n11674_, new_n11675_, new_n11676_, new_n11677_,
    new_n11678_, new_n11679_, new_n11680_, new_n11681_, new_n11682_,
    new_n11683_, new_n11684_, new_n11685_, new_n11686_, new_n11687_,
    new_n11688_, new_n11689_, new_n11690_, new_n11691_, new_n11692_,
    new_n11693_, new_n11694_, new_n11695_, new_n11696_, new_n11697_,
    new_n11698_, new_n11699_, new_n11700_, new_n11701_, new_n11702_,
    new_n11703_, new_n11704_, new_n11705_, new_n11706_, new_n11707_,
    new_n11708_, new_n11709_, new_n11710_, new_n11711_, new_n11712_,
    new_n11713_, new_n11714_, new_n11715_, new_n11716_, new_n11717_,
    new_n11718_, new_n11720_, new_n11721_, new_n11722_, new_n11723_,
    new_n11724_, new_n11725_, new_n11726_, new_n11727_, new_n11728_,
    new_n11729_, new_n11730_, new_n11731_, new_n11732_, new_n11733_,
    new_n11734_, new_n11735_, new_n11736_, new_n11737_, new_n11738_,
    new_n11739_, new_n11740_, new_n11741_, new_n11742_, new_n11743_,
    new_n11744_, new_n11745_, new_n11746_, new_n11747_, new_n11748_,
    new_n11749_, new_n11750_, new_n11751_, new_n11752_, new_n11753_,
    new_n11754_, new_n11755_, new_n11756_, new_n11757_, new_n11758_,
    new_n11759_, new_n11760_, new_n11761_, new_n11762_, new_n11763_,
    new_n11764_, new_n11765_, new_n11766_, new_n11767_, new_n11768_,
    new_n11769_, new_n11770_, new_n11771_, new_n11772_, new_n11774_,
    new_n11775_, new_n11776_, new_n11777_, new_n11778_, new_n11779_,
    new_n11780_, new_n11781_, new_n11783_, new_n11784_, new_n11785_,
    new_n11786_, new_n11787_, new_n11788_, new_n11789_, new_n11790_,
    new_n11791_, new_n11792_, new_n11793_, new_n11794_, new_n11795_,
    new_n11796_, new_n11797_, new_n11798_, new_n11799_, new_n11800_,
    new_n11801_, new_n11802_, new_n11803_, new_n11804_, new_n11805_,
    new_n11806_, new_n11807_, new_n11808_, new_n11809_, new_n11810_,
    new_n11811_, new_n11812_, new_n11813_, new_n11814_, new_n11815_,
    new_n11816_, new_n11817_, new_n11818_, new_n11819_, new_n11820_,
    new_n11821_, new_n11822_, new_n11823_, new_n11824_, new_n11825_,
    new_n11826_, new_n11827_, new_n11828_, new_n11829_, new_n11830_,
    new_n11831_, new_n11832_, new_n11833_, new_n11834_, new_n11835_,
    new_n11836_, new_n11837_, new_n11838_, new_n11839_, new_n11840_,
    new_n11841_, new_n11842_, new_n11843_, new_n11844_, new_n11845_,
    new_n11846_, new_n11847_, new_n11849_, new_n11850_, new_n11851_,
    new_n11852_, new_n11853_, new_n11854_, new_n11855_, new_n11856_,
    new_n11857_, new_n11858_, new_n11859_, new_n11860_, new_n11861_,
    new_n11862_, new_n11863_, new_n11864_, new_n11865_, new_n11866_,
    new_n11867_, new_n11868_, new_n11869_, new_n11870_, new_n11871_,
    new_n11872_, new_n11873_, new_n11874_, new_n11875_, new_n11876_,
    new_n11877_, new_n11878_, new_n11879_, new_n11880_, new_n11882_,
    new_n11883_, new_n11884_, new_n11885_, new_n11886_, new_n11887_,
    new_n11888_, new_n11889_, new_n11890_, new_n11891_, new_n11892_,
    new_n11893_, new_n11894_, new_n11895_, new_n11896_, new_n11897_,
    new_n11898_, new_n11899_, new_n11900_, new_n11901_, new_n11902_,
    new_n11903_, new_n11904_, new_n11905_, new_n11906_, new_n11907_,
    new_n11908_, new_n11909_, new_n11910_, new_n11911_, new_n11912_,
    new_n11913_, new_n11914_, new_n11915_, new_n11916_, new_n11917_,
    new_n11918_, new_n11919_, new_n11920_, new_n11921_, new_n11922_,
    new_n11923_, new_n11925_, new_n11926_, new_n11927_, new_n11928_,
    new_n11929_, new_n11930_, new_n11931_, new_n11932_, new_n11933_,
    new_n11934_, new_n11935_, new_n11936_, new_n11937_, new_n11938_,
    new_n11939_, new_n11940_, new_n11941_, new_n11942_, new_n11943_,
    new_n11944_, new_n11945_, new_n11946_, new_n11947_, new_n11948_,
    new_n11949_, new_n11950_, new_n11951_, new_n11952_, new_n11953_,
    new_n11954_, new_n11955_, new_n11956_, new_n11957_, new_n11958_,
    new_n11959_, new_n11960_, new_n11961_, new_n11962_, new_n11963_,
    new_n11964_, new_n11965_, new_n11966_, new_n11967_, new_n11968_,
    new_n11969_, new_n11970_, new_n11971_, new_n11972_, new_n11973_,
    new_n11974_, new_n11975_, new_n11976_, new_n11977_, new_n11978_,
    new_n11979_, new_n11980_, new_n11981_, new_n11982_, new_n11983_,
    new_n11984_, new_n11985_, new_n11986_, new_n11987_, new_n11988_,
    new_n11989_, new_n11990_, new_n11991_, new_n11992_, new_n11993_,
    new_n11994_, new_n11995_, new_n11996_, new_n11997_, new_n11998_,
    new_n11999_, new_n12000_, new_n12001_, new_n12002_, new_n12003_,
    new_n12004_, new_n12005_, new_n12006_, new_n12007_, new_n12008_,
    new_n12009_, new_n12010_, new_n12011_, new_n12012_, new_n12013_,
    new_n12014_, new_n12015_, new_n12016_, new_n12017_, new_n12018_,
    new_n12019_, new_n12020_, new_n12021_, new_n12022_, new_n12023_,
    new_n12024_, new_n12025_, new_n12026_, new_n12027_, new_n12028_,
    new_n12029_, new_n12030_, new_n12031_, new_n12032_, new_n12033_,
    new_n12034_, new_n12035_, new_n12036_, new_n12037_, new_n12038_,
    new_n12039_, new_n12040_, new_n12041_, new_n12042_, new_n12043_,
    new_n12044_, new_n12045_, new_n12046_, new_n12047_, new_n12048_,
    new_n12049_, new_n12050_, new_n12051_, new_n12052_, new_n12053_,
    new_n12054_, new_n12055_, new_n12056_, new_n12057_, new_n12058_,
    new_n12059_, new_n12060_, new_n12061_, new_n12062_, new_n12063_,
    new_n12064_, new_n12065_, new_n12066_, new_n12067_, new_n12068_,
    new_n12069_, new_n12070_, new_n12071_, new_n12072_, new_n12073_,
    new_n12074_, new_n12075_, new_n12076_, new_n12077_, new_n12078_,
    new_n12079_, new_n12080_, new_n12081_, new_n12082_, new_n12083_,
    new_n12084_, new_n12085_, new_n12086_, new_n12087_, new_n12088_,
    new_n12089_, new_n12090_, new_n12091_, new_n12092_, new_n12093_,
    new_n12094_, new_n12095_, new_n12096_, new_n12097_, new_n12098_,
    new_n12099_, new_n12100_, new_n12101_, new_n12102_, new_n12103_,
    new_n12104_, new_n12105_, new_n12106_, new_n12107_, new_n12108_,
    new_n12109_, new_n12110_, new_n12111_, new_n12112_, new_n12113_,
    new_n12114_, new_n12115_, new_n12116_, new_n12117_, new_n12118_,
    new_n12119_, new_n12120_, new_n12121_, new_n12122_, new_n12123_,
    new_n12124_, new_n12125_, new_n12126_, new_n12127_, new_n12128_,
    new_n12129_, new_n12130_, new_n12131_, new_n12132_, new_n12133_,
    new_n12134_, new_n12135_, new_n12136_, new_n12137_, new_n12138_,
    new_n12139_, new_n12140_, new_n12141_, new_n12142_, new_n12143_,
    new_n12144_, new_n12145_, new_n12146_, new_n12147_, new_n12148_,
    new_n12149_, new_n12150_, new_n12151_, new_n12152_, new_n12153_,
    new_n12154_, new_n12155_, new_n12156_, new_n12157_, new_n12158_,
    new_n12159_, new_n12160_, new_n12161_, new_n12162_, new_n12163_,
    new_n12164_, new_n12165_, new_n12166_, new_n12167_, new_n12168_,
    new_n12169_, new_n12170_, new_n12171_, new_n12172_, new_n12173_,
    new_n12174_, new_n12175_, new_n12176_, new_n12177_, new_n12178_,
    new_n12179_, new_n12180_, new_n12181_, new_n12182_, new_n12183_,
    new_n12184_, new_n12185_, new_n12186_, new_n12187_, new_n12188_,
    new_n12189_, new_n12190_, new_n12191_, new_n12192_, new_n12193_,
    new_n12194_, new_n12195_, new_n12196_, new_n12197_, new_n12198_,
    new_n12199_, new_n12200_, new_n12201_, new_n12202_, new_n12203_,
    new_n12204_, new_n12205_, new_n12206_, new_n12207_, new_n12208_,
    new_n12209_, new_n12210_, new_n12211_, new_n12212_, new_n12213_,
    new_n12214_, new_n12215_, new_n12216_, new_n12217_, new_n12218_,
    new_n12219_, new_n12220_, new_n12221_, new_n12222_, new_n12223_,
    new_n12224_, new_n12225_, new_n12226_, new_n12227_, new_n12228_,
    new_n12229_, new_n12230_, new_n12231_, new_n12232_, new_n12233_,
    new_n12234_, new_n12235_, new_n12236_, new_n12237_, new_n12238_,
    new_n12239_, new_n12240_, new_n12241_, new_n12242_, new_n12243_,
    new_n12244_, new_n12245_, new_n12246_, new_n12247_, new_n12248_,
    new_n12249_, new_n12250_, new_n12251_, new_n12252_, new_n12253_,
    new_n12254_, new_n12255_, new_n12256_, new_n12257_, new_n12258_,
    new_n12259_, new_n12260_, new_n12261_, new_n12262_, new_n12263_,
    new_n12264_, new_n12265_, new_n12266_, new_n12267_, new_n12268_,
    new_n12269_, new_n12270_, new_n12271_, new_n12272_, new_n12273_,
    new_n12274_, new_n12275_, new_n12276_, new_n12277_, new_n12278_,
    new_n12279_, new_n12280_, new_n12281_, new_n12282_, new_n12283_,
    new_n12284_, new_n12285_, new_n12286_, new_n12287_, new_n12288_,
    new_n12289_, new_n12290_, new_n12291_, new_n12292_, new_n12293_,
    new_n12294_, new_n12295_, new_n12296_, new_n12297_, new_n12298_,
    new_n12299_, new_n12300_, new_n12301_, new_n12302_, new_n12303_,
    new_n12304_, new_n12305_, new_n12306_, new_n12307_, new_n12308_,
    new_n12309_, new_n12310_, new_n12311_, new_n12312_, new_n12313_,
    new_n12314_, new_n12315_, new_n12316_, new_n12317_, new_n12318_,
    new_n12319_, new_n12320_, new_n12321_, new_n12322_, new_n12323_,
    new_n12324_, new_n12325_, new_n12326_, new_n12327_, new_n12328_,
    new_n12329_, new_n12330_, new_n12331_, new_n12332_, new_n12333_,
    new_n12334_, new_n12335_, new_n12336_, new_n12337_, new_n12338_,
    new_n12339_, new_n12340_, new_n12341_, new_n12342_, new_n12343_,
    new_n12344_, new_n12345_, new_n12346_, new_n12347_, new_n12348_,
    new_n12349_, new_n12350_, new_n12351_, new_n12352_, new_n12353_,
    new_n12354_, new_n12355_, new_n12356_, new_n12357_, new_n12358_,
    new_n12359_, new_n12360_, new_n12361_, new_n12362_, new_n12363_,
    new_n12364_, new_n12365_, new_n12366_, new_n12367_, new_n12368_,
    new_n12369_, new_n12370_, new_n12371_, new_n12372_, new_n12373_,
    new_n12374_, new_n12375_, new_n12376_, new_n12377_, new_n12378_,
    new_n12379_, new_n12380_, new_n12381_, new_n12382_, new_n12383_,
    new_n12384_, new_n12385_, new_n12386_, new_n12387_, new_n12388_,
    new_n12389_, new_n12390_, new_n12391_, new_n12392_, new_n12393_,
    new_n12394_, new_n12395_, new_n12396_, new_n12397_, new_n12398_,
    new_n12399_, new_n12400_, new_n12401_, new_n12402_, new_n12403_,
    new_n12404_, new_n12405_, new_n12406_, new_n12407_, new_n12408_,
    new_n12409_, new_n12410_, new_n12411_, new_n12412_, new_n12413_,
    new_n12414_, new_n12415_, new_n12416_, new_n12417_, new_n12418_,
    new_n12419_, new_n12420_, new_n12421_, new_n12422_, new_n12423_,
    new_n12424_, new_n12425_, new_n12426_, new_n12427_, new_n12428_,
    new_n12429_, new_n12430_, new_n12431_, new_n12432_, new_n12433_,
    new_n12434_, new_n12435_, new_n12436_, new_n12437_, new_n12438_,
    new_n12439_, new_n12440_, new_n12441_, new_n12442_, new_n12443_,
    new_n12444_, new_n12445_, new_n12446_, new_n12447_, new_n12448_,
    new_n12449_, new_n12450_, new_n12451_, new_n12452_, new_n12453_,
    new_n12454_, new_n12455_, new_n12456_, new_n12457_, new_n12458_,
    new_n12459_, new_n12460_, new_n12461_, new_n12462_, new_n12463_,
    new_n12464_, new_n12465_, new_n12466_, new_n12467_, new_n12468_,
    new_n12469_, new_n12470_, new_n12471_, new_n12472_, new_n12473_,
    new_n12474_, new_n12475_, new_n12476_, new_n12477_, new_n12478_,
    new_n12479_, new_n12480_, new_n12481_, new_n12482_, new_n12483_,
    new_n12484_, new_n12485_, new_n12486_, new_n12487_, new_n12488_,
    new_n12489_, new_n12490_, new_n12491_, new_n12492_, new_n12493_,
    new_n12494_, new_n12495_, new_n12496_, new_n12497_, new_n12498_,
    new_n12499_, new_n12500_, new_n12501_, new_n12502_, new_n12503_,
    new_n12504_, new_n12505_, new_n12506_, new_n12507_, new_n12508_,
    new_n12509_, new_n12510_, new_n12511_, new_n12512_, new_n12513_,
    new_n12514_, new_n12515_, new_n12516_, new_n12517_, new_n12518_,
    new_n12519_, new_n12520_, new_n12521_, new_n12522_, new_n12523_,
    new_n12524_, new_n12525_, new_n12526_, new_n12527_, new_n12528_,
    new_n12529_, new_n12530_, new_n12531_, new_n12532_, new_n12533_,
    new_n12534_, new_n12535_, new_n12536_, new_n12537_, new_n12538_,
    new_n12539_, new_n12540_, new_n12541_, new_n12542_, new_n12543_,
    new_n12544_, new_n12545_, new_n12546_, new_n12547_, new_n12548_,
    new_n12549_, new_n12550_, new_n12551_, new_n12552_, new_n12553_,
    new_n12554_, new_n12555_, new_n12556_, new_n12557_, new_n12558_,
    new_n12559_, new_n12560_, new_n12561_, new_n12562_, new_n12563_,
    new_n12564_, new_n12565_, new_n12566_, new_n12567_, new_n12568_,
    new_n12569_, new_n12570_, new_n12571_, new_n12572_, new_n12573_,
    new_n12574_, new_n12575_, new_n12576_, new_n12577_, new_n12578_,
    new_n12579_, new_n12580_, new_n12581_, new_n12582_, new_n12583_,
    new_n12584_, new_n12585_, new_n12586_, new_n12587_, new_n12588_,
    new_n12589_, new_n12590_, new_n12591_, new_n12592_, new_n12593_,
    new_n12594_, new_n12595_, new_n12596_, new_n12597_, new_n12598_,
    new_n12599_, new_n12600_, new_n12601_, new_n12602_, new_n12603_,
    new_n12604_, new_n12605_, new_n12606_, new_n12607_, new_n12608_,
    new_n12609_, new_n12610_, new_n12611_, new_n12612_, new_n12613_,
    new_n12614_, new_n12615_, new_n12616_, new_n12617_, new_n12618_,
    new_n12619_, new_n12620_, new_n12621_, new_n12622_, new_n12623_,
    new_n12624_, new_n12625_, new_n12626_, new_n12627_, new_n12628_,
    new_n12629_, new_n12630_, new_n12631_, new_n12632_, new_n12633_,
    new_n12634_, new_n12635_, new_n12636_, new_n12637_, new_n12638_,
    new_n12639_, new_n12640_, new_n12641_, new_n12642_, new_n12643_,
    new_n12644_, new_n12645_, new_n12646_, new_n12647_, new_n12648_,
    new_n12649_, new_n12650_, new_n12651_, new_n12652_, new_n12653_,
    new_n12654_, new_n12655_, new_n12656_, new_n12657_, new_n12658_,
    new_n12659_, new_n12660_, new_n12661_, new_n12662_, new_n12663_,
    new_n12664_, new_n12665_, new_n12666_, new_n12667_, new_n12668_,
    new_n12669_, new_n12670_, new_n12671_, new_n12672_, new_n12673_,
    new_n12674_, new_n12675_, new_n12676_, new_n12677_, new_n12678_,
    new_n12679_, new_n12680_, new_n12681_, new_n12682_, new_n12683_,
    new_n12684_, new_n12685_, new_n12686_, new_n12687_, new_n12688_,
    new_n12689_, new_n12690_, new_n12691_, new_n12692_, new_n12693_,
    new_n12694_, new_n12695_, new_n12696_, new_n12697_, new_n12698_,
    new_n12699_, new_n12700_, new_n12701_, new_n12702_, new_n12703_,
    new_n12704_, new_n12705_, new_n12706_, new_n12707_, new_n12708_,
    new_n12709_, new_n12710_, new_n12711_, new_n12712_, new_n12713_,
    new_n12714_, new_n12715_, new_n12716_, new_n12717_, new_n12718_,
    new_n12719_, new_n12720_, new_n12721_, new_n12722_, new_n12723_,
    new_n12724_, new_n12725_, new_n12726_, new_n12727_, new_n12728_,
    new_n12729_, new_n12730_, new_n12731_, new_n12732_, new_n12733_,
    new_n12734_, new_n12735_, new_n12736_, new_n12737_, new_n12738_,
    new_n12739_, new_n12740_, new_n12741_, new_n12742_, new_n12743_,
    new_n12744_, new_n12745_, new_n12746_, new_n12747_, new_n12748_,
    new_n12749_, new_n12750_, new_n12751_, new_n12752_, new_n12753_,
    new_n12754_, new_n12755_, new_n12756_, new_n12757_, new_n12758_,
    new_n12759_, new_n12760_, new_n12761_, new_n12762_, new_n12763_,
    new_n12764_, new_n12765_, new_n12766_, new_n12767_, new_n12768_,
    new_n12769_, new_n12770_, new_n12771_, new_n12772_, new_n12773_,
    new_n12774_, new_n12775_, new_n12776_, new_n12777_, new_n12778_,
    new_n12779_, new_n12780_, new_n12781_, new_n12782_, new_n12783_,
    new_n12784_, new_n12785_, new_n12786_, new_n12787_, new_n12788_,
    new_n12789_, new_n12790_, new_n12791_, new_n12792_, new_n12793_,
    new_n12794_, new_n12795_, new_n12796_, new_n12797_, new_n12798_,
    new_n12799_, new_n12800_, new_n12801_, new_n12802_, new_n12803_,
    new_n12804_, new_n12805_, new_n12806_, new_n12807_, new_n12808_,
    new_n12809_, new_n12810_, new_n12811_, new_n12812_, new_n12813_,
    new_n12814_, new_n12815_, new_n12816_, new_n12817_, new_n12818_,
    new_n12819_, new_n12820_, new_n12821_, new_n12822_, new_n12823_,
    new_n12824_, new_n12825_, new_n12826_, new_n12827_, new_n12828_,
    new_n12829_, new_n12830_, new_n12831_, new_n12832_, new_n12833_,
    new_n12834_, new_n12835_, new_n12836_, new_n12837_, new_n12838_,
    new_n12839_, new_n12840_, new_n12841_, new_n12842_, new_n12843_,
    new_n12844_, new_n12845_, new_n12846_, new_n12847_, new_n12848_,
    new_n12849_, new_n12850_, new_n12851_, new_n12852_, new_n12853_,
    new_n12854_, new_n12855_, new_n12856_, new_n12857_, new_n12858_,
    new_n12859_, new_n12860_, new_n12861_, new_n12862_, new_n12863_,
    new_n12864_, new_n12865_, new_n12866_, new_n12867_, new_n12868_,
    new_n12869_, new_n12870_, new_n12871_, new_n12872_, new_n12873_,
    new_n12874_, new_n12875_, new_n12876_, new_n12877_, new_n12878_,
    new_n12879_, new_n12880_, new_n12881_, new_n12882_, new_n12883_,
    new_n12884_, new_n12885_, new_n12886_, new_n12887_, new_n12888_,
    new_n12889_, new_n12890_, new_n12891_, new_n12892_, new_n12893_,
    new_n12894_, new_n12895_, new_n12896_, new_n12897_, new_n12898_,
    new_n12899_, new_n12901_, new_n12902_, new_n12903_, new_n12904_,
    new_n12905_, new_n12906_, new_n12907_, new_n12908_, new_n12909_,
    new_n12910_, new_n12911_, new_n12912_, new_n12913_, new_n12914_,
    new_n12915_, new_n12916_, new_n12917_, new_n12918_, new_n12919_,
    new_n12920_, new_n12921_, new_n12922_, new_n12923_, new_n12924_,
    new_n12925_, new_n12926_, new_n12927_, new_n12928_, new_n12929_,
    new_n12930_, new_n12931_, new_n12932_, new_n12933_, new_n12934_,
    new_n12935_, new_n12936_, new_n12937_, new_n12938_, new_n12939_,
    new_n12940_, new_n12941_, new_n12942_, new_n12943_, new_n12944_,
    new_n12945_, new_n12946_, new_n12947_, new_n12948_, new_n12949_,
    new_n12950_, new_n12951_, new_n12952_, new_n12953_, new_n12954_,
    new_n12955_, new_n12956_, new_n12957_, new_n12958_, new_n12959_,
    new_n12960_, new_n12961_, new_n12962_, new_n12963_, new_n12964_,
    new_n12965_, new_n12966_, new_n12967_, new_n12968_, new_n12969_,
    new_n12970_, new_n12971_, new_n12972_, new_n12973_, new_n12974_,
    new_n12975_, new_n12976_, new_n12977_, new_n12978_, new_n12979_,
    new_n12980_, new_n12981_, new_n12982_, new_n12983_, new_n12984_,
    new_n12985_, new_n12986_, new_n12987_, new_n12988_, new_n12989_,
    new_n12990_, new_n12991_, new_n12992_, new_n12993_, new_n12994_,
    new_n12995_, new_n12996_, new_n12997_, new_n12998_, new_n12999_,
    new_n13000_, new_n13001_, new_n13002_, new_n13003_, new_n13004_,
    new_n13005_, new_n13006_, new_n13007_, new_n13008_, new_n13009_,
    new_n13010_, new_n13011_, new_n13012_, new_n13013_, new_n13014_,
    new_n13015_, new_n13016_, new_n13017_, new_n13018_, new_n13019_,
    new_n13020_, new_n13021_, new_n13022_, new_n13023_, new_n13024_,
    new_n13025_, new_n13026_, new_n13027_, new_n13028_, new_n13029_,
    new_n13030_, new_n13031_, new_n13032_, new_n13033_, new_n13034_,
    new_n13035_, new_n13036_, new_n13037_, new_n13038_, new_n13039_,
    new_n13040_, new_n13041_, new_n13042_, new_n13043_, new_n13044_,
    new_n13045_, new_n13046_, new_n13047_, new_n13048_, new_n13049_,
    new_n13050_, new_n13051_, new_n13052_, new_n13053_, new_n13054_,
    new_n13055_, new_n13056_, new_n13057_, new_n13058_, new_n13059_,
    new_n13060_, new_n13061_, new_n13062_, new_n13063_, new_n13064_,
    new_n13065_, new_n13066_, new_n13067_, new_n13068_, new_n13069_,
    new_n13070_, new_n13071_, new_n13072_, new_n13073_, new_n13074_,
    new_n13075_, new_n13076_, new_n13077_, new_n13078_, new_n13079_,
    new_n13080_, new_n13081_, new_n13082_, new_n13083_, new_n13084_,
    new_n13085_, new_n13086_, new_n13087_, new_n13088_, new_n13089_,
    new_n13090_, new_n13091_, new_n13092_, new_n13093_, new_n13094_,
    new_n13095_, new_n13096_, new_n13097_, new_n13098_, new_n13099_,
    new_n13100_, new_n13101_, new_n13102_, new_n13103_, new_n13104_,
    new_n13105_, new_n13106_, new_n13107_, new_n13108_, new_n13109_,
    new_n13110_, new_n13111_, new_n13112_, new_n13113_, new_n13114_,
    new_n13115_, new_n13116_, new_n13117_, new_n13118_, new_n13119_,
    new_n13120_, new_n13121_, new_n13122_, new_n13123_, new_n13124_,
    new_n13125_, new_n13126_, new_n13127_, new_n13128_, new_n13129_,
    new_n13130_, new_n13131_, new_n13132_, new_n13133_, new_n13134_,
    new_n13135_, new_n13136_, new_n13137_, new_n13138_, new_n13139_,
    new_n13140_, new_n13141_, new_n13142_, new_n13143_, new_n13144_,
    new_n13145_, new_n13146_, new_n13147_, new_n13148_, new_n13149_,
    new_n13150_, new_n13151_, new_n13152_, new_n13153_, new_n13154_,
    new_n13155_, new_n13156_, new_n13157_, new_n13158_, new_n13159_,
    new_n13160_, new_n13161_, new_n13162_, new_n13163_, new_n13164_,
    new_n13165_, new_n13166_, new_n13167_, new_n13168_, new_n13169_,
    new_n13170_, new_n13171_, new_n13172_, new_n13173_, new_n13174_,
    new_n13175_, new_n13176_, new_n13177_, new_n13178_, new_n13179_,
    new_n13180_, new_n13181_, new_n13182_, new_n13183_, new_n13184_,
    new_n13185_, new_n13186_, new_n13187_, new_n13188_, new_n13189_,
    new_n13190_, new_n13191_, new_n13192_, new_n13193_, new_n13194_,
    new_n13195_, new_n13196_, new_n13197_, new_n13198_, new_n13199_,
    new_n13200_, new_n13201_, new_n13202_, new_n13203_, new_n13204_,
    new_n13205_, new_n13206_, new_n13207_, new_n13208_, new_n13209_,
    new_n13210_, new_n13211_, new_n13212_, new_n13213_, new_n13214_,
    new_n13215_, new_n13216_, new_n13217_, new_n13219_, new_n13220_,
    new_n13221_, new_n13222_, new_n13223_, new_n13224_, new_n13225_,
    new_n13226_, new_n13227_, new_n13228_, new_n13229_, new_n13230_,
    new_n13231_, new_n13232_, new_n13233_, new_n13234_, new_n13235_,
    new_n13236_, new_n13237_, new_n13238_, new_n13239_, new_n13240_,
    new_n13241_, new_n13242_, new_n13243_, new_n13244_, new_n13245_,
    new_n13246_, new_n13247_, new_n13248_, new_n13249_, new_n13250_,
    new_n13251_, new_n13252_, new_n13253_, new_n13254_, new_n13255_,
    new_n13256_, new_n13257_, new_n13258_, new_n13259_, new_n13260_,
    new_n13261_, new_n13262_, new_n13263_, new_n13264_, new_n13265_,
    new_n13266_, new_n13267_, new_n13268_, new_n13269_, new_n13270_,
    new_n13271_, new_n13272_, new_n13273_, new_n13274_, new_n13275_,
    new_n13276_, new_n13277_, new_n13278_, new_n13279_, new_n13280_,
    new_n13281_, new_n13282_, new_n13283_, new_n13284_, new_n13285_,
    new_n13286_, new_n13287_, new_n13288_, new_n13289_, new_n13290_,
    new_n13291_, new_n13292_, new_n13293_, new_n13294_, new_n13295_,
    new_n13296_, new_n13297_, new_n13298_, new_n13299_, new_n13300_,
    new_n13301_, new_n13302_, new_n13303_, new_n13304_, new_n13305_,
    new_n13306_, new_n13307_, new_n13308_, new_n13309_, new_n13310_,
    new_n13311_, new_n13312_, new_n13313_, new_n13314_, new_n13315_,
    new_n13316_, new_n13317_, new_n13318_, new_n13319_, new_n13320_,
    new_n13321_, new_n13322_, new_n13323_, new_n13324_, new_n13325_,
    new_n13326_, new_n13327_, new_n13328_, new_n13329_, new_n13330_,
    new_n13331_, new_n13332_, new_n13333_, new_n13334_, new_n13335_,
    new_n13336_, new_n13337_, new_n13338_, new_n13339_, new_n13340_,
    new_n13341_, new_n13342_, new_n13343_, new_n13344_, new_n13345_,
    new_n13346_, new_n13347_, new_n13348_, new_n13349_, new_n13350_,
    new_n13351_, new_n13352_, new_n13353_, new_n13354_, new_n13355_,
    new_n13356_, new_n13357_, new_n13358_, new_n13359_, new_n13360_,
    new_n13361_, new_n13362_, new_n13363_, new_n13364_, new_n13365_,
    new_n13366_, new_n13367_, new_n13368_, new_n13369_, new_n13370_,
    new_n13371_, new_n13372_, new_n13373_, new_n13374_, new_n13375_,
    new_n13376_, new_n13377_, new_n13378_, new_n13379_, new_n13380_,
    new_n13381_, new_n13382_, new_n13383_, new_n13384_, new_n13385_,
    new_n13386_, new_n13387_, new_n13388_, new_n13389_, new_n13390_,
    new_n13391_, new_n13392_, new_n13393_, new_n13394_, new_n13395_,
    new_n13396_, new_n13397_, new_n13398_, new_n13399_, new_n13400_,
    new_n13401_, new_n13402_, new_n13403_, new_n13404_, new_n13405_,
    new_n13406_, new_n13407_, new_n13408_, new_n13409_, new_n13410_,
    new_n13411_, new_n13412_, new_n13413_, new_n13414_, new_n13415_,
    new_n13416_, new_n13417_, new_n13418_, new_n13419_, new_n13420_,
    new_n13421_, new_n13422_, new_n13423_, new_n13424_, new_n13425_,
    new_n13426_, new_n13427_, new_n13428_, new_n13429_, new_n13430_,
    new_n13431_, new_n13432_, new_n13433_, new_n13434_, new_n13435_,
    new_n13436_, new_n13437_, new_n13438_, new_n13439_, new_n13440_,
    new_n13441_, new_n13442_, new_n13443_, new_n13444_, new_n13445_,
    new_n13446_, new_n13447_, new_n13448_, new_n13449_, new_n13450_,
    new_n13451_, new_n13452_, new_n13453_, new_n13454_, new_n13455_,
    new_n13456_, new_n13457_, new_n13458_, new_n13459_, new_n13460_,
    new_n13461_, new_n13462_, new_n13463_, new_n13464_, new_n13465_,
    new_n13466_, new_n13467_, new_n13468_, new_n13469_, new_n13470_,
    new_n13471_, new_n13472_, new_n13473_, new_n13474_, new_n13475_,
    new_n13476_, new_n13477_, new_n13478_, new_n13479_, new_n13480_,
    new_n13481_, new_n13482_, new_n13483_, new_n13484_, new_n13485_,
    new_n13486_, new_n13487_, new_n13488_, new_n13489_, new_n13490_,
    new_n13491_, new_n13492_, new_n13493_, new_n13494_, new_n13495_,
    new_n13496_, new_n13497_, new_n13498_, new_n13499_, new_n13500_,
    new_n13501_, new_n13502_, new_n13503_, new_n13504_, new_n13505_,
    new_n13506_, new_n13507_, new_n13508_, new_n13509_, new_n13510_,
    new_n13511_, new_n13512_, new_n13513_, new_n13514_, new_n13515_,
    new_n13516_, new_n13517_, new_n13518_, new_n13519_, new_n13520_,
    new_n13521_, new_n13522_, new_n13523_, new_n13524_, new_n13525_,
    new_n13526_, new_n13527_, new_n13528_, new_n13529_, new_n13530_,
    new_n13531_, new_n13532_, new_n13533_, new_n13534_, new_n13535_,
    new_n13536_, new_n13537_, new_n13538_, new_n13539_, new_n13540_,
    new_n13541_, new_n13542_, new_n13543_, new_n13544_, new_n13545_,
    new_n13546_, new_n13547_, new_n13548_, new_n13549_, new_n13550_,
    new_n13551_, new_n13552_, new_n13553_, new_n13554_, new_n13555_,
    new_n13556_, new_n13557_, new_n13558_, new_n13559_, new_n13560_,
    new_n13561_, new_n13562_, new_n13563_, new_n13564_, new_n13565_,
    new_n13566_, new_n13567_, new_n13568_, new_n13569_, new_n13570_,
    new_n13571_, new_n13572_, new_n13573_, new_n13574_, new_n13575_,
    new_n13576_, new_n13577_, new_n13578_, new_n13579_, new_n13580_,
    new_n13581_, new_n13582_, new_n13583_, new_n13584_, new_n13585_,
    new_n13586_, new_n13587_, new_n13588_, new_n13589_, new_n13590_,
    new_n13591_, new_n13592_, new_n13593_, new_n13594_, new_n13595_,
    new_n13596_, new_n13597_, new_n13598_, new_n13599_, new_n13600_,
    new_n13601_, new_n13602_, new_n13603_, new_n13604_, new_n13605_,
    new_n13606_, new_n13607_, new_n13608_, new_n13609_, new_n13610_,
    new_n13611_, new_n13612_, new_n13613_, new_n13614_, new_n13615_,
    new_n13616_, new_n13617_, new_n13618_, new_n13619_, new_n13620_,
    new_n13621_, new_n13622_, new_n13623_, new_n13624_, new_n13625_,
    new_n13626_, new_n13627_, new_n13628_, new_n13629_, new_n13630_,
    new_n13631_, new_n13632_, new_n13633_, new_n13634_, new_n13635_,
    new_n13636_, new_n13637_, new_n13638_, new_n13639_, new_n13640_,
    new_n13641_, new_n13642_, new_n13643_, new_n13644_, new_n13645_,
    new_n13646_, new_n13647_, new_n13648_, new_n13649_, new_n13650_,
    new_n13651_, new_n13652_, new_n13653_, new_n13654_, new_n13655_,
    new_n13656_, new_n13657_, new_n13658_, new_n13659_, new_n13660_,
    new_n13661_, new_n13662_, new_n13663_, new_n13664_, new_n13665_,
    new_n13666_, new_n13667_, new_n13669_, new_n13670_, new_n13671_,
    new_n13672_, new_n13673_, new_n13674_, new_n13675_, new_n13676_,
    new_n13677_, new_n13678_, new_n13679_, new_n13680_, new_n13681_,
    new_n13682_, new_n13683_, new_n13684_, new_n13685_, new_n13686_,
    new_n13687_, new_n13688_, new_n13689_, new_n13690_, new_n13691_,
    new_n13692_, new_n13693_, new_n13694_, new_n13695_, new_n13696_,
    new_n13697_, new_n13698_, new_n13699_, new_n13700_, new_n13701_,
    new_n13702_, new_n13703_, new_n13704_, new_n13705_, new_n13706_,
    new_n13707_, new_n13708_, new_n13709_, new_n13710_, new_n13711_,
    new_n13712_, new_n13713_, new_n13714_, new_n13715_, new_n13716_,
    new_n13717_, new_n13718_, new_n13719_, new_n13720_, new_n13721_,
    new_n13722_, new_n13723_, new_n13724_, new_n13725_, new_n13726_,
    new_n13727_, new_n13728_, new_n13729_, new_n13730_, new_n13731_,
    new_n13732_, new_n13733_, new_n13734_, new_n13735_, new_n13736_,
    new_n13737_, new_n13738_, new_n13739_, new_n13740_, new_n13741_,
    new_n13742_, new_n13743_, new_n13744_, new_n13745_, new_n13746_,
    new_n13747_, new_n13748_, new_n13749_, new_n13750_, new_n13751_,
    new_n13752_, new_n13753_, new_n13754_, new_n13755_, new_n13756_,
    new_n13757_, new_n13758_, new_n13759_, new_n13760_, new_n13761_,
    new_n13762_, new_n13763_, new_n13764_, new_n13765_, new_n13766_,
    new_n13767_, new_n13768_, new_n13769_, new_n13770_, new_n13771_,
    new_n13772_, new_n13773_, new_n13774_, new_n13775_, new_n13776_,
    new_n13777_, new_n13778_, new_n13779_, new_n13780_, new_n13781_,
    new_n13782_, new_n13783_, new_n13784_, new_n13785_, new_n13786_,
    new_n13787_, new_n13788_, new_n13789_, new_n13790_, new_n13791_,
    new_n13792_, new_n13793_, new_n13794_, new_n13795_, new_n13796_,
    new_n13797_, new_n13798_, new_n13799_, new_n13800_, new_n13801_,
    new_n13802_, new_n13803_, new_n13804_, new_n13805_, new_n13806_,
    new_n13807_, new_n13808_, new_n13809_, new_n13810_, new_n13811_,
    new_n13812_, new_n13813_, new_n13814_, new_n13815_, new_n13816_,
    new_n13817_, new_n13818_, new_n13819_, new_n13820_, new_n13821_,
    new_n13822_, new_n13823_, new_n13824_, new_n13825_, new_n13826_,
    new_n13827_, new_n13828_, new_n13829_, new_n13830_, new_n13831_,
    new_n13832_, new_n13833_, new_n13834_, new_n13835_, new_n13836_,
    new_n13837_, new_n13838_, new_n13839_, new_n13840_, new_n13841_,
    new_n13842_, new_n13843_, new_n13844_, new_n13845_, new_n13846_,
    new_n13847_, new_n13848_, new_n13849_, new_n13850_, new_n13851_,
    new_n13852_, new_n13853_, new_n13854_, new_n13855_, new_n13856_,
    new_n13857_, new_n13858_, new_n13859_, new_n13860_, new_n13861_,
    new_n13862_, new_n13863_, new_n13864_, new_n13865_, new_n13866_,
    new_n13867_, new_n13868_, new_n13869_, new_n13870_, new_n13871_,
    new_n13872_, new_n13873_, new_n13874_, new_n13875_, new_n13876_,
    new_n13877_, new_n13878_, new_n13879_, new_n13880_, new_n13881_,
    new_n13882_, new_n13883_, new_n13884_, new_n13885_, new_n13886_,
    new_n13887_, new_n13888_, new_n13889_, new_n13890_, new_n13891_,
    new_n13892_, new_n13893_, new_n13894_, new_n13895_, new_n13896_,
    new_n13897_, new_n13898_, new_n13899_, new_n13900_, new_n13901_,
    new_n13902_, new_n13903_, new_n13904_, new_n13905_, new_n13906_,
    new_n13907_, new_n13908_, new_n13909_, new_n13910_, new_n13911_,
    new_n13912_, new_n13913_, new_n13914_, new_n13915_, new_n13916_,
    new_n13917_, new_n13918_, new_n13919_, new_n13920_, new_n13921_,
    new_n13922_, new_n13923_, new_n13924_, new_n13925_, new_n13926_,
    new_n13927_, new_n13928_, new_n13929_, new_n13930_, new_n13931_,
    new_n13932_, new_n13933_, new_n13934_, new_n13935_, new_n13936_,
    new_n13937_, new_n13938_, new_n13939_, new_n13940_, new_n13941_,
    new_n13942_, new_n13943_, new_n13944_, new_n13945_, new_n13946_,
    new_n13947_, new_n13948_, new_n13949_, new_n13950_, new_n13951_,
    new_n13952_, new_n13953_, new_n13954_, new_n13955_, new_n13956_,
    new_n13957_, new_n13958_, new_n13959_, new_n13960_, new_n13961_,
    new_n13962_, new_n13963_, new_n13964_, new_n13965_, new_n13966_,
    new_n13967_, new_n13969_, new_n13970_, new_n13971_, new_n13972_,
    new_n13973_, new_n13974_, new_n13975_, new_n13976_, new_n13977_,
    new_n13978_, new_n13979_, new_n13980_, new_n13981_, new_n13982_,
    new_n13983_, new_n13984_, new_n13985_, new_n13986_, new_n13987_,
    new_n13988_, new_n13989_, new_n13990_, new_n13991_, new_n13992_,
    new_n13993_, new_n13994_, new_n13995_, new_n13996_, new_n13997_,
    new_n13998_, new_n13999_, new_n14000_, new_n14001_, new_n14002_,
    new_n14003_, new_n14004_, new_n14005_, new_n14006_, new_n14007_,
    new_n14008_, new_n14009_, new_n14010_, new_n14011_, new_n14012_,
    new_n14013_, new_n14014_, new_n14015_, new_n14016_, new_n14017_,
    new_n14018_, new_n14019_, new_n14020_, new_n14021_, new_n14022_,
    new_n14023_, new_n14024_, new_n14025_, new_n14026_, new_n14027_,
    new_n14028_, new_n14029_, new_n14030_, new_n14031_, new_n14032_,
    new_n14033_, new_n14034_, new_n14035_, new_n14036_, new_n14037_,
    new_n14038_, new_n14039_, new_n14040_, new_n14041_, new_n14042_,
    new_n14043_, new_n14044_, new_n14045_, new_n14046_, new_n14047_,
    new_n14048_, new_n14049_, new_n14050_, new_n14051_, new_n14052_,
    new_n14053_, new_n14054_, new_n14055_, new_n14056_, new_n14057_,
    new_n14058_, new_n14059_, new_n14060_, new_n14061_, new_n14062_,
    new_n14063_, new_n14064_, new_n14065_, new_n14066_, new_n14067_,
    new_n14068_, new_n14069_, new_n14070_, new_n14071_, new_n14072_,
    new_n14073_, new_n14074_, new_n14075_, new_n14076_, new_n14077_,
    new_n14078_, new_n14079_, new_n14080_, new_n14081_, new_n14082_,
    new_n14083_, new_n14084_, new_n14085_, new_n14086_, new_n14087_,
    new_n14088_, new_n14089_, new_n14090_, new_n14091_, new_n14092_,
    new_n14093_, new_n14094_, new_n14095_, new_n14096_, new_n14097_,
    new_n14098_, new_n14099_, new_n14100_, new_n14101_, new_n14102_,
    new_n14103_, new_n14104_, new_n14105_, new_n14106_, new_n14107_,
    new_n14108_, new_n14109_, new_n14110_, new_n14111_, new_n14112_,
    new_n14113_, new_n14114_, new_n14115_, new_n14116_, new_n14117_,
    new_n14118_, new_n14119_, new_n14120_, new_n14121_, new_n14122_,
    new_n14123_, new_n14124_, new_n14125_, new_n14126_, new_n14127_,
    new_n14128_, new_n14129_, new_n14130_, new_n14131_, new_n14132_,
    new_n14133_, new_n14134_, new_n14135_, new_n14136_, new_n14137_,
    new_n14138_, new_n14139_, new_n14140_, new_n14141_, new_n14142_,
    new_n14143_, new_n14144_, new_n14145_, new_n14146_, new_n14147_,
    new_n14148_, new_n14149_, new_n14150_, new_n14151_, new_n14152_,
    new_n14153_, new_n14154_, new_n14155_, new_n14156_, new_n14157_,
    new_n14158_, new_n14159_, new_n14160_, new_n14161_, new_n14162_,
    new_n14163_, new_n14164_, new_n14165_, new_n14166_, new_n14167_,
    new_n14168_, new_n14169_, new_n14170_, new_n14171_, new_n14172_,
    new_n14173_, new_n14174_, new_n14175_, new_n14176_, new_n14177_,
    new_n14178_, new_n14179_, new_n14180_, new_n14181_, new_n14182_,
    new_n14183_, new_n14184_, new_n14185_, new_n14186_, new_n14187_,
    new_n14188_, new_n14189_, new_n14190_, new_n14191_, new_n14192_,
    new_n14193_, new_n14194_, new_n14195_, new_n14196_, new_n14197_,
    new_n14198_, new_n14199_, new_n14200_, new_n14201_, new_n14202_,
    new_n14203_, new_n14204_, new_n14205_, new_n14206_, new_n14207_,
    new_n14208_, new_n14209_, new_n14210_, new_n14211_, new_n14212_,
    new_n14213_, new_n14214_, new_n14215_, new_n14216_, new_n14217_,
    new_n14218_, new_n14219_, new_n14220_, new_n14221_, new_n14222_,
    new_n14223_, new_n14224_, new_n14225_, new_n14226_, new_n14227_,
    new_n14228_, new_n14229_, new_n14230_, new_n14231_, new_n14232_,
    new_n14233_, new_n14234_, new_n14235_, new_n14236_, new_n14237_,
    new_n14238_, new_n14239_, new_n14240_, new_n14241_, new_n14242_,
    new_n14243_, new_n14244_, new_n14245_, new_n14246_, new_n14247_,
    new_n14248_, new_n14249_, new_n14250_, new_n14251_, new_n14252_,
    new_n14253_, new_n14254_, new_n14255_, new_n14256_, new_n14257_,
    new_n14258_, new_n14259_, new_n14260_, new_n14261_, new_n14262_,
    new_n14263_, new_n14264_, new_n14265_, new_n14266_, new_n14267_,
    new_n14268_, new_n14269_, new_n14270_, new_n14271_, new_n14272_,
    new_n14273_, new_n14274_, new_n14275_, new_n14276_, new_n14277_,
    new_n14278_, new_n14279_, new_n14280_, new_n14281_, new_n14282_,
    new_n14283_, new_n14284_, new_n14285_, new_n14286_, new_n14287_,
    new_n14288_, new_n14289_, new_n14290_, new_n14291_, new_n14292_,
    new_n14293_, new_n14294_, new_n14295_, new_n14296_, new_n14297_,
    new_n14298_, new_n14299_, new_n14300_, new_n14301_, new_n14303_,
    new_n14304_, new_n14305_, new_n14306_, new_n14307_, new_n14308_,
    new_n14309_, new_n14310_, new_n14311_, new_n14312_, new_n14313_,
    new_n14314_, new_n14315_, new_n14316_, new_n14317_, new_n14318_,
    new_n14319_, new_n14320_, new_n14321_, new_n14322_, new_n14323_,
    new_n14324_, new_n14325_, new_n14326_, new_n14327_, new_n14328_,
    new_n14329_, new_n14330_, new_n14331_, new_n14332_, new_n14333_,
    new_n14334_, new_n14335_, new_n14336_, new_n14337_, new_n14338_,
    new_n14339_, new_n14340_, new_n14341_, new_n14342_, new_n14343_,
    new_n14344_, new_n14345_, new_n14346_, new_n14347_, new_n14348_,
    new_n14349_, new_n14350_, new_n14351_, new_n14352_, new_n14353_,
    new_n14354_, new_n14355_, new_n14356_, new_n14357_, new_n14358_,
    new_n14359_, new_n14360_, new_n14361_, new_n14362_, new_n14363_,
    new_n14364_, new_n14365_, new_n14366_, new_n14367_, new_n14368_,
    new_n14369_, new_n14370_, new_n14371_, new_n14372_, new_n14373_,
    new_n14374_, new_n14375_, new_n14376_, new_n14377_, new_n14378_,
    new_n14379_, new_n14380_, new_n14381_, new_n14382_, new_n14383_,
    new_n14384_, new_n14385_, new_n14386_, new_n14387_, new_n14388_,
    new_n14389_, new_n14390_, new_n14391_, new_n14392_, new_n14393_,
    new_n14394_, new_n14395_, new_n14396_, new_n14397_, new_n14398_,
    new_n14399_, new_n14400_, new_n14401_, new_n14402_, new_n14403_,
    new_n14404_, new_n14405_, new_n14406_, new_n14407_, new_n14408_,
    new_n14409_, new_n14410_, new_n14411_, new_n14412_, new_n14413_,
    new_n14414_, new_n14415_, new_n14416_, new_n14417_, new_n14418_,
    new_n14419_, new_n14420_, new_n14421_, new_n14422_, new_n14423_,
    new_n14424_, new_n14425_, new_n14426_, new_n14427_, new_n14428_,
    new_n14429_, new_n14430_, new_n14431_, new_n14432_, new_n14433_,
    new_n14434_, new_n14435_, new_n14436_, new_n14437_, new_n14438_,
    new_n14439_, new_n14440_, new_n14441_, new_n14442_, new_n14443_,
    new_n14444_, new_n14445_, new_n14446_, new_n14447_, new_n14448_,
    new_n14449_, new_n14450_, new_n14451_, new_n14452_, new_n14453_,
    new_n14454_, new_n14455_, new_n14456_, new_n14457_, new_n14458_,
    new_n14459_, new_n14460_, new_n14461_, new_n14462_, new_n14463_,
    new_n14464_, new_n14465_, new_n14466_, new_n14467_, new_n14468_,
    new_n14469_, new_n14470_, new_n14471_, new_n14472_, new_n14473_,
    new_n14474_, new_n14475_, new_n14476_, new_n14477_, new_n14478_,
    new_n14479_, new_n14480_, new_n14481_, new_n14482_, new_n14483_,
    new_n14484_, new_n14485_, new_n14486_, new_n14487_, new_n14488_,
    new_n14489_, new_n14490_, new_n14491_, new_n14492_, new_n14493_,
    new_n14494_, new_n14495_, new_n14496_, new_n14497_, new_n14498_,
    new_n14499_, new_n14500_, new_n14501_, new_n14502_, new_n14503_,
    new_n14504_, new_n14505_, new_n14506_, new_n14507_, new_n14508_,
    new_n14509_, new_n14510_, new_n14511_, new_n14512_, new_n14513_,
    new_n14514_, new_n14515_, new_n14516_, new_n14517_, new_n14518_,
    new_n14519_, new_n14520_, new_n14521_, new_n14522_, new_n14523_,
    new_n14524_, new_n14525_, new_n14526_, new_n14527_, new_n14528_,
    new_n14529_, new_n14530_, new_n14531_, new_n14532_, new_n14533_,
    new_n14534_, new_n14535_, new_n14536_, new_n14537_, new_n14538_,
    new_n14539_, new_n14540_, new_n14541_, new_n14542_, new_n14543_,
    new_n14544_, new_n14545_, new_n14546_, new_n14547_, new_n14548_,
    new_n14549_, new_n14550_, new_n14551_, new_n14552_, new_n14553_,
    new_n14554_, new_n14555_, new_n14556_, new_n14557_, new_n14558_,
    new_n14559_, new_n14560_, new_n14561_, new_n14562_, new_n14563_,
    new_n14564_, new_n14565_, new_n14566_, new_n14567_, new_n14568_,
    new_n14569_, new_n14570_, new_n14571_, new_n14572_, new_n14573_,
    new_n14574_, new_n14575_, new_n14576_, new_n14577_, new_n14578_,
    new_n14579_, new_n14580_, new_n14581_, new_n14582_, new_n14583_,
    new_n14584_, new_n14585_, new_n14586_, new_n14587_, new_n14588_,
    new_n14590_, new_n14591_, new_n14592_, new_n14593_, new_n14594_,
    new_n14595_, new_n14596_, new_n14597_, new_n14598_, new_n14599_,
    new_n14600_, new_n14601_, new_n14602_, new_n14603_, new_n14604_,
    new_n14605_, new_n14606_, new_n14607_, new_n14608_, new_n14609_,
    new_n14610_, new_n14611_, new_n14612_, new_n14613_, new_n14614_,
    new_n14615_, new_n14616_, new_n14617_, new_n14618_, new_n14619_,
    new_n14620_, new_n14621_, new_n14622_, new_n14623_, new_n14624_,
    new_n14625_, new_n14626_, new_n14627_, new_n14628_, new_n14629_,
    new_n14630_, new_n14631_, new_n14632_, new_n14633_, new_n14634_,
    new_n14635_, new_n14637_, new_n14638_, new_n14639_, new_n14640_,
    new_n14641_, new_n14642_, new_n14643_, new_n14644_, new_n14645_,
    new_n14646_, new_n14647_, new_n14648_, new_n14649_, new_n14650_,
    new_n14651_, new_n14652_, new_n14653_, new_n14654_, new_n14655_,
    new_n14656_, new_n14657_, new_n14658_, new_n14659_, new_n14660_,
    new_n14661_, new_n14662_, new_n14663_, new_n14664_, new_n14665_,
    new_n14666_, new_n14667_, new_n14668_, new_n14669_, new_n14670_,
    new_n14671_, new_n14672_, new_n14673_, new_n14674_, new_n14675_,
    new_n14676_, new_n14677_, new_n14678_, new_n14679_, new_n14680_,
    new_n14681_, new_n14682_, new_n14683_, new_n14684_, new_n14685_,
    new_n14686_, new_n14687_, new_n14688_, new_n14689_, new_n14690_,
    new_n14691_, new_n14692_, new_n14693_, new_n14694_, new_n14695_,
    new_n14696_, new_n14697_, new_n14698_, new_n14699_, new_n14700_,
    new_n14701_, new_n14702_, new_n14703_, new_n14704_, new_n14705_,
    new_n14706_, new_n14707_, new_n14708_, new_n14709_, new_n14710_,
    new_n14711_, new_n14712_, new_n14713_, new_n14714_, new_n14715_,
    new_n14716_, new_n14717_, new_n14718_, new_n14719_, new_n14720_,
    new_n14721_, new_n14722_, new_n14723_, new_n14724_, new_n14725_,
    new_n14726_, new_n14727_, new_n14728_, new_n14729_, new_n14730_,
    new_n14731_, new_n14732_, new_n14733_, new_n14734_, new_n14735_,
    new_n14736_, new_n14737_, new_n14738_, new_n14740_, new_n14741_,
    new_n14742_, new_n14743_, new_n14744_, new_n14745_, new_n14746_,
    new_n14747_, new_n14748_, new_n14749_, new_n14750_, new_n14751_,
    new_n14752_, new_n14753_, new_n14754_, new_n14755_, new_n14756_,
    new_n14757_, new_n14758_, new_n14759_, new_n14760_, new_n14761_,
    new_n14762_, new_n14763_, new_n14764_, new_n14765_, new_n14766_,
    new_n14767_, new_n14768_, new_n14769_, new_n14770_, new_n14771_,
    new_n14772_, new_n14773_, new_n14774_, new_n14775_, new_n14776_,
    new_n14777_, new_n14778_, new_n14779_, new_n14780_, new_n14782_,
    new_n14783_, new_n14784_, new_n14785_, new_n14786_, new_n14787_,
    new_n14788_, new_n14789_, new_n14790_, new_n14791_, new_n14792_,
    new_n14793_, new_n14794_, new_n14795_, new_n14796_, new_n14797_,
    new_n14798_, new_n14799_, new_n14800_, new_n14801_, new_n14802_,
    new_n14803_, new_n14804_, new_n14805_, new_n14806_, new_n14807_,
    new_n14808_, new_n14809_, new_n14810_, new_n14811_, new_n14812_,
    new_n14813_, new_n14814_, new_n14815_, new_n14816_, new_n14817_,
    new_n14819_, new_n14820_, new_n14821_, new_n14822_, new_n14823_,
    new_n14824_, new_n14825_, new_n14826_, new_n14827_, new_n14828_,
    new_n14829_, new_n14830_, new_n14831_, new_n14832_, new_n14833_,
    new_n14834_, new_n14835_, new_n14836_, new_n14837_, new_n14838_,
    new_n14839_, new_n14840_, new_n14841_, new_n14842_, new_n14843_,
    new_n14844_, new_n14845_, new_n14846_, new_n14847_, new_n14848_,
    new_n14849_, new_n14850_, new_n14852_, new_n14853_, new_n14854_,
    new_n14855_, new_n14856_, new_n14857_, new_n14858_, new_n14859_,
    new_n14860_, new_n14861_, new_n14862_, new_n14863_, new_n14864_,
    new_n14865_, new_n14866_, new_n14867_, new_n14868_, new_n14869_,
    new_n14870_, new_n14871_, new_n14872_, new_n14873_, new_n14874_,
    new_n14875_, new_n14876_, new_n14877_, new_n14878_, new_n14879_,
    new_n14880_, new_n14881_, new_n14882_, new_n14883_, new_n14884_,
    new_n14885_, new_n14886_, new_n14887_, new_n14888_, new_n14889_,
    new_n14890_, new_n14891_, new_n14892_, new_n14893_, new_n14894_,
    new_n14895_, new_n14896_, new_n14897_, new_n14898_, new_n14899_,
    new_n14900_, new_n14901_, new_n14902_, new_n14903_, new_n14904_,
    new_n14905_, new_n14906_, new_n14908_, new_n14909_, new_n14910_,
    new_n14911_, new_n14912_, new_n14913_, new_n14914_, new_n14915_,
    new_n14916_, new_n14917_, new_n14918_, new_n14919_, new_n14920_,
    new_n14921_, new_n14922_, new_n14923_, new_n14924_, new_n14925_,
    new_n14926_, new_n14927_, new_n14928_, new_n14929_, new_n14930_,
    new_n14931_, new_n14932_, new_n14933_, new_n14934_, new_n14935_,
    new_n14936_, new_n14937_, new_n14938_, new_n14939_, new_n14940_,
    new_n14941_, new_n14942_, new_n14943_, new_n14944_, new_n14945_,
    new_n14946_, new_n14947_, new_n14948_, new_n14949_, new_n14950_,
    new_n14951_, new_n14952_, new_n14953_, new_n14954_, new_n14955_,
    new_n14956_, new_n14957_, new_n14958_, new_n14959_, new_n14960_,
    new_n14961_, new_n14962_, new_n14963_, new_n14964_, new_n14965_,
    new_n14966_, new_n14967_, new_n14968_, new_n14969_, new_n14970_,
    new_n14971_, new_n14972_, new_n14973_, new_n14974_, new_n14975_,
    new_n14977_, new_n14978_, new_n14979_, new_n14980_, new_n14981_,
    new_n14982_, new_n14983_, new_n14984_, new_n14985_, new_n14986_,
    new_n14987_, new_n14988_, new_n14989_, new_n14990_, new_n14991_,
    new_n14992_, new_n14993_, new_n14994_, new_n14995_, new_n14996_,
    new_n14997_, new_n14998_, new_n14999_, new_n15000_, new_n15001_,
    new_n15002_, new_n15003_, new_n15004_, new_n15005_, new_n15006_,
    new_n15007_, new_n15008_, new_n15009_, new_n15010_, new_n15011_,
    new_n15012_, new_n15013_, new_n15014_, new_n15015_, new_n15016_,
    new_n15017_, new_n15018_, new_n15019_, new_n15020_, new_n15021_,
    new_n15022_, new_n15023_, new_n15024_, new_n15025_, new_n15026_,
    new_n15027_, new_n15028_, new_n15029_, new_n15030_, new_n15032_,
    new_n15033_, new_n15034_, new_n15035_, new_n15036_, new_n15037_,
    new_n15038_, new_n15039_, new_n15040_, new_n15041_, new_n15042_,
    new_n15043_, new_n15044_, new_n15045_, new_n15046_, new_n15047_,
    new_n15048_, new_n15049_, new_n15050_, new_n15051_, new_n15052_,
    new_n15053_, new_n15054_, new_n15055_, new_n15056_, new_n15057_,
    new_n15058_, new_n15059_, new_n15060_, new_n15061_, new_n15062_,
    new_n15064_, new_n15065_, new_n15066_, new_n15067_, new_n15068_,
    new_n15069_, new_n15070_, new_n15071_, new_n15072_, new_n15073_,
    new_n15074_, new_n15075_, new_n15076_, new_n15077_, new_n15078_,
    new_n15079_, new_n15080_, new_n15081_, new_n15082_, new_n15083_,
    new_n15084_, new_n15085_, new_n15086_, new_n15088_, new_n15089_,
    new_n15090_, new_n15091_, new_n15092_, new_n15093_, new_n15094_,
    new_n15095_, new_n15096_, new_n15097_, new_n15098_, new_n15099_,
    new_n15100_, new_n15101_, new_n15102_, new_n15103_, new_n15104_,
    new_n15106_, new_n15107_, new_n15108_, new_n15109_, new_n15110_,
    new_n15111_, new_n15112_, new_n15113_, new_n15114_, new_n15115_,
    new_n15116_, new_n15117_, new_n15118_, new_n15119_, new_n15120_,
    new_n15121_, new_n15122_, new_n15123_, new_n15124_, new_n15125_,
    new_n15126_, new_n15127_, new_n15128_, new_n15129_, new_n15130_,
    new_n15131_, new_n15132_, new_n15133_, new_n15134_, new_n15135_,
    new_n15136_, new_n15137_, new_n15138_, new_n15139_, new_n15141_,
    new_n15142_, new_n15143_, new_n15144_, new_n15145_, new_n15146_,
    new_n15147_, new_n15148_, new_n15149_, new_n15150_, new_n15151_,
    new_n15152_, new_n15153_, new_n15154_, new_n15155_, new_n15156_,
    new_n15157_, new_n15158_, new_n15159_, new_n15160_, new_n15161_,
    new_n15162_, new_n15163_, new_n15164_, new_n15165_, new_n15166_,
    new_n15167_, new_n15168_, new_n15169_, new_n15170_, new_n15172_,
    new_n15173_, new_n15174_, new_n15175_, new_n15176_, new_n15177_,
    new_n15178_, new_n15179_, new_n15180_, new_n15181_, new_n15182_,
    new_n15183_, new_n15184_, new_n15185_, new_n15186_, new_n15187_,
    new_n15188_, new_n15189_, new_n15190_, new_n15191_, new_n15192_,
    new_n15193_, new_n15194_, new_n15195_, new_n15196_, new_n15197_,
    new_n15198_, new_n15199_, new_n15200_, new_n15201_, new_n15203_,
    new_n15204_, new_n15205_, new_n15206_, new_n15207_, new_n15208_,
    new_n15209_, new_n15210_, new_n15211_, new_n15212_, new_n15213_,
    new_n15214_, new_n15215_, new_n15216_, new_n15217_, new_n15218_,
    new_n15219_, new_n15220_, new_n15221_, new_n15222_, new_n15223_,
    new_n15224_, new_n15225_, new_n15226_, new_n15227_, new_n15228_,
    new_n15229_, new_n15230_, new_n15231_, new_n15232_, new_n15233_,
    new_n15234_, new_n15235_, new_n15236_, new_n15238_, new_n15239_,
    new_n15240_, new_n15241_, new_n15242_, new_n15243_, new_n15244_,
    new_n15245_, new_n15246_, new_n15247_, new_n15248_, new_n15249_,
    new_n15250_, new_n15251_, new_n15252_, new_n15253_, new_n15254_,
    new_n15255_, new_n15256_, new_n15257_, new_n15258_, new_n15259_,
    new_n15260_, new_n15261_, new_n15262_, new_n15263_, new_n15264_,
    new_n15265_, new_n15266_, new_n15267_, new_n15268_, new_n15269_,
    new_n15270_, new_n15271_, new_n15272_, new_n15273_, new_n15274_,
    new_n15275_, new_n15276_, new_n15277_, new_n15278_, new_n15279_,
    new_n15280_, new_n15281_, new_n15282_, new_n15283_, new_n15284_,
    new_n15285_, new_n15286_, new_n15287_, new_n15288_, new_n15289_,
    new_n15290_, new_n15291_, new_n15292_, new_n15293_, new_n15294_,
    new_n15296_, new_n15297_, new_n15298_, new_n15299_, new_n15300_,
    new_n15301_, new_n15302_, new_n15303_, new_n15304_, new_n15305_,
    new_n15306_, new_n15307_, new_n15308_, new_n15309_, new_n15310_,
    new_n15311_, new_n15312_, new_n15313_, new_n15314_, new_n15315_,
    new_n15316_, new_n15317_, new_n15318_, new_n15319_, new_n15320_,
    new_n15321_, new_n15322_, new_n15323_, new_n15324_, new_n15325_,
    new_n15326_, new_n15327_, new_n15329_, new_n15330_, new_n15331_,
    new_n15332_, new_n15333_, new_n15334_, new_n15335_, new_n15336_,
    new_n15337_, new_n15338_, new_n15339_, new_n15340_, new_n15341_,
    new_n15342_, new_n15343_, new_n15344_, new_n15345_, new_n15346_,
    new_n15347_, new_n15348_, new_n15349_, new_n15350_, new_n15351_,
    new_n15352_, new_n15353_, new_n15354_, new_n15355_, new_n15356_,
    new_n15357_, new_n15358_, new_n15359_, new_n15360_, new_n15361_,
    new_n15362_, new_n15364_, new_n15365_, new_n15366_, new_n15367_,
    new_n15368_, new_n15369_, new_n15370_, new_n15371_, new_n15372_,
    new_n15373_, new_n15374_, new_n15375_, new_n15376_, new_n15377_,
    new_n15378_, new_n15379_, new_n15380_, new_n15381_, new_n15382_,
    new_n15383_, new_n15384_, new_n15385_, new_n15387_, new_n15388_,
    new_n15389_, new_n15390_, new_n15391_, new_n15392_, new_n15393_,
    new_n15394_, new_n15395_, new_n15396_, new_n15397_, new_n15398_,
    new_n15399_, new_n15400_, new_n15401_, new_n15402_, new_n15403_,
    new_n15404_, new_n15405_, new_n15406_, new_n15408_, new_n15409_,
    new_n15410_, new_n15411_, new_n15412_, new_n15413_, new_n15414_,
    new_n15415_, new_n15416_, new_n15417_, new_n15418_, new_n15419_,
    new_n15420_, new_n15421_, new_n15422_, new_n15423_, new_n15424_,
    new_n15425_, new_n15426_, new_n15427_, new_n15428_, new_n15429_,
    new_n15430_, new_n15431_, new_n15432_, new_n15433_, new_n15434_,
    new_n15435_, new_n15436_, new_n15437_, new_n15438_, new_n15439_,
    new_n15440_, new_n15441_, new_n15442_, new_n15443_, new_n15444_,
    new_n15445_, new_n15446_, new_n15447_, new_n15448_, new_n15449_,
    new_n15450_, new_n15451_, new_n15452_, new_n15453_, new_n15454_,
    new_n15455_, new_n15456_, new_n15457_, new_n15458_, new_n15459_,
    new_n15460_, new_n15461_, new_n15462_, new_n15463_, new_n15464_,
    new_n15465_, new_n15466_, new_n15467_, new_n15468_, new_n15470_,
    new_n15471_, new_n15472_, new_n15473_, new_n15474_, new_n15475_,
    new_n15476_, new_n15477_, new_n15478_, new_n15479_, new_n15480_,
    new_n15481_, new_n15482_, new_n15483_, new_n15484_, new_n15485_,
    new_n15486_, new_n15487_, new_n15488_, new_n15489_, new_n15490_,
    new_n15491_, new_n15492_, new_n15493_, new_n15495_, new_n15496_,
    new_n15497_, new_n15498_, new_n15499_, new_n15500_, new_n15501_,
    new_n15502_, new_n15503_, new_n15504_, new_n15505_, new_n15506_,
    new_n15507_, new_n15508_, new_n15509_, new_n15510_, new_n15511_,
    new_n15512_, new_n15513_, new_n15514_, new_n15515_, new_n15516_,
    new_n15517_, new_n15518_, new_n15519_, new_n15520_, new_n15521_,
    new_n15522_, new_n15523_, new_n15524_, new_n15525_, new_n15526_,
    new_n15527_, new_n15528_, new_n15529_, new_n15530_, new_n15531_,
    new_n15532_, new_n15533_, new_n15534_, new_n15535_, new_n15536_,
    new_n15537_, new_n15538_, new_n15539_, new_n15540_, new_n15541_,
    new_n15542_, new_n15543_, new_n15545_, new_n15546_, new_n15547_,
    new_n15548_, new_n15549_, new_n15550_, new_n15551_, new_n15552_,
    new_n15553_, new_n15554_, new_n15555_, new_n15556_, new_n15557_,
    new_n15558_, new_n15559_, new_n15560_, new_n15561_, new_n15562_,
    new_n15563_, new_n15564_, new_n15565_, new_n15566_, new_n15567_,
    new_n15568_, new_n15569_, new_n15570_, new_n15571_, new_n15572_,
    new_n15573_, new_n15574_, new_n15575_, new_n15576_, new_n15577_,
    new_n15578_, new_n15579_, new_n15580_, new_n15581_, new_n15582_,
    new_n15583_, new_n15584_, new_n15585_, new_n15586_, new_n15587_,
    new_n15588_, new_n15589_, new_n15590_, new_n15591_, new_n15592_,
    new_n15593_, new_n15595_, new_n15596_, new_n15597_, new_n15598_,
    new_n15599_, new_n15600_, new_n15601_, new_n15602_, new_n15603_,
    new_n15604_, new_n15605_, new_n15606_, new_n15607_, new_n15608_,
    new_n15609_, new_n15610_, new_n15611_, new_n15612_, new_n15613_,
    new_n15614_, new_n15615_, new_n15616_, new_n15617_, new_n15618_,
    new_n15619_, new_n15620_, new_n15621_, new_n15622_, new_n15623_,
    new_n15624_, new_n15625_, new_n15626_, new_n15627_, new_n15628_,
    new_n15629_, new_n15630_, new_n15631_, new_n15632_, new_n15633_,
    new_n15634_, new_n15635_, new_n15636_, new_n15637_, new_n15638_,
    new_n15639_, new_n15641_, new_n15642_, new_n15643_, new_n15644_,
    new_n15645_, new_n15646_, new_n15647_, new_n15648_, new_n15649_,
    new_n15650_, new_n15651_, new_n15652_, new_n15653_, new_n15654_,
    new_n15655_, new_n15656_, new_n15657_, new_n15658_, new_n15659_,
    new_n15660_, new_n15661_, new_n15662_, new_n15663_, new_n15664_,
    new_n15665_, new_n15666_, new_n15667_, new_n15668_, new_n15669_,
    new_n15670_, new_n15671_, new_n15672_, new_n15673_, new_n15674_,
    new_n15675_, new_n15676_, new_n15677_, new_n15678_, new_n15679_,
    new_n15680_, new_n15681_, new_n15682_, new_n15683_, new_n15684_,
    new_n15685_, new_n15686_, new_n15687_, new_n15688_, new_n15689_,
    new_n15691_, new_n15692_, new_n15693_, new_n15694_, new_n15695_,
    new_n15696_, new_n15697_, new_n15698_, new_n15699_, new_n15700_,
    new_n15701_, new_n15702_, new_n15703_, new_n15704_, new_n15705_,
    new_n15706_, new_n15707_, new_n15708_, new_n15709_, new_n15710_,
    new_n15711_, new_n15712_, new_n15713_, new_n15714_, new_n15715_,
    new_n15716_, new_n15717_, new_n15718_, new_n15719_, new_n15720_,
    new_n15721_, new_n15722_, new_n15723_, new_n15724_, new_n15725_,
    new_n15726_, new_n15727_, new_n15728_, new_n15729_, new_n15730_,
    new_n15731_, new_n15732_, new_n15733_, new_n15734_, new_n15735_,
    new_n15736_, new_n15737_, new_n15738_, new_n15739_, new_n15740_,
    new_n15742_, new_n15743_, new_n15744_, new_n15745_, new_n15746_,
    new_n15747_, new_n15748_, new_n15749_, new_n15750_, new_n15751_,
    new_n15752_, new_n15753_, new_n15754_, new_n15755_, new_n15756_,
    new_n15757_, new_n15758_, new_n15759_, new_n15760_, new_n15761_,
    new_n15762_, new_n15763_, new_n15764_, new_n15765_, new_n15766_,
    new_n15767_, new_n15768_, new_n15769_, new_n15770_, new_n15771_,
    new_n15772_, new_n15773_, new_n15774_, new_n15775_, new_n15776_,
    new_n15777_, new_n15778_, new_n15779_, new_n15780_, new_n15781_,
    new_n15782_, new_n15783_, new_n15784_, new_n15785_, new_n15786_,
    new_n15787_, new_n15788_, new_n15789_, new_n15790_, new_n15791_,
    new_n15792_, new_n15793_, new_n15794_, new_n15795_, new_n15796_,
    new_n15797_, new_n15798_, new_n15799_, new_n15800_, new_n15801_,
    new_n15802_, new_n15803_, new_n15804_, new_n15805_, new_n15806_,
    new_n15807_, new_n15808_, new_n15809_, new_n15810_, new_n15811_,
    new_n15812_, new_n15813_, new_n15814_, new_n15815_, new_n15816_,
    new_n15817_, new_n15818_, new_n15819_, new_n15820_, new_n15821_,
    new_n15822_, new_n15823_, new_n15824_, new_n15825_, new_n15826_,
    new_n15827_, new_n15828_, new_n15829_, new_n15830_, new_n15831_,
    new_n15832_, new_n15833_, new_n15834_, new_n15835_, new_n15836_,
    new_n15837_, new_n15838_, new_n15839_, new_n15840_, new_n15841_,
    new_n15842_, new_n15843_, new_n15844_, new_n15845_, new_n15846_,
    new_n15847_, new_n15848_, new_n15849_, new_n15850_, new_n15851_,
    new_n15852_, new_n15853_, new_n15854_, new_n15855_, new_n15856_,
    new_n15857_, new_n15858_, new_n15859_, new_n15860_, new_n15861_,
    new_n15862_, new_n15863_, new_n15864_, new_n15865_, new_n15866_,
    new_n15867_, new_n15868_, new_n15869_, new_n15870_, new_n15871_,
    new_n15872_, new_n15873_, new_n15874_, new_n15875_, new_n15876_,
    new_n15877_, new_n15878_, new_n15879_, new_n15880_, new_n15881_,
    new_n15882_, new_n15883_, new_n15884_, new_n15885_, new_n15886_,
    new_n15887_, new_n15888_, new_n15889_, new_n15890_, new_n15891_,
    new_n15892_, new_n15893_, new_n15894_, new_n15895_, new_n15896_,
    new_n15897_, new_n15898_, new_n15899_, new_n15900_, new_n15901_,
    new_n15902_, new_n15903_, new_n15904_, new_n15905_, new_n15906_,
    new_n15907_, new_n15908_, new_n15909_, new_n15910_, new_n15911_,
    new_n15912_, new_n15913_, new_n15914_, new_n15915_, new_n15916_,
    new_n15917_, new_n15918_, new_n15919_, new_n15920_, new_n15921_,
    new_n15922_, new_n15923_, new_n15924_, new_n15925_, new_n15926_,
    new_n15927_, new_n15928_, new_n15929_, new_n15930_, new_n15931_,
    new_n15932_, new_n15933_, new_n15934_, new_n15935_, new_n15936_,
    new_n15937_, new_n15938_, new_n15939_, new_n15940_, new_n15941_,
    new_n15942_, new_n15943_, new_n15944_, new_n15945_, new_n15946_,
    new_n15947_, new_n15948_, new_n15949_, new_n15950_, new_n15951_,
    new_n15952_, new_n15953_, new_n15954_, new_n15955_, new_n15956_,
    new_n15957_, new_n15958_, new_n15959_, new_n15960_, new_n15961_,
    new_n15962_, new_n15963_, new_n15964_, new_n15965_, new_n15966_,
    new_n15967_, new_n15968_, new_n15969_, new_n15970_, new_n15971_,
    new_n15972_, new_n15973_, new_n15974_, new_n15975_, new_n15976_,
    new_n15977_, new_n15978_, new_n15979_, new_n15980_, new_n15981_,
    new_n15982_, new_n15983_, new_n15984_, new_n15985_, new_n15986_,
    new_n15987_, new_n15988_, new_n15989_, new_n15990_, new_n15991_,
    new_n15992_, new_n15993_, new_n15994_, new_n15995_, new_n15996_,
    new_n15997_, new_n15998_, new_n15999_, new_n16000_, new_n16001_,
    new_n16002_, new_n16003_, new_n16004_, new_n16005_, new_n16006_,
    new_n16007_, new_n16008_, new_n16009_, new_n16010_, new_n16011_,
    new_n16012_, new_n16013_, new_n16015_, new_n16016_, new_n16017_,
    new_n16018_, new_n16019_, new_n16020_, new_n16021_, new_n16022_,
    new_n16023_, new_n16024_, new_n16025_, new_n16026_, new_n16027_,
    new_n16028_, new_n16029_, new_n16030_, new_n16031_, new_n16032_,
    new_n16033_, new_n16034_, new_n16035_, new_n16036_, new_n16037_,
    new_n16038_, new_n16039_, new_n16040_, new_n16041_, new_n16042_,
    new_n16043_, new_n16044_, new_n16045_, new_n16046_, new_n16047_,
    new_n16048_, new_n16049_, new_n16050_, new_n16051_, new_n16052_,
    new_n16053_, new_n16054_, new_n16055_, new_n16056_, new_n16057_,
    new_n16058_, new_n16059_, new_n16060_, new_n16061_, new_n16062_,
    new_n16063_, new_n16064_, new_n16065_, new_n16066_, new_n16067_,
    new_n16068_, new_n16069_, new_n16070_, new_n16071_, new_n16072_,
    new_n16073_, new_n16074_, new_n16075_, new_n16076_, new_n16077_,
    new_n16078_, new_n16079_, new_n16080_, new_n16081_, new_n16082_,
    new_n16083_, new_n16084_, new_n16085_, new_n16086_, new_n16087_,
    new_n16088_, new_n16089_, new_n16090_, new_n16091_, new_n16092_,
    new_n16093_, new_n16094_, new_n16095_, new_n16096_, new_n16097_,
    new_n16098_, new_n16099_, new_n16100_, new_n16101_, new_n16102_,
    new_n16103_, new_n16104_, new_n16105_, new_n16106_, new_n16107_,
    new_n16108_, new_n16109_, new_n16110_, new_n16111_, new_n16112_,
    new_n16113_, new_n16114_, new_n16115_, new_n16116_, new_n16117_,
    new_n16118_, new_n16119_, new_n16120_, new_n16121_, new_n16122_,
    new_n16123_, new_n16124_, new_n16125_, new_n16126_, new_n16127_,
    new_n16128_, new_n16129_, new_n16130_, new_n16131_, new_n16132_,
    new_n16133_, new_n16134_, new_n16135_, new_n16136_, new_n16137_,
    new_n16138_, new_n16139_, new_n16140_, new_n16141_, new_n16142_,
    new_n16143_, new_n16144_, new_n16145_, new_n16146_, new_n16147_,
    new_n16148_, new_n16149_, new_n16150_, new_n16151_, new_n16152_,
    new_n16153_, new_n16154_, new_n16155_, new_n16156_, new_n16157_,
    new_n16158_, new_n16159_, new_n16160_, new_n16161_, new_n16162_,
    new_n16163_, new_n16164_, new_n16165_, new_n16166_, new_n16167_,
    new_n16168_, new_n16169_, new_n16170_, new_n16171_, new_n16172_,
    new_n16173_, new_n16174_, new_n16175_, new_n16176_, new_n16177_,
    new_n16178_, new_n16179_, new_n16180_, new_n16181_, new_n16182_,
    new_n16183_, new_n16184_, new_n16185_, new_n16186_, new_n16187_,
    new_n16188_, new_n16189_, new_n16190_, new_n16191_, new_n16192_,
    new_n16193_, new_n16194_, new_n16195_, new_n16196_, new_n16197_,
    new_n16198_, new_n16199_, new_n16200_, new_n16201_, new_n16202_,
    new_n16203_, new_n16204_, new_n16205_, new_n16206_, new_n16207_,
    new_n16208_, new_n16209_, new_n16210_, new_n16211_, new_n16212_,
    new_n16213_, new_n16214_, new_n16215_, new_n16216_, new_n16217_,
    new_n16218_, new_n16219_, new_n16220_, new_n16221_, new_n16222_,
    new_n16223_, new_n16224_, new_n16225_, new_n16226_, new_n16227_,
    new_n16228_, new_n16229_, new_n16230_, new_n16231_, new_n16232_,
    new_n16233_, new_n16234_, new_n16235_, new_n16236_, new_n16237_,
    new_n16238_, new_n16239_, new_n16240_, new_n16241_, new_n16242_,
    new_n16243_, new_n16244_, new_n16245_, new_n16246_, new_n16247_,
    new_n16248_, new_n16249_, new_n16250_, new_n16251_, new_n16252_,
    new_n16253_, new_n16254_, new_n16255_, new_n16256_, new_n16257_,
    new_n16258_, new_n16259_, new_n16260_, new_n16261_, new_n16262_,
    new_n16263_, new_n16264_, new_n16265_, new_n16266_, new_n16267_,
    new_n16268_, new_n16269_, new_n16270_, new_n16271_, new_n16272_,
    new_n16273_, new_n16274_, new_n16275_, new_n16276_, new_n16277_,
    new_n16278_, new_n16279_, new_n16280_, new_n16281_, new_n16282_,
    new_n16283_, new_n16284_, new_n16285_, new_n16286_, new_n16287_,
    new_n16288_, new_n16289_, new_n16290_, new_n16291_, new_n16292_,
    new_n16293_, new_n16294_, new_n16295_, new_n16296_, new_n16297_,
    new_n16298_, new_n16299_, new_n16300_, new_n16301_, new_n16302_,
    new_n16303_, new_n16304_, new_n16305_, new_n16307_, new_n16308_,
    new_n16309_, new_n16310_, new_n16311_, new_n16312_, new_n16313_,
    new_n16314_, new_n16315_, new_n16316_, new_n16317_, new_n16318_,
    new_n16319_, new_n16320_, new_n16321_, new_n16322_, new_n16323_,
    new_n16324_, new_n16325_, new_n16326_, new_n16327_, new_n16328_,
    new_n16329_, new_n16330_, new_n16331_, new_n16332_, new_n16333_,
    new_n16334_, new_n16335_, new_n16336_, new_n16337_, new_n16338_,
    new_n16339_, new_n16340_, new_n16341_, new_n16342_, new_n16343_,
    new_n16344_, new_n16345_, new_n16346_, new_n16347_, new_n16348_,
    new_n16349_, new_n16350_, new_n16351_, new_n16352_, new_n16353_,
    new_n16354_, new_n16355_, new_n16356_, new_n16357_, new_n16358_,
    new_n16359_, new_n16360_, new_n16361_, new_n16362_, new_n16363_,
    new_n16364_, new_n16365_, new_n16366_, new_n16367_, new_n16368_,
    new_n16369_, new_n16370_, new_n16371_, new_n16372_, new_n16373_,
    new_n16374_, new_n16375_, new_n16376_, new_n16377_, new_n16378_,
    new_n16379_, new_n16380_, new_n16381_, new_n16382_, new_n16383_,
    new_n16384_, new_n16385_, new_n16386_, new_n16387_, new_n16388_,
    new_n16389_, new_n16390_, new_n16391_, new_n16392_, new_n16393_,
    new_n16394_, new_n16395_, new_n16396_, new_n16397_, new_n16398_,
    new_n16399_, new_n16400_, new_n16401_, new_n16402_, new_n16403_,
    new_n16404_, new_n16405_, new_n16406_, new_n16407_, new_n16408_,
    new_n16409_, new_n16410_, new_n16411_, new_n16412_, new_n16413_,
    new_n16414_, new_n16415_, new_n16416_, new_n16417_, new_n16418_,
    new_n16419_, new_n16420_, new_n16421_, new_n16422_, new_n16423_,
    new_n16424_, new_n16425_, new_n16426_, new_n16427_, new_n16428_,
    new_n16429_, new_n16430_, new_n16431_, new_n16432_, new_n16433_,
    new_n16434_, new_n16435_, new_n16436_, new_n16437_, new_n16438_,
    new_n16439_, new_n16440_, new_n16441_, new_n16442_, new_n16443_,
    new_n16444_, new_n16445_, new_n16446_, new_n16447_, new_n16448_,
    new_n16449_, new_n16450_, new_n16451_, new_n16452_, new_n16453_,
    new_n16454_, new_n16455_, new_n16456_, new_n16457_, new_n16458_,
    new_n16459_, new_n16460_, new_n16461_, new_n16462_, new_n16463_,
    new_n16464_, new_n16465_, new_n16466_, new_n16467_, new_n16468_,
    new_n16469_, new_n16470_, new_n16471_, new_n16472_, new_n16473_,
    new_n16474_, new_n16475_, new_n16476_, new_n16477_, new_n16478_,
    new_n16479_, new_n16480_, new_n16481_, new_n16482_, new_n16483_,
    new_n16484_, new_n16485_, new_n16486_, new_n16487_, new_n16488_,
    new_n16489_, new_n16490_, new_n16491_, new_n16492_, new_n16493_,
    new_n16494_, new_n16495_, new_n16496_, new_n16497_, new_n16498_,
    new_n16499_, new_n16500_, new_n16501_, new_n16502_, new_n16503_,
    new_n16504_, new_n16505_, new_n16506_, new_n16507_, new_n16508_,
    new_n16509_, new_n16510_, new_n16511_, new_n16512_, new_n16513_,
    new_n16514_, new_n16515_, new_n16516_, new_n16517_, new_n16518_,
    new_n16519_, new_n16520_, new_n16521_, new_n16522_, new_n16523_,
    new_n16524_, new_n16525_, new_n16526_, new_n16527_, new_n16528_,
    new_n16529_, new_n16530_, new_n16531_, new_n16532_, new_n16533_,
    new_n16534_, new_n16535_, new_n16536_, new_n16537_, new_n16538_,
    new_n16539_, new_n16540_, new_n16541_, new_n16542_, new_n16543_,
    new_n16544_, new_n16545_, new_n16546_, new_n16547_, new_n16548_,
    new_n16549_, new_n16550_, new_n16551_, new_n16552_, new_n16553_,
    new_n16554_, new_n16555_, new_n16556_, new_n16557_, new_n16558_,
    new_n16559_, new_n16560_, new_n16561_, new_n16562_, new_n16563_,
    new_n16564_, new_n16565_, new_n16566_, new_n16567_, new_n16568_,
    new_n16569_, new_n16570_, new_n16571_, new_n16572_, new_n16573_,
    new_n16574_, new_n16575_, new_n16576_, new_n16577_, new_n16578_,
    new_n16579_, new_n16580_, new_n16581_, new_n16582_, new_n16583_,
    new_n16584_, new_n16585_, new_n16586_, new_n16587_, new_n16588_,
    new_n16589_, new_n16591_, new_n16592_, new_n16593_, new_n16594_,
    new_n16595_, new_n16596_, new_n16597_, new_n16598_, new_n16599_,
    new_n16600_, new_n16601_, new_n16602_, new_n16603_, new_n16604_,
    new_n16605_, new_n16606_, new_n16607_, new_n16608_, new_n16609_,
    new_n16610_, new_n16611_, new_n16612_, new_n16613_, new_n16614_,
    new_n16615_, new_n16616_, new_n16617_, new_n16618_, new_n16619_,
    new_n16620_, new_n16621_, new_n16622_, new_n16623_, new_n16624_,
    new_n16625_, new_n16626_, new_n16627_, new_n16628_, new_n16629_,
    new_n16630_, new_n16631_, new_n16632_, new_n16633_, new_n16634_,
    new_n16635_, new_n16636_, new_n16637_, new_n16638_, new_n16639_,
    new_n16640_, new_n16641_, new_n16642_, new_n16643_, new_n16644_,
    new_n16645_, new_n16646_, new_n16647_, new_n16648_, new_n16649_,
    new_n16650_, new_n16651_, new_n16652_, new_n16653_, new_n16654_,
    new_n16655_, new_n16656_, new_n16657_, new_n16658_, new_n16659_,
    new_n16660_, new_n16661_, new_n16662_, new_n16663_, new_n16664_,
    new_n16665_, new_n16666_, new_n16667_, new_n16668_, new_n16669_,
    new_n16670_, new_n16671_, new_n16672_, new_n16673_, new_n16674_,
    new_n16675_, new_n16676_, new_n16677_, new_n16678_, new_n16679_,
    new_n16680_, new_n16681_, new_n16682_, new_n16683_, new_n16684_,
    new_n16685_, new_n16686_, new_n16687_, new_n16688_, new_n16689_,
    new_n16690_, new_n16691_, new_n16692_, new_n16693_, new_n16694_,
    new_n16695_, new_n16696_, new_n16697_, new_n16698_, new_n16699_,
    new_n16700_, new_n16701_, new_n16702_, new_n16703_, new_n16704_,
    new_n16705_, new_n16706_, new_n16707_, new_n16708_, new_n16709_,
    new_n16710_, new_n16711_, new_n16712_, new_n16713_, new_n16714_,
    new_n16715_, new_n16716_, new_n16717_, new_n16718_, new_n16719_,
    new_n16720_, new_n16721_, new_n16722_, new_n16723_, new_n16724_,
    new_n16725_, new_n16726_, new_n16727_, new_n16728_, new_n16729_,
    new_n16730_, new_n16731_, new_n16732_, new_n16733_, new_n16734_,
    new_n16735_, new_n16736_, new_n16737_, new_n16738_, new_n16739_,
    new_n16740_, new_n16741_, new_n16742_, new_n16743_, new_n16744_,
    new_n16745_, new_n16746_, new_n16747_, new_n16748_, new_n16749_,
    new_n16750_, new_n16751_, new_n16752_, new_n16753_, new_n16754_,
    new_n16755_, new_n16756_, new_n16757_, new_n16758_, new_n16759_,
    new_n16760_, new_n16761_, new_n16762_, new_n16763_, new_n16764_,
    new_n16765_, new_n16766_, new_n16767_, new_n16768_, new_n16769_,
    new_n16770_, new_n16771_, new_n16772_, new_n16773_, new_n16774_,
    new_n16775_, new_n16776_, new_n16777_, new_n16778_, new_n16779_,
    new_n16780_, new_n16781_, new_n16782_, new_n16783_, new_n16784_,
    new_n16785_, new_n16786_, new_n16787_, new_n16788_, new_n16789_,
    new_n16790_, new_n16791_, new_n16792_, new_n16793_, new_n16794_,
    new_n16795_, new_n16796_, new_n16797_, new_n16798_, new_n16799_,
    new_n16800_, new_n16801_, new_n16802_, new_n16803_, new_n16804_,
    new_n16805_, new_n16806_, new_n16807_, new_n16808_, new_n16809_,
    new_n16810_, new_n16811_, new_n16812_, new_n16813_, new_n16814_,
    new_n16815_, new_n16816_, new_n16817_, new_n16818_, new_n16819_,
    new_n16820_, new_n16821_, new_n16822_, new_n16823_, new_n16824_,
    new_n16825_, new_n16826_, new_n16827_, new_n16828_, new_n16829_,
    new_n16830_, new_n16831_, new_n16832_, new_n16833_, new_n16834_,
    new_n16835_, new_n16836_, new_n16837_, new_n16838_, new_n16839_,
    new_n16840_, new_n16841_, new_n16842_, new_n16843_, new_n16844_,
    new_n16845_, new_n16846_, new_n16847_, new_n16848_, new_n16849_,
    new_n16850_, new_n16851_, new_n16853_, new_n16854_, new_n16855_,
    new_n16856_, new_n16857_, new_n16858_, new_n16859_, new_n16860_,
    new_n16861_, new_n16862_, new_n16863_, new_n16864_, new_n16865_,
    new_n16866_, new_n16867_, new_n16868_, new_n16869_, new_n16870_,
    new_n16871_, new_n16872_, new_n16873_, new_n16874_, new_n16875_,
    new_n16876_, new_n16877_, new_n16878_, new_n16879_, new_n16880_,
    new_n16881_, new_n16882_, new_n16883_, new_n16884_, new_n16885_,
    new_n16886_, new_n16887_, new_n16888_, new_n16889_, new_n16890_,
    new_n16891_, new_n16892_, new_n16893_, new_n16894_, new_n16895_,
    new_n16896_, new_n16897_, new_n16898_, new_n16899_, new_n16900_,
    new_n16901_, new_n16902_, new_n16903_, new_n16904_, new_n16905_,
    new_n16906_, new_n16907_, new_n16908_, new_n16909_, new_n16910_,
    new_n16911_, new_n16912_, new_n16913_, new_n16914_, new_n16915_,
    new_n16916_, new_n16917_, new_n16918_, new_n16919_, new_n16920_,
    new_n16921_, new_n16922_, new_n16923_, new_n16924_, new_n16925_,
    new_n16926_, new_n16927_, new_n16928_, new_n16929_, new_n16930_,
    new_n16931_, new_n16932_, new_n16933_, new_n16934_, new_n16935_,
    new_n16936_, new_n16937_, new_n16938_, new_n16939_, new_n16940_,
    new_n16941_, new_n16942_, new_n16943_, new_n16944_, new_n16945_,
    new_n16946_, new_n16947_, new_n16948_, new_n16949_, new_n16950_,
    new_n16951_, new_n16952_, new_n16953_, new_n16954_, new_n16955_,
    new_n16956_, new_n16957_, new_n16958_, new_n16959_, new_n16960_,
    new_n16961_, new_n16962_, new_n16963_, new_n16964_, new_n16965_,
    new_n16966_, new_n16967_, new_n16968_, new_n16969_, new_n16970_,
    new_n16971_, new_n16972_, new_n16973_, new_n16974_, new_n16975_,
    new_n16976_, new_n16977_, new_n16978_, new_n16979_, new_n16980_,
    new_n16981_, new_n16982_, new_n16983_, new_n16984_, new_n16985_,
    new_n16986_, new_n16987_, new_n16988_, new_n16989_, new_n16990_,
    new_n16991_, new_n16992_, new_n16993_, new_n16994_, new_n16995_,
    new_n16996_, new_n16997_, new_n16998_, new_n16999_, new_n17000_,
    new_n17001_, new_n17002_, new_n17003_, new_n17004_, new_n17005_,
    new_n17006_, new_n17007_, new_n17008_, new_n17009_, new_n17010_,
    new_n17011_, new_n17012_, new_n17013_, new_n17014_, new_n17015_,
    new_n17016_, new_n17017_, new_n17018_, new_n17019_, new_n17020_,
    new_n17021_, new_n17022_, new_n17023_, new_n17024_, new_n17025_,
    new_n17026_, new_n17027_, new_n17028_, new_n17029_, new_n17030_,
    new_n17031_, new_n17032_, new_n17033_, new_n17034_, new_n17035_,
    new_n17036_, new_n17037_, new_n17038_, new_n17039_, new_n17040_,
    new_n17041_, new_n17042_, new_n17043_, new_n17044_, new_n17045_,
    new_n17046_, new_n17047_, new_n17048_, new_n17049_, new_n17050_,
    new_n17051_, new_n17052_, new_n17053_, new_n17054_, new_n17055_,
    new_n17056_, new_n17057_, new_n17058_, new_n17059_, new_n17060_,
    new_n17061_, new_n17062_, new_n17063_, new_n17064_, new_n17065_,
    new_n17066_, new_n17067_, new_n17068_, new_n17069_, new_n17070_,
    new_n17071_, new_n17072_, new_n17073_, new_n17074_, new_n17075_,
    new_n17076_, new_n17077_, new_n17078_, new_n17079_, new_n17080_,
    new_n17081_, new_n17082_, new_n17083_, new_n17084_, new_n17085_,
    new_n17086_, new_n17087_, new_n17088_, new_n17089_, new_n17090_,
    new_n17091_, new_n17092_, new_n17093_, new_n17094_, new_n17095_,
    new_n17096_, new_n17097_, new_n17098_, new_n17099_, new_n17100_,
    new_n17101_, new_n17102_, new_n17103_, new_n17104_, new_n17105_,
    new_n17106_, new_n17107_, new_n17108_, new_n17109_, new_n17110_,
    new_n17111_, new_n17112_, new_n17113_, new_n17114_, new_n17115_,
    new_n17116_, new_n17117_, new_n17118_, new_n17119_, new_n17120_,
    new_n17121_, new_n17122_, new_n17123_, new_n17124_, new_n17125_,
    new_n17126_, new_n17127_, new_n17128_, new_n17129_, new_n17131_,
    new_n17132_, new_n17133_, new_n17134_, new_n17135_, new_n17136_,
    new_n17137_, new_n17138_, new_n17139_, new_n17140_, new_n17141_,
    new_n17142_, new_n17143_, new_n17144_, new_n17145_, new_n17146_,
    new_n17147_, new_n17148_, new_n17149_, new_n17150_, new_n17151_,
    new_n17152_, new_n17153_, new_n17154_, new_n17155_, new_n17156_,
    new_n17157_, new_n17158_, new_n17159_, new_n17160_, new_n17161_,
    new_n17162_, new_n17163_, new_n17164_, new_n17165_, new_n17166_,
    new_n17167_, new_n17168_, new_n17169_, new_n17170_, new_n17171_,
    new_n17172_, new_n17173_, new_n17174_, new_n17175_, new_n17176_,
    new_n17177_, new_n17178_, new_n17179_, new_n17180_, new_n17181_,
    new_n17182_, new_n17183_, new_n17184_, new_n17185_, new_n17186_,
    new_n17187_, new_n17188_, new_n17189_, new_n17190_, new_n17191_,
    new_n17192_, new_n17193_, new_n17194_, new_n17195_, new_n17196_,
    new_n17197_, new_n17198_, new_n17199_, new_n17200_, new_n17201_,
    new_n17202_, new_n17203_, new_n17204_, new_n17205_, new_n17206_,
    new_n17207_, new_n17208_, new_n17209_, new_n17210_, new_n17211_,
    new_n17212_, new_n17213_, new_n17214_, new_n17215_, new_n17216_,
    new_n17217_, new_n17218_, new_n17219_, new_n17220_, new_n17221_,
    new_n17222_, new_n17223_, new_n17224_, new_n17225_, new_n17226_,
    new_n17227_, new_n17228_, new_n17229_, new_n17230_, new_n17231_,
    new_n17232_, new_n17233_, new_n17234_, new_n17235_, new_n17236_,
    new_n17237_, new_n17238_, new_n17239_, new_n17240_, new_n17241_,
    new_n17242_, new_n17243_, new_n17244_, new_n17245_, new_n17246_,
    new_n17247_, new_n17248_, new_n17249_, new_n17250_, new_n17251_,
    new_n17252_, new_n17253_, new_n17254_, new_n17255_, new_n17256_,
    new_n17257_, new_n17258_, new_n17259_, new_n17260_, new_n17261_,
    new_n17262_, new_n17263_, new_n17264_, new_n17265_, new_n17266_,
    new_n17267_, new_n17268_, new_n17269_, new_n17270_, new_n17271_,
    new_n17272_, new_n17273_, new_n17274_, new_n17275_, new_n17276_,
    new_n17277_, new_n17278_, new_n17279_, new_n17280_, new_n17281_,
    new_n17282_, new_n17283_, new_n17284_, new_n17285_, new_n17286_,
    new_n17287_, new_n17288_, new_n17289_, new_n17290_, new_n17291_,
    new_n17292_, new_n17293_, new_n17294_, new_n17295_, new_n17296_,
    new_n17297_, new_n17298_, new_n17299_, new_n17300_, new_n17301_,
    new_n17302_, new_n17303_, new_n17304_, new_n17305_, new_n17306_,
    new_n17307_, new_n17308_, new_n17309_, new_n17310_, new_n17311_,
    new_n17312_, new_n17313_, new_n17314_, new_n17315_, new_n17316_,
    new_n17317_, new_n17318_, new_n17319_, new_n17320_, new_n17321_,
    new_n17322_, new_n17323_, new_n17324_, new_n17325_, new_n17326_,
    new_n17327_, new_n17328_, new_n17329_, new_n17330_, new_n17331_,
    new_n17332_, new_n17333_, new_n17334_, new_n17335_, new_n17336_,
    new_n17337_, new_n17338_, new_n17339_, new_n17340_, new_n17341_,
    new_n17342_, new_n17343_, new_n17344_, new_n17345_, new_n17346_,
    new_n17347_, new_n17348_, new_n17349_, new_n17350_, new_n17351_,
    new_n17352_, new_n17353_, new_n17354_, new_n17355_, new_n17356_,
    new_n17357_, new_n17358_, new_n17359_, new_n17360_, new_n17361_,
    new_n17362_, new_n17363_, new_n17364_, new_n17365_, new_n17366_,
    new_n17367_, new_n17368_, new_n17369_, new_n17370_, new_n17371_,
    new_n17372_, new_n17373_, new_n17374_, new_n17375_, new_n17376_,
    new_n17377_, new_n17378_, new_n17379_, new_n17380_, new_n17381_,
    new_n17382_, new_n17383_, new_n17384_, new_n17385_, new_n17386_,
    new_n17387_, new_n17388_, new_n17389_, new_n17390_, new_n17391_,
    new_n17392_, new_n17393_, new_n17394_, new_n17395_, new_n17396_,
    new_n17397_, new_n17398_, new_n17399_, new_n17400_, new_n17402_,
    new_n17403_, new_n17404_, new_n17405_, new_n17406_, new_n17407_,
    new_n17408_, new_n17409_, new_n17410_, new_n17411_, new_n17412_,
    new_n17413_, new_n17414_, new_n17415_, new_n17416_, new_n17417_,
    new_n17418_, new_n17419_, new_n17420_, new_n17421_, new_n17422_,
    new_n17423_, new_n17424_, new_n17425_, new_n17426_, new_n17427_,
    new_n17428_, new_n17429_, new_n17430_, new_n17431_, new_n17432_,
    new_n17433_, new_n17434_, new_n17435_, new_n17436_, new_n17437_,
    new_n17438_, new_n17439_, new_n17440_, new_n17441_, new_n17442_,
    new_n17443_, new_n17444_, new_n17445_, new_n17446_, new_n17447_,
    new_n17448_, new_n17449_, new_n17450_, new_n17451_, new_n17452_,
    new_n17453_, new_n17454_, new_n17455_, new_n17456_, new_n17457_,
    new_n17458_, new_n17459_, new_n17460_, new_n17461_, new_n17462_,
    new_n17463_, new_n17464_, new_n17465_, new_n17466_, new_n17467_,
    new_n17468_, new_n17469_, new_n17470_, new_n17471_, new_n17472_,
    new_n17473_, new_n17474_, new_n17475_, new_n17476_, new_n17477_,
    new_n17478_, new_n17479_, new_n17480_, new_n17481_, new_n17482_,
    new_n17483_, new_n17484_, new_n17485_, new_n17486_, new_n17487_,
    new_n17488_, new_n17489_, new_n17490_, new_n17491_, new_n17492_,
    new_n17493_, new_n17494_, new_n17495_, new_n17496_, new_n17497_,
    new_n17498_, new_n17499_, new_n17500_, new_n17501_, new_n17502_,
    new_n17503_, new_n17504_, new_n17505_, new_n17506_, new_n17507_,
    new_n17508_, new_n17509_, new_n17510_, new_n17511_, new_n17512_,
    new_n17513_, new_n17514_, new_n17515_, new_n17516_, new_n17517_,
    new_n17518_, new_n17519_, new_n17520_, new_n17521_, new_n17522_,
    new_n17523_, new_n17524_, new_n17525_, new_n17526_, new_n17527_,
    new_n17528_, new_n17529_, new_n17530_, new_n17531_, new_n17532_,
    new_n17533_, new_n17534_, new_n17535_, new_n17536_, new_n17537_,
    new_n17538_, new_n17539_, new_n17540_, new_n17541_, new_n17542_,
    new_n17543_, new_n17544_, new_n17545_, new_n17546_, new_n17547_,
    new_n17548_, new_n17549_, new_n17550_, new_n17551_, new_n17552_,
    new_n17553_, new_n17554_, new_n17555_, new_n17556_, new_n17557_,
    new_n17558_, new_n17559_, new_n17560_, new_n17561_, new_n17562_,
    new_n17563_, new_n17564_, new_n17565_, new_n17566_, new_n17567_,
    new_n17568_, new_n17569_, new_n17570_, new_n17571_, new_n17572_,
    new_n17573_, new_n17574_, new_n17575_, new_n17576_, new_n17577_,
    new_n17578_, new_n17579_, new_n17580_, new_n17581_, new_n17582_,
    new_n17583_, new_n17584_, new_n17585_, new_n17586_, new_n17587_,
    new_n17588_, new_n17589_, new_n17590_, new_n17591_, new_n17592_,
    new_n17593_, new_n17594_, new_n17595_, new_n17596_, new_n17597_,
    new_n17598_, new_n17599_, new_n17600_, new_n17601_, new_n17602_,
    new_n17603_, new_n17604_, new_n17605_, new_n17606_, new_n17607_,
    new_n17608_, new_n17609_, new_n17610_, new_n17611_, new_n17612_,
    new_n17613_, new_n17614_, new_n17615_, new_n17616_, new_n17617_,
    new_n17618_, new_n17619_, new_n17620_, new_n17621_, new_n17622_,
    new_n17623_, new_n17624_, new_n17625_, new_n17626_, new_n17627_,
    new_n17628_, new_n17629_, new_n17630_, new_n17631_, new_n17632_,
    new_n17633_, new_n17634_, new_n17635_, new_n17636_, new_n17637_,
    new_n17638_, new_n17639_, new_n17640_, new_n17641_, new_n17642_,
    new_n17643_, new_n17644_, new_n17645_, new_n17646_, new_n17647_,
    new_n17648_, new_n17649_, new_n17650_, new_n17651_, new_n17652_,
    new_n17653_, new_n17654_, new_n17655_, new_n17656_, new_n17657_,
    new_n17658_, new_n17659_, new_n17660_, new_n17661_, new_n17662_,
    new_n17663_, new_n17664_, new_n17665_, new_n17666_, new_n17667_,
    new_n17668_, new_n17669_, new_n17670_, new_n17672_, new_n17673_,
    new_n17674_, new_n17675_, new_n17676_, new_n17677_, new_n17678_,
    new_n17679_, new_n17680_, new_n17681_, new_n17682_, new_n17683_,
    new_n17684_, new_n17685_, new_n17686_, new_n17687_, new_n17688_,
    new_n17689_, new_n17690_, new_n17691_, new_n17692_, new_n17693_,
    new_n17694_, new_n17695_, new_n17696_, new_n17697_, new_n17698_,
    new_n17699_, new_n17700_, new_n17701_, new_n17702_, new_n17703_,
    new_n17704_, new_n17705_, new_n17706_, new_n17707_, new_n17708_,
    new_n17709_, new_n17710_, new_n17711_, new_n17712_, new_n17713_,
    new_n17714_, new_n17715_, new_n17716_, new_n17717_, new_n17718_,
    new_n17719_, new_n17720_, new_n17721_, new_n17722_, new_n17723_,
    new_n17724_, new_n17725_, new_n17726_, new_n17727_, new_n17728_,
    new_n17729_, new_n17730_, new_n17731_, new_n17732_, new_n17733_,
    new_n17734_, new_n17735_, new_n17736_, new_n17737_, new_n17738_,
    new_n17739_, new_n17740_, new_n17741_, new_n17742_, new_n17743_,
    new_n17744_, new_n17745_, new_n17746_, new_n17747_, new_n17748_,
    new_n17749_, new_n17750_, new_n17751_, new_n17752_, new_n17753_,
    new_n17754_, new_n17755_, new_n17756_, new_n17757_, new_n17758_,
    new_n17759_, new_n17760_, new_n17761_, new_n17762_, new_n17763_,
    new_n17764_, new_n17765_, new_n17766_, new_n17767_, new_n17768_,
    new_n17769_, new_n17770_, new_n17771_, new_n17772_, new_n17773_,
    new_n17774_, new_n17775_, new_n17776_, new_n17777_, new_n17778_,
    new_n17779_, new_n17780_, new_n17781_, new_n17782_, new_n17783_,
    new_n17784_, new_n17785_, new_n17786_, new_n17787_, new_n17788_,
    new_n17789_, new_n17790_, new_n17791_, new_n17792_, new_n17793_,
    new_n17794_, new_n17795_, new_n17796_, new_n17797_, new_n17798_,
    new_n17799_, new_n17800_, new_n17801_, new_n17802_, new_n17803_,
    new_n17804_, new_n17805_, new_n17806_, new_n17807_, new_n17808_,
    new_n17809_, new_n17810_, new_n17811_, new_n17812_, new_n17813_,
    new_n17814_, new_n17815_, new_n17816_, new_n17817_, new_n17818_,
    new_n17819_, new_n17820_, new_n17821_, new_n17822_, new_n17823_,
    new_n17824_, new_n17825_, new_n17826_, new_n17827_, new_n17828_,
    new_n17829_, new_n17830_, new_n17831_, new_n17832_, new_n17833_,
    new_n17834_, new_n17835_, new_n17836_, new_n17837_, new_n17838_,
    new_n17839_, new_n17840_, new_n17841_, new_n17842_, new_n17843_,
    new_n17844_, new_n17845_, new_n17846_, new_n17847_, new_n17848_,
    new_n17849_, new_n17850_, new_n17851_, new_n17852_, new_n17853_,
    new_n17854_, new_n17855_, new_n17856_, new_n17857_, new_n17858_,
    new_n17859_, new_n17860_, new_n17861_, new_n17862_, new_n17863_,
    new_n17864_, new_n17865_, new_n17866_, new_n17867_, new_n17868_,
    new_n17869_, new_n17870_, new_n17871_, new_n17872_, new_n17873_,
    new_n17874_, new_n17875_, new_n17876_, new_n17877_, new_n17878_,
    new_n17879_, new_n17880_, new_n17881_, new_n17882_, new_n17883_,
    new_n17884_, new_n17885_, new_n17886_, new_n17887_, new_n17888_,
    new_n17889_, new_n17890_, new_n17891_, new_n17892_, new_n17893_,
    new_n17894_, new_n17895_, new_n17896_, new_n17897_, new_n17898_,
    new_n17899_, new_n17900_, new_n17901_, new_n17902_, new_n17903_,
    new_n17904_, new_n17905_, new_n17906_, new_n17907_, new_n17908_,
    new_n17909_, new_n17910_, new_n17911_, new_n17912_, new_n17913_,
    new_n17914_, new_n17915_, new_n17916_, new_n17917_, new_n17918_,
    new_n17919_, new_n17920_, new_n17921_, new_n17922_, new_n17923_,
    new_n17924_, new_n17925_, new_n17926_, new_n17927_, new_n17928_,
    new_n17929_, new_n17930_, new_n17931_, new_n17932_, new_n17933_,
    new_n17934_, new_n17935_, new_n17936_, new_n17937_, new_n17938_,
    new_n17939_, new_n17940_, new_n17941_, new_n17942_, new_n17943_,
    new_n17945_, new_n17946_, new_n17947_, new_n17948_, new_n17949_,
    new_n17950_, new_n17951_, new_n17952_, new_n17953_, new_n17954_,
    new_n17955_, new_n17956_, new_n17957_, new_n17958_, new_n17959_,
    new_n17960_, new_n17961_, new_n17962_, new_n17963_, new_n17964_,
    new_n17965_, new_n17966_, new_n17967_, new_n17968_, new_n17969_,
    new_n17970_, new_n17971_, new_n17972_, new_n17973_, new_n17974_,
    new_n17975_, new_n17976_, new_n17977_, new_n17978_, new_n17979_,
    new_n17980_, new_n17981_, new_n17982_, new_n17983_, new_n17984_,
    new_n17985_, new_n17986_, new_n17987_, new_n17988_, new_n17989_,
    new_n17990_, new_n17991_, new_n17992_, new_n17993_, new_n17994_,
    new_n17995_, new_n17996_, new_n17997_, new_n17998_, new_n17999_,
    new_n18000_, new_n18001_, new_n18002_, new_n18003_, new_n18004_,
    new_n18005_, new_n18006_, new_n18007_, new_n18008_, new_n18009_,
    new_n18010_, new_n18011_, new_n18012_, new_n18013_, new_n18014_,
    new_n18015_, new_n18016_, new_n18017_, new_n18018_, new_n18019_,
    new_n18020_, new_n18021_, new_n18022_, new_n18023_, new_n18024_,
    new_n18025_, new_n18026_, new_n18027_, new_n18028_, new_n18029_,
    new_n18030_, new_n18031_, new_n18032_, new_n18033_, new_n18034_,
    new_n18035_, new_n18036_, new_n18037_, new_n18038_, new_n18039_,
    new_n18040_, new_n18041_, new_n18042_, new_n18043_, new_n18044_,
    new_n18045_, new_n18046_, new_n18047_, new_n18048_, new_n18049_,
    new_n18050_, new_n18051_, new_n18052_, new_n18053_, new_n18054_,
    new_n18055_, new_n18056_, new_n18057_, new_n18058_, new_n18059_,
    new_n18060_, new_n18061_, new_n18062_, new_n18063_, new_n18064_,
    new_n18065_, new_n18066_, new_n18067_, new_n18068_, new_n18069_,
    new_n18070_, new_n18071_, new_n18072_, new_n18073_, new_n18074_,
    new_n18075_, new_n18076_, new_n18077_, new_n18078_, new_n18079_,
    new_n18080_, new_n18081_, new_n18082_, new_n18083_, new_n18084_,
    new_n18085_, new_n18086_, new_n18087_, new_n18088_, new_n18089_,
    new_n18090_, new_n18091_, new_n18092_, new_n18093_, new_n18094_,
    new_n18095_, new_n18096_, new_n18097_, new_n18098_, new_n18099_,
    new_n18100_, new_n18101_, new_n18102_, new_n18103_, new_n18104_,
    new_n18105_, new_n18106_, new_n18107_, new_n18108_, new_n18109_,
    new_n18110_, new_n18111_, new_n18112_, new_n18113_, new_n18114_,
    new_n18115_, new_n18116_, new_n18117_, new_n18118_, new_n18119_,
    new_n18120_, new_n18121_, new_n18122_, new_n18123_, new_n18124_,
    new_n18125_, new_n18126_, new_n18127_, new_n18128_, new_n18129_,
    new_n18130_, new_n18131_, new_n18132_, new_n18133_, new_n18134_,
    new_n18135_, new_n18136_, new_n18137_, new_n18138_, new_n18139_,
    new_n18140_, new_n18141_, new_n18142_, new_n18143_, new_n18144_,
    new_n18145_, new_n18146_, new_n18147_, new_n18148_, new_n18149_,
    new_n18150_, new_n18151_, new_n18152_, new_n18153_, new_n18154_,
    new_n18155_, new_n18156_, new_n18157_, new_n18158_, new_n18159_,
    new_n18160_, new_n18161_, new_n18162_, new_n18163_, new_n18164_,
    new_n18165_, new_n18166_, new_n18167_, new_n18168_, new_n18169_,
    new_n18170_, new_n18171_, new_n18172_, new_n18173_, new_n18174_,
    new_n18175_, new_n18176_, new_n18177_, new_n18178_, new_n18179_,
    new_n18180_, new_n18181_, new_n18182_, new_n18183_, new_n18184_,
    new_n18185_, new_n18186_, new_n18187_, new_n18188_, new_n18189_,
    new_n18190_, new_n18191_, new_n18192_, new_n18193_, new_n18194_,
    new_n18195_, new_n18196_, new_n18197_, new_n18198_, new_n18199_,
    new_n18200_, new_n18201_, new_n18202_, new_n18203_, new_n18204_,
    new_n18205_, new_n18206_, new_n18207_, new_n18208_, new_n18209_,
    new_n18210_, new_n18211_, new_n18212_, new_n18213_, new_n18214_,
    new_n18215_, new_n18216_, new_n18218_, new_n18219_, new_n18220_,
    new_n18221_, new_n18222_, new_n18223_, new_n18224_, new_n18225_,
    new_n18226_, new_n18227_, new_n18228_, new_n18229_, new_n18230_,
    new_n18231_, new_n18232_, new_n18233_, new_n18234_, new_n18235_,
    new_n18236_, new_n18237_, new_n18238_, new_n18239_, new_n18240_,
    new_n18241_, new_n18242_, new_n18243_, new_n18244_, new_n18245_,
    new_n18246_, new_n18247_, new_n18248_, new_n18249_, new_n18250_,
    new_n18251_, new_n18252_, new_n18253_, new_n18254_, new_n18255_,
    new_n18256_, new_n18257_, new_n18258_, new_n18259_, new_n18260_,
    new_n18261_, new_n18262_, new_n18263_, new_n18264_, new_n18265_,
    new_n18266_, new_n18267_, new_n18268_, new_n18269_, new_n18270_,
    new_n18271_, new_n18272_, new_n18273_, new_n18274_, new_n18275_,
    new_n18276_, new_n18277_, new_n18278_, new_n18279_, new_n18280_,
    new_n18281_, new_n18282_, new_n18283_, new_n18284_, new_n18285_,
    new_n18286_, new_n18287_, new_n18288_, new_n18289_, new_n18290_,
    new_n18291_, new_n18292_, new_n18293_, new_n18294_, new_n18295_,
    new_n18296_, new_n18297_, new_n18298_, new_n18299_, new_n18300_,
    new_n18301_, new_n18302_, new_n18303_, new_n18304_, new_n18305_,
    new_n18306_, new_n18307_, new_n18308_, new_n18309_, new_n18310_,
    new_n18311_, new_n18312_, new_n18313_, new_n18314_, new_n18315_,
    new_n18316_, new_n18317_, new_n18318_, new_n18319_, new_n18320_,
    new_n18321_, new_n18322_, new_n18323_, new_n18324_, new_n18325_,
    new_n18326_, new_n18327_, new_n18328_, new_n18329_, new_n18330_,
    new_n18331_, new_n18332_, new_n18333_, new_n18334_, new_n18335_,
    new_n18336_, new_n18337_, new_n18338_, new_n18339_, new_n18340_,
    new_n18341_, new_n18342_, new_n18343_, new_n18344_, new_n18345_,
    new_n18346_, new_n18347_, new_n18348_, new_n18349_, new_n18350_,
    new_n18351_, new_n18352_, new_n18353_, new_n18354_, new_n18355_,
    new_n18356_, new_n18357_, new_n18358_, new_n18359_, new_n18360_,
    new_n18361_, new_n18362_, new_n18363_, new_n18364_, new_n18365_,
    new_n18366_, new_n18367_, new_n18368_, new_n18369_, new_n18370_,
    new_n18371_, new_n18372_, new_n18373_, new_n18374_, new_n18375_,
    new_n18376_, new_n18377_, new_n18378_, new_n18379_, new_n18380_,
    new_n18381_, new_n18382_, new_n18383_, new_n18384_, new_n18385_,
    new_n18386_, new_n18387_, new_n18388_, new_n18389_, new_n18390_,
    new_n18391_, new_n18392_, new_n18393_, new_n18394_, new_n18395_,
    new_n18396_, new_n18397_, new_n18398_, new_n18399_, new_n18400_,
    new_n18401_, new_n18402_, new_n18403_, new_n18404_, new_n18405_,
    new_n18406_, new_n18407_, new_n18408_, new_n18409_, new_n18410_,
    new_n18411_, new_n18412_, new_n18413_, new_n18414_, new_n18415_,
    new_n18416_, new_n18417_, new_n18418_, new_n18419_, new_n18420_,
    new_n18421_, new_n18422_, new_n18423_, new_n18424_, new_n18425_,
    new_n18426_, new_n18427_, new_n18428_, new_n18429_, new_n18430_,
    new_n18431_, new_n18432_, new_n18433_, new_n18434_, new_n18435_,
    new_n18436_, new_n18437_, new_n18438_, new_n18439_, new_n18440_,
    new_n18441_, new_n18442_, new_n18443_, new_n18444_, new_n18445_,
    new_n18446_, new_n18447_, new_n18448_, new_n18449_, new_n18450_,
    new_n18451_, new_n18452_, new_n18453_, new_n18454_, new_n18455_,
    new_n18456_, new_n18457_, new_n18458_, new_n18459_, new_n18460_,
    new_n18461_, new_n18462_, new_n18463_, new_n18464_, new_n18465_,
    new_n18466_, new_n18467_, new_n18468_, new_n18469_, new_n18470_,
    new_n18471_, new_n18472_, new_n18473_, new_n18474_, new_n18475_,
    new_n18476_, new_n18477_, new_n18478_, new_n18479_, new_n18480_,
    new_n18481_, new_n18482_, new_n18483_, new_n18484_, new_n18485_,
    new_n18486_, new_n18488_, new_n18489_, new_n18490_, new_n18491_,
    new_n18492_, new_n18493_, new_n18494_, new_n18495_, new_n18496_,
    new_n18497_, new_n18498_, new_n18499_, new_n18500_, new_n18501_,
    new_n18502_, new_n18503_, new_n18504_, new_n18505_, new_n18506_,
    new_n18507_, new_n18508_, new_n18509_, new_n18510_, new_n18511_,
    new_n18512_, new_n18513_, new_n18514_, new_n18515_, new_n18516_,
    new_n18517_, new_n18518_, new_n18519_, new_n18520_, new_n18521_,
    new_n18522_, new_n18523_, new_n18524_, new_n18525_, new_n18526_,
    new_n18527_, new_n18528_, new_n18529_, new_n18530_, new_n18531_,
    new_n18532_, new_n18533_, new_n18534_, new_n18535_, new_n18536_,
    new_n18537_, new_n18538_, new_n18539_, new_n18540_, new_n18541_,
    new_n18542_, new_n18543_, new_n18544_, new_n18545_, new_n18546_,
    new_n18547_, new_n18548_, new_n18549_, new_n18550_, new_n18551_,
    new_n18552_, new_n18553_, new_n18554_, new_n18555_, new_n18556_,
    new_n18557_, new_n18558_, new_n18559_, new_n18560_, new_n18561_,
    new_n18562_, new_n18563_, new_n18564_, new_n18565_, new_n18566_,
    new_n18567_, new_n18568_, new_n18569_, new_n18570_, new_n18571_,
    new_n18572_, new_n18573_, new_n18574_, new_n18575_, new_n18576_,
    new_n18577_, new_n18578_, new_n18579_, new_n18580_, new_n18581_,
    new_n18582_, new_n18583_, new_n18584_, new_n18585_, new_n18586_,
    new_n18587_, new_n18588_, new_n18589_, new_n18590_, new_n18591_,
    new_n18592_, new_n18593_, new_n18594_, new_n18595_, new_n18596_,
    new_n18597_, new_n18598_, new_n18599_, new_n18600_, new_n18601_,
    new_n18602_, new_n18603_, new_n18604_, new_n18605_, new_n18606_,
    new_n18607_, new_n18608_, new_n18609_, new_n18610_, new_n18611_,
    new_n18612_, new_n18613_, new_n18614_, new_n18615_, new_n18616_,
    new_n18617_, new_n18618_, new_n18619_, new_n18620_, new_n18621_,
    new_n18622_, new_n18623_, new_n18624_, new_n18625_, new_n18626_,
    new_n18627_, new_n18628_, new_n18629_, new_n18630_, new_n18631_,
    new_n18632_, new_n18633_, new_n18634_, new_n18635_, new_n18636_,
    new_n18637_, new_n18638_, new_n18639_, new_n18640_, new_n18641_,
    new_n18642_, new_n18643_, new_n18644_, new_n18645_, new_n18646_,
    new_n18647_, new_n18648_, new_n18649_, new_n18650_, new_n18651_,
    new_n18652_, new_n18653_, new_n18654_, new_n18655_, new_n18656_,
    new_n18657_, new_n18658_, new_n18659_, new_n18660_, new_n18661_,
    new_n18662_, new_n18663_, new_n18664_, new_n18665_, new_n18666_,
    new_n18667_, new_n18668_, new_n18669_, new_n18670_, new_n18671_,
    new_n18672_, new_n18673_, new_n18674_, new_n18675_, new_n18676_,
    new_n18677_, new_n18678_, new_n18679_, new_n18680_, new_n18681_,
    new_n18682_, new_n18683_, new_n18684_, new_n18685_, new_n18686_,
    new_n18687_, new_n18688_, new_n18689_, new_n18690_, new_n18691_,
    new_n18692_, new_n18693_, new_n18694_, new_n18695_, new_n18696_,
    new_n18697_, new_n18698_, new_n18699_, new_n18700_, new_n18701_,
    new_n18702_, new_n18703_, new_n18704_, new_n18705_, new_n18706_,
    new_n18707_, new_n18708_, new_n18709_, new_n18710_, new_n18711_,
    new_n18712_, new_n18713_, new_n18714_, new_n18715_, new_n18716_,
    new_n18717_, new_n18718_, new_n18719_, new_n18720_, new_n18721_,
    new_n18722_, new_n18723_, new_n18724_, new_n18725_, new_n18726_,
    new_n18727_, new_n18728_, new_n18729_, new_n18730_, new_n18731_,
    new_n18732_, new_n18733_, new_n18734_, new_n18735_, new_n18736_,
    new_n18737_, new_n18738_, new_n18739_, new_n18740_, new_n18741_,
    new_n18742_, new_n18743_, new_n18744_, new_n18745_, new_n18746_,
    new_n18747_, new_n18748_, new_n18749_, new_n18750_, new_n18751_,
    new_n18752_, new_n18753_, new_n18754_, new_n18755_, new_n18756_,
    new_n18758_, new_n18759_, new_n18760_, new_n18761_, new_n18762_,
    new_n18763_, new_n18764_, new_n18765_, new_n18766_, new_n18767_,
    new_n18768_, new_n18769_, new_n18770_, new_n18771_, new_n18772_,
    new_n18773_, new_n18774_, new_n18775_, new_n18776_, new_n18777_,
    new_n18778_, new_n18779_, new_n18780_, new_n18781_, new_n18782_,
    new_n18783_, new_n18784_, new_n18785_, new_n18786_, new_n18787_,
    new_n18788_, new_n18789_, new_n18790_, new_n18791_, new_n18792_,
    new_n18793_, new_n18794_, new_n18795_, new_n18796_, new_n18797_,
    new_n18798_, new_n18799_, new_n18800_, new_n18801_, new_n18802_,
    new_n18803_, new_n18804_, new_n18805_, new_n18806_, new_n18807_,
    new_n18808_, new_n18809_, new_n18810_, new_n18811_, new_n18812_,
    new_n18813_, new_n18814_, new_n18815_, new_n18816_, new_n18817_,
    new_n18818_, new_n18819_, new_n18820_, new_n18821_, new_n18822_,
    new_n18823_, new_n18824_, new_n18825_, new_n18826_, new_n18827_,
    new_n18828_, new_n18829_, new_n18830_, new_n18831_, new_n18832_,
    new_n18833_, new_n18834_, new_n18835_, new_n18836_, new_n18837_,
    new_n18838_, new_n18839_, new_n18840_, new_n18841_, new_n18842_,
    new_n18843_, new_n18844_, new_n18845_, new_n18846_, new_n18847_,
    new_n18848_, new_n18849_, new_n18850_, new_n18851_, new_n18852_,
    new_n18853_, new_n18854_, new_n18855_, new_n18856_, new_n18857_,
    new_n18858_, new_n18859_, new_n18860_, new_n18861_, new_n18862_,
    new_n18863_, new_n18864_, new_n18865_, new_n18866_, new_n18867_,
    new_n18868_, new_n18869_, new_n18870_, new_n18871_, new_n18872_,
    new_n18873_, new_n18874_, new_n18875_, new_n18876_, new_n18877_,
    new_n18878_, new_n18879_, new_n18880_, new_n18881_, new_n18882_,
    new_n18883_, new_n18884_, new_n18885_, new_n18886_, new_n18887_,
    new_n18888_, new_n18889_, new_n18890_, new_n18891_, new_n18892_,
    new_n18893_, new_n18894_, new_n18895_, new_n18896_, new_n18897_,
    new_n18898_, new_n18899_, new_n18900_, new_n18901_, new_n18902_,
    new_n18903_, new_n18904_, new_n18905_, new_n18906_, new_n18907_,
    new_n18908_, new_n18909_, new_n18910_, new_n18911_, new_n18912_,
    new_n18913_, new_n18914_, new_n18915_, new_n18916_, new_n18917_,
    new_n18918_, new_n18919_, new_n18920_, new_n18921_, new_n18922_,
    new_n18923_, new_n18924_, new_n18925_, new_n18926_, new_n18927_,
    new_n18928_, new_n18929_, new_n18930_, new_n18931_, new_n18932_,
    new_n18933_, new_n18934_, new_n18935_, new_n18936_, new_n18937_,
    new_n18938_, new_n18939_, new_n18940_, new_n18941_, new_n18942_,
    new_n18943_, new_n18944_, new_n18945_, new_n18946_, new_n18947_,
    new_n18948_, new_n18949_, new_n18950_, new_n18951_, new_n18952_,
    new_n18953_, new_n18954_, new_n18955_, new_n18956_, new_n18957_,
    new_n18958_, new_n18959_, new_n18960_, new_n18961_, new_n18962_,
    new_n18963_, new_n18964_, new_n18965_, new_n18966_, new_n18967_,
    new_n18968_, new_n18969_, new_n18970_, new_n18971_, new_n18972_,
    new_n18973_, new_n18974_, new_n18975_, new_n18976_, new_n18977_,
    new_n18978_, new_n18979_, new_n18980_, new_n18981_, new_n18982_,
    new_n18983_, new_n18984_, new_n18985_, new_n18986_, new_n18987_,
    new_n18988_, new_n18989_, new_n18990_, new_n18991_, new_n18992_,
    new_n18993_, new_n18994_, new_n18995_, new_n18996_, new_n18997_,
    new_n18998_, new_n18999_, new_n19000_, new_n19001_, new_n19002_,
    new_n19003_, new_n19004_, new_n19005_, new_n19006_, new_n19007_,
    new_n19008_, new_n19009_, new_n19010_, new_n19011_, new_n19012_,
    new_n19013_, new_n19014_, new_n19015_, new_n19016_, new_n19017_,
    new_n19018_, new_n19019_, new_n19020_, new_n19021_, new_n19022_,
    new_n19023_, new_n19024_, new_n19025_, new_n19026_, new_n19028_,
    new_n19029_, new_n19030_, new_n19031_, new_n19032_, new_n19033_,
    new_n19034_, new_n19035_, new_n19036_, new_n19037_, new_n19038_,
    new_n19039_, new_n19040_, new_n19041_, new_n19042_, new_n19043_,
    new_n19044_, new_n19045_, new_n19046_, new_n19047_, new_n19048_,
    new_n19049_, new_n19050_, new_n19051_, new_n19052_, new_n19053_,
    new_n19054_, new_n19055_, new_n19056_, new_n19057_, new_n19058_,
    new_n19059_, new_n19060_, new_n19061_, new_n19062_, new_n19063_,
    new_n19064_, new_n19065_, new_n19066_, new_n19067_, new_n19068_,
    new_n19069_, new_n19070_, new_n19071_, new_n19072_, new_n19073_,
    new_n19074_, new_n19075_, new_n19076_, new_n19077_, new_n19078_,
    new_n19079_, new_n19080_, new_n19081_, new_n19082_, new_n19083_,
    new_n19084_, new_n19085_, new_n19086_, new_n19087_, new_n19088_,
    new_n19089_, new_n19090_, new_n19091_, new_n19092_, new_n19093_,
    new_n19094_, new_n19095_, new_n19096_, new_n19097_, new_n19098_,
    new_n19099_, new_n19100_, new_n19101_, new_n19102_, new_n19103_,
    new_n19104_, new_n19105_, new_n19106_, new_n19107_, new_n19108_,
    new_n19109_, new_n19110_, new_n19111_, new_n19112_, new_n19113_,
    new_n19114_, new_n19115_, new_n19116_, new_n19117_, new_n19118_,
    new_n19119_, new_n19120_, new_n19121_, new_n19122_, new_n19123_,
    new_n19124_, new_n19125_, new_n19126_, new_n19127_, new_n19128_,
    new_n19129_, new_n19130_, new_n19131_, new_n19132_, new_n19133_,
    new_n19134_, new_n19135_, new_n19136_, new_n19137_, new_n19138_,
    new_n19139_, new_n19140_, new_n19141_, new_n19142_, new_n19143_,
    new_n19144_, new_n19145_, new_n19146_, new_n19147_, new_n19148_,
    new_n19149_, new_n19150_, new_n19151_, new_n19152_, new_n19153_,
    new_n19154_, new_n19155_, new_n19156_, new_n19157_, new_n19158_,
    new_n19159_, new_n19160_, new_n19161_, new_n19162_, new_n19163_,
    new_n19164_, new_n19165_, new_n19166_, new_n19167_, new_n19168_,
    new_n19169_, new_n19170_, new_n19171_, new_n19172_, new_n19173_,
    new_n19174_, new_n19175_, new_n19176_, new_n19177_, new_n19178_,
    new_n19179_, new_n19180_, new_n19181_, new_n19182_, new_n19183_,
    new_n19184_, new_n19185_, new_n19186_, new_n19187_, new_n19188_,
    new_n19189_, new_n19190_, new_n19191_, new_n19192_, new_n19193_,
    new_n19194_, new_n19195_, new_n19196_, new_n19197_, new_n19198_,
    new_n19199_, new_n19200_, new_n19201_, new_n19202_, new_n19203_,
    new_n19204_, new_n19205_, new_n19206_, new_n19207_, new_n19208_,
    new_n19209_, new_n19210_, new_n19211_, new_n19212_, new_n19213_,
    new_n19214_, new_n19215_, new_n19216_, new_n19217_, new_n19218_,
    new_n19219_, new_n19220_, new_n19221_, new_n19222_, new_n19223_,
    new_n19224_, new_n19225_, new_n19226_, new_n19227_, new_n19228_,
    new_n19229_, new_n19230_, new_n19231_, new_n19232_, new_n19233_,
    new_n19234_, new_n19235_, new_n19236_, new_n19237_, new_n19238_,
    new_n19239_, new_n19240_, new_n19241_, new_n19242_, new_n19243_,
    new_n19244_, new_n19245_, new_n19246_, new_n19247_, new_n19248_,
    new_n19249_, new_n19250_, new_n19251_, new_n19252_, new_n19253_,
    new_n19254_, new_n19255_, new_n19256_, new_n19257_, new_n19258_,
    new_n19259_, new_n19260_, new_n19261_, new_n19262_, new_n19263_,
    new_n19264_, new_n19265_, new_n19266_, new_n19267_, new_n19268_,
    new_n19269_, new_n19270_, new_n19271_, new_n19272_, new_n19273_,
    new_n19274_, new_n19275_, new_n19276_, new_n19277_, new_n19278_,
    new_n19279_, new_n19280_, new_n19281_, new_n19282_, new_n19283_,
    new_n19284_, new_n19285_, new_n19286_, new_n19287_, new_n19288_,
    new_n19289_, new_n19290_, new_n19291_, new_n19292_, new_n19293_,
    new_n19294_, new_n19295_, new_n19296_, new_n19297_, new_n19298_,
    new_n19299_, new_n19301_, new_n19302_, new_n19303_, new_n19304_,
    new_n19305_, new_n19306_, new_n19307_, new_n19308_, new_n19309_,
    new_n19310_, new_n19311_, new_n19312_, new_n19313_, new_n19314_,
    new_n19315_, new_n19316_, new_n19317_, new_n19318_, new_n19319_,
    new_n19320_, new_n19321_, new_n19322_, new_n19323_, new_n19324_,
    new_n19325_, new_n19326_, new_n19327_, new_n19328_, new_n19329_,
    new_n19330_, new_n19331_, new_n19332_, new_n19333_, new_n19334_,
    new_n19335_, new_n19336_, new_n19337_, new_n19338_, new_n19339_,
    new_n19340_, new_n19341_, new_n19342_, new_n19343_, new_n19344_,
    new_n19345_, new_n19346_, new_n19347_, new_n19348_, new_n19349_,
    new_n19350_, new_n19351_, new_n19352_, new_n19353_, new_n19354_,
    new_n19355_, new_n19356_, new_n19357_, new_n19358_, new_n19359_,
    new_n19360_, new_n19361_, new_n19362_, new_n19363_, new_n19364_,
    new_n19365_, new_n19366_, new_n19367_, new_n19368_, new_n19369_,
    new_n19370_, new_n19371_, new_n19372_, new_n19373_, new_n19374_,
    new_n19375_, new_n19376_, new_n19377_, new_n19378_, new_n19379_,
    new_n19380_, new_n19381_, new_n19382_, new_n19383_, new_n19384_,
    new_n19385_, new_n19386_, new_n19387_, new_n19388_, new_n19389_,
    new_n19390_, new_n19391_, new_n19392_, new_n19393_, new_n19394_,
    new_n19395_, new_n19396_, new_n19397_, new_n19398_, new_n19399_,
    new_n19400_, new_n19401_, new_n19402_, new_n19403_, new_n19404_,
    new_n19405_, new_n19406_, new_n19407_, new_n19408_, new_n19409_,
    new_n19410_, new_n19411_, new_n19412_, new_n19413_, new_n19414_,
    new_n19415_, new_n19416_, new_n19417_, new_n19418_, new_n19419_,
    new_n19420_, new_n19421_, new_n19422_, new_n19423_, new_n19424_,
    new_n19425_, new_n19426_, new_n19427_, new_n19428_, new_n19429_,
    new_n19430_, new_n19431_, new_n19432_, new_n19433_, new_n19434_,
    new_n19435_, new_n19436_, new_n19437_, new_n19438_, new_n19439_,
    new_n19440_, new_n19441_, new_n19442_, new_n19443_, new_n19444_,
    new_n19445_, new_n19446_, new_n19447_, new_n19448_, new_n19449_,
    new_n19450_, new_n19451_, new_n19452_, new_n19453_, new_n19454_,
    new_n19455_, new_n19456_, new_n19457_, new_n19458_, new_n19459_,
    new_n19460_, new_n19461_, new_n19462_, new_n19463_, new_n19464_,
    new_n19465_, new_n19466_, new_n19467_, new_n19468_, new_n19469_,
    new_n19470_, new_n19471_, new_n19472_, new_n19473_, new_n19474_,
    new_n19475_, new_n19476_, new_n19477_, new_n19478_, new_n19479_,
    new_n19480_, new_n19481_, new_n19482_, new_n19483_, new_n19484_,
    new_n19485_, new_n19486_, new_n19487_, new_n19488_, new_n19489_,
    new_n19490_, new_n19491_, new_n19492_, new_n19493_, new_n19494_,
    new_n19495_, new_n19496_, new_n19497_, new_n19498_, new_n19499_,
    new_n19500_, new_n19501_, new_n19502_, new_n19503_, new_n19504_,
    new_n19505_, new_n19506_, new_n19507_, new_n19508_, new_n19509_,
    new_n19510_, new_n19511_, new_n19512_, new_n19513_, new_n19514_,
    new_n19515_, new_n19516_, new_n19517_, new_n19518_, new_n19519_,
    new_n19520_, new_n19521_, new_n19522_, new_n19523_, new_n19524_,
    new_n19525_, new_n19526_, new_n19527_, new_n19528_, new_n19529_,
    new_n19530_, new_n19531_, new_n19532_, new_n19533_, new_n19534_,
    new_n19535_, new_n19536_, new_n19537_, new_n19538_, new_n19539_,
    new_n19540_, new_n19541_, new_n19542_, new_n19543_, new_n19544_,
    new_n19545_, new_n19546_, new_n19547_, new_n19548_, new_n19549_,
    new_n19550_, new_n19551_, new_n19552_, new_n19553_, new_n19554_,
    new_n19555_, new_n19556_, new_n19557_, new_n19558_, new_n19559_,
    new_n19560_, new_n19561_, new_n19562_, new_n19563_, new_n19564_,
    new_n19565_, new_n19566_, new_n19567_, new_n19568_, new_n19569_,
    new_n19570_, new_n19572_, new_n19573_, new_n19574_, new_n19575_,
    new_n19576_, new_n19577_, new_n19578_, new_n19579_, new_n19580_,
    new_n19581_, new_n19582_, new_n19583_, new_n19584_, new_n19585_,
    new_n19586_, new_n19587_, new_n19588_, new_n19589_, new_n19590_,
    new_n19591_, new_n19592_, new_n19593_, new_n19594_, new_n19595_,
    new_n19596_, new_n19597_, new_n19598_, new_n19599_, new_n19600_,
    new_n19601_, new_n19602_, new_n19603_, new_n19604_, new_n19605_,
    new_n19606_, new_n19607_, new_n19608_, new_n19609_, new_n19610_,
    new_n19611_, new_n19612_, new_n19613_, new_n19614_, new_n19615_,
    new_n19616_, new_n19617_, new_n19618_, new_n19619_, new_n19620_,
    new_n19621_, new_n19622_, new_n19623_, new_n19624_, new_n19625_,
    new_n19626_, new_n19627_, new_n19628_, new_n19629_, new_n19630_,
    new_n19631_, new_n19632_, new_n19633_, new_n19634_, new_n19635_,
    new_n19636_, new_n19637_, new_n19638_, new_n19639_, new_n19640_,
    new_n19641_, new_n19642_, new_n19643_, new_n19644_, new_n19645_,
    new_n19646_, new_n19647_, new_n19648_, new_n19649_, new_n19650_,
    new_n19651_, new_n19652_, new_n19653_, new_n19654_, new_n19655_,
    new_n19656_, new_n19657_, new_n19658_, new_n19659_, new_n19660_,
    new_n19661_, new_n19662_, new_n19663_, new_n19664_, new_n19665_,
    new_n19666_, new_n19667_, new_n19668_, new_n19669_, new_n19670_,
    new_n19671_, new_n19672_, new_n19673_, new_n19674_, new_n19675_,
    new_n19676_, new_n19677_, new_n19678_, new_n19679_, new_n19680_,
    new_n19681_, new_n19682_, new_n19683_, new_n19684_, new_n19685_,
    new_n19686_, new_n19687_, new_n19688_, new_n19689_, new_n19690_,
    new_n19691_, new_n19692_, new_n19693_, new_n19694_, new_n19695_,
    new_n19696_, new_n19697_, new_n19698_, new_n19699_, new_n19700_,
    new_n19701_, new_n19702_, new_n19703_, new_n19704_, new_n19705_,
    new_n19706_, new_n19707_, new_n19708_, new_n19709_, new_n19710_,
    new_n19711_, new_n19712_, new_n19713_, new_n19714_, new_n19715_,
    new_n19716_, new_n19717_, new_n19718_, new_n19719_, new_n19720_,
    new_n19721_, new_n19722_, new_n19723_, new_n19724_, new_n19725_,
    new_n19726_, new_n19727_, new_n19728_, new_n19729_, new_n19730_,
    new_n19731_, new_n19732_, new_n19733_, new_n19734_, new_n19735_,
    new_n19736_, new_n19737_, new_n19738_, new_n19739_, new_n19740_,
    new_n19741_, new_n19742_, new_n19743_, new_n19744_, new_n19745_,
    new_n19746_, new_n19747_, new_n19748_, new_n19749_, new_n19750_,
    new_n19751_, new_n19752_, new_n19753_, new_n19754_, new_n19755_,
    new_n19756_, new_n19757_, new_n19758_, new_n19759_, new_n19760_,
    new_n19761_, new_n19762_, new_n19763_, new_n19764_, new_n19765_,
    new_n19766_, new_n19767_, new_n19768_, new_n19769_, new_n19770_,
    new_n19771_, new_n19772_, new_n19773_, new_n19774_, new_n19775_,
    new_n19776_, new_n19777_, new_n19778_, new_n19779_, new_n19780_,
    new_n19781_, new_n19782_, new_n19783_, new_n19784_, new_n19785_,
    new_n19786_, new_n19787_, new_n19788_, new_n19789_, new_n19790_,
    new_n19791_, new_n19792_, new_n19793_, new_n19794_, new_n19795_,
    new_n19796_, new_n19797_, new_n19798_, new_n19799_, new_n19800_,
    new_n19801_, new_n19802_, new_n19803_, new_n19804_, new_n19805_,
    new_n19806_, new_n19807_, new_n19808_, new_n19809_, new_n19810_,
    new_n19811_, new_n19812_, new_n19813_, new_n19814_, new_n19815_,
    new_n19816_, new_n19817_, new_n19818_, new_n19819_, new_n19820_,
    new_n19821_, new_n19822_, new_n19823_, new_n19824_, new_n19825_,
    new_n19826_, new_n19827_, new_n19828_, new_n19829_, new_n19830_,
    new_n19831_, new_n19832_, new_n19833_, new_n19834_, new_n19835_,
    new_n19836_, new_n19837_, new_n19838_, new_n19839_, new_n19840_,
    new_n19841_, new_n19842_, new_n19843_, new_n19844_, new_n19845_,
    new_n19846_, new_n19847_, new_n19848_, new_n19850_, new_n19851_,
    new_n19852_, new_n19853_, new_n19854_, new_n19855_, new_n19856_,
    new_n19857_, new_n19858_, new_n19859_, new_n19860_, new_n19861_,
    new_n19862_, new_n19863_, new_n19864_, new_n19865_, new_n19866_,
    new_n19867_, new_n19868_, new_n19869_, new_n19870_, new_n19871_,
    new_n19872_, new_n19873_, new_n19874_, new_n19875_, new_n19876_,
    new_n19877_, new_n19878_, new_n19879_, new_n19880_, new_n19881_,
    new_n19882_, new_n19883_, new_n19884_, new_n19885_, new_n19886_,
    new_n19887_, new_n19888_, new_n19889_, new_n19890_, new_n19891_,
    new_n19892_, new_n19893_, new_n19894_, new_n19895_, new_n19896_,
    new_n19897_, new_n19898_, new_n19899_, new_n19900_, new_n19901_,
    new_n19902_, new_n19903_, new_n19904_, new_n19905_, new_n19906_,
    new_n19907_, new_n19908_, new_n19909_, new_n19910_, new_n19911_,
    new_n19912_, new_n19913_, new_n19914_, new_n19915_, new_n19916_,
    new_n19917_, new_n19918_, new_n19919_, new_n19920_, new_n19921_,
    new_n19922_, new_n19923_, new_n19924_, new_n19925_, new_n19926_,
    new_n19927_, new_n19928_, new_n19929_, new_n19930_, new_n19931_,
    new_n19932_, new_n19933_, new_n19934_, new_n19935_, new_n19936_,
    new_n19937_, new_n19938_, new_n19939_, new_n19940_, new_n19941_,
    new_n19942_, new_n19943_, new_n19944_, new_n19945_, new_n19946_,
    new_n19947_, new_n19948_, new_n19949_, new_n19950_, new_n19951_,
    new_n19952_, new_n19953_, new_n19954_, new_n19955_, new_n19956_,
    new_n19957_, new_n19958_, new_n19959_, new_n19960_, new_n19961_,
    new_n19962_, new_n19963_, new_n19964_, new_n19965_, new_n19966_,
    new_n19967_, new_n19968_, new_n19969_, new_n19970_, new_n19971_,
    new_n19972_, new_n19973_, new_n19974_, new_n19975_, new_n19976_,
    new_n19977_, new_n19978_, new_n19979_, new_n19980_, new_n19981_,
    new_n19982_, new_n19983_, new_n19984_, new_n19985_, new_n19986_,
    new_n19987_, new_n19988_, new_n19989_, new_n19990_, new_n19991_,
    new_n19992_, new_n19993_, new_n19994_, new_n19995_, new_n19996_,
    new_n19997_, new_n19998_, new_n19999_, new_n20000_, new_n20001_,
    new_n20002_, new_n20003_, new_n20004_, new_n20005_, new_n20006_,
    new_n20007_, new_n20008_, new_n20009_, new_n20010_, new_n20011_,
    new_n20012_, new_n20013_, new_n20014_, new_n20015_, new_n20016_,
    new_n20017_, new_n20018_, new_n20019_, new_n20020_, new_n20021_,
    new_n20022_, new_n20023_, new_n20024_, new_n20025_, new_n20026_,
    new_n20027_, new_n20028_, new_n20029_, new_n20030_, new_n20031_,
    new_n20032_, new_n20033_, new_n20034_, new_n20035_, new_n20036_,
    new_n20037_, new_n20038_, new_n20039_, new_n20040_, new_n20041_,
    new_n20042_, new_n20043_, new_n20044_, new_n20045_, new_n20046_,
    new_n20047_, new_n20048_, new_n20049_, new_n20050_, new_n20051_,
    new_n20052_, new_n20053_, new_n20054_, new_n20055_, new_n20056_,
    new_n20057_, new_n20058_, new_n20059_, new_n20060_, new_n20061_,
    new_n20062_, new_n20063_, new_n20064_, new_n20065_, new_n20066_,
    new_n20067_, new_n20068_, new_n20069_, new_n20070_, new_n20071_,
    new_n20072_, new_n20073_, new_n20074_, new_n20075_, new_n20076_,
    new_n20077_, new_n20078_, new_n20079_, new_n20080_, new_n20081_,
    new_n20082_, new_n20083_, new_n20084_, new_n20085_, new_n20086_,
    new_n20087_, new_n20088_, new_n20089_, new_n20090_, new_n20091_,
    new_n20092_, new_n20093_, new_n20094_, new_n20095_, new_n20096_,
    new_n20097_, new_n20098_, new_n20099_, new_n20100_, new_n20101_,
    new_n20102_, new_n20103_, new_n20104_, new_n20105_, new_n20106_,
    new_n20107_, new_n20108_, new_n20109_, new_n20110_, new_n20111_,
    new_n20112_, new_n20113_, new_n20114_, new_n20115_, new_n20116_,
    new_n20117_, new_n20118_, new_n20119_, new_n20120_, new_n20121_,
    new_n20122_, new_n20123_, new_n20124_, new_n20125_, new_n20126_,
    new_n20128_, new_n20129_, new_n20130_, new_n20131_, new_n20132_,
    new_n20133_, new_n20134_, new_n20135_, new_n20136_, new_n20137_,
    new_n20138_, new_n20139_, new_n20140_, new_n20141_, new_n20142_,
    new_n20143_, new_n20144_, new_n20145_, new_n20146_, new_n20147_,
    new_n20148_, new_n20149_, new_n20150_, new_n20151_, new_n20152_,
    new_n20153_, new_n20154_, new_n20155_, new_n20156_, new_n20157_,
    new_n20158_, new_n20159_, new_n20160_, new_n20161_, new_n20162_,
    new_n20163_, new_n20164_, new_n20165_, new_n20166_, new_n20167_,
    new_n20168_, new_n20169_, new_n20170_, new_n20171_, new_n20172_,
    new_n20173_, new_n20174_, new_n20175_, new_n20176_, new_n20177_,
    new_n20178_, new_n20179_, new_n20180_, new_n20181_, new_n20182_,
    new_n20183_, new_n20184_, new_n20185_, new_n20186_, new_n20187_,
    new_n20188_, new_n20189_, new_n20190_, new_n20191_, new_n20192_,
    new_n20193_, new_n20194_, new_n20195_, new_n20196_, new_n20197_,
    new_n20198_, new_n20199_, new_n20200_, new_n20201_, new_n20202_,
    new_n20203_, new_n20204_, new_n20205_, new_n20206_, new_n20207_,
    new_n20208_, new_n20209_, new_n20210_, new_n20211_, new_n20212_,
    new_n20213_, new_n20214_, new_n20215_, new_n20216_, new_n20217_,
    new_n20218_, new_n20219_, new_n20220_, new_n20221_, new_n20222_,
    new_n20223_, new_n20224_, new_n20225_, new_n20226_, new_n20227_,
    new_n20228_, new_n20229_, new_n20230_, new_n20231_, new_n20232_,
    new_n20233_, new_n20234_, new_n20235_, new_n20236_, new_n20237_,
    new_n20238_, new_n20239_, new_n20240_, new_n20241_, new_n20242_,
    new_n20243_, new_n20244_, new_n20245_, new_n20246_, new_n20247_,
    new_n20248_, new_n20249_, new_n20250_, new_n20251_, new_n20252_,
    new_n20253_, new_n20254_, new_n20255_, new_n20256_, new_n20257_,
    new_n20258_, new_n20259_, new_n20260_, new_n20261_, new_n20262_,
    new_n20263_, new_n20264_, new_n20265_, new_n20266_, new_n20267_,
    new_n20268_, new_n20269_, new_n20270_, new_n20271_, new_n20272_,
    new_n20273_, new_n20274_, new_n20275_, new_n20276_, new_n20277_,
    new_n20278_, new_n20279_, new_n20280_, new_n20281_, new_n20282_,
    new_n20283_, new_n20284_, new_n20285_, new_n20286_, new_n20287_,
    new_n20288_, new_n20289_, new_n20290_, new_n20291_, new_n20292_,
    new_n20293_, new_n20294_, new_n20295_, new_n20296_, new_n20297_,
    new_n20298_, new_n20299_, new_n20300_, new_n20301_, new_n20302_,
    new_n20303_, new_n20304_, new_n20305_, new_n20306_, new_n20307_,
    new_n20308_, new_n20309_, new_n20310_, new_n20311_, new_n20312_,
    new_n20313_, new_n20314_, new_n20315_, new_n20316_, new_n20317_,
    new_n20318_, new_n20319_, new_n20320_, new_n20321_, new_n20322_,
    new_n20323_, new_n20324_, new_n20325_, new_n20326_, new_n20327_,
    new_n20328_, new_n20329_, new_n20330_, new_n20331_, new_n20332_,
    new_n20333_, new_n20334_, new_n20335_, new_n20336_, new_n20337_,
    new_n20338_, new_n20339_, new_n20340_, new_n20341_, new_n20342_,
    new_n20343_, new_n20344_, new_n20345_, new_n20346_, new_n20347_,
    new_n20348_, new_n20349_, new_n20350_, new_n20351_, new_n20352_,
    new_n20353_, new_n20354_, new_n20355_, new_n20356_, new_n20357_,
    new_n20358_, new_n20359_, new_n20360_, new_n20361_, new_n20362_,
    new_n20363_, new_n20364_, new_n20365_, new_n20366_, new_n20367_,
    new_n20368_, new_n20369_, new_n20370_, new_n20371_, new_n20372_,
    new_n20373_, new_n20374_, new_n20375_, new_n20376_, new_n20377_,
    new_n20378_, new_n20379_, new_n20380_, new_n20381_, new_n20382_,
    new_n20383_, new_n20384_, new_n20385_, new_n20386_, new_n20387_,
    new_n20388_, new_n20389_, new_n20390_, new_n20391_, new_n20392_,
    new_n20393_, new_n20394_, new_n20395_, new_n20396_, new_n20397_,
    new_n20398_, new_n20399_, new_n20400_, new_n20401_, new_n20402_,
    new_n20403_, new_n20404_, new_n20405_, new_n20406_, new_n20407_,
    new_n20409_, new_n20410_, new_n20411_, new_n20412_, new_n20413_,
    new_n20414_, new_n20415_, new_n20416_, new_n20417_, new_n20418_,
    new_n20419_, new_n20420_, new_n20421_, new_n20422_, new_n20423_,
    new_n20424_, new_n20425_, new_n20426_, new_n20427_, new_n20428_,
    new_n20429_, new_n20430_, new_n20431_, new_n20432_, new_n20433_,
    new_n20434_, new_n20435_, new_n20436_, new_n20437_, new_n20438_,
    new_n20439_, new_n20440_, new_n20441_, new_n20442_, new_n20443_,
    new_n20444_, new_n20445_, new_n20446_, new_n20447_, new_n20448_,
    new_n20449_, new_n20450_, new_n20451_, new_n20452_, new_n20453_,
    new_n20454_, new_n20455_, new_n20456_, new_n20457_, new_n20458_,
    new_n20459_, new_n20460_, new_n20461_, new_n20462_, new_n20463_,
    new_n20464_, new_n20465_, new_n20466_, new_n20467_, new_n20468_,
    new_n20469_, new_n20470_, new_n20471_, new_n20472_, new_n20473_,
    new_n20474_, new_n20475_, new_n20476_, new_n20477_, new_n20478_,
    new_n20479_, new_n20480_, new_n20481_, new_n20482_, new_n20483_,
    new_n20484_, new_n20485_, new_n20486_, new_n20487_, new_n20488_,
    new_n20489_, new_n20490_, new_n20491_, new_n20492_, new_n20493_,
    new_n20494_, new_n20495_, new_n20496_, new_n20497_, new_n20498_,
    new_n20499_, new_n20500_, new_n20501_, new_n20502_, new_n20503_,
    new_n20504_, new_n20505_, new_n20506_, new_n20507_, new_n20508_,
    new_n20509_, new_n20510_, new_n20511_, new_n20512_, new_n20513_,
    new_n20514_, new_n20515_, new_n20516_, new_n20517_, new_n20518_,
    new_n20519_, new_n20520_, new_n20521_, new_n20522_, new_n20523_,
    new_n20524_, new_n20525_, new_n20526_, new_n20527_, new_n20528_,
    new_n20529_, new_n20530_, new_n20531_, new_n20532_, new_n20533_,
    new_n20534_, new_n20535_, new_n20536_, new_n20537_, new_n20538_,
    new_n20539_, new_n20540_, new_n20541_, new_n20542_, new_n20543_,
    new_n20544_, new_n20545_, new_n20546_, new_n20547_, new_n20548_,
    new_n20549_, new_n20550_, new_n20551_, new_n20552_, new_n20553_,
    new_n20554_, new_n20555_, new_n20556_, new_n20557_, new_n20558_,
    new_n20559_, new_n20560_, new_n20561_, new_n20562_, new_n20563_,
    new_n20564_, new_n20565_, new_n20566_, new_n20567_, new_n20568_,
    new_n20569_, new_n20570_, new_n20571_, new_n20572_, new_n20573_,
    new_n20574_, new_n20575_, new_n20576_, new_n20577_, new_n20578_,
    new_n20579_, new_n20580_, new_n20581_, new_n20582_, new_n20583_,
    new_n20584_, new_n20585_, new_n20586_, new_n20587_, new_n20588_,
    new_n20589_, new_n20590_, new_n20591_, new_n20592_, new_n20593_,
    new_n20594_, new_n20595_, new_n20596_, new_n20597_, new_n20598_,
    new_n20599_, new_n20600_, new_n20601_, new_n20602_, new_n20603_,
    new_n20604_, new_n20605_, new_n20606_, new_n20607_, new_n20608_,
    new_n20609_, new_n20610_, new_n20611_, new_n20612_, new_n20613_,
    new_n20614_, new_n20615_, new_n20616_, new_n20617_, new_n20618_,
    new_n20619_, new_n20620_, new_n20621_, new_n20622_, new_n20623_,
    new_n20624_, new_n20625_, new_n20626_, new_n20627_, new_n20628_,
    new_n20629_, new_n20630_, new_n20631_, new_n20632_, new_n20633_,
    new_n20634_, new_n20635_, new_n20636_, new_n20637_, new_n20638_,
    new_n20639_, new_n20640_, new_n20641_, new_n20642_, new_n20643_,
    new_n20644_, new_n20645_, new_n20646_, new_n20647_, new_n20648_,
    new_n20649_, new_n20650_, new_n20651_, new_n20652_, new_n20653_,
    new_n20654_, new_n20655_, new_n20656_, new_n20657_, new_n20658_,
    new_n20659_, new_n20660_, new_n20661_, new_n20662_, new_n20663_,
    new_n20664_, new_n20665_, new_n20666_, new_n20667_, new_n20668_,
    new_n20669_, new_n20670_, new_n20671_, new_n20672_, new_n20673_,
    new_n20674_, new_n20675_, new_n20676_, new_n20677_, new_n20678_,
    new_n20679_, new_n20680_, new_n20681_, new_n20682_, new_n20683_,
    new_n20685_, new_n20686_, new_n20687_, new_n20688_, new_n20689_,
    new_n20690_, new_n20691_, new_n20692_, new_n20693_, new_n20694_,
    new_n20695_, new_n20696_, new_n20697_, new_n20698_, new_n20699_,
    new_n20700_, new_n20701_, new_n20702_, new_n20703_, new_n20704_,
    new_n20705_, new_n20706_, new_n20707_, new_n20708_, new_n20709_,
    new_n20710_, new_n20711_, new_n20712_, new_n20713_, new_n20714_,
    new_n20715_, new_n20716_, new_n20717_, new_n20718_, new_n20719_,
    new_n20720_, new_n20721_, new_n20722_, new_n20723_, new_n20724_,
    new_n20725_, new_n20726_, new_n20727_, new_n20728_, new_n20729_,
    new_n20730_, new_n20731_, new_n20732_, new_n20733_, new_n20734_,
    new_n20735_, new_n20736_, new_n20737_, new_n20738_, new_n20739_,
    new_n20740_, new_n20741_, new_n20742_, new_n20743_, new_n20744_,
    new_n20745_, new_n20746_, new_n20747_, new_n20748_, new_n20749_,
    new_n20750_, new_n20751_, new_n20752_, new_n20753_, new_n20754_,
    new_n20755_, new_n20756_, new_n20757_, new_n20758_, new_n20759_,
    new_n20760_, new_n20761_, new_n20762_, new_n20763_, new_n20764_,
    new_n20765_, new_n20766_, new_n20767_, new_n20768_, new_n20769_,
    new_n20770_, new_n20771_, new_n20772_, new_n20773_, new_n20774_,
    new_n20775_, new_n20776_, new_n20777_, new_n20778_, new_n20779_,
    new_n20780_, new_n20781_, new_n20782_, new_n20783_, new_n20784_,
    new_n20785_, new_n20786_, new_n20787_, new_n20788_, new_n20789_,
    new_n20790_, new_n20791_, new_n20792_, new_n20793_, new_n20794_,
    new_n20795_, new_n20796_, new_n20797_, new_n20798_, new_n20799_,
    new_n20800_, new_n20801_, new_n20802_, new_n20803_, new_n20804_,
    new_n20805_, new_n20806_, new_n20807_, new_n20808_, new_n20809_,
    new_n20810_, new_n20811_, new_n20812_, new_n20813_, new_n20814_,
    new_n20815_, new_n20816_, new_n20817_, new_n20818_, new_n20819_,
    new_n20820_, new_n20821_, new_n20822_, new_n20823_, new_n20824_,
    new_n20825_, new_n20826_, new_n20827_, new_n20828_, new_n20829_,
    new_n20830_, new_n20831_, new_n20832_, new_n20833_, new_n20834_,
    new_n20835_, new_n20836_, new_n20837_, new_n20838_, new_n20839_,
    new_n20840_, new_n20841_, new_n20842_, new_n20843_, new_n20844_,
    new_n20845_, new_n20846_, new_n20847_, new_n20848_, new_n20849_,
    new_n20850_, new_n20851_, new_n20852_, new_n20853_, new_n20854_,
    new_n20855_, new_n20856_, new_n20857_, new_n20858_, new_n20859_,
    new_n20860_, new_n20861_, new_n20862_, new_n20863_, new_n20864_,
    new_n20865_, new_n20866_, new_n20867_, new_n20868_, new_n20869_,
    new_n20870_, new_n20871_, new_n20872_, new_n20873_, new_n20874_,
    new_n20875_, new_n20876_, new_n20877_, new_n20878_, new_n20879_,
    new_n20880_, new_n20881_, new_n20882_, new_n20883_, new_n20884_,
    new_n20885_, new_n20886_, new_n20887_, new_n20888_, new_n20889_,
    new_n20890_, new_n20891_, new_n20892_, new_n20893_, new_n20894_,
    new_n20895_, new_n20896_, new_n20897_, new_n20898_, new_n20899_,
    new_n20900_, new_n20901_, new_n20902_, new_n20903_, new_n20904_,
    new_n20905_, new_n20906_, new_n20907_, new_n20908_, new_n20909_,
    new_n20910_, new_n20911_, new_n20912_, new_n20913_, new_n20914_,
    new_n20915_, new_n20916_, new_n20917_, new_n20918_, new_n20919_,
    new_n20920_, new_n20921_, new_n20922_, new_n20923_, new_n20924_,
    new_n20925_, new_n20926_, new_n20927_, new_n20928_, new_n20929_,
    new_n20930_, new_n20931_, new_n20932_, new_n20933_, new_n20934_,
    new_n20935_, new_n20936_, new_n20937_, new_n20938_, new_n20939_,
    new_n20940_, new_n20941_, new_n20942_, new_n20943_, new_n20944_,
    new_n20945_, new_n20946_, new_n20947_, new_n20948_, new_n20949_,
    new_n20950_, new_n20951_, new_n20952_, new_n20953_, new_n20954_,
    new_n20955_, new_n20956_, new_n20957_, new_n20958_, new_n20959_,
    new_n20961_, new_n20962_, new_n20963_, new_n20964_, new_n20965_,
    new_n20966_, new_n20967_, new_n20968_, new_n20969_, new_n20970_,
    new_n20971_, new_n20972_, new_n20973_, new_n20974_, new_n20975_,
    new_n20976_, new_n20977_, new_n20978_, new_n20979_, new_n20980_,
    new_n20981_, new_n20982_, new_n20983_, new_n20984_, new_n20985_,
    new_n20986_, new_n20987_, new_n20988_, new_n20989_, new_n20990_,
    new_n20991_, new_n20992_, new_n20993_, new_n20994_, new_n20995_,
    new_n20996_, new_n20997_, new_n20998_, new_n20999_, new_n21000_,
    new_n21001_, new_n21002_, new_n21003_, new_n21004_, new_n21005_,
    new_n21006_, new_n21007_, new_n21008_, new_n21009_, new_n21010_,
    new_n21011_, new_n21012_, new_n21013_, new_n21014_, new_n21015_,
    new_n21016_, new_n21017_, new_n21018_, new_n21019_, new_n21020_,
    new_n21021_, new_n21022_, new_n21023_, new_n21024_, new_n21025_,
    new_n21026_, new_n21027_, new_n21028_, new_n21029_, new_n21030_,
    new_n21031_, new_n21032_, new_n21033_, new_n21034_, new_n21035_,
    new_n21036_, new_n21037_, new_n21038_, new_n21039_, new_n21040_,
    new_n21041_, new_n21042_, new_n21043_, new_n21044_, new_n21045_,
    new_n21046_, new_n21047_, new_n21048_, new_n21049_, new_n21050_,
    new_n21051_, new_n21052_, new_n21053_, new_n21054_, new_n21055_,
    new_n21056_, new_n21057_, new_n21058_, new_n21059_, new_n21060_,
    new_n21061_, new_n21062_, new_n21063_, new_n21064_, new_n21065_,
    new_n21066_, new_n21067_, new_n21068_, new_n21069_, new_n21070_,
    new_n21071_, new_n21072_, new_n21073_, new_n21074_, new_n21075_,
    new_n21076_, new_n21077_, new_n21078_, new_n21079_, new_n21080_,
    new_n21081_, new_n21082_, new_n21083_, new_n21084_, new_n21085_,
    new_n21086_, new_n21087_, new_n21088_, new_n21089_, new_n21090_,
    new_n21091_, new_n21092_, new_n21093_, new_n21094_, new_n21095_,
    new_n21096_, new_n21097_, new_n21098_, new_n21099_, new_n21100_,
    new_n21101_, new_n21102_, new_n21103_, new_n21104_, new_n21105_,
    new_n21106_, new_n21107_, new_n21108_, new_n21109_, new_n21110_,
    new_n21111_, new_n21112_, new_n21113_, new_n21114_, new_n21115_,
    new_n21116_, new_n21117_, new_n21118_, new_n21119_, new_n21120_,
    new_n21121_, new_n21122_, new_n21123_, new_n21124_, new_n21125_,
    new_n21126_, new_n21127_, new_n21128_, new_n21129_, new_n21130_,
    new_n21131_, new_n21132_, new_n21133_, new_n21134_, new_n21135_,
    new_n21136_, new_n21137_, new_n21138_, new_n21139_, new_n21140_,
    new_n21141_, new_n21142_, new_n21143_, new_n21144_, new_n21145_,
    new_n21146_, new_n21147_, new_n21148_, new_n21149_, new_n21150_,
    new_n21151_, new_n21152_, new_n21153_, new_n21154_, new_n21155_,
    new_n21156_, new_n21157_, new_n21158_, new_n21159_, new_n21160_,
    new_n21161_, new_n21162_, new_n21163_, new_n21164_, new_n21165_,
    new_n21166_, new_n21167_, new_n21168_, new_n21169_, new_n21170_,
    new_n21171_, new_n21172_, new_n21173_, new_n21174_, new_n21175_,
    new_n21176_, new_n21177_, new_n21178_, new_n21179_, new_n21180_,
    new_n21181_, new_n21182_, new_n21183_, new_n21184_, new_n21185_,
    new_n21186_, new_n21187_, new_n21188_, new_n21189_, new_n21190_,
    new_n21191_, new_n21192_, new_n21193_, new_n21194_, new_n21195_,
    new_n21196_, new_n21197_, new_n21198_, new_n21199_, new_n21200_,
    new_n21201_, new_n21202_, new_n21203_, new_n21204_, new_n21205_,
    new_n21206_, new_n21207_, new_n21208_, new_n21209_, new_n21210_,
    new_n21211_, new_n21212_, new_n21213_, new_n21214_, new_n21215_,
    new_n21216_, new_n21217_, new_n21218_, new_n21219_, new_n21220_,
    new_n21221_, new_n21222_, new_n21223_, new_n21224_, new_n21225_,
    new_n21226_, new_n21227_, new_n21228_, new_n21229_, new_n21230_,
    new_n21231_, new_n21232_, new_n21233_, new_n21234_, new_n21235_,
    new_n21237_, new_n21238_, new_n21239_, new_n21240_, new_n21241_,
    new_n21242_, new_n21243_, new_n21244_, new_n21245_, new_n21246_,
    new_n21247_, new_n21248_, new_n21249_, new_n21250_, new_n21251_,
    new_n21252_, new_n21253_, new_n21254_, new_n21255_, new_n21256_,
    new_n21257_, new_n21258_, new_n21259_, new_n21260_, new_n21261_,
    new_n21262_, new_n21263_, new_n21264_, new_n21265_, new_n21266_,
    new_n21267_, new_n21268_, new_n21269_, new_n21270_, new_n21271_,
    new_n21272_, new_n21273_, new_n21274_, new_n21275_, new_n21276_,
    new_n21277_, new_n21278_, new_n21279_, new_n21280_, new_n21281_,
    new_n21282_, new_n21283_, new_n21284_, new_n21285_, new_n21286_,
    new_n21287_, new_n21288_, new_n21289_, new_n21290_, new_n21291_,
    new_n21292_, new_n21293_, new_n21294_, new_n21295_, new_n21296_,
    new_n21297_, new_n21298_, new_n21299_, new_n21300_, new_n21301_,
    new_n21302_, new_n21303_, new_n21304_, new_n21305_, new_n21306_,
    new_n21307_, new_n21308_, new_n21309_, new_n21310_, new_n21311_,
    new_n21312_, new_n21313_, new_n21314_, new_n21315_, new_n21316_,
    new_n21317_, new_n21318_, new_n21319_, new_n21320_, new_n21321_,
    new_n21322_, new_n21323_, new_n21324_, new_n21325_, new_n21326_,
    new_n21327_, new_n21328_, new_n21329_, new_n21330_, new_n21331_,
    new_n21332_, new_n21333_, new_n21334_, new_n21335_, new_n21336_,
    new_n21337_, new_n21338_, new_n21339_, new_n21340_, new_n21341_,
    new_n21342_, new_n21343_, new_n21344_, new_n21345_, new_n21346_,
    new_n21347_, new_n21348_, new_n21349_, new_n21350_, new_n21351_,
    new_n21352_, new_n21353_, new_n21354_, new_n21355_, new_n21356_,
    new_n21357_, new_n21358_, new_n21359_, new_n21360_, new_n21361_,
    new_n21362_, new_n21363_, new_n21364_, new_n21365_, new_n21366_,
    new_n21367_, new_n21368_, new_n21369_, new_n21370_, new_n21371_,
    new_n21372_, new_n21373_, new_n21374_, new_n21375_, new_n21376_,
    new_n21377_, new_n21378_, new_n21379_, new_n21380_, new_n21381_,
    new_n21382_, new_n21383_, new_n21384_, new_n21385_, new_n21386_,
    new_n21387_, new_n21388_, new_n21389_, new_n21390_, new_n21391_,
    new_n21392_, new_n21393_, new_n21394_, new_n21395_, new_n21396_,
    new_n21397_, new_n21398_, new_n21399_, new_n21400_, new_n21401_,
    new_n21402_, new_n21403_, new_n21404_, new_n21405_, new_n21406_,
    new_n21407_, new_n21408_, new_n21409_, new_n21410_, new_n21411_,
    new_n21412_, new_n21413_, new_n21414_, new_n21415_, new_n21416_,
    new_n21417_, new_n21418_, new_n21419_, new_n21420_, new_n21421_,
    new_n21422_, new_n21423_, new_n21424_, new_n21425_, new_n21426_,
    new_n21427_, new_n21428_, new_n21429_, new_n21430_, new_n21431_,
    new_n21432_, new_n21433_, new_n21434_, new_n21435_, new_n21436_,
    new_n21437_, new_n21438_, new_n21439_, new_n21440_, new_n21441_,
    new_n21442_, new_n21443_, new_n21444_, new_n21445_, new_n21446_,
    new_n21447_, new_n21448_, new_n21449_, new_n21450_, new_n21451_,
    new_n21452_, new_n21453_, new_n21454_, new_n21455_, new_n21456_,
    new_n21457_, new_n21458_, new_n21459_, new_n21460_, new_n21461_,
    new_n21462_, new_n21463_, new_n21464_, new_n21465_, new_n21466_,
    new_n21467_, new_n21468_, new_n21469_, new_n21470_, new_n21471_,
    new_n21472_, new_n21473_, new_n21474_, new_n21475_, new_n21476_,
    new_n21477_, new_n21478_, new_n21479_, new_n21480_, new_n21481_,
    new_n21482_, new_n21483_, new_n21484_, new_n21485_, new_n21486_,
    new_n21487_, new_n21488_, new_n21489_, new_n21490_, new_n21491_,
    new_n21492_, new_n21493_, new_n21494_, new_n21495_, new_n21496_,
    new_n21497_, new_n21498_, new_n21499_, new_n21500_, new_n21501_,
    new_n21502_, new_n21503_, new_n21504_, new_n21505_, new_n21507_,
    new_n21508_, new_n21509_, new_n21510_, new_n21511_, new_n21512_,
    new_n21513_, new_n21514_, new_n21515_, new_n21516_, new_n21517_,
    new_n21518_, new_n21519_, new_n21520_, new_n21521_, new_n21522_,
    new_n21523_, new_n21524_, new_n21525_, new_n21526_, new_n21527_,
    new_n21528_, new_n21529_, new_n21530_, new_n21531_, new_n21532_,
    new_n21533_, new_n21534_, new_n21535_, new_n21536_, new_n21537_,
    new_n21538_, new_n21539_, new_n21540_, new_n21541_, new_n21542_,
    new_n21543_, new_n21544_, new_n21545_, new_n21546_, new_n21547_,
    new_n21548_, new_n21549_, new_n21550_, new_n21551_, new_n21552_,
    new_n21553_, new_n21554_, new_n21555_, new_n21556_, new_n21557_,
    new_n21558_, new_n21559_, new_n21560_, new_n21561_, new_n21562_,
    new_n21563_, new_n21564_, new_n21565_, new_n21566_, new_n21567_,
    new_n21568_, new_n21569_, new_n21570_, new_n21571_, new_n21572_,
    new_n21573_, new_n21574_, new_n21575_, new_n21576_, new_n21577_,
    new_n21578_, new_n21579_, new_n21580_, new_n21581_, new_n21582_,
    new_n21583_, new_n21584_, new_n21585_, new_n21586_, new_n21587_,
    new_n21588_, new_n21589_, new_n21590_, new_n21591_, new_n21592_,
    new_n21593_, new_n21594_, new_n21595_, new_n21596_, new_n21597_,
    new_n21598_, new_n21599_, new_n21600_, new_n21601_, new_n21602_,
    new_n21603_, new_n21604_, new_n21605_, new_n21606_, new_n21607_,
    new_n21608_, new_n21609_, new_n21610_, new_n21611_, new_n21612_,
    new_n21613_, new_n21614_, new_n21615_, new_n21616_, new_n21617_,
    new_n21618_, new_n21619_, new_n21620_, new_n21621_, new_n21622_,
    new_n21623_, new_n21624_, new_n21625_, new_n21626_, new_n21627_,
    new_n21628_, new_n21629_, new_n21630_, new_n21631_, new_n21632_,
    new_n21633_, new_n21634_, new_n21635_, new_n21636_, new_n21637_,
    new_n21638_, new_n21639_, new_n21640_, new_n21641_, new_n21642_,
    new_n21643_, new_n21644_, new_n21645_, new_n21646_, new_n21647_,
    new_n21648_, new_n21649_, new_n21650_, new_n21651_, new_n21652_,
    new_n21653_, new_n21654_, new_n21655_, new_n21656_, new_n21657_,
    new_n21658_, new_n21659_, new_n21660_, new_n21661_, new_n21662_,
    new_n21663_, new_n21664_, new_n21665_, new_n21666_, new_n21667_,
    new_n21668_, new_n21669_, new_n21670_, new_n21671_, new_n21672_,
    new_n21673_, new_n21674_, new_n21675_, new_n21676_, new_n21677_,
    new_n21678_, new_n21679_, new_n21680_, new_n21681_, new_n21682_,
    new_n21683_, new_n21684_, new_n21685_, new_n21686_, new_n21687_,
    new_n21688_, new_n21689_, new_n21690_, new_n21691_, new_n21692_,
    new_n21693_, new_n21694_, new_n21695_, new_n21696_, new_n21697_,
    new_n21698_, new_n21699_, new_n21700_, new_n21701_, new_n21702_,
    new_n21703_, new_n21704_, new_n21705_, new_n21706_, new_n21707_,
    new_n21708_, new_n21709_, new_n21710_, new_n21711_, new_n21712_,
    new_n21713_, new_n21714_, new_n21715_, new_n21716_, new_n21717_,
    new_n21718_, new_n21719_, new_n21720_, new_n21721_, new_n21722_,
    new_n21723_, new_n21724_, new_n21725_, new_n21726_, new_n21727_,
    new_n21728_, new_n21729_, new_n21730_, new_n21731_, new_n21732_,
    new_n21733_, new_n21734_, new_n21735_, new_n21736_, new_n21737_,
    new_n21738_, new_n21739_, new_n21740_, new_n21741_, new_n21742_,
    new_n21743_, new_n21744_, new_n21745_, new_n21746_, new_n21747_,
    new_n21748_, new_n21749_, new_n21750_, new_n21751_, new_n21752_,
    new_n21753_, new_n21754_, new_n21755_, new_n21756_, new_n21757_,
    new_n21758_, new_n21759_, new_n21760_, new_n21761_, new_n21762_,
    new_n21763_, new_n21764_, new_n21765_, new_n21766_, new_n21767_,
    new_n21768_, new_n21769_, new_n21771_, new_n21772_, new_n21773_,
    new_n21774_, new_n21775_, new_n21776_, new_n21777_, new_n21778_,
    new_n21779_, new_n21780_, new_n21781_, new_n21782_, new_n21783_,
    new_n21784_, new_n21785_, new_n21786_, new_n21787_, new_n21788_,
    new_n21789_, new_n21790_, new_n21791_, new_n21792_, new_n21793_,
    new_n21794_, new_n21795_, new_n21796_, new_n21797_, new_n21798_,
    new_n21799_, new_n21800_, new_n21801_, new_n21802_, new_n21804_,
    new_n21805_, new_n21806_, new_n21807_, new_n21808_, new_n21809_,
    new_n21810_, new_n21811_, new_n21812_, new_n21813_, new_n21814_,
    new_n21815_, new_n21816_, new_n21817_, new_n21818_, new_n21819_,
    new_n21820_, new_n21821_, new_n21822_, new_n21823_, new_n21824_,
    new_n21825_, new_n21826_, new_n21827_, new_n21828_, new_n21829_,
    new_n21830_, new_n21831_, new_n21832_, new_n21833_, new_n21834_,
    new_n21835_, new_n21836_, new_n21837_, new_n21838_, new_n21839_,
    new_n21840_, new_n21841_, new_n21842_, new_n21843_, new_n21844_,
    new_n21846_, new_n21847_, new_n21848_, new_n21849_, new_n21850_,
    new_n21851_, new_n21852_, new_n21853_, new_n21854_, new_n21855_,
    new_n21856_, new_n21857_, new_n21858_, new_n21859_, new_n21860_,
    new_n21861_, new_n21862_, new_n21863_, new_n21864_, new_n21865_,
    new_n21866_, new_n21867_, new_n21868_, new_n21869_, new_n21870_,
    new_n21871_, new_n21872_, new_n21873_, new_n21874_, new_n21875_,
    new_n21876_, new_n21877_, new_n21878_, new_n21879_, new_n21881_,
    new_n21882_, new_n21883_, new_n21884_, new_n21885_, new_n21886_,
    new_n21887_, new_n21888_, new_n21889_, new_n21890_, new_n21891_,
    new_n21892_, new_n21893_, new_n21894_, new_n21895_, new_n21896_,
    new_n21897_, new_n21898_, new_n21899_, new_n21900_, new_n21901_,
    new_n21902_, new_n21903_, new_n21904_, new_n21905_, new_n21906_,
    new_n21907_, new_n21908_, new_n21909_, new_n21910_, new_n21911_,
    new_n21912_, new_n21913_, new_n21914_, new_n21915_, new_n21916_,
    new_n21917_, new_n21918_, new_n21919_, new_n21920_, new_n21921_,
    new_n21922_, new_n21923_, new_n21924_, new_n21925_, new_n21926_,
    new_n21927_, new_n21928_, new_n21929_, new_n21930_, new_n21931_,
    new_n21932_, new_n21933_, new_n21934_, new_n21935_, new_n21936_,
    new_n21937_, new_n21938_, new_n21939_, new_n21940_, new_n21941_,
    new_n21942_, new_n21943_, new_n21944_, new_n21945_, new_n21946_,
    new_n21947_, new_n21948_, new_n21949_, new_n21950_, new_n21951_,
    new_n21952_, new_n21953_, new_n21954_, new_n21955_, new_n21956_,
    new_n21957_, new_n21958_, new_n21959_, new_n21960_, new_n21961_,
    new_n21962_, new_n21963_, new_n21964_, new_n21965_, new_n21966_,
    new_n21967_, new_n21968_, new_n21969_, new_n21970_, new_n21971_,
    new_n21972_, new_n21973_, new_n21974_, new_n21975_, new_n21976_,
    new_n21977_, new_n21978_, new_n21979_, new_n21980_, new_n21981_,
    new_n21982_, new_n21983_, new_n21984_, new_n21985_, new_n21986_,
    new_n21987_, new_n21988_, new_n21989_, new_n21990_, new_n21991_,
    new_n21992_, new_n21993_, new_n21994_, new_n21995_, new_n21996_,
    new_n21997_, new_n21998_, new_n21999_, new_n22000_, new_n22001_,
    new_n22002_, new_n22003_, new_n22004_, new_n22005_, new_n22006_,
    new_n22007_, new_n22008_, new_n22009_, new_n22010_, new_n22011_,
    new_n22012_, new_n22013_, new_n22014_, new_n22015_, new_n22016_,
    new_n22017_, new_n22018_, new_n22019_, new_n22020_, new_n22021_,
    new_n22022_, new_n22023_, new_n22024_, new_n22025_, new_n22026_,
    new_n22027_, new_n22028_, new_n22029_, new_n22030_, new_n22031_,
    new_n22032_, new_n22033_, new_n22034_, new_n22035_, new_n22036_,
    new_n22037_, new_n22038_, new_n22039_, new_n22040_, new_n22041_,
    new_n22042_, new_n22043_, new_n22044_, new_n22045_, new_n22046_,
    new_n22047_, new_n22048_, new_n22049_, new_n22050_, new_n22051_,
    new_n22052_, new_n22053_, new_n22054_, new_n22055_, new_n22056_,
    new_n22057_, new_n22058_, new_n22059_, new_n22060_, new_n22061_,
    new_n22062_, new_n22063_, new_n22064_, new_n22065_, new_n22066_,
    new_n22067_, new_n22068_, new_n22069_, new_n22070_, new_n22071_,
    new_n22072_, new_n22073_, new_n22074_, new_n22075_, new_n22076_,
    new_n22077_, new_n22078_, new_n22079_, new_n22080_, new_n22081_,
    new_n22082_, new_n22083_, new_n22084_, new_n22085_, new_n22086_,
    new_n22087_, new_n22088_, new_n22089_, new_n22090_, new_n22091_,
    new_n22092_, new_n22093_, new_n22094_, new_n22095_, new_n22096_,
    new_n22097_, new_n22098_, new_n22099_, new_n22100_, new_n22101_,
    new_n22102_, new_n22103_, new_n22104_, new_n22105_, new_n22106_,
    new_n22107_, new_n22108_, new_n22109_, new_n22110_, new_n22111_,
    new_n22112_, new_n22113_, new_n22114_, new_n22115_, new_n22116_,
    new_n22117_, new_n22118_, new_n22119_, new_n22120_, new_n22121_,
    new_n22122_, new_n22123_, new_n22124_, new_n22125_, new_n22126_,
    new_n22127_, new_n22128_, new_n22129_, new_n22130_, new_n22131_,
    new_n22132_, new_n22133_, new_n22134_, new_n22135_, new_n22136_,
    new_n22137_, new_n22138_, new_n22139_, new_n22140_, new_n22141_,
    new_n22142_, new_n22143_, new_n22144_, new_n22145_, new_n22146_,
    new_n22147_, new_n22148_, new_n22149_, new_n22150_, new_n22151_,
    new_n22152_, new_n22153_, new_n22154_, new_n22155_, new_n22156_,
    new_n22157_, new_n22158_, new_n22159_, new_n22160_, new_n22161_,
    new_n22162_, new_n22163_, new_n22164_, new_n22165_, new_n22166_,
    new_n22167_, new_n22168_, new_n22169_, new_n22170_, new_n22171_,
    new_n22172_, new_n22173_, new_n22174_, new_n22175_, new_n22176_,
    new_n22177_, new_n22178_, new_n22179_, new_n22180_, new_n22181_,
    new_n22182_, new_n22183_, new_n22184_, new_n22185_, new_n22186_,
    new_n22187_, new_n22188_, new_n22189_, new_n22190_, new_n22191_,
    new_n22192_, new_n22193_, new_n22194_, new_n22195_, new_n22196_,
    new_n22197_, new_n22198_, new_n22199_, new_n22200_, new_n22201_,
    new_n22202_, new_n22203_, new_n22204_, new_n22205_, new_n22206_,
    new_n22207_, new_n22208_, new_n22209_, new_n22210_, new_n22211_,
    new_n22212_, new_n22213_, new_n22214_, new_n22215_, new_n22216_,
    new_n22217_, new_n22218_, new_n22219_, new_n22220_, new_n22221_,
    new_n22222_, new_n22223_, new_n22224_, new_n22225_, new_n22226_,
    new_n22227_, new_n22228_, new_n22229_, new_n22230_, new_n22231_,
    new_n22232_, new_n22233_, new_n22234_, new_n22235_, new_n22236_,
    new_n22237_, new_n22238_, new_n22239_, new_n22240_, new_n22241_,
    new_n22242_, new_n22243_, new_n22244_, new_n22245_, new_n22246_,
    new_n22247_, new_n22248_, new_n22249_, new_n22250_, new_n22251_,
    new_n22252_, new_n22253_, new_n22254_, new_n22255_, new_n22256_,
    new_n22257_, new_n22258_, new_n22259_, new_n22260_, new_n22261_,
    new_n22262_, new_n22263_, new_n22264_, new_n22265_, new_n22266_,
    new_n22267_, new_n22268_, new_n22270_, new_n22271_, new_n22272_,
    new_n22273_, new_n22274_, new_n22275_, new_n22276_, new_n22277_,
    new_n22278_, new_n22279_, new_n22280_, new_n22281_, new_n22282_,
    new_n22283_, new_n22284_, new_n22285_, new_n22286_, new_n22287_,
    new_n22288_, new_n22289_, new_n22290_, new_n22291_, new_n22292_,
    new_n22293_, new_n22294_, new_n22295_, new_n22296_, new_n22297_,
    new_n22298_, new_n22299_, new_n22300_, new_n22301_, new_n22302_,
    new_n22303_, new_n22304_, new_n22305_, new_n22306_, new_n22307_,
    new_n22308_, new_n22309_, new_n22310_, new_n22311_, new_n22312_,
    new_n22313_, new_n22314_, new_n22315_, new_n22316_, new_n22317_,
    new_n22318_, new_n22319_, new_n22320_, new_n22321_, new_n22322_,
    new_n22323_, new_n22324_, new_n22325_, new_n22326_, new_n22327_,
    new_n22328_, new_n22329_, new_n22330_, new_n22331_, new_n22332_,
    new_n22333_, new_n22334_, new_n22335_, new_n22336_, new_n22337_,
    new_n22338_, new_n22339_, new_n22340_, new_n22341_, new_n22342_,
    new_n22343_, new_n22344_, new_n22345_, new_n22346_, new_n22347_,
    new_n22348_, new_n22349_, new_n22350_, new_n22351_, new_n22352_,
    new_n22353_, new_n22354_, new_n22355_, new_n22356_, new_n22357_,
    new_n22358_, new_n22359_, new_n22360_, new_n22361_, new_n22362_,
    new_n22363_, new_n22364_, new_n22365_, new_n22366_, new_n22367_,
    new_n22368_, new_n22369_, new_n22370_, new_n22371_, new_n22372_,
    new_n22373_, new_n22374_, new_n22375_, new_n22376_, new_n22377_,
    new_n22378_, new_n22379_, new_n22380_, new_n22381_, new_n22382_,
    new_n22383_, new_n22384_, new_n22385_, new_n22386_, new_n22387_,
    new_n22388_, new_n22389_, new_n22390_, new_n22391_, new_n22392_,
    new_n22393_, new_n22394_, new_n22395_, new_n22396_, new_n22397_,
    new_n22398_, new_n22399_, new_n22400_, new_n22401_, new_n22402_,
    new_n22403_, new_n22404_, new_n22405_, new_n22406_, new_n22407_,
    new_n22408_, new_n22409_, new_n22410_, new_n22411_, new_n22412_,
    new_n22413_, new_n22414_, new_n22415_, new_n22416_, new_n22417_,
    new_n22418_, new_n22419_, new_n22420_, new_n22421_, new_n22422_,
    new_n22423_, new_n22424_, new_n22425_, new_n22426_, new_n22427_,
    new_n22428_, new_n22430_, new_n22431_, new_n22432_, new_n22433_,
    new_n22434_, new_n22435_, new_n22436_, new_n22437_, new_n22438_,
    new_n22439_, new_n22440_, new_n22441_, new_n22442_, new_n22443_,
    new_n22444_, new_n22445_, new_n22446_, new_n22447_, new_n22448_,
    new_n22449_, new_n22450_, new_n22451_, new_n22452_, new_n22453_,
    new_n22454_, new_n22455_, new_n22456_, new_n22457_, new_n22458_,
    new_n22459_, new_n22460_, new_n22461_, new_n22462_, new_n22463_,
    new_n22464_, new_n22465_, new_n22466_, new_n22467_, new_n22468_,
    new_n22469_, new_n22470_, new_n22471_, new_n22472_, new_n22473_,
    new_n22474_, new_n22475_, new_n22476_, new_n22477_, new_n22478_,
    new_n22479_, new_n22480_, new_n22481_, new_n22482_, new_n22483_,
    new_n22484_, new_n22485_, new_n22486_, new_n22487_, new_n22488_,
    new_n22489_, new_n22490_, new_n22491_, new_n22492_, new_n22493_,
    new_n22494_, new_n22495_, new_n22496_, new_n22497_, new_n22498_,
    new_n22499_, new_n22500_, new_n22501_, new_n22502_, new_n22503_,
    new_n22504_, new_n22505_, new_n22506_, new_n22507_, new_n22508_,
    new_n22509_, new_n22510_, new_n22511_, new_n22512_, new_n22513_,
    new_n22514_, new_n22515_, new_n22516_, new_n22517_, new_n22518_,
    new_n22519_, new_n22520_, new_n22521_, new_n22522_, new_n22523_,
    new_n22524_, new_n22525_, new_n22526_, new_n22527_, new_n22528_,
    new_n22529_, new_n22530_, new_n22531_, new_n22532_, new_n22533_,
    new_n22534_, new_n22535_, new_n22536_, new_n22537_, new_n22538_,
    new_n22539_, new_n22540_, new_n22541_, new_n22542_, new_n22543_,
    new_n22544_, new_n22545_, new_n22546_, new_n22547_, new_n22548_,
    new_n22549_, new_n22550_, new_n22551_, new_n22552_, new_n22553_,
    new_n22554_, new_n22555_, new_n22556_, new_n22557_, new_n22558_,
    new_n22559_, new_n22560_, new_n22561_, new_n22562_, new_n22563_,
    new_n22564_, new_n22565_, new_n22566_, new_n22567_, new_n22568_,
    new_n22569_, new_n22570_, new_n22571_, new_n22572_, new_n22573_,
    new_n22574_, new_n22575_, new_n22576_, new_n22577_, new_n22578_,
    new_n22579_, new_n22580_, new_n22581_, new_n22582_, new_n22583_,
    new_n22584_, new_n22585_, new_n22586_, new_n22588_, new_n22589_,
    new_n22590_, new_n22591_, new_n22592_, new_n22593_, new_n22594_,
    new_n22595_, new_n22596_, new_n22597_, new_n22598_, new_n22599_,
    new_n22600_, new_n22601_, new_n22602_, new_n22603_, new_n22604_,
    new_n22605_, new_n22606_, new_n22607_, new_n22608_, new_n22609_,
    new_n22610_, new_n22611_, new_n22612_, new_n22613_, new_n22614_,
    new_n22615_, new_n22616_, new_n22617_, new_n22618_, new_n22619_,
    new_n22620_, new_n22621_, new_n22622_, new_n22623_, new_n22624_,
    new_n22625_, new_n22626_, new_n22627_, new_n22628_, new_n22629_,
    new_n22630_, new_n22631_, new_n22632_, new_n22633_, new_n22634_,
    new_n22635_, new_n22636_, new_n22637_, new_n22638_, new_n22639_,
    new_n22640_, new_n22641_, new_n22642_, new_n22643_, new_n22644_,
    new_n22645_, new_n22646_, new_n22647_, new_n22648_, new_n22649_,
    new_n22650_, new_n22651_, new_n22652_, new_n22653_, new_n22654_,
    new_n22655_, new_n22656_, new_n22657_, new_n22658_, new_n22659_,
    new_n22660_, new_n22661_, new_n22662_, new_n22663_, new_n22664_,
    new_n22665_, new_n22666_, new_n22667_, new_n22668_, new_n22669_,
    new_n22670_, new_n22671_, new_n22672_, new_n22673_, new_n22674_,
    new_n22675_, new_n22676_, new_n22677_, new_n22678_, new_n22679_,
    new_n22680_, new_n22681_, new_n22682_, new_n22683_, new_n22684_,
    new_n22685_, new_n22686_, new_n22687_, new_n22688_, new_n22689_,
    new_n22690_, new_n22691_, new_n22692_, new_n22693_, new_n22694_,
    new_n22695_, new_n22696_, new_n22697_, new_n22698_, new_n22699_,
    new_n22700_, new_n22701_, new_n22702_, new_n22703_, new_n22704_,
    new_n22705_, new_n22706_, new_n22707_, new_n22708_, new_n22709_,
    new_n22710_, new_n22711_, new_n22712_, new_n22713_, new_n22714_,
    new_n22715_, new_n22717_, new_n22718_, new_n22719_, new_n22720_,
    new_n22721_, new_n22722_, new_n22724_, new_n22725_, new_n22726_,
    new_n22727_, new_n22728_, new_n22730_, new_n22731_, new_n22732_,
    new_n22733_, new_n22734_, new_n22735_, new_n22736_, new_n22737_,
    new_n22738_, new_n22739_, new_n22740_, new_n22741_, new_n22742_,
    new_n22743_, new_n22744_, new_n22745_, new_n22746_, new_n22747_,
    new_n22748_, new_n22749_, new_n22750_, new_n22751_, new_n22752_,
    new_n22753_, new_n22754_, new_n22755_, new_n22756_, new_n22757_,
    new_n22758_, new_n22759_, new_n22760_, new_n22761_, new_n22762_,
    new_n22763_, new_n22764_, new_n22765_, new_n22766_, new_n22767_,
    new_n22768_, new_n22769_, new_n22770_, new_n22771_, new_n22772_,
    new_n22773_, new_n22774_, new_n22775_, new_n22776_, new_n22777_,
    new_n22778_, new_n22779_, new_n22780_, new_n22781_, new_n22782_,
    new_n22783_, new_n22784_, new_n22785_, new_n22786_, new_n22787_,
    new_n22788_, new_n22789_, new_n22790_, new_n22791_, new_n22792_,
    new_n22794_, new_n22795_, new_n22797_, new_n22798_, new_n22799_,
    new_n22800_, new_n22801_, new_n22803_, new_n22804_, new_n22805_,
    new_n22806_, new_n22807_, new_n22808_, new_n22809_, new_n22810_,
    new_n22811_, new_n22812_, new_n22813_, new_n22814_, new_n22815_,
    new_n22816_, new_n22817_, new_n22818_, new_n22819_, new_n22820_,
    new_n22821_, new_n22822_, new_n22823_, new_n22824_, new_n22825_,
    new_n22826_, new_n22827_, new_n22828_, new_n22829_, new_n22830_,
    new_n22831_, new_n22832_, new_n22833_, new_n22834_, new_n22835_,
    new_n22836_, new_n22837_, new_n22838_, new_n22839_, new_n22840_,
    new_n22841_, new_n22842_, new_n22843_, new_n22844_, new_n22845_,
    new_n22846_, new_n22847_, new_n22848_, new_n22849_, new_n22850_,
    new_n22851_, new_n22852_, new_n22853_, new_n22854_, new_n22855_,
    new_n22856_, new_n22857_, new_n22858_, new_n22859_, new_n22860_,
    new_n22861_, new_n22862_, new_n22863_, new_n22864_, new_n22865_,
    new_n22866_, new_n22867_, new_n22868_, new_n22869_, new_n22870_,
    new_n22871_, new_n22872_, new_n22873_, new_n22874_, new_n22875_,
    new_n22876_, new_n22877_, new_n22878_, new_n22879_, new_n22880_,
    new_n22881_, new_n22882_, new_n22883_, new_n22884_, new_n22885_,
    new_n22886_, new_n22887_, new_n22888_, new_n22889_, new_n22890_,
    new_n22891_, new_n22892_, new_n22893_, new_n22894_, new_n22895_,
    new_n22896_, new_n22897_, new_n22898_, new_n22899_, new_n22900_,
    new_n22901_, new_n22902_, new_n22903_, new_n22904_, new_n22905_,
    new_n22906_, new_n22907_, new_n22908_, new_n22909_, new_n22910_,
    new_n22911_, new_n22912_, new_n22913_, new_n22914_, new_n22915_,
    new_n22916_, new_n22917_, new_n22918_, new_n22919_, new_n22920_,
    new_n22921_, new_n22922_, new_n22923_, new_n22924_, new_n22925_,
    new_n22926_, new_n22927_, new_n22928_, new_n22929_, new_n22930_,
    new_n22931_, new_n22932_, new_n22933_, new_n22934_, new_n22935_,
    new_n22936_, new_n22937_, new_n22938_, new_n22939_, new_n22940_,
    new_n22941_, new_n22942_, new_n22943_, new_n22944_, new_n22945_,
    new_n22946_, new_n22947_, new_n22948_, new_n22949_, new_n22950_,
    new_n22951_, new_n22952_, new_n22953_, new_n22954_, new_n22955_,
    new_n22956_, new_n22957_, new_n22958_, new_n22959_, new_n22960_,
    new_n22961_, new_n22962_, new_n22963_, new_n22964_, new_n22965_,
    new_n22966_, new_n22967_, new_n22968_, new_n22969_, new_n22970_,
    new_n22971_, new_n22972_, new_n22973_, new_n22974_, new_n22975_,
    new_n22976_, new_n22977_, new_n22978_, new_n22979_, new_n22980_,
    new_n22981_, new_n22982_, new_n22983_, new_n22984_, new_n22985_,
    new_n22986_, new_n22987_, new_n22988_, new_n22989_, new_n22990_,
    new_n22991_, new_n22992_, new_n22993_, new_n22994_, new_n22995_,
    new_n22996_, new_n22997_, new_n22998_, new_n22999_, new_n23000_,
    new_n23001_, new_n23002_, new_n23003_, new_n23004_, new_n23005_,
    new_n23006_, new_n23007_, new_n23008_, new_n23009_, new_n23010_,
    new_n23011_, new_n23012_, new_n23013_, new_n23014_, new_n23015_,
    new_n23016_, new_n23017_, new_n23018_, new_n23019_, new_n23020_,
    new_n23021_, new_n23022_, new_n23023_, new_n23024_, new_n23025_,
    new_n23026_, new_n23027_, new_n23028_, new_n23029_, new_n23030_,
    new_n23031_, new_n23032_, new_n23033_, new_n23034_, new_n23035_,
    new_n23036_, new_n23037_, new_n23038_, new_n23039_, new_n23040_,
    new_n23041_, new_n23042_, new_n23043_, new_n23044_, new_n23045_,
    new_n23046_, new_n23047_, new_n23048_, new_n23049_, new_n23050_,
    new_n23051_, new_n23052_, new_n23053_, new_n23054_, new_n23055_,
    new_n23056_, new_n23057_, new_n23058_, new_n23059_, new_n23060_,
    new_n23061_, new_n23062_, new_n23063_, new_n23064_, new_n23065_,
    new_n23066_, new_n23067_, new_n23068_, new_n23069_, new_n23070_,
    new_n23071_, new_n23072_, new_n23073_, new_n23074_, new_n23075_,
    new_n23076_, new_n23077_, new_n23078_, new_n23079_, new_n23080_,
    new_n23081_, new_n23082_, new_n23083_, new_n23084_, new_n23085_,
    new_n23086_, new_n23087_, new_n23088_, new_n23089_, new_n23090_,
    new_n23091_, new_n23092_, new_n23093_, new_n23094_, new_n23095_,
    new_n23096_, new_n23097_, new_n23098_, new_n23099_, new_n23100_,
    new_n23101_, new_n23102_, new_n23103_, new_n23104_, new_n23105_,
    new_n23106_, new_n23107_, new_n23109_, new_n23110_, new_n23111_,
    new_n23112_, new_n23113_, new_n23114_, new_n23115_, new_n23116_,
    new_n23117_, new_n23118_, new_n23119_, new_n23120_, new_n23121_,
    new_n23122_, new_n23123_, new_n23124_, new_n23125_, new_n23126_,
    new_n23127_, new_n23128_, new_n23129_, new_n23130_, new_n23131_,
    new_n23132_, new_n23133_, new_n23134_, new_n23135_, new_n23136_,
    new_n23137_, new_n23138_, new_n23139_, new_n23140_, new_n23141_,
    new_n23142_, new_n23143_, new_n23144_, new_n23145_, new_n23146_,
    new_n23147_, new_n23148_, new_n23149_, new_n23151_, new_n23152_,
    new_n23153_, new_n23154_, new_n23155_, new_n23156_, new_n23157_,
    new_n23158_, new_n23159_, new_n23160_, new_n23161_, new_n23162_,
    new_n23163_, new_n23164_, new_n23165_, new_n23166_, new_n23167_,
    new_n23168_, new_n23169_, new_n23170_, new_n23171_, new_n23172_,
    new_n23173_, new_n23174_, new_n23175_, new_n23176_, new_n23177_,
    new_n23178_, new_n23179_, new_n23180_, new_n23181_, new_n23182_,
    new_n23183_, new_n23184_, new_n23185_, new_n23186_, new_n23187_,
    new_n23188_, new_n23189_, new_n23190_, new_n23191_, new_n23192_,
    new_n23193_, new_n23194_, new_n23195_, new_n23196_, new_n23197_,
    new_n23198_, new_n23199_, new_n23200_, new_n23201_, new_n23202_,
    new_n23203_, new_n23204_, new_n23205_, new_n23206_, new_n23207_,
    new_n23208_, new_n23209_, new_n23210_, new_n23211_, new_n23212_,
    new_n23213_, new_n23214_, new_n23215_, new_n23216_, new_n23217_,
    new_n23218_, new_n23219_, new_n23220_, new_n23221_, new_n23222_,
    new_n23223_, new_n23224_, new_n23225_, new_n23226_, new_n23227_,
    new_n23228_, new_n23229_, new_n23230_, new_n23231_, new_n23232_,
    new_n23233_, new_n23234_, new_n23235_, new_n23236_, new_n23237_,
    new_n23238_, new_n23239_, new_n23240_, new_n23241_, new_n23242_,
    new_n23243_, new_n23244_, new_n23245_, new_n23246_, new_n23247_,
    new_n23248_, new_n23249_, new_n23250_, new_n23251_, new_n23253_,
    new_n23254_, new_n23255_, new_n23256_, new_n23257_, new_n23258_,
    new_n23259_, new_n23260_, new_n23261_, new_n23262_, new_n23263_,
    new_n23264_, new_n23265_, new_n23266_, new_n23267_, new_n23268_,
    new_n23269_, new_n23270_, new_n23271_, new_n23272_, new_n23273_,
    new_n23274_, new_n23275_, new_n23276_, new_n23277_, new_n23278_,
    new_n23279_, new_n23280_, new_n23281_, new_n23282_, new_n23283_,
    new_n23284_, new_n23285_, new_n23286_, new_n23287_, new_n23288_,
    new_n23289_, new_n23290_, new_n23291_, new_n23292_, new_n23293_,
    new_n23294_, new_n23295_, new_n23296_, new_n23297_, new_n23298_,
    new_n23299_, new_n23300_, new_n23301_, new_n23302_, new_n23303_,
    new_n23304_, new_n23305_, new_n23306_, new_n23307_, new_n23308_,
    new_n23309_, new_n23310_, new_n23311_, new_n23312_, new_n23313_,
    new_n23314_, new_n23315_, new_n23316_, new_n23317_, new_n23318_,
    new_n23319_, new_n23320_, new_n23321_, new_n23322_, new_n23323_,
    new_n23324_, new_n23325_, new_n23326_, new_n23328_, new_n23329_,
    new_n23330_, new_n23331_, new_n23332_, new_n23333_, new_n23334_,
    new_n23335_, new_n23336_, new_n23337_, new_n23338_, new_n23339_,
    new_n23340_, new_n23341_, new_n23342_, new_n23344_, new_n23345_,
    new_n23346_, new_n23347_, new_n23348_, new_n23349_, new_n23350_,
    new_n23351_, new_n23352_, new_n23353_, new_n23355_, new_n23356_,
    new_n23357_, new_n23358_, new_n23359_, new_n23360_, new_n23361_,
    new_n23362_, new_n23363_, new_n23364_, new_n23365_, new_n23367_,
    new_n23368_, new_n23369_, new_n23370_, new_n23371_, new_n23372_,
    new_n23373_, new_n23374_, new_n23375_, new_n23376_, new_n23378_,
    new_n23379_, new_n23380_, new_n23381_, new_n23382_, new_n23383_,
    new_n23384_, new_n23385_, new_n23386_, new_n23387_, new_n23388_,
    new_n23389_, new_n23390_, new_n23391_, new_n23392_, new_n23393_,
    new_n23394_, new_n23395_, new_n23396_, new_n23397_, new_n23398_,
    new_n23399_, new_n23400_, new_n23401_, new_n23402_, new_n23403_,
    new_n23404_, new_n23405_, new_n23406_, new_n23407_, new_n23408_,
    new_n23409_, new_n23410_, new_n23411_, new_n23412_, new_n23413_,
    new_n23414_, new_n23415_, new_n23416_, new_n23417_, new_n23418_,
    new_n23419_, new_n23420_, new_n23421_, new_n23422_, new_n23423_,
    new_n23424_, new_n23425_, new_n23426_, new_n23427_, new_n23428_,
    new_n23429_, new_n23430_, new_n23431_, new_n23432_, new_n23433_,
    new_n23434_, new_n23435_, new_n23436_, new_n23437_, new_n23438_,
    new_n23439_, new_n23440_, new_n23441_, new_n23442_, new_n23443_,
    new_n23444_, new_n23445_, new_n23446_, new_n23447_, new_n23448_,
    new_n23449_, new_n23450_, new_n23452_, new_n23453_, new_n23454_,
    new_n23455_, new_n23456_, new_n23457_, new_n23458_, new_n23459_,
    new_n23460_, new_n23461_, new_n23462_, new_n23463_, new_n23464_,
    new_n23465_, new_n23466_, new_n23467_, new_n23468_, new_n23469_,
    new_n23470_, new_n23471_, new_n23472_, new_n23473_, new_n23474_,
    new_n23475_, new_n23476_, new_n23477_, new_n23478_, new_n23479_,
    new_n23480_, new_n23481_, new_n23482_, new_n23483_, new_n23484_,
    new_n23485_, new_n23486_, new_n23487_, new_n23488_, new_n23489_,
    new_n23490_, new_n23491_, new_n23492_, new_n23493_, new_n23494_,
    new_n23495_, new_n23496_, new_n23497_, new_n23498_, new_n23499_,
    new_n23500_, new_n23501_, new_n23502_, new_n23503_, new_n23504_,
    new_n23505_, new_n23506_, new_n23507_, new_n23508_, new_n23509_,
    new_n23510_, new_n23511_, new_n23512_, new_n23513_, new_n23514_,
    new_n23515_, new_n23516_, new_n23517_, new_n23518_, new_n23519_,
    new_n23520_, new_n23521_, new_n23523_, new_n23524_, new_n23525_,
    new_n23526_, new_n23527_, new_n23528_, new_n23529_, new_n23530_,
    new_n23531_, new_n23532_, new_n23533_, new_n23534_, new_n23536_,
    new_n23537_, new_n23539_, new_n23540_, new_n23541_, new_n23542_,
    new_n23543_, new_n23544_, new_n23545_, new_n23546_, new_n23547_,
    new_n23548_, new_n23549_, new_n23551_, new_n23552_, new_n23553_,
    new_n23555_, new_n23556_, new_n23557_, new_n23558_, new_n23559_,
    new_n23560_, new_n23561_, new_n23562_, new_n23563_, new_n23564_,
    new_n23565_, new_n23566_, new_n23567_, new_n23568_, new_n23569_,
    new_n23570_, new_n23571_, new_n23572_, new_n23573_, new_n23574_,
    new_n23575_, new_n23576_, new_n23577_, new_n23578_, new_n23579_,
    new_n23580_, new_n23581_, new_n23582_, new_n23583_, new_n23584_,
    new_n23585_, new_n23586_, new_n23587_, new_n23588_, new_n23589_,
    new_n23590_, new_n23591_, new_n23592_, new_n23593_, new_n23594_,
    new_n23595_, new_n23596_, new_n23597_, new_n23598_, new_n23599_,
    new_n23600_, new_n23601_, new_n23602_, new_n23603_, new_n23604_,
    new_n23605_, new_n23606_, new_n23607_, new_n23608_, new_n23609_,
    new_n23610_, new_n23611_, new_n23612_, new_n23613_, new_n23614_,
    new_n23615_, new_n23616_, new_n23617_, new_n23618_, new_n23619_,
    new_n23620_, new_n23622_, new_n23623_, new_n23624_, new_n23625_,
    new_n23626_, new_n23627_, new_n23628_, new_n23629_, new_n23630_,
    new_n23631_, new_n23632_, new_n23633_, new_n23634_, new_n23635_,
    new_n23636_, new_n23637_, new_n23638_, new_n23639_, new_n23640_,
    new_n23641_, new_n23642_, new_n23643_, new_n23644_, new_n23645_,
    new_n23646_, new_n23647_, new_n23648_, new_n23649_, new_n23650_,
    new_n23651_, new_n23652_, new_n23653_, new_n23654_, new_n23655_,
    new_n23656_, new_n23657_, new_n23658_, new_n23659_, new_n23660_,
    new_n23661_, new_n23662_, new_n23663_, new_n23664_, new_n23665_,
    new_n23666_, new_n23667_, new_n23668_, new_n23669_, new_n23670_,
    new_n23671_, new_n23672_, new_n23673_, new_n23674_, new_n23675_,
    new_n23676_, new_n23677_, new_n23678_, new_n23679_, new_n23680_,
    new_n23681_, new_n23682_, new_n23683_, new_n23684_, new_n23685_,
    new_n23686_, new_n23687_, new_n23688_, new_n23689_, new_n23690_,
    new_n23691_, new_n23692_, new_n23693_, new_n23694_, new_n23695_,
    new_n23696_, new_n23697_, new_n23698_, new_n23699_, new_n23700_,
    new_n23701_, new_n23702_, new_n23703_, new_n23704_, new_n23705_,
    new_n23706_, new_n23707_, new_n23708_, new_n23709_, new_n23710_,
    new_n23711_, new_n23712_, new_n23713_, new_n23714_, new_n23715_,
    new_n23716_, new_n23717_, new_n23718_, new_n23719_, new_n23720_,
    new_n23721_, new_n23722_, new_n23723_, new_n23724_, new_n23725_,
    new_n23726_, new_n23727_, new_n23728_, new_n23729_, new_n23730_,
    new_n23731_, new_n23732_, new_n23733_, new_n23734_, new_n23735_,
    new_n23736_, new_n23737_, new_n23738_, new_n23739_, new_n23740_,
    new_n23741_, new_n23742_, new_n23743_, new_n23744_, new_n23745_,
    new_n23746_, new_n23747_, new_n23748_, new_n23749_, new_n23750_,
    new_n23751_, new_n23752_, new_n23753_, new_n23754_, new_n23755_,
    new_n23756_, new_n23757_, new_n23758_, new_n23759_, new_n23760_,
    new_n23761_, new_n23762_, new_n23763_, new_n23764_, new_n23765_,
    new_n23766_, new_n23767_, new_n23768_, new_n23769_, new_n23770_,
    new_n23771_, new_n23772_, new_n23773_, new_n23774_, new_n23775_,
    new_n23776_, new_n23777_, new_n23778_, new_n23779_, new_n23780_,
    new_n23781_, new_n23782_, new_n23783_, new_n23784_, new_n23785_,
    new_n23786_, new_n23787_, new_n23788_, new_n23789_, new_n23790_,
    new_n23791_, new_n23792_, new_n23793_, new_n23794_, new_n23795_,
    new_n23796_, new_n23797_, new_n23798_, new_n23799_, new_n23800_,
    new_n23801_, new_n23802_, new_n23803_, new_n23804_, new_n23805_,
    new_n23806_, new_n23807_, new_n23808_, new_n23809_, new_n23810_,
    new_n23811_, new_n23812_, new_n23813_, new_n23814_, new_n23815_,
    new_n23816_, new_n23817_, new_n23818_, new_n23819_, new_n23820_,
    new_n23821_, new_n23822_, new_n23823_, new_n23824_, new_n23825_,
    new_n23826_, new_n23827_, new_n23828_, new_n23829_, new_n23830_,
    new_n23831_, new_n23832_, new_n23833_, new_n23834_, new_n23835_,
    new_n23836_, new_n23837_, new_n23838_, new_n23839_, new_n23840_,
    new_n23841_, new_n23842_, new_n23843_, new_n23844_, new_n23845_,
    new_n23846_, new_n23847_, new_n23848_, new_n23849_, new_n23850_,
    new_n23851_, new_n23852_, new_n23853_, new_n23854_, new_n23855_,
    new_n23856_, new_n23857_, new_n23858_, new_n23859_, new_n23860_,
    new_n23861_, new_n23862_, new_n23863_, new_n23864_, new_n23865_,
    new_n23866_, new_n23867_, new_n23868_, new_n23869_, new_n23870_,
    new_n23871_, new_n23872_, new_n23873_, new_n23874_, new_n23875_,
    new_n23876_, new_n23877_, new_n23878_, new_n23879_, new_n23880_,
    new_n23881_, new_n23882_, new_n23883_, new_n23884_, new_n23885_,
    new_n23886_, new_n23887_, new_n23888_, new_n23889_, new_n23890_,
    new_n23891_, new_n23892_, new_n23893_, new_n23894_, new_n23895_,
    new_n23896_, new_n23897_, new_n23898_, new_n23899_, new_n23900_,
    new_n23901_, new_n23902_, new_n23903_, new_n23904_, new_n23905_,
    new_n23906_, new_n23907_, new_n23908_, new_n23909_, new_n23910_,
    new_n23911_, new_n23912_, new_n23913_, new_n23914_, new_n23915_,
    new_n23916_, new_n23917_, new_n23918_, new_n23919_, new_n23920_,
    new_n23921_, new_n23922_, new_n23923_, new_n23924_, new_n23925_,
    new_n23926_, new_n23927_, new_n23928_, new_n23929_, new_n23930_,
    new_n23931_, new_n23932_, new_n23933_, new_n23934_, new_n23935_,
    new_n23936_, new_n23937_, new_n23938_, new_n23939_, new_n23940_,
    new_n23941_, new_n23942_, new_n23943_, new_n23944_, new_n23945_,
    new_n23946_, new_n23947_, new_n23948_, new_n23949_, new_n23950_,
    new_n23951_, new_n23952_, new_n23953_, new_n23954_, new_n23955_,
    new_n23956_, new_n23957_, new_n23958_, new_n23959_, new_n23960_,
    new_n23961_, new_n23962_, new_n23963_, new_n23964_, new_n23965_,
    new_n23966_, new_n23967_, new_n23968_, new_n23969_, new_n23970_,
    new_n23971_, new_n23972_, new_n23973_, new_n23974_, new_n23975_,
    new_n23976_, new_n23977_, new_n23978_, new_n23979_, new_n23980_,
    new_n23981_, new_n23982_, new_n23983_, new_n23984_, new_n23985_,
    new_n23986_, new_n23987_, new_n23988_, new_n23989_, new_n23990_,
    new_n23991_, new_n23992_, new_n23993_, new_n23994_, new_n23995_,
    new_n23996_, new_n23997_, new_n23998_, new_n23999_, new_n24000_,
    new_n24001_, new_n24002_, new_n24003_, new_n24004_, new_n24005_,
    new_n24006_, new_n24007_, new_n24008_, new_n24009_, new_n24010_,
    new_n24011_, new_n24012_, new_n24013_, new_n24014_, new_n24015_,
    new_n24016_, new_n24017_, new_n24018_, new_n24019_, new_n24020_,
    new_n24021_, new_n24022_, new_n24024_, new_n24025_, new_n24026_,
    new_n24027_, new_n24028_, new_n24029_, new_n24030_, new_n24031_,
    new_n24032_, new_n24033_, new_n24034_, new_n24035_, new_n24036_,
    new_n24037_, new_n24038_, new_n24039_, new_n24040_, new_n24041_,
    new_n24042_, new_n24043_, new_n24044_, new_n24045_, new_n24046_,
    new_n24047_, new_n24048_, new_n24049_, new_n24050_, new_n24051_,
    new_n24052_, new_n24053_, new_n24054_, new_n24055_, new_n24056_,
    new_n24057_, new_n24058_, new_n24059_, new_n24060_, new_n24061_,
    new_n24062_, new_n24063_, new_n24064_, new_n24065_, new_n24066_,
    new_n24067_, new_n24068_, new_n24069_, new_n24070_, new_n24071_,
    new_n24072_, new_n24073_, new_n24074_, new_n24075_, new_n24076_,
    new_n24077_, new_n24078_, new_n24079_, new_n24080_, new_n24081_,
    new_n24082_, new_n24083_, new_n24084_, new_n24085_, new_n24086_,
    new_n24087_, new_n24088_, new_n24089_, new_n24090_, new_n24091_,
    new_n24092_, new_n24093_, new_n24094_, new_n24095_, new_n24096_,
    new_n24097_, new_n24098_, new_n24099_, new_n24100_, new_n24101_,
    new_n24102_, new_n24103_, new_n24104_, new_n24105_, new_n24106_,
    new_n24107_, new_n24108_, new_n24109_, new_n24110_, new_n24111_,
    new_n24112_, new_n24113_, new_n24114_, new_n24115_, new_n24116_,
    new_n24117_, new_n24118_, new_n24119_, new_n24120_, new_n24121_,
    new_n24122_, new_n24123_, new_n24124_, new_n24125_, new_n24126_,
    new_n24127_, new_n24128_, new_n24129_, new_n24130_, new_n24131_,
    new_n24132_, new_n24133_, new_n24134_, new_n24135_, new_n24136_,
    new_n24137_, new_n24138_, new_n24139_, new_n24140_, new_n24141_,
    new_n24142_, new_n24143_, new_n24144_, new_n24145_, new_n24146_,
    new_n24147_, new_n24148_, new_n24149_, new_n24150_, new_n24151_,
    new_n24152_, new_n24153_, new_n24154_, new_n24155_, new_n24156_,
    new_n24157_, new_n24158_, new_n24159_, new_n24160_, new_n24161_,
    new_n24162_, new_n24163_, new_n24164_, new_n24165_, new_n24166_,
    new_n24167_, new_n24168_, new_n24169_, new_n24170_, new_n24171_,
    new_n24172_, new_n24173_, new_n24174_, new_n24175_, new_n24176_,
    new_n24177_, new_n24178_, new_n24179_, new_n24180_, new_n24181_,
    new_n24182_, new_n24183_, new_n24184_, new_n24185_, new_n24186_,
    new_n24187_, new_n24188_, new_n24189_, new_n24190_, new_n24191_,
    new_n24192_, new_n24193_, new_n24194_, new_n24195_, new_n24196_,
    new_n24197_, new_n24198_, new_n24199_, new_n24200_, new_n24201_,
    new_n24202_, new_n24203_, new_n24204_, new_n24205_, new_n24206_,
    new_n24207_, new_n24208_, new_n24209_, new_n24210_, new_n24211_,
    new_n24212_, new_n24213_, new_n24214_, new_n24215_, new_n24216_,
    new_n24217_, new_n24218_, new_n24219_, new_n24220_, new_n24221_,
    new_n24222_, new_n24223_, new_n24224_, new_n24225_, new_n24226_,
    new_n24227_, new_n24228_, new_n24229_, new_n24230_, new_n24231_,
    new_n24232_, new_n24233_, new_n24234_, new_n24235_, new_n24236_,
    new_n24237_, new_n24238_, new_n24239_, new_n24240_, new_n24241_,
    new_n24242_, new_n24243_, new_n24244_, new_n24245_, new_n24246_,
    new_n24247_, new_n24248_, new_n24249_, new_n24250_, new_n24251_,
    new_n24252_, new_n24253_, new_n24254_, new_n24255_, new_n24256_,
    new_n24257_, new_n24258_, new_n24259_, new_n24260_, new_n24261_,
    new_n24262_, new_n24263_, new_n24264_, new_n24265_, new_n24266_,
    new_n24267_, new_n24268_, new_n24269_, new_n24270_, new_n24271_,
    new_n24272_, new_n24273_, new_n24274_, new_n24275_, new_n24276_,
    new_n24277_, new_n24278_, new_n24279_, new_n24280_, new_n24281_,
    new_n24282_, new_n24283_, new_n24284_, new_n24285_, new_n24286_,
    new_n24287_, new_n24288_, new_n24289_, new_n24290_, new_n24291_,
    new_n24292_, new_n24293_, new_n24294_, new_n24295_, new_n24296_,
    new_n24297_, new_n24298_, new_n24299_, new_n24300_, new_n24301_,
    new_n24302_, new_n24303_, new_n24304_, new_n24305_, new_n24306_,
    new_n24307_, new_n24308_, new_n24309_, new_n24310_, new_n24311_,
    new_n24312_, new_n24313_, new_n24314_, new_n24315_, new_n24316_,
    new_n24317_, new_n24318_, new_n24319_, new_n24320_, new_n24321_,
    new_n24322_, new_n24323_, new_n24324_, new_n24325_, new_n24326_,
    new_n24327_, new_n24328_, new_n24329_, new_n24330_, new_n24331_,
    new_n24332_, new_n24333_, new_n24334_, new_n24335_, new_n24336_,
    new_n24337_, new_n24338_, new_n24339_, new_n24340_, new_n24341_,
    new_n24342_, new_n24343_, new_n24344_, new_n24345_, new_n24346_,
    new_n24347_, new_n24348_, new_n24349_, new_n24350_, new_n24351_,
    new_n24352_, new_n24353_, new_n24354_, new_n24355_, new_n24356_,
    new_n24357_, new_n24358_, new_n24359_, new_n24360_, new_n24361_,
    new_n24362_, new_n24363_, new_n24364_, new_n24365_, new_n24366_,
    new_n24367_, new_n24368_, new_n24369_, new_n24370_, new_n24371_,
    new_n24372_, new_n24373_, new_n24374_, new_n24375_, new_n24376_,
    new_n24377_, new_n24378_, new_n24379_, new_n24380_, new_n24381_,
    new_n24383_, new_n24384_, new_n24385_, new_n24386_, new_n24387_,
    new_n24388_, new_n24389_, new_n24390_, new_n24391_, new_n24392_,
    new_n24393_, new_n24394_, new_n24395_, new_n24396_, new_n24397_,
    new_n24398_, new_n24399_, new_n24400_, new_n24401_, new_n24402_,
    new_n24403_, new_n24404_, new_n24405_, new_n24406_, new_n24407_,
    new_n24408_, new_n24409_, new_n24410_, new_n24411_, new_n24412_,
    new_n24413_, new_n24414_, new_n24415_, new_n24416_, new_n24417_,
    new_n24418_, new_n24419_, new_n24420_, new_n24421_, new_n24422_,
    new_n24423_, new_n24424_, new_n24425_, new_n24426_, new_n24427_,
    new_n24428_, new_n24429_, new_n24430_, new_n24431_, new_n24432_,
    new_n24433_, new_n24434_, new_n24435_, new_n24436_, new_n24437_,
    new_n24438_, new_n24439_, new_n24440_, new_n24441_, new_n24442_,
    new_n24443_, new_n24444_, new_n24445_, new_n24446_, new_n24447_,
    new_n24448_, new_n24449_, new_n24450_, new_n24451_, new_n24452_,
    new_n24453_, new_n24454_, new_n24455_, new_n24456_, new_n24457_,
    new_n24458_, new_n24459_, new_n24460_, new_n24461_, new_n24462_,
    new_n24463_, new_n24464_, new_n24465_, new_n24466_, new_n24467_,
    new_n24468_, new_n24469_, new_n24470_, new_n24471_, new_n24472_,
    new_n24473_, new_n24474_, new_n24475_, new_n24476_, new_n24477_,
    new_n24478_, new_n24479_, new_n24480_, new_n24481_, new_n24482_,
    new_n24483_, new_n24484_, new_n24485_, new_n24486_, new_n24487_,
    new_n24488_, new_n24489_, new_n24490_, new_n24491_, new_n24492_,
    new_n24493_, new_n24494_, new_n24495_, new_n24496_, new_n24497_,
    new_n24498_, new_n24499_, new_n24500_, new_n24501_, new_n24502_,
    new_n24503_, new_n24504_, new_n24505_, new_n24506_, new_n24507_,
    new_n24508_, new_n24509_, new_n24510_, new_n24511_, new_n24512_,
    new_n24513_, new_n24514_, new_n24515_, new_n24516_, new_n24517_,
    new_n24518_, new_n24519_, new_n24520_, new_n24521_, new_n24522_,
    new_n24523_, new_n24524_, new_n24525_, new_n24526_, new_n24527_,
    new_n24528_, new_n24529_, new_n24530_, new_n24531_, new_n24532_,
    new_n24533_, new_n24534_, new_n24535_, new_n24536_, new_n24537_,
    new_n24538_, new_n24539_, new_n24540_, new_n24541_, new_n24542_,
    new_n24543_, new_n24544_, new_n24545_, new_n24546_, new_n24547_,
    new_n24548_, new_n24549_, new_n24550_, new_n24551_, new_n24552_,
    new_n24553_, new_n24554_, new_n24555_, new_n24556_, new_n24557_,
    new_n24558_, new_n24559_, new_n24560_, new_n24561_, new_n24562_,
    new_n24563_, new_n24564_, new_n24565_, new_n24566_, new_n24567_,
    new_n24568_, new_n24569_, new_n24570_, new_n24571_, new_n24572_,
    new_n24573_, new_n24574_, new_n24575_, new_n24576_, new_n24577_,
    new_n24578_, new_n24579_, new_n24580_, new_n24581_, new_n24582_,
    new_n24583_, new_n24584_, new_n24585_, new_n24586_, new_n24587_,
    new_n24588_, new_n24589_, new_n24590_, new_n24591_, new_n24592_,
    new_n24593_, new_n24594_, new_n24595_, new_n24596_, new_n24597_,
    new_n24598_, new_n24599_, new_n24600_, new_n24601_, new_n24602_,
    new_n24603_, new_n24604_, new_n24605_, new_n24606_, new_n24607_,
    new_n24608_, new_n24609_, new_n24610_, new_n24611_, new_n24612_,
    new_n24613_, new_n24614_, new_n24615_, new_n24616_, new_n24617_,
    new_n24618_, new_n24619_, new_n24620_, new_n24621_, new_n24622_,
    new_n24623_, new_n24624_, new_n24625_, new_n24626_, new_n24627_,
    new_n24628_, new_n24629_, new_n24630_, new_n24631_, new_n24632_,
    new_n24633_, new_n24634_, new_n24635_, new_n24636_, new_n24637_,
    new_n24638_, new_n24639_, new_n24640_, new_n24641_, new_n24642_,
    new_n24643_, new_n24644_, new_n24645_, new_n24646_, new_n24647_,
    new_n24648_, new_n24649_, new_n24650_, new_n24651_, new_n24652_,
    new_n24653_, new_n24654_, new_n24655_, new_n24656_, new_n24657_,
    new_n24658_, new_n24659_, new_n24660_, new_n24661_, new_n24662_,
    new_n24663_, new_n24664_, new_n24665_, new_n24666_, new_n24667_,
    new_n24668_, new_n24669_, new_n24670_, new_n24671_, new_n24672_,
    new_n24673_, new_n24674_, new_n24675_, new_n24676_, new_n24677_,
    new_n24678_, new_n24679_, new_n24680_, new_n24681_, new_n24682_,
    new_n24683_, new_n24684_, new_n24685_, new_n24686_, new_n24687_,
    new_n24688_, new_n24689_, new_n24690_, new_n24691_, new_n24692_,
    new_n24693_, new_n24694_, new_n24695_, new_n24696_, new_n24697_,
    new_n24698_, new_n24699_, new_n24700_, new_n24701_, new_n24702_,
    new_n24703_, new_n24704_, new_n24705_, new_n24706_, new_n24707_,
    new_n24708_, new_n24709_, new_n24710_, new_n24711_, new_n24712_,
    new_n24713_, new_n24714_, new_n24715_, new_n24716_, new_n24717_,
    new_n24718_, new_n24719_, new_n24720_, new_n24721_, new_n24722_,
    new_n24723_, new_n24725_, new_n24726_, new_n24727_, new_n24728_,
    new_n24729_, new_n24730_, new_n24731_, new_n24732_, new_n24733_,
    new_n24734_, new_n24735_, new_n24736_, new_n24737_, new_n24738_,
    new_n24739_, new_n24740_, new_n24741_, new_n24742_, new_n24743_,
    new_n24744_, new_n24745_, new_n24746_, new_n24747_, new_n24748_,
    new_n24749_, new_n24750_, new_n24751_, new_n24752_, new_n24753_,
    new_n24754_, new_n24755_, new_n24756_, new_n24757_, new_n24758_,
    new_n24759_, new_n24760_, new_n24761_, new_n24762_, new_n24763_,
    new_n24764_, new_n24765_, new_n24766_, new_n24767_, new_n24768_,
    new_n24769_, new_n24770_, new_n24771_, new_n24772_, new_n24773_,
    new_n24774_, new_n24775_, new_n24776_, new_n24777_, new_n24778_,
    new_n24779_, new_n24780_, new_n24781_, new_n24782_, new_n24783_,
    new_n24784_, new_n24785_, new_n24786_, new_n24787_, new_n24788_,
    new_n24789_, new_n24790_, new_n24791_, new_n24792_, new_n24793_,
    new_n24794_, new_n24795_, new_n24796_, new_n24797_, new_n24798_,
    new_n24799_, new_n24800_, new_n24801_, new_n24803_, new_n24804_,
    new_n24805_, new_n24806_, new_n24807_, new_n24808_, new_n24809_,
    new_n24810_, new_n24811_, new_n24812_, new_n24813_, new_n24814_,
    new_n24815_, new_n24816_, new_n24817_, new_n24818_, new_n24819_,
    new_n24820_, new_n24821_, new_n24822_, new_n24823_, new_n24824_,
    new_n24825_, new_n24826_, new_n24827_, new_n24828_, new_n24829_,
    new_n24830_, new_n24831_, new_n24833_, new_n24834_, new_n24835_,
    new_n24836_, new_n24837_, new_n24838_, new_n24839_, new_n24840_,
    new_n24841_, new_n24842_, new_n24843_, new_n24844_, new_n24845_,
    new_n24846_, new_n24847_, new_n24848_, new_n24849_, new_n24850_,
    new_n24851_, new_n24852_, new_n24853_, new_n24854_, new_n24856_,
    new_n24857_, new_n24858_, new_n24859_, new_n24860_, new_n24861_,
    new_n24863_, new_n24864_, new_n24865_, new_n24866_, new_n24867_,
    new_n24868_, new_n24869_, new_n24870_, new_n24871_, new_n24872_,
    new_n24873_, new_n24874_, new_n24875_, new_n24876_, new_n24877_,
    new_n24878_, new_n24879_, new_n24880_, new_n24881_, new_n24882_,
    new_n24883_, new_n24884_, new_n24885_, new_n24886_, new_n24887_,
    new_n24888_, new_n24889_, new_n24890_, new_n24891_, new_n24892_,
    new_n24893_, new_n24894_, new_n24895_, new_n24896_, new_n24897_,
    new_n24898_, new_n24899_, new_n24900_, new_n24901_, new_n24902_,
    new_n24903_, new_n24904_, new_n24905_, new_n24906_, new_n24907_,
    new_n24908_, new_n24909_, new_n24910_, new_n24911_, new_n24912_,
    new_n24913_, new_n24914_, new_n24915_, new_n24917_, new_n24918_,
    new_n24919_, new_n24920_, new_n24921_, new_n24922_, new_n24923_,
    new_n24924_, new_n24925_, new_n24926_, new_n24927_, new_n24928_,
    new_n24929_, new_n24930_, new_n24931_, new_n24932_, new_n24933_,
    new_n24934_, new_n24935_, new_n24936_, new_n24937_, new_n24938_,
    new_n24940_, new_n24941_, new_n24942_, new_n24943_, new_n24944_,
    new_n24945_, new_n24946_, new_n24947_, new_n24948_, new_n24949_,
    new_n24950_, new_n24951_, new_n24952_, new_n24954_, new_n24955_,
    new_n24956_, new_n24957_, new_n24958_, new_n24959_, new_n24960_,
    new_n24961_, new_n24962_, new_n24963_, new_n24964_, new_n24965_,
    new_n24966_, new_n24967_, new_n24968_, new_n24969_, new_n24970_,
    new_n24971_, new_n24972_, new_n24973_, new_n24974_, new_n24975_,
    new_n24976_, new_n24977_, new_n24978_, new_n24979_, new_n24980_,
    new_n24981_, new_n24982_, new_n24983_, new_n24984_, new_n24985_,
    new_n24986_, new_n24987_, new_n24988_, new_n24989_, new_n24990_,
    new_n24991_, new_n24992_, new_n24993_, new_n24994_, new_n24995_,
    new_n24996_, new_n24997_, new_n24998_, new_n24999_, new_n25000_,
    new_n25001_, new_n25002_, new_n25003_, new_n25004_, new_n25005_,
    new_n25006_, new_n25007_, new_n25008_, new_n25009_, new_n25010_,
    new_n25011_, new_n25012_, new_n25013_, new_n25014_, new_n25015_,
    new_n25016_, new_n25017_, new_n25018_, new_n25019_, new_n25020_,
    new_n25021_, new_n25022_, new_n25023_, new_n25024_, new_n25025_,
    new_n25026_, new_n25027_, new_n25028_, new_n25029_, new_n25030_,
    new_n25031_, new_n25032_, new_n25033_, new_n25034_, new_n25035_,
    new_n25036_, new_n25037_, new_n25038_, new_n25039_, new_n25040_,
    new_n25041_, new_n25042_, new_n25043_, new_n25044_, new_n25045_,
    new_n25046_, new_n25047_, new_n25048_, new_n25049_, new_n25050_,
    new_n25051_, new_n25052_, new_n25053_, new_n25054_, new_n25055_,
    new_n25056_, new_n25057_, new_n25058_, new_n25059_, new_n25060_,
    new_n25061_, new_n25062_, new_n25063_, new_n25064_, new_n25065_,
    new_n25066_, new_n25067_, new_n25068_, new_n25069_, new_n25070_,
    new_n25071_, new_n25072_, new_n25073_, new_n25074_, new_n25075_,
    new_n25076_, new_n25077_, new_n25078_, new_n25079_, new_n25080_,
    new_n25081_, new_n25082_, new_n25083_, new_n25084_, new_n25085_,
    new_n25086_, new_n25087_, new_n25088_, new_n25089_, new_n25090_,
    new_n25091_, new_n25092_, new_n25093_, new_n25094_, new_n25095_,
    new_n25096_, new_n25097_, new_n25098_, new_n25099_, new_n25100_,
    new_n25101_, new_n25102_, new_n25103_, new_n25104_, new_n25105_,
    new_n25106_, new_n25107_, new_n25108_, new_n25109_, new_n25110_,
    new_n25111_, new_n25112_, new_n25113_, new_n25114_, new_n25115_,
    new_n25116_, new_n25117_, new_n25118_, new_n25119_, new_n25120_,
    new_n25121_, new_n25122_, new_n25123_, new_n25124_, new_n25125_,
    new_n25126_, new_n25127_, new_n25128_, new_n25129_, new_n25130_,
    new_n25131_, new_n25132_, new_n25133_, new_n25134_, new_n25135_,
    new_n25136_, new_n25137_, new_n25138_, new_n25139_, new_n25140_,
    new_n25141_, new_n25142_, new_n25143_, new_n25144_, new_n25145_,
    new_n25146_, new_n25147_, new_n25148_, new_n25149_, new_n25150_,
    new_n25151_, new_n25152_, new_n25153_, new_n25154_, new_n25155_,
    new_n25156_, new_n25157_, new_n25158_, new_n25159_, new_n25160_,
    new_n25161_, new_n25162_, new_n25163_, new_n25164_, new_n25165_,
    new_n25166_, new_n25167_, new_n25168_, new_n25169_, new_n25170_,
    new_n25171_, new_n25172_, new_n25173_, new_n25174_, new_n25175_,
    new_n25176_, new_n25177_, new_n25178_, new_n25179_, new_n25180_,
    new_n25181_, new_n25182_, new_n25183_, new_n25184_, new_n25185_,
    new_n25186_, new_n25187_, new_n25188_, new_n25189_, new_n25190_,
    new_n25191_, new_n25192_, new_n25193_, new_n25194_, new_n25195_,
    new_n25196_, new_n25197_, new_n25198_, new_n25199_, new_n25200_,
    new_n25201_, new_n25202_, new_n25203_, new_n25204_, new_n25205_,
    new_n25206_, new_n25207_, new_n25208_, new_n25209_, new_n25210_,
    new_n25211_, new_n25212_, new_n25213_, new_n25214_, new_n25215_,
    new_n25216_, new_n25217_, new_n25218_, new_n25219_, new_n25220_,
    new_n25221_, new_n25222_, new_n25223_, new_n25224_, new_n25225_,
    new_n25226_, new_n25227_, new_n25228_, new_n25229_, new_n25230_,
    new_n25231_, new_n25232_, new_n25233_, new_n25234_, new_n25235_,
    new_n25236_, new_n25237_, new_n25238_, new_n25239_, new_n25240_,
    new_n25241_, new_n25242_, new_n25243_, new_n25244_, new_n25245_,
    new_n25246_, new_n25247_, new_n25248_, new_n25249_, new_n25250_,
    new_n25251_, new_n25253_, new_n25254_, new_n25255_, new_n25256_,
    new_n25257_, new_n25258_, new_n25259_, new_n25260_, new_n25261_,
    new_n25262_, new_n25263_, new_n25264_, new_n25265_, new_n25266_,
    new_n25267_, new_n25268_, new_n25269_, new_n25270_, new_n25271_,
    new_n25272_, new_n25273_, new_n25274_, new_n25275_, new_n25276_,
    new_n25277_, new_n25278_, new_n25279_, new_n25280_, new_n25281_,
    new_n25282_, new_n25283_, new_n25284_, new_n25285_, new_n25286_,
    new_n25287_, new_n25288_, new_n25289_, new_n25290_, new_n25291_,
    new_n25292_, new_n25293_, new_n25294_, new_n25295_, new_n25296_,
    new_n25297_, new_n25298_, new_n25299_, new_n25300_, new_n25301_,
    new_n25302_, new_n25303_, new_n25304_, new_n25305_, new_n25306_,
    new_n25307_, new_n25308_, new_n25309_, new_n25310_, new_n25311_,
    new_n25312_, new_n25313_, new_n25314_, new_n25315_, new_n25316_,
    new_n25317_, new_n25318_, new_n25319_, new_n25320_, new_n25321_,
    new_n25322_, new_n25323_, new_n25324_, new_n25325_, new_n25326_,
    new_n25327_, new_n25328_, new_n25329_, new_n25330_, new_n25331_,
    new_n25332_, new_n25333_, new_n25334_, new_n25335_, new_n25336_,
    new_n25337_, new_n25338_, new_n25339_, new_n25340_, new_n25341_,
    new_n25342_, new_n25343_, new_n25344_, new_n25345_, new_n25346_,
    new_n25347_, new_n25348_, new_n25349_, new_n25350_, new_n25351_,
    new_n25352_, new_n25353_, new_n25354_, new_n25355_, new_n25356_,
    new_n25357_, new_n25358_, new_n25359_, new_n25360_, new_n25361_,
    new_n25362_, new_n25363_, new_n25364_, new_n25365_, new_n25366_,
    new_n25367_, new_n25368_, new_n25369_, new_n25370_, new_n25371_,
    new_n25372_, new_n25373_, new_n25374_, new_n25375_, new_n25376_,
    new_n25377_, new_n25378_, new_n25379_, new_n25380_, new_n25381_,
    new_n25382_, new_n25383_, new_n25384_, new_n25385_, new_n25386_,
    new_n25387_, new_n25388_, new_n25389_, new_n25390_, new_n25391_,
    new_n25392_, new_n25393_, new_n25394_, new_n25395_, new_n25396_,
    new_n25397_, new_n25398_, new_n25399_, new_n25400_, new_n25401_,
    new_n25402_, new_n25403_, new_n25404_, new_n25405_, new_n25406_,
    new_n25407_, new_n25408_, new_n25409_, new_n25410_, new_n25411_,
    new_n25412_, new_n25413_, new_n25414_, new_n25415_, new_n25416_,
    new_n25417_, new_n25418_, new_n25419_, new_n25420_, new_n25421_,
    new_n25422_, new_n25423_, new_n25424_, new_n25425_, new_n25426_,
    new_n25427_, new_n25428_, new_n25429_, new_n25430_, new_n25431_,
    new_n25432_, new_n25433_, new_n25434_, new_n25435_, new_n25436_,
    new_n25437_, new_n25438_, new_n25439_, new_n25440_, new_n25441_,
    new_n25442_, new_n25443_, new_n25444_, new_n25445_, new_n25446_,
    new_n25447_, new_n25448_, new_n25449_, new_n25450_, new_n25451_,
    new_n25452_, new_n25453_, new_n25454_, new_n25455_, new_n25456_,
    new_n25457_, new_n25458_, new_n25459_, new_n25460_, new_n25461_,
    new_n25462_, new_n25463_, new_n25464_, new_n25465_, new_n25466_,
    new_n25467_, new_n25468_, new_n25469_, new_n25470_, new_n25471_,
    new_n25472_, new_n25473_, new_n25474_, new_n25475_, new_n25476_,
    new_n25478_, new_n25479_, new_n25480_, new_n25481_, new_n25482_,
    new_n25483_, new_n25484_, new_n25485_, new_n25486_, new_n25487_,
    new_n25488_, new_n25489_, new_n25490_, new_n25491_, new_n25492_,
    new_n25493_, new_n25494_, new_n25495_, new_n25496_, new_n25497_,
    new_n25498_, new_n25499_, new_n25500_, new_n25501_, new_n25502_,
    new_n25503_, new_n25504_, new_n25505_, new_n25506_, new_n25507_,
    new_n25508_, new_n25509_, new_n25510_, new_n25511_, new_n25512_,
    new_n25513_, new_n25514_, new_n25515_, new_n25516_, new_n25517_,
    new_n25518_, new_n25519_, new_n25520_, new_n25521_, new_n25522_,
    new_n25523_, new_n25524_, new_n25525_, new_n25526_, new_n25527_,
    new_n25528_, new_n25529_, new_n25530_, new_n25531_, new_n25532_,
    new_n25533_, new_n25534_, new_n25535_, new_n25536_, new_n25537_,
    new_n25538_, new_n25539_, new_n25540_, new_n25541_, new_n25542_,
    new_n25543_, new_n25544_, new_n25545_, new_n25546_, new_n25547_,
    new_n25548_, new_n25549_, new_n25550_, new_n25551_, new_n25552_,
    new_n25553_, new_n25554_, new_n25555_, new_n25556_, new_n25557_,
    new_n25558_, new_n25559_, new_n25560_, new_n25561_, new_n25562_,
    new_n25563_, new_n25564_, new_n25565_, new_n25566_, new_n25567_,
    new_n25568_, new_n25569_, new_n25570_, new_n25571_, new_n25572_,
    new_n25573_, new_n25574_, new_n25575_, new_n25576_, new_n25577_,
    new_n25578_, new_n25579_, new_n25580_, new_n25581_, new_n25582_,
    new_n25583_, new_n25584_, new_n25585_, new_n25586_, new_n25587_,
    new_n25588_, new_n25589_, new_n25590_, new_n25591_, new_n25592_,
    new_n25593_, new_n25594_, new_n25595_, new_n25596_, new_n25597_,
    new_n25598_, new_n25599_, new_n25600_, new_n25601_, new_n25602_,
    new_n25603_, new_n25604_, new_n25605_, new_n25606_, new_n25607_,
    new_n25608_, new_n25609_, new_n25610_, new_n25611_, new_n25612_,
    new_n25613_, new_n25615_, new_n25616_, new_n25617_, new_n25618_,
    new_n25619_, new_n25620_, new_n25622_, new_n25623_, new_n25624_,
    new_n25625_, new_n25626_, new_n25627_, new_n25628_, new_n25629_,
    new_n25630_, new_n25631_, new_n25632_, new_n25633_, new_n25634_,
    new_n25635_, new_n25636_, new_n25637_, new_n25638_, new_n25639_,
    new_n25640_, new_n25641_, new_n25642_, new_n25643_, new_n25644_,
    new_n25645_, new_n25646_, new_n25647_, new_n25648_, new_n25649_,
    new_n25650_, new_n25651_, new_n25652_, new_n25653_, new_n25654_,
    new_n25655_, new_n25656_, new_n25657_, new_n25658_, new_n25659_,
    new_n25660_, new_n25661_, new_n25662_, new_n25663_, new_n25664_,
    new_n25665_, new_n25666_, new_n25667_, new_n25668_, new_n25669_,
    new_n25670_, new_n25671_, new_n25672_, new_n25673_, new_n25674_,
    new_n25675_, new_n25676_, new_n25677_, new_n25678_, new_n25679_,
    new_n25680_, new_n25681_, new_n25682_, new_n25683_, new_n25684_,
    new_n25685_, new_n25686_, new_n25687_, new_n25688_, new_n25689_,
    new_n25690_, new_n25691_, new_n25692_, new_n25693_, new_n25694_,
    new_n25695_, new_n25696_, new_n25697_, new_n25698_, new_n25699_,
    new_n25700_, new_n25701_, new_n25702_, new_n25703_, new_n25704_,
    new_n25705_, new_n25706_, new_n25707_, new_n25708_, new_n25709_,
    new_n25710_, new_n25711_, new_n25712_, new_n25713_, new_n25714_,
    new_n25715_, new_n25716_, new_n25717_, new_n25718_, new_n25719_,
    new_n25720_, new_n25721_, new_n25722_, new_n25723_, new_n25724_,
    new_n25725_, new_n25726_, new_n25727_, new_n25728_, new_n25729_,
    new_n25730_, new_n25731_, new_n25732_, new_n25733_, new_n25734_,
    new_n25735_, new_n25736_, new_n25737_, new_n25738_, new_n25739_,
    new_n25740_, new_n25741_, new_n25742_, new_n25743_, new_n25744_,
    new_n25745_, new_n25746_, new_n25747_, new_n25748_, new_n25749_,
    new_n25750_, new_n25751_, new_n25752_, new_n25753_, new_n25754_,
    new_n25755_, new_n25756_, new_n25757_, new_n25758_, new_n25759_,
    new_n25760_, new_n25761_, new_n25762_, new_n25763_, new_n25764_,
    new_n25765_, new_n25766_, new_n25767_, new_n25768_, new_n25769_,
    new_n25770_, new_n25771_, new_n25772_, new_n25773_, new_n25774_,
    new_n25775_, new_n25776_, new_n25777_, new_n25778_, new_n25779_,
    new_n25780_, new_n25781_, new_n25782_, new_n25783_, new_n25784_,
    new_n25785_, new_n25786_, new_n25787_, new_n25788_, new_n25789_,
    new_n25790_, new_n25791_, new_n25792_, new_n25793_, new_n25794_,
    new_n25796_, new_n25797_, new_n25798_, new_n25799_, new_n25800_,
    new_n25801_, new_n25802_, new_n25803_, new_n25804_, new_n25805_,
    new_n25806_, new_n25807_, new_n25808_, new_n25809_, new_n25810_,
    new_n25811_, new_n25812_, new_n25813_, new_n25814_, new_n25815_,
    new_n25816_, new_n25817_, new_n25818_, new_n25819_, new_n25820_,
    new_n25821_, new_n25822_, new_n25823_, new_n25824_, new_n25825_,
    new_n25826_, new_n25827_, new_n25828_, new_n25829_, new_n25830_,
    new_n25831_, new_n25832_, new_n25833_, new_n25834_, new_n25835_,
    new_n25836_, new_n25837_, new_n25838_, new_n25839_, new_n25840_,
    new_n25841_, new_n25842_, new_n25843_, new_n25844_, new_n25845_,
    new_n25846_, new_n25847_, new_n25848_, new_n25849_, new_n25850_,
    new_n25851_, new_n25852_, new_n25853_, new_n25854_, new_n25855_,
    new_n25856_, new_n25857_, new_n25858_, new_n25859_, new_n25860_,
    new_n25861_, new_n25862_, new_n25863_, new_n25864_, new_n25865_,
    new_n25866_, new_n25867_, new_n25868_, new_n25869_, new_n25870_,
    new_n25871_, new_n25872_, new_n25873_, new_n25874_, new_n25875_,
    new_n25876_, new_n25877_, new_n25878_, new_n25879_, new_n25880_,
    new_n25881_, new_n25882_, new_n25883_, new_n25884_, new_n25885_,
    new_n25886_, new_n25887_, new_n25888_, new_n25889_, new_n25890_,
    new_n25891_, new_n25892_, new_n25893_, new_n25894_, new_n25895_,
    new_n25896_, new_n25897_, new_n25898_, new_n25899_, new_n25900_,
    new_n25901_, new_n25902_, new_n25903_, new_n25904_, new_n25905_,
    new_n25906_, new_n25907_, new_n25908_, new_n25909_, new_n25910_,
    new_n25911_, new_n25912_, new_n25913_, new_n25914_, new_n25915_,
    new_n25916_, new_n25917_, new_n25918_, new_n25919_, new_n25920_,
    new_n25921_, new_n25922_, new_n25923_, new_n25924_, new_n25925_,
    new_n25926_, new_n25927_, new_n25928_, new_n25929_, new_n25930_,
    new_n25931_, new_n25932_, new_n25933_, new_n25934_, new_n25935_,
    new_n25936_, new_n25937_, new_n25938_, new_n25939_, new_n25940_,
    new_n25941_, new_n25942_, new_n25943_, new_n25944_, new_n25945_,
    new_n25946_, new_n25947_, new_n25948_, new_n25949_, new_n25950_,
    new_n25951_, new_n25952_, new_n25953_, new_n25954_, new_n25955_,
    new_n25956_, new_n25957_, new_n25958_, new_n25959_, new_n25960_,
    new_n25961_, new_n25962_, new_n25963_, new_n25964_, new_n25965_,
    new_n25966_, new_n25967_, new_n25968_, new_n25969_, new_n25970_,
    new_n25971_, new_n25972_, new_n25973_, new_n25974_, new_n25975_,
    new_n25976_, new_n25977_, new_n25978_, new_n25979_, new_n25980_,
    new_n25981_, new_n25982_, new_n25983_, new_n25984_, new_n25985_,
    new_n25986_, new_n25987_, new_n25988_, new_n25989_, new_n25990_,
    new_n25991_, new_n25992_, new_n25993_, new_n25994_, new_n25995_,
    new_n25996_, new_n25997_, new_n25998_, new_n25999_, new_n26000_,
    new_n26001_, new_n26002_, new_n26003_, new_n26004_, new_n26005_,
    new_n26006_, new_n26007_, new_n26008_, new_n26009_, new_n26010_,
    new_n26011_, new_n26012_, new_n26013_, new_n26014_, new_n26015_,
    new_n26016_, new_n26017_, new_n26018_, new_n26019_, new_n26020_,
    new_n26021_, new_n26022_, new_n26023_, new_n26024_, new_n26025_,
    new_n26026_, new_n26028_, new_n26029_, new_n26030_, new_n26031_,
    new_n26032_, new_n26033_, new_n26034_, new_n26035_, new_n26036_,
    new_n26037_, new_n26038_, new_n26039_, new_n26040_, new_n26041_,
    new_n26042_, new_n26043_, new_n26044_, new_n26045_, new_n26046_,
    new_n26047_, new_n26048_, new_n26049_, new_n26050_, new_n26051_,
    new_n26052_, new_n26053_, new_n26054_, new_n26055_, new_n26056_,
    new_n26057_, new_n26058_, new_n26059_, new_n26060_, new_n26061_,
    new_n26062_, new_n26063_, new_n26064_, new_n26065_, new_n26066_,
    new_n26067_, new_n26068_, new_n26069_, new_n26070_, new_n26071_,
    new_n26072_, new_n26073_, new_n26074_, new_n26075_, new_n26076_,
    new_n26077_, new_n26078_, new_n26079_, new_n26080_, new_n26081_,
    new_n26082_, new_n26083_, new_n26084_, new_n26085_, new_n26086_,
    new_n26087_, new_n26088_, new_n26089_, new_n26091_, new_n26092_,
    new_n26093_, new_n26094_, new_n26095_, new_n26096_, new_n26097_,
    new_n26098_, new_n26099_, new_n26100_, new_n26101_, new_n26102_,
    new_n26103_, new_n26104_, new_n26105_, new_n26106_, new_n26107_,
    new_n26108_, new_n26109_, new_n26110_, new_n26111_, new_n26112_,
    new_n26113_, new_n26114_, new_n26115_, new_n26116_, new_n26117_,
    new_n26118_, new_n26119_, new_n26120_, new_n26121_, new_n26122_,
    new_n26123_, new_n26124_, new_n26125_, new_n26126_, new_n26127_,
    new_n26128_, new_n26129_, new_n26130_, new_n26131_, new_n26132_,
    new_n26133_, new_n26134_, new_n26135_, new_n26136_, new_n26137_,
    new_n26138_, new_n26139_, new_n26140_, new_n26141_, new_n26142_,
    new_n26143_, new_n26144_, new_n26145_, new_n26146_, new_n26147_,
    new_n26148_, new_n26149_, new_n26150_, new_n26151_, new_n26152_,
    new_n26153_, new_n26154_, new_n26155_, new_n26156_, new_n26157_,
    new_n26158_, new_n26159_, new_n26160_, new_n26161_, new_n26162_,
    new_n26163_, new_n26164_, new_n26165_, new_n26166_, new_n26167_,
    new_n26168_, new_n26169_, new_n26170_, new_n26171_, new_n26172_,
    new_n26173_, new_n26174_, new_n26175_, new_n26176_, new_n26177_,
    new_n26178_, new_n26179_, new_n26180_, new_n26181_, new_n26182_,
    new_n26183_, new_n26184_, new_n26185_, new_n26186_, new_n26187_,
    new_n26188_, new_n26189_, new_n26190_, new_n26191_, new_n26192_,
    new_n26193_, new_n26194_, new_n26195_, new_n26196_, new_n26197_,
    new_n26198_, new_n26199_, new_n26200_, new_n26201_, new_n26202_,
    new_n26203_, new_n26204_, new_n26205_, new_n26206_, new_n26207_,
    new_n26208_, new_n26209_, new_n26210_, new_n26211_, new_n26212_,
    new_n26213_, new_n26214_, new_n26215_, new_n26216_, new_n26217_,
    new_n26218_, new_n26219_, new_n26220_, new_n26221_, new_n26222_,
    new_n26223_, new_n26224_, new_n26225_, new_n26226_, new_n26227_,
    new_n26228_, new_n26229_, new_n26230_, new_n26231_, new_n26232_,
    new_n26233_, new_n26234_, new_n26235_, new_n26236_, new_n26237_,
    new_n26238_, new_n26239_, new_n26240_, new_n26241_, new_n26242_,
    new_n26243_, new_n26244_, new_n26245_, new_n26246_, new_n26247_,
    new_n26248_, new_n26249_, new_n26250_, new_n26251_, new_n26252_,
    new_n26253_, new_n26254_, new_n26255_, new_n26256_, new_n26257_,
    new_n26258_, new_n26259_, new_n26260_, new_n26261_, new_n26262_,
    new_n26263_, new_n26264_, new_n26265_, new_n26266_, new_n26267_,
    new_n26268_, new_n26269_, new_n26270_, new_n26271_, new_n26272_,
    new_n26273_, new_n26274_, new_n26275_, new_n26276_, new_n26277_,
    new_n26278_, new_n26279_, new_n26280_, new_n26281_, new_n26282_,
    new_n26283_, new_n26284_, new_n26285_, new_n26286_, new_n26287_,
    new_n26288_, new_n26289_, new_n26290_, new_n26291_, new_n26292_,
    new_n26293_, new_n26294_, new_n26295_, new_n26296_, new_n26297_,
    new_n26298_, new_n26299_, new_n26300_, new_n26301_, new_n26302_,
    new_n26303_, new_n26304_, new_n26305_, new_n26306_, new_n26307_,
    new_n26308_, new_n26309_, new_n26310_, new_n26311_, new_n26312_,
    new_n26313_, new_n26314_, new_n26315_, new_n26316_, new_n26317_,
    new_n26318_, new_n26319_, new_n26320_, new_n26321_, new_n26322_,
    new_n26323_, new_n26324_, new_n26325_, new_n26326_, new_n26327_,
    new_n26328_, new_n26329_, new_n26330_, new_n26331_, new_n26332_,
    new_n26333_, new_n26334_, new_n26335_, new_n26336_, new_n26337_,
    new_n26338_, new_n26339_, new_n26340_, new_n26341_, new_n26342_,
    new_n26343_, new_n26344_, new_n26345_, new_n26346_, new_n26347_,
    new_n26348_, new_n26349_, new_n26350_, new_n26351_, new_n26352_,
    new_n26353_, new_n26354_, new_n26355_, new_n26356_, new_n26357_,
    new_n26358_, new_n26359_, new_n26360_, new_n26361_, new_n26362_,
    new_n26363_, new_n26364_, new_n26365_, new_n26366_, new_n26367_,
    new_n26368_, new_n26369_, new_n26370_, new_n26371_, new_n26372_,
    new_n26373_, new_n26374_, new_n26375_, new_n26376_, new_n26377_,
    new_n26378_, new_n26379_, new_n26380_, new_n26381_, new_n26382_,
    new_n26383_, new_n26384_, new_n26385_, new_n26386_, new_n26387_,
    new_n26388_, new_n26389_, new_n26390_, new_n26391_, new_n26392_,
    new_n26393_, new_n26394_, new_n26395_, new_n26396_, new_n26397_,
    new_n26398_, new_n26399_, new_n26400_, new_n26401_, new_n26402_,
    new_n26403_, new_n26404_, new_n26405_, new_n26406_, new_n26407_,
    new_n26408_, new_n26409_, new_n26410_, new_n26411_, new_n26412_,
    new_n26413_, new_n26414_, new_n26416_, new_n26417_, new_n26418_,
    new_n26419_, new_n26420_, new_n26421_, new_n26422_, new_n26423_,
    new_n26424_, new_n26425_, new_n26426_, new_n26427_, new_n26428_,
    new_n26429_, new_n26430_, new_n26431_, new_n26432_, new_n26433_,
    new_n26434_, new_n26435_, new_n26436_, new_n26437_, new_n26438_,
    new_n26439_, new_n26440_, new_n26441_, new_n26442_, new_n26443_,
    new_n26444_, new_n26445_, new_n26446_, new_n26447_, new_n26448_,
    new_n26449_, new_n26450_, new_n26451_, new_n26452_, new_n26453_,
    new_n26454_, new_n26455_, new_n26456_, new_n26457_, new_n26458_,
    new_n26459_, new_n26460_, new_n26461_, new_n26462_, new_n26463_,
    new_n26464_, new_n26465_, new_n26466_, new_n26467_, new_n26468_,
    new_n26469_, new_n26470_, new_n26471_, new_n26472_, new_n26473_,
    new_n26474_, new_n26475_, new_n26476_, new_n26477_, new_n26478_,
    new_n26479_, new_n26480_, new_n26481_, new_n26482_, new_n26483_,
    new_n26484_, new_n26485_, new_n26486_, new_n26487_, new_n26488_,
    new_n26489_, new_n26490_, new_n26491_, new_n26492_, new_n26493_,
    new_n26494_, new_n26495_, new_n26496_, new_n26497_, new_n26498_,
    new_n26499_, new_n26500_, new_n26501_, new_n26502_, new_n26503_,
    new_n26504_, new_n26505_, new_n26506_, new_n26507_, new_n26508_,
    new_n26509_, new_n26510_, new_n26511_, new_n26512_, new_n26513_,
    new_n26514_, new_n26515_, new_n26516_, new_n26517_, new_n26518_,
    new_n26519_, new_n26520_, new_n26521_, new_n26522_, new_n26523_,
    new_n26524_, new_n26525_, new_n26526_, new_n26527_, new_n26528_,
    new_n26529_, new_n26530_, new_n26531_, new_n26532_, new_n26533_,
    new_n26534_, new_n26535_, new_n26536_, new_n26537_, new_n26538_,
    new_n26539_, new_n26540_, new_n26541_, new_n26542_, new_n26543_,
    new_n26544_, new_n26545_, new_n26546_, new_n26547_, new_n26548_,
    new_n26549_, new_n26550_, new_n26551_, new_n26552_, new_n26553_,
    new_n26554_, new_n26555_, new_n26556_, new_n26557_, new_n26558_,
    new_n26559_, new_n26560_, new_n26561_, new_n26562_, new_n26563_,
    new_n26564_, new_n26565_, new_n26566_, new_n26567_, new_n26568_,
    new_n26569_, new_n26570_, new_n26571_, new_n26572_, new_n26573_,
    new_n26574_, new_n26575_, new_n26576_, new_n26577_, new_n26578_,
    new_n26579_, new_n26580_, new_n26581_, new_n26582_, new_n26583_,
    new_n26584_, new_n26585_, new_n26586_, new_n26587_, new_n26588_,
    new_n26589_, new_n26590_, new_n26591_, new_n26592_, new_n26593_,
    new_n26594_, new_n26595_, new_n26596_, new_n26597_, new_n26598_,
    new_n26599_, new_n26600_, new_n26601_, new_n26602_, new_n26603_,
    new_n26604_, new_n26605_, new_n26606_, new_n26607_, new_n26608_,
    new_n26609_, new_n26610_, new_n26611_, new_n26612_, new_n26613_,
    new_n26615_, new_n26616_, new_n26617_, new_n26618_, new_n26619_,
    new_n26620_, new_n26621_, new_n26622_, new_n26623_, new_n26624_,
    new_n26625_, new_n26626_, new_n26627_, new_n26628_, new_n26629_,
    new_n26630_, new_n26631_, new_n26632_, new_n26633_, new_n26634_,
    new_n26635_, new_n26636_, new_n26637_, new_n26638_, new_n26639_,
    new_n26640_, new_n26641_, new_n26642_, new_n26643_, new_n26644_,
    new_n26645_, new_n26646_, new_n26647_, new_n26648_, new_n26649_,
    new_n26650_, new_n26651_, new_n26652_, new_n26653_, new_n26654_,
    new_n26655_, new_n26656_, new_n26657_, new_n26658_, new_n26659_,
    new_n26660_, new_n26661_, new_n26662_, new_n26663_, new_n26664_,
    new_n26665_, new_n26666_, new_n26667_, new_n26668_, new_n26669_,
    new_n26670_, new_n26671_, new_n26673_, new_n26674_, new_n26675_,
    new_n26676_, new_n26677_, new_n26678_, new_n26679_, new_n26680_,
    new_n26681_, new_n26682_, new_n26683_, new_n26684_, new_n26685_,
    new_n26686_, new_n26687_, new_n26688_, new_n26689_, new_n26690_,
    new_n26691_, new_n26692_, new_n26693_, new_n26694_, new_n26695_,
    new_n26696_, new_n26697_, new_n26698_, new_n26699_, new_n26700_,
    new_n26701_, new_n26702_, new_n26703_, new_n26704_, new_n26705_,
    new_n26706_, new_n26707_, new_n26708_, new_n26709_, new_n26710_,
    new_n26711_, new_n26712_, new_n26713_, new_n26714_, new_n26715_,
    new_n26716_, new_n26717_, new_n26718_, new_n26719_, new_n26720_,
    new_n26721_, new_n26722_, new_n26723_, new_n26724_, new_n26725_,
    new_n26726_, new_n26727_, new_n26728_, new_n26729_, new_n26730_,
    new_n26731_, new_n26732_, new_n26733_, new_n26734_, new_n26735_,
    new_n26736_, new_n26737_, new_n26738_, new_n26739_, new_n26740_,
    new_n26741_, new_n26742_, new_n26743_, new_n26744_, new_n26745_,
    new_n26746_, new_n26747_, new_n26748_, new_n26749_, new_n26750_,
    new_n26751_, new_n26752_, new_n26753_, new_n26754_, new_n26755_,
    new_n26756_, new_n26757_, new_n26758_, new_n26759_, new_n26760_,
    new_n26761_, new_n26762_, new_n26763_, new_n26764_, new_n26765_,
    new_n26766_, new_n26767_, new_n26768_, new_n26769_, new_n26770_,
    new_n26771_, new_n26772_, new_n26773_, new_n26774_, new_n26775_,
    new_n26776_, new_n26777_, new_n26778_, new_n26779_, new_n26780_,
    new_n26781_, new_n26782_, new_n26783_, new_n26784_, new_n26785_,
    new_n26786_, new_n26787_, new_n26788_, new_n26789_, new_n26790_,
    new_n26791_, new_n26792_, new_n26793_, new_n26794_, new_n26795_,
    new_n26796_, new_n26797_, new_n26798_, new_n26799_, new_n26800_,
    new_n26801_, new_n26802_, new_n26803_, new_n26804_, new_n26805_,
    new_n26806_, new_n26807_, new_n26808_, new_n26809_, new_n26810_,
    new_n26811_, new_n26812_, new_n26813_, new_n26814_, new_n26815_,
    new_n26816_, new_n26817_, new_n26818_, new_n26819_, new_n26820_,
    new_n26821_, new_n26822_, new_n26823_, new_n26824_, new_n26825_,
    new_n26826_, new_n26827_, new_n26828_, new_n26829_, new_n26830_,
    new_n26831_, new_n26832_, new_n26833_, new_n26834_, new_n26835_,
    new_n26836_, new_n26837_, new_n26838_, new_n26839_, new_n26840_,
    new_n26841_, new_n26842_, new_n26843_, new_n26844_, new_n26845_,
    new_n26846_, new_n26847_, new_n26848_, new_n26849_, new_n26850_,
    new_n26851_, new_n26852_, new_n26853_, new_n26854_, new_n26855_,
    new_n26856_, new_n26857_, new_n26858_, new_n26859_, new_n26860_,
    new_n26861_, new_n26862_, new_n26863_, new_n26864_, new_n26865_,
    new_n26866_, new_n26867_, new_n26868_, new_n26869_, new_n26870_,
    new_n26871_, new_n26872_, new_n26873_, new_n26874_, new_n26875_,
    new_n26876_, new_n26877_, new_n26878_, new_n26879_, new_n26880_,
    new_n26881_, new_n26882_, new_n26883_, new_n26884_, new_n26885_,
    new_n26886_, new_n26887_, new_n26888_, new_n26889_, new_n26890_,
    new_n26891_, new_n26892_, new_n26893_, new_n26894_, new_n26895_,
    new_n26896_, new_n26897_, new_n26898_, new_n26899_, new_n26900_,
    new_n26901_, new_n26902_, new_n26903_, new_n26904_, new_n26905_,
    new_n26906_, new_n26907_, new_n26908_, new_n26910_, new_n26911_,
    new_n26912_, new_n26913_, new_n26914_, new_n26915_, new_n26916_,
    new_n26917_, new_n26918_, new_n26919_, new_n26920_, new_n26921_,
    new_n26922_, new_n26923_, new_n26924_, new_n26925_, new_n26926_,
    new_n26927_, new_n26928_, new_n26929_, new_n26930_, new_n26931_,
    new_n26932_, new_n26933_, new_n26934_, new_n26935_, new_n26936_,
    new_n26937_, new_n26938_, new_n26939_, new_n26940_, new_n26941_,
    new_n26943_, new_n26944_, new_n26945_, new_n26946_, new_n26947_,
    new_n26948_, new_n26949_, new_n26950_, new_n26951_, new_n26952_,
    new_n26953_, new_n26954_, new_n26955_, new_n26956_, new_n26957_,
    new_n26958_, new_n26959_, new_n26960_, new_n26961_, new_n26962_,
    new_n26963_, new_n26964_, new_n26965_, new_n26966_, new_n26967_,
    new_n26968_, new_n26969_, new_n26970_, new_n26971_, new_n26972_,
    new_n26973_, new_n26974_, new_n26975_, new_n26976_, new_n26977_,
    new_n26978_, new_n26979_, new_n26980_, new_n26981_, new_n26982_,
    new_n26983_, new_n26984_, new_n26985_, new_n26986_, new_n26987_,
    new_n26988_, new_n26989_, new_n26990_, new_n26991_, new_n26992_,
    new_n26993_, new_n26994_, new_n26995_, new_n26996_, new_n26997_,
    new_n26998_, new_n26999_, new_n27000_, new_n27001_, new_n27002_,
    new_n27003_, new_n27004_, new_n27005_, new_n27006_, new_n27007_,
    new_n27008_, new_n27009_, new_n27010_, new_n27011_, new_n27012_,
    new_n27013_, new_n27014_, new_n27015_, new_n27016_, new_n27017_,
    new_n27018_, new_n27019_, new_n27020_, new_n27021_, new_n27022_,
    new_n27023_, new_n27024_, new_n27025_, new_n27026_, new_n27027_,
    new_n27028_, new_n27029_, new_n27030_, new_n27031_, new_n27032_,
    new_n27033_, new_n27034_, new_n27035_, new_n27036_, new_n27037_,
    new_n27038_, new_n27039_, new_n27040_, new_n27041_, new_n27042_,
    new_n27043_, new_n27044_, new_n27045_, new_n27046_, new_n27047_,
    new_n27048_, new_n27049_, new_n27050_, new_n27051_, new_n27052_,
    new_n27053_, new_n27054_, new_n27055_, new_n27056_, new_n27057_,
    new_n27058_, new_n27059_, new_n27060_, new_n27061_, new_n27062_,
    new_n27063_, new_n27064_, new_n27065_, new_n27066_, new_n27067_,
    new_n27068_, new_n27069_, new_n27070_, new_n27071_, new_n27072_,
    new_n27073_, new_n27074_, new_n27075_, new_n27076_, new_n27077_,
    new_n27078_, new_n27079_, new_n27080_, new_n27081_, new_n27082_,
    new_n27083_, new_n27084_, new_n27085_, new_n27086_, new_n27087_,
    new_n27088_, new_n27089_, new_n27090_, new_n27091_, new_n27092_,
    new_n27093_, new_n27094_, new_n27095_, new_n27096_, new_n27097_,
    new_n27098_, new_n27099_, new_n27100_, new_n27101_, new_n27102_,
    new_n27103_, new_n27104_, new_n27105_, new_n27106_, new_n27107_,
    new_n27108_, new_n27109_, new_n27110_, new_n27111_, new_n27112_,
    new_n27113_, new_n27114_, new_n27115_, new_n27116_, new_n27117_,
    new_n27119_, new_n27120_, new_n27121_, new_n27122_, new_n27123_,
    new_n27124_, new_n27125_, new_n27126_, new_n27127_, new_n27128_,
    new_n27129_, new_n27130_, new_n27131_, new_n27132_, new_n27133_,
    new_n27134_, new_n27135_, new_n27136_, new_n27137_, new_n27138_,
    new_n27139_, new_n27140_, new_n27141_, new_n27142_, new_n27143_,
    new_n27144_, new_n27145_, new_n27146_, new_n27147_, new_n27148_,
    new_n27149_, new_n27150_, new_n27151_, new_n27152_, new_n27153_,
    new_n27154_, new_n27155_, new_n27156_, new_n27157_, new_n27158_,
    new_n27159_, new_n27160_, new_n27161_, new_n27162_, new_n27163_,
    new_n27164_, new_n27165_, new_n27166_, new_n27167_, new_n27168_,
    new_n27169_, new_n27170_, new_n27171_, new_n27172_, new_n27173_,
    new_n27174_, new_n27175_, new_n27176_, new_n27177_, new_n27178_,
    new_n27179_, new_n27180_, new_n27181_, new_n27182_, new_n27183_,
    new_n27184_, new_n27185_, new_n27186_, new_n27187_, new_n27188_,
    new_n27189_, new_n27190_, new_n27191_, new_n27192_, new_n27193_,
    new_n27194_, new_n27195_, new_n27196_, new_n27197_, new_n27198_,
    new_n27199_, new_n27200_, new_n27201_, new_n27202_, new_n27203_,
    new_n27204_, new_n27205_, new_n27206_, new_n27207_, new_n27208_,
    new_n27209_, new_n27210_, new_n27211_, new_n27212_, new_n27213_,
    new_n27214_, new_n27215_, new_n27216_, new_n27217_, new_n27218_,
    new_n27219_, new_n27220_, new_n27221_, new_n27222_, new_n27223_,
    new_n27224_, new_n27225_, new_n27226_, new_n27227_, new_n27228_,
    new_n27229_, new_n27230_, new_n27231_, new_n27232_, new_n27233_,
    new_n27234_, new_n27235_, new_n27236_, new_n27237_, new_n27238_,
    new_n27239_, new_n27240_, new_n27241_, new_n27242_, new_n27243_,
    new_n27244_, new_n27245_, new_n27246_, new_n27247_, new_n27248_,
    new_n27249_, new_n27250_, new_n27251_, new_n27252_, new_n27253_,
    new_n27254_, new_n27255_, new_n27256_, new_n27257_, new_n27258_,
    new_n27259_, new_n27260_, new_n27261_, new_n27262_, new_n27263_,
    new_n27264_, new_n27265_, new_n27266_, new_n27267_, new_n27268_,
    new_n27269_, new_n27270_, new_n27271_, new_n27272_, new_n27273_,
    new_n27274_, new_n27275_, new_n27276_, new_n27277_, new_n27278_,
    new_n27279_, new_n27280_, new_n27281_, new_n27282_, new_n27283_,
    new_n27284_, new_n27285_, new_n27286_, new_n27287_, new_n27288_,
    new_n27289_, new_n27290_, new_n27291_, new_n27292_, new_n27293_,
    new_n27294_, new_n27296_, new_n27297_, new_n27298_, new_n27299_,
    new_n27300_, new_n27301_, new_n27302_, new_n27303_, new_n27304_,
    new_n27305_, new_n27306_, new_n27307_, new_n27308_, new_n27309_,
    new_n27310_, new_n27311_, new_n27312_, new_n27313_, new_n27314_,
    new_n27315_, new_n27316_, new_n27317_, new_n27318_, new_n27319_,
    new_n27320_, new_n27321_, new_n27322_, new_n27323_, new_n27324_,
    new_n27325_, new_n27326_, new_n27327_, new_n27328_, new_n27329_,
    new_n27330_, new_n27331_, new_n27332_, new_n27333_, new_n27334_,
    new_n27335_, new_n27336_, new_n27337_, new_n27338_, new_n27339_,
    new_n27340_, new_n27341_, new_n27342_, new_n27343_, new_n27344_,
    new_n27345_, new_n27346_, new_n27347_, new_n27348_, new_n27349_,
    new_n27350_, new_n27351_, new_n27352_, new_n27353_, new_n27354_,
    new_n27355_, new_n27356_, new_n27357_, new_n27358_, new_n27359_,
    new_n27360_, new_n27361_, new_n27362_, new_n27363_, new_n27364_,
    new_n27365_, new_n27366_, new_n27367_, new_n27368_, new_n27369_,
    new_n27370_, new_n27371_, new_n27372_, new_n27373_, new_n27374_,
    new_n27375_, new_n27376_, new_n27377_, new_n27378_, new_n27379_,
    new_n27380_, new_n27381_, new_n27382_, new_n27383_, new_n27384_,
    new_n27385_, new_n27386_, new_n27387_, new_n27388_, new_n27389_,
    new_n27390_, new_n27391_, new_n27392_, new_n27393_, new_n27394_,
    new_n27395_, new_n27396_, new_n27397_, new_n27398_, new_n27399_,
    new_n27400_, new_n27401_, new_n27402_, new_n27403_, new_n27404_,
    new_n27405_, new_n27406_, new_n27407_, new_n27408_, new_n27409_,
    new_n27410_, new_n27411_, new_n27412_, new_n27413_, new_n27414_,
    new_n27415_, new_n27416_, new_n27417_, new_n27418_, new_n27419_,
    new_n27420_, new_n27421_, new_n27422_, new_n27423_, new_n27424_,
    new_n27425_, new_n27426_, new_n27427_, new_n27428_, new_n27429_,
    new_n27430_, new_n27431_, new_n27432_, new_n27433_, new_n27434_,
    new_n27435_, new_n27436_, new_n27437_, new_n27438_, new_n27439_,
    new_n27440_, new_n27441_, new_n27442_, new_n27443_, new_n27444_,
    new_n27445_, new_n27446_, new_n27447_, new_n27448_, new_n27449_,
    new_n27450_, new_n27451_, new_n27452_, new_n27453_, new_n27454_,
    new_n27456_, new_n27457_, new_n27458_, new_n27459_, new_n27460_,
    new_n27461_, new_n27462_, new_n27463_, new_n27464_, new_n27465_,
    new_n27466_, new_n27467_, new_n27468_, new_n27469_, new_n27470_,
    new_n27471_, new_n27472_, new_n27473_, new_n27474_, new_n27475_,
    new_n27476_, new_n27477_, new_n27478_, new_n27479_, new_n27480_,
    new_n27481_, new_n27482_, new_n27483_, new_n27484_, new_n27485_,
    new_n27486_, new_n27487_, new_n27488_, new_n27489_, new_n27490_,
    new_n27491_, new_n27492_, new_n27493_, new_n27494_, new_n27495_,
    new_n27496_, new_n27497_, new_n27498_, new_n27499_, new_n27500_,
    new_n27501_, new_n27502_, new_n27503_, new_n27504_, new_n27505_,
    new_n27506_, new_n27507_, new_n27508_, new_n27509_, new_n27510_,
    new_n27511_, new_n27512_, new_n27513_, new_n27514_, new_n27515_,
    new_n27516_, new_n27517_, new_n27518_, new_n27519_, new_n27520_,
    new_n27521_, new_n27522_, new_n27523_, new_n27524_, new_n27525_,
    new_n27526_, new_n27527_, new_n27528_, new_n27529_, new_n27530_,
    new_n27531_, new_n27532_, new_n27533_, new_n27534_, new_n27535_,
    new_n27536_, new_n27537_, new_n27538_, new_n27539_, new_n27540_,
    new_n27541_, new_n27542_, new_n27543_, new_n27544_, new_n27545_,
    new_n27546_, new_n27547_, new_n27548_, new_n27549_, new_n27550_,
    new_n27551_, new_n27552_, new_n27553_, new_n27554_, new_n27555_,
    new_n27556_, new_n27557_, new_n27558_, new_n27559_, new_n27560_,
    new_n27561_, new_n27562_, new_n27563_, new_n27564_, new_n27565_,
    new_n27566_, new_n27567_, new_n27568_, new_n27570_, new_n27571_,
    new_n27572_, new_n27573_, new_n27574_, new_n27575_, new_n27576_,
    new_n27577_, new_n27578_, new_n27579_, new_n27580_, new_n27581_,
    new_n27582_, new_n27583_, new_n27584_, new_n27585_, new_n27586_,
    new_n27587_, new_n27588_, new_n27589_, new_n27590_, new_n27591_,
    new_n27592_, new_n27593_, new_n27594_, new_n27595_, new_n27596_,
    new_n27597_, new_n27598_, new_n27599_, new_n27600_, new_n27601_,
    new_n27602_, new_n27603_, new_n27604_, new_n27605_, new_n27606_,
    new_n27607_, new_n27608_, new_n27609_, new_n27610_, new_n27611_,
    new_n27612_, new_n27613_, new_n27614_, new_n27615_, new_n27616_,
    new_n27617_, new_n27618_, new_n27619_, new_n27620_, new_n27621_,
    new_n27622_, new_n27623_, new_n27624_, new_n27625_, new_n27626_,
    new_n27627_, new_n27628_, new_n27629_, new_n27630_, new_n27631_,
    new_n27632_, new_n27633_, new_n27634_, new_n27635_, new_n27636_,
    new_n27637_, new_n27638_, new_n27639_, new_n27640_, new_n27641_,
    new_n27642_, new_n27643_, new_n27644_, new_n27645_, new_n27646_,
    new_n27647_, new_n27648_, new_n27649_, new_n27650_, new_n27651_,
    new_n27652_, new_n27653_, new_n27654_, new_n27655_, new_n27656_,
    new_n27657_, new_n27658_, new_n27659_, new_n27660_, new_n27661_,
    new_n27662_, new_n27663_, new_n27664_, new_n27665_, new_n27666_,
    new_n27667_, new_n27668_, new_n27669_, new_n27670_, new_n27671_,
    new_n27672_, new_n27673_, new_n27674_, new_n27675_, new_n27676_,
    new_n27677_, new_n27678_, new_n27679_, new_n27680_, new_n27681_,
    new_n27682_, new_n27683_, new_n27684_, new_n27685_, new_n27686_,
    new_n27688_, new_n27689_, new_n27690_, new_n27691_, new_n27693_,
    new_n27694_, new_n27695_, new_n27696_, new_n27697_, new_n27699_,
    new_n27700_, new_n27701_, new_n27702_, new_n27703_, new_n27704_,
    new_n27705_, new_n27706_, new_n27707_, new_n27708_, new_n27709_,
    new_n27710_, new_n27711_, new_n27712_, new_n27713_, new_n27714_,
    new_n27715_, new_n27716_, new_n27717_, new_n27718_, new_n27719_,
    new_n27720_, new_n27722_, new_n27723_, new_n27724_, new_n27725_,
    new_n27726_, new_n27727_, new_n27728_, new_n27729_, new_n27730_,
    new_n27731_, new_n27732_, new_n27733_, new_n27734_, new_n27735_,
    new_n27736_, new_n27737_, new_n27738_, new_n27739_, new_n27740_,
    new_n27741_, new_n27742_, new_n27743_, new_n27744_, new_n27745_,
    new_n27746_, new_n27747_, new_n27748_, new_n27749_, new_n27750_,
    new_n27751_, new_n27752_, new_n27753_, new_n27754_, new_n27755_,
    new_n27756_, new_n27757_, new_n27758_, new_n27759_, new_n27760_,
    new_n27761_, new_n27762_, new_n27763_, new_n27764_, new_n27765_,
    new_n27766_, new_n27767_, new_n27768_, new_n27769_, new_n27770_,
    new_n27771_, new_n27772_, new_n27773_, new_n27774_, new_n27775_,
    new_n27776_, new_n27777_, new_n27778_, new_n27779_, new_n27780_,
    new_n27781_, new_n27782_, new_n27783_, new_n27784_, new_n27785_,
    new_n27786_, new_n27787_, new_n27788_, new_n27789_, new_n27790_,
    new_n27791_, new_n27792_, new_n27793_, new_n27794_, new_n27795_,
    new_n27796_, new_n27797_, new_n27798_, new_n27799_, new_n27800_,
    new_n27801_, new_n27802_, new_n27803_, new_n27804_, new_n27805_,
    new_n27806_, new_n27807_, new_n27808_, new_n27809_, new_n27810_,
    new_n27811_, new_n27812_, new_n27813_, new_n27814_, new_n27815_,
    new_n27816_, new_n27817_, new_n27818_, new_n27819_, new_n27820_,
    new_n27821_, new_n27822_, new_n27823_, new_n27824_, new_n27825_,
    new_n27826_, new_n27827_, new_n27828_, new_n27829_, new_n27830_,
    new_n27831_, new_n27832_, new_n27833_, new_n27834_, new_n27835_,
    new_n27836_, new_n27837_, new_n27838_, new_n27839_, new_n27840_,
    new_n27841_, new_n27842_, new_n27843_, new_n27844_, new_n27845_,
    new_n27846_, new_n27847_, new_n27848_, new_n27849_, new_n27850_,
    new_n27851_, new_n27852_, new_n27853_, new_n27854_, new_n27855_,
    new_n27856_, new_n27857_, new_n27858_, new_n27859_, new_n27860_,
    new_n27861_, new_n27862_, new_n27863_, new_n27864_, new_n27865_,
    new_n27866_, new_n27867_, new_n27868_, new_n27869_, new_n27870_,
    new_n27871_, new_n27872_, new_n27873_, new_n27874_, new_n27875_,
    new_n27876_, new_n27877_, new_n27878_, new_n27879_, new_n27880_,
    new_n27881_, new_n27882_, new_n27883_, new_n27884_, new_n27885_,
    new_n27886_, new_n27887_, new_n27888_, new_n27889_, new_n27890_,
    new_n27891_, new_n27892_, new_n27893_, new_n27894_, new_n27895_,
    new_n27896_, new_n27897_, new_n27899_, new_n27900_, new_n27901_,
    new_n27902_, new_n27903_, new_n27904_, new_n27905_, new_n27906_,
    new_n27907_, new_n27908_, new_n27909_, new_n27910_, new_n27911_,
    new_n27912_, new_n27913_, new_n27914_, new_n27915_, new_n27916_,
    new_n27917_, new_n27918_, new_n27919_, new_n27920_, new_n27921_,
    new_n27922_, new_n27923_, new_n27924_, new_n27925_, new_n27926_,
    new_n27927_, new_n27928_, new_n27929_, new_n27930_, new_n27931_,
    new_n27932_, new_n27933_, new_n27934_, new_n27935_, new_n27936_,
    new_n27937_, new_n27938_, new_n27939_, new_n27940_, new_n27941_,
    new_n27942_, new_n27943_, new_n27944_, new_n27945_, new_n27946_,
    new_n27947_, new_n27948_, new_n27949_, new_n27950_, new_n27951_,
    new_n27952_, new_n27953_, new_n27954_, new_n27955_, new_n27956_,
    new_n27957_, new_n27958_, new_n27959_, new_n27960_, new_n27961_,
    new_n27962_, new_n27963_, new_n27964_, new_n27965_, new_n27966_,
    new_n27967_, new_n27968_, new_n27969_, new_n27970_, new_n27971_,
    new_n27972_, new_n27973_, new_n27974_, new_n27975_, new_n27976_,
    new_n27977_, new_n27978_, new_n27979_, new_n27980_, new_n27981_,
    new_n27982_, new_n27983_, new_n27984_, new_n27985_, new_n27986_,
    new_n27987_, new_n27988_, new_n27989_, new_n27990_, new_n27991_,
    new_n27992_, new_n27993_, new_n27994_, new_n27995_, new_n27996_,
    new_n27997_, new_n27998_, new_n27999_, new_n28000_, new_n28001_,
    new_n28002_, new_n28003_, new_n28004_, new_n28005_, new_n28006_,
    new_n28007_, new_n28008_, new_n28009_, new_n28010_, new_n28011_,
    new_n28012_, new_n28013_, new_n28014_, new_n28015_, new_n28016_,
    new_n28017_, new_n28018_, new_n28019_, new_n28020_, new_n28021_,
    new_n28022_, new_n28023_, new_n28024_, new_n28025_, new_n28026_,
    new_n28027_, new_n28028_, new_n28029_, new_n28030_, new_n28031_,
    new_n28032_, new_n28033_, new_n28034_, new_n28035_, new_n28036_,
    new_n28037_, new_n28038_, new_n28039_, new_n28040_, new_n28041_,
    new_n28043_, new_n28045_, new_n28047_, new_n28049_, new_n28051_,
    new_n28053_, new_n28054_, new_n28055_, new_n28057_, new_n28058_,
    new_n28059_, new_n28061_, new_n28062_, new_n28063_, new_n28064_,
    new_n28065_, new_n28066_, new_n28067_, new_n28068_, new_n28069_,
    new_n28070_, new_n28071_, new_n28072_, new_n28073_, new_n28074_,
    new_n28075_, new_n28076_, new_n28077_, new_n28078_, new_n28079_,
    new_n28080_, new_n28081_, new_n28082_, new_n28084_, new_n28085_,
    new_n28086_, new_n28087_, new_n28088_, new_n28089_, new_n28090_,
    new_n28091_, new_n28092_, new_n28093_, new_n28094_, new_n28095_,
    new_n28096_, new_n28097_, new_n28098_, new_n28099_, new_n28100_,
    new_n28101_, new_n28102_, new_n28103_, new_n28104_, new_n28105_,
    new_n28106_, new_n28107_, new_n28108_, new_n28109_, new_n28110_,
    new_n28111_, new_n28112_, new_n28113_, new_n28114_, new_n28115_,
    new_n28116_, new_n28117_, new_n28118_, new_n28119_, new_n28120_,
    new_n28121_, new_n28122_, new_n28123_, new_n28124_, new_n28125_,
    new_n28126_, new_n28127_, new_n28128_, new_n28129_, new_n28130_,
    new_n28131_, new_n28132_, new_n28133_, new_n28134_, new_n28135_,
    new_n28136_, new_n28137_, new_n28138_, new_n28139_, new_n28140_,
    new_n28141_, new_n28142_, new_n28143_, new_n28144_, new_n28145_,
    new_n28146_, new_n28147_, new_n28148_, new_n28149_, new_n28150_,
    new_n28151_, new_n28152_, new_n28153_, new_n28154_, new_n28155_,
    new_n28156_, new_n28157_, new_n28158_, new_n28159_, new_n28160_,
    new_n28161_, new_n28162_, new_n28163_, new_n28164_, new_n28165_,
    new_n28166_, new_n28167_, new_n28168_, new_n28169_, new_n28170_,
    new_n28171_, new_n28172_, new_n28173_, new_n28174_, new_n28175_,
    new_n28176_, new_n28177_, new_n28178_, new_n28179_, new_n28180_,
    new_n28181_, new_n28182_, new_n28183_, new_n28184_, new_n28185_,
    new_n28186_, new_n28187_, new_n28188_, new_n28189_, new_n28190_,
    new_n28191_, new_n28192_, new_n28193_, new_n28194_, new_n28195_,
    new_n28196_, new_n28197_, new_n28198_, new_n28199_, new_n28200_,
    new_n28201_, new_n28202_, new_n28203_, new_n28204_, new_n28205_,
    new_n28206_, new_n28207_, new_n28208_, new_n28209_, new_n28210_,
    new_n28211_, new_n28212_, new_n28213_, new_n28214_, new_n28215_,
    new_n28216_, new_n28217_, new_n28218_, new_n28219_, new_n28220_,
    new_n28221_, new_n28222_, new_n28223_, new_n28224_, new_n28225_,
    new_n28226_, new_n28227_, new_n28228_, new_n28229_, new_n28230_,
    new_n28231_, new_n28232_, new_n28233_, new_n28234_, new_n28235_,
    new_n28236_, new_n28237_, new_n28238_, new_n28239_, new_n28241_,
    new_n28242_, new_n28243_, new_n28244_, new_n28245_, new_n28246_,
    new_n28247_, new_n28248_, new_n28249_, new_n28250_, new_n28251_,
    new_n28252_, new_n28253_, new_n28254_, new_n28255_, new_n28256_,
    new_n28257_, new_n28258_, new_n28259_, new_n28260_, new_n28261_,
    new_n28262_, new_n28263_, new_n28264_, new_n28265_, new_n28266_,
    new_n28267_, new_n28268_, new_n28270_, new_n28271_, new_n28272_,
    new_n28273_, new_n28274_, new_n28275_, new_n28276_, new_n28277_,
    new_n28278_, new_n28279_, new_n28280_, new_n28281_, new_n28282_,
    new_n28283_, new_n28284_, new_n28285_, new_n28286_, new_n28287_,
    new_n28288_, new_n28289_, new_n28290_, new_n28291_, new_n28292_,
    new_n28293_, new_n28295_, new_n28296_, new_n28297_, new_n28298_,
    new_n28299_, new_n28300_, new_n28301_, new_n28302_, new_n28303_,
    new_n28304_, new_n28305_, new_n28306_, new_n28307_, new_n28308_,
    new_n28309_, new_n28310_, new_n28311_, new_n28312_, new_n28313_,
    new_n28314_, new_n28315_, new_n28316_, new_n28317_, new_n28318_,
    new_n28319_, new_n28320_, new_n28321_, new_n28322_, new_n28323_,
    new_n28324_, new_n28325_, new_n28326_, new_n28327_, new_n28328_,
    new_n28329_, new_n28330_, new_n28331_, new_n28332_, new_n28333_,
    new_n28334_, new_n28335_, new_n28336_, new_n28338_, new_n28339_,
    new_n28340_, new_n28341_, new_n28342_, new_n28343_, new_n28344_,
    new_n28345_, new_n28346_, new_n28347_, new_n28348_, new_n28349_,
    new_n28350_, new_n28351_, new_n28352_, new_n28353_, new_n28354_,
    new_n28355_, new_n28356_, new_n28357_, new_n28358_, new_n28359_,
    new_n28360_, new_n28361_, new_n28362_, new_n28363_, new_n28364_,
    new_n28365_, new_n28366_, new_n28367_, new_n28368_, new_n28369_,
    new_n28370_, new_n28371_, new_n28372_, new_n28373_, new_n28374_,
    new_n28375_, new_n28376_, new_n28377_, new_n28378_, new_n28379_,
    new_n28380_, new_n28381_, new_n28382_, new_n28383_, new_n28384_,
    new_n28385_, new_n28386_, new_n28387_, new_n28388_, new_n28389_,
    new_n28390_, new_n28391_, new_n28392_, new_n28393_, new_n28394_,
    new_n28395_, new_n28396_, new_n28397_, new_n28398_, new_n28399_,
    new_n28400_, new_n28401_, new_n28402_, new_n28403_, new_n28404_,
    new_n28405_, new_n28406_, new_n28407_, new_n28408_, new_n28409_,
    new_n28410_, new_n28411_, new_n28412_, new_n28413_, new_n28414_,
    new_n28415_, new_n28416_, new_n28417_, new_n28418_, new_n28419_,
    new_n28420_, new_n28421_, new_n28422_, new_n28423_, new_n28424_,
    new_n28425_, new_n28426_, new_n28427_, new_n28428_, new_n28429_,
    new_n28430_, new_n28431_, new_n28432_, new_n28433_, new_n28434_,
    new_n28435_, new_n28436_, new_n28437_, new_n28438_, new_n28439_,
    new_n28440_, new_n28441_, new_n28442_, new_n28443_, new_n28444_,
    new_n28445_, new_n28446_, new_n28447_, new_n28448_, new_n28449_,
    new_n28450_, new_n28451_, new_n28452_, new_n28453_, new_n28454_,
    new_n28455_, new_n28456_, new_n28457_, new_n28458_, new_n28459_,
    new_n28460_, new_n28461_, new_n28462_, new_n28463_, new_n28464_,
    new_n28465_, new_n28466_, new_n28467_, new_n28468_, new_n28469_,
    new_n28471_, new_n28472_, new_n28473_, new_n28474_, new_n28475_,
    new_n28476_, new_n28477_, new_n28478_, new_n28479_, new_n28480_,
    new_n28481_, new_n28482_, new_n28483_, new_n28484_, new_n28485_,
    new_n28486_, new_n28487_, new_n28488_, new_n28489_, new_n28490_,
    new_n28491_, new_n28492_, new_n28493_, new_n28494_, new_n28495_,
    new_n28496_, new_n28497_, new_n28498_, new_n28499_, new_n28500_,
    new_n28501_, new_n28502_, new_n28503_, new_n28504_, new_n28505_,
    new_n28506_, new_n28507_, new_n28508_, new_n28509_, new_n28510_,
    new_n28511_, new_n28512_, new_n28513_, new_n28514_, new_n28515_,
    new_n28516_, new_n28517_, new_n28518_, new_n28519_, new_n28520_,
    new_n28521_, new_n28522_, new_n28523_, new_n28524_, new_n28525_,
    new_n28526_, new_n28527_, new_n28528_, new_n28529_, new_n28530_,
    new_n28531_, new_n28532_, new_n28533_, new_n28534_, new_n28535_,
    new_n28536_, new_n28537_, new_n28538_, new_n28539_, new_n28540_,
    new_n28541_, new_n28542_, new_n28543_, new_n28544_, new_n28545_,
    new_n28546_, new_n28547_, new_n28548_, new_n28549_, new_n28550_,
    new_n28551_, new_n28552_, new_n28553_, new_n28554_, new_n28555_,
    new_n28556_, new_n28557_, new_n28558_, new_n28559_, new_n28560_,
    new_n28561_, new_n28562_, new_n28563_, new_n28564_, new_n28565_,
    new_n28566_, new_n28567_, new_n28568_, new_n28569_, new_n28570_,
    new_n28571_, new_n28572_, new_n28573_, new_n28574_, new_n28575_,
    new_n28576_, new_n28577_, new_n28578_, new_n28580_, new_n28581_,
    new_n28582_, new_n28583_, new_n28584_, new_n28585_, new_n28586_,
    new_n28587_, new_n28588_, new_n28589_, new_n28590_, new_n28591_,
    new_n28592_, new_n28593_, new_n28594_, new_n28595_, new_n28596_,
    new_n28597_, new_n28598_, new_n28599_, new_n28600_, new_n28601_,
    new_n28602_, new_n28603_, new_n28605_, new_n28606_, new_n28607_,
    new_n28608_, new_n28609_, new_n28610_, new_n28611_, new_n28612_,
    new_n28613_, new_n28614_, new_n28615_, new_n28616_, new_n28617_,
    new_n28618_, new_n28619_, new_n28620_, new_n28621_, new_n28622_,
    new_n28623_, new_n28624_, new_n28625_, new_n28626_, new_n28627_,
    new_n28628_, new_n28629_, new_n28631_, new_n28632_, new_n28633_,
    new_n28634_, new_n28635_, new_n28636_, new_n28637_, new_n28638_,
    new_n28639_, new_n28640_, new_n28641_, new_n28642_, new_n28643_,
    new_n28644_, new_n28645_, new_n28646_, new_n28647_, new_n28648_,
    new_n28649_, new_n28650_, new_n28651_, new_n28652_, new_n28653_,
    new_n28654_, new_n28655_, new_n28656_, new_n28657_, new_n28659_,
    new_n28660_, new_n28661_, new_n28662_, new_n28663_, new_n28664_,
    new_n28665_, new_n28666_, new_n28667_, new_n28668_, new_n28669_,
    new_n28670_, new_n28671_, new_n28672_, new_n28673_, new_n28674_,
    new_n28675_, new_n28676_, new_n28677_, new_n28678_, new_n28679_,
    new_n28680_, new_n28681_, new_n28682_, new_n28683_, new_n28684_,
    new_n28685_, new_n28686_, new_n28687_, new_n28688_, new_n28689_,
    new_n28690_, new_n28691_, new_n28692_, new_n28693_, new_n28694_,
    new_n28695_, new_n28696_, new_n28697_, new_n28698_, new_n28699_,
    new_n28700_, new_n28701_, new_n28702_, new_n28703_, new_n28704_,
    new_n28705_, new_n28706_, new_n28707_, new_n28708_, new_n28709_,
    new_n28710_, new_n28711_, new_n28712_, new_n28713_, new_n28714_,
    new_n28715_, new_n28716_, new_n28717_, new_n28719_, new_n28720_,
    new_n28721_, new_n28722_, new_n28723_, new_n28724_, new_n28725_,
    new_n28726_, new_n28727_, new_n28728_, new_n28729_, new_n28730_,
    new_n28731_, new_n28732_, new_n28733_, new_n28734_, new_n28735_,
    new_n28736_, new_n28737_, new_n28738_, new_n28739_, new_n28740_,
    new_n28741_, new_n28742_, new_n28743_, new_n28744_, new_n28745_,
    new_n28746_, new_n28747_, new_n28748_, new_n28749_, new_n28750_,
    new_n28751_, new_n28752_, new_n28753_, new_n28754_, new_n28755_,
    new_n28756_, new_n28757_, new_n28759_, new_n28760_, new_n28761_,
    new_n28762_, new_n28763_, new_n28764_, new_n28765_, new_n28766_,
    new_n28767_, new_n28768_, new_n28769_, new_n28770_, new_n28771_,
    new_n28772_, new_n28773_, new_n28774_, new_n28775_, new_n28776_,
    new_n28777_, new_n28778_, new_n28779_, new_n28780_, new_n28781_,
    new_n28782_, new_n28783_, new_n28784_, new_n28785_, new_n28787_,
    new_n28788_, new_n28789_, new_n28790_, new_n28791_, new_n28792_,
    new_n28793_, new_n28794_, new_n28795_, new_n28796_, new_n28797_,
    new_n28798_, new_n28799_, new_n28800_, new_n28801_, new_n28802_,
    new_n28803_, new_n28804_, new_n28805_, new_n28806_, new_n28807_,
    new_n28808_, new_n28809_, new_n28810_, new_n28811_, new_n28812_,
    new_n28813_, new_n28814_, new_n28815_, new_n28816_, new_n28817_,
    new_n28818_, new_n28819_, new_n28820_, new_n28821_, new_n28822_,
    new_n28823_, new_n28824_, new_n28825_, new_n28826_, new_n28827_,
    new_n28828_, new_n28829_, new_n28830_, new_n28831_, new_n28833_,
    new_n28834_, new_n28835_, new_n28836_, new_n28837_, new_n28838_,
    new_n28839_, new_n28840_, new_n28841_, new_n28842_, new_n28843_,
    new_n28844_, new_n28845_, new_n28846_, new_n28848_, new_n28849_,
    new_n28850_, new_n28851_, new_n28852_, new_n28853_, new_n28854_,
    new_n28855_, new_n28856_, new_n28857_, new_n28858_, new_n28859_,
    new_n28860_, new_n28861_, new_n28862_, new_n28863_, new_n28864_,
    new_n28865_, new_n28866_, new_n28867_, new_n28868_, new_n28869_,
    new_n28870_, new_n28873_, new_n28874_, new_n28875_, new_n28876_,
    new_n28877_, new_n28878_, new_n28879_, new_n28880_, new_n28881_,
    new_n28882_, new_n28883_, new_n28884_, new_n28885_, new_n28886_,
    new_n28887_, new_n28888_, new_n28889_, new_n28890_, new_n28891_,
    new_n28892_, new_n28893_, new_n28894_, new_n28895_, new_n28896_,
    new_n28897_, new_n28898_, new_n28899_, new_n28900_, new_n28901_,
    new_n28902_, new_n28903_, new_n28904_, new_n28905_, new_n28906_,
    new_n28907_, new_n28908_, new_n28909_, new_n28910_, new_n28911_,
    new_n28912_, new_n28913_, new_n28915_, new_n28916_, new_n28917_,
    new_n28918_, new_n28919_, new_n28920_, new_n28921_, new_n28922_,
    new_n28923_, new_n28924_, new_n28925_, new_n28926_, new_n28927_,
    new_n28928_, new_n28929_, new_n28930_, new_n28931_, new_n28932_,
    new_n28933_, new_n28934_, new_n28935_, new_n28936_, new_n28937_,
    new_n28938_, new_n28939_, new_n28940_, new_n28941_, new_n28942_,
    new_n28943_, new_n28944_, new_n28946_, new_n28947_, new_n28948_,
    new_n28949_, new_n28950_, new_n28951_, new_n28952_, new_n28953_,
    new_n28954_, new_n28955_, new_n28956_, new_n28957_, new_n28958_,
    new_n28959_, new_n28960_, new_n28961_, new_n28962_, new_n28963_,
    new_n28964_, new_n28965_, new_n28966_, new_n28967_, new_n28968_,
    new_n28969_, new_n28970_, new_n28972_, new_n28973_, new_n28974_,
    new_n28975_, new_n28976_, new_n28977_, new_n28978_, new_n28979_,
    new_n28980_, new_n28981_, new_n28982_, new_n28983_, new_n28984_,
    new_n28985_, new_n28986_, new_n28987_, new_n28988_, new_n28989_,
    new_n28990_, new_n28992_, new_n28993_, new_n28994_, new_n28995_,
    new_n28996_, new_n28997_, new_n28998_, new_n28999_, new_n29000_,
    new_n29001_, new_n29002_, new_n29003_, new_n29004_, new_n29005_,
    new_n29006_, new_n29007_, new_n29008_, new_n29009_, new_n29010_,
    new_n29012_, new_n29013_, new_n29014_, new_n29015_, new_n29016_,
    new_n29017_, new_n29018_, new_n29019_, new_n29020_, new_n29021_,
    new_n29022_, new_n29023_, new_n29024_, new_n29025_, new_n29026_,
    new_n29027_, new_n29028_, new_n29029_, new_n29030_, new_n29031_,
    new_n29032_, new_n29033_, new_n29034_, new_n29035_, new_n29036_,
    new_n29037_, new_n29038_, new_n29039_, new_n29040_, new_n29041_,
    new_n29042_, new_n29043_, new_n29044_, new_n29045_, new_n29047_,
    new_n29049_, new_n29050_, new_n29051_, new_n29052_, new_n29053_,
    new_n29054_, new_n29055_, new_n29056_, new_n29057_, new_n29058_,
    new_n29059_, new_n29060_, new_n29061_, new_n29062_, new_n29063_,
    new_n29065_, new_n29066_, new_n29067_, new_n29068_, new_n29069_,
    new_n29070_, new_n29071_, new_n29072_, new_n29073_, new_n29074_,
    new_n29075_, new_n29076_, new_n29077_, new_n29078_, new_n29081_,
    new_n29083_, new_n29085_, new_n29086_, new_n29087_, new_n29088_,
    new_n29089_, new_n29090_, new_n29091_, new_n29092_, new_n29093_,
    new_n29094_, new_n29105_, new_n29106_, new_n29107_, new_n29108_,
    new_n29110_, new_n29111_, new_n29112_, new_n29113_, new_n29114_,
    new_n29116_, new_n29117_, new_n29118_, new_n29119_, new_n29121_,
    new_n29122_, new_n29123_, new_n29124_, new_n29125_, new_n29126_,
    new_n29127_, new_n29128_, new_n29129_, new_n29130_, new_n29131_,
    new_n29132_, new_n29133_, new_n29134_, new_n29135_, new_n29144_,
    new_n29145_, new_n29146_, new_n29147_, new_n29148_, new_n29149_,
    new_n29150_, new_n29151_, new_n29152_, new_n29153_, new_n29154_,
    new_n29155_, new_n29156_, new_n29157_, new_n29158_, new_n29160_,
    new_n29162_, new_n29164_, new_n29165_, new_n29166_, new_n29167_,
    new_n29169_, new_n29170_, new_n29171_, new_n29172_, new_n29173_,
    new_n29174_, new_n29175_, new_n29177_, new_n29180_, new_n29182_,
    new_n29195_, new_n29196_, new_n29197_, new_n29198_, new_n29199_,
    new_n29201_, new_n29203_, new_n29204_, new_n29205_, new_n29206_,
    new_n29207_, new_n29208_, new_n29217_, new_n29218_, new_n29219_,
    new_n29221_, new_n29295_, new_n29339_, new_n29340_, new_n29341_,
    new_n29342_, new_n29343_, new_n29344_, new_n29345_, new_n29346_,
    new_n29347_, new_n29348_, new_n29349_, new_n29350_, new_n29351_,
    new_n29352_, new_n29353_, new_n29354_, new_n29355_, new_n29356_,
    new_n29357_, new_n29358_, new_n29359_, new_n29360_, new_n29369_,
    new_n29370_, new_n29371_, new_n29372_, new_n29373_, new_n29374_,
    new_n29375_, new_n29376_, new_n29377_, new_n29378_, new_n29379_,
    new_n29380_, new_n29381_, new_n29383_, new_n29384_, new_n29385_,
    new_n29386_, new_n29387_, new_n29388_, new_n29389_, new_n29390_,
    new_n29391_, new_n29392_, new_n29393_, new_n29395_, new_n29396_,
    new_n29397_, new_n29398_, new_n29399_, new_n29400_, new_n29401_,
    new_n29402_, new_n29403_, new_n29404_, new_n29405_, new_n29406_,
    new_n29407_, new_n29408_, new_n29409_, new_n29410_, new_n29412_,
    new_n29414_, new_n29415_, new_n29416_, new_n29417_, new_n29418_,
    new_n29419_, new_n29420_, new_n29421_, new_n29422_, new_n29423_,
    new_n29425_, new_n29426_, new_n29427_, new_n29428_, new_n29429_,
    new_n29430_, new_n29431_, new_n29432_, new_n29433_, new_n29434_,
    new_n29436_, new_n29437_, new_n29438_, new_n29439_, new_n29440_,
    new_n29441_, new_n29442_, new_n29443_, new_n29444_, new_n29445_,
    new_n29447_, new_n29448_, new_n29449_, new_n29450_, new_n29451_,
    new_n29452_, new_n29453_, new_n29454_, new_n29455_, new_n29456_,
    new_n29458_, new_n29459_, new_n29460_, new_n29461_, new_n29462_,
    new_n29463_, new_n29465_, new_n29466_, new_n29467_, new_n29468_,
    new_n29469_, new_n29470_, new_n29472_, new_n29473_, new_n29474_,
    new_n29475_, new_n29476_, new_n29477_, new_n29479_, new_n29480_,
    new_n29481_, new_n29482_, new_n29483_, new_n29484_, new_n29495_,
    new_n29502_, new_n29506_, new_n29515_, new_n29516_, new_n29517_,
    new_n29518_, new_n29519_, new_n29520_, new_n29527_, new_n29528_,
    new_n29529_, new_n29537_, new_n29538_, new_n29539_, new_n29540_,
    new_n29542_, new_n29547_, new_n29548_, new_n29549_, new_n29551_,
    new_n29562_, new_n29573_, new_n29574_, new_n29575_, new_n29582_,
    new_n29590_, new_n29591_, new_n29592_, new_n29603_, new_n29604_,
    new_n29605_, new_n29606_, new_n29607_, new_n29608_, new_n29609_,
    new_n29610_, new_n29611_, new_n29612_, new_n29613_, new_n29614_,
    new_n29615_, new_n29616_, new_n29617_, new_n29618_, new_n29619_,
    new_n29620_, new_n29621_, new_n29622_, new_n29623_, new_n29624_,
    new_n29625_, new_n29626_, new_n29627_, new_n29628_, new_n29629_,
    new_n29630_, new_n29631_, new_n29632_, new_n29633_, new_n29634_,
    new_n29635_, new_n29636_, new_n29637_, new_n29638_, new_n29639_,
    new_n29640_, new_n29641_, new_n29642_, new_n29643_, new_n29644_,
    new_n29645_, new_n29646_, new_n29647_, new_n29648_, new_n29649_,
    new_n29650_, new_n29651_, new_n29652_, new_n29653_, new_n29654_,
    new_n29655_, new_n29656_, new_n29657_, new_n29658_, new_n29659_,
    new_n29660_, new_n29661_, new_n29662_, new_n29663_, new_n29666_,
    new_n29668_, new_n29669_, new_n29670_, new_n29687_, new_n29688_,
    new_n29690_, new_n29691_, new_n29693_, new_n29694_, new_n29695_,
    new_n29696_, new_n29697_, new_n29698_, new_n29699_, new_n29700_,
    new_n29701_, new_n29702_, new_n29703_, new_n29704_, new_n29706_,
    new_n29707_, new_n29709_, new_n29711_, new_n29713_, new_n29714_,
    new_n29715_, new_n29716_, new_n29717_, new_n29718_, new_n29719_,
    new_n29720_, new_n29721_, new_n29722_, new_n29723_, new_n29724_,
    new_n29725_, new_n29726_, new_n29727_, new_n29728_, new_n29729_,
    new_n29730_, new_n29731_, new_n29732_, new_n29733_, new_n29734_,
    new_n29735_, new_n29736_, new_n29737_, new_n29738_, new_n29739_,
    new_n29740_, new_n29741_, new_n29742_, new_n29743_, new_n29744_,
    new_n29745_, new_n29746_, new_n29747_, new_n29748_, new_n29749_,
    new_n29750_, new_n29751_, new_n29752_, new_n29753_, new_n29754_,
    new_n29755_, new_n29756_, new_n29757_, new_n29758_, new_n29759_,
    new_n29760_, new_n29761_, new_n29762_, new_n29763_, new_n29764_,
    new_n29765_, new_n29766_, new_n29767_, new_n29768_, new_n29769_,
    new_n29770_, new_n29771_, new_n29772_, new_n29773_, new_n29774_,
    new_n29775_, new_n29776_, new_n29777_, new_n29778_, new_n29779_,
    new_n29780_, new_n29781_, new_n29782_, new_n29783_, new_n29784_,
    new_n29785_, new_n29786_, new_n29787_, new_n29788_, new_n29789_,
    new_n29790_, new_n29791_, new_n29792_, new_n29793_, new_n29794_,
    new_n29795_, new_n29796_, new_n29797_, new_n29798_, new_n29799_,
    new_n29800_, new_n29801_, new_n29802_, new_n29803_, new_n29804_,
    new_n29805_, new_n29806_, new_n29807_, new_n29808_, new_n29809_,
    new_n29810_, new_n29811_, new_n29812_, new_n29813_, new_n29814_,
    new_n29815_, new_n29816_, new_n29817_, new_n29818_, new_n29819_,
    new_n29820_, new_n29821_, new_n29822_, new_n29823_, new_n29824_,
    new_n29825_, new_n29826_, new_n29827_, new_n29828_, new_n29829_,
    new_n29830_, new_n29831_, new_n29832_, new_n29833_, new_n29834_,
    new_n29835_, new_n29836_, new_n29837_, new_n29838_, new_n29839_,
    new_n29840_, new_n29841_, new_n29842_, new_n29843_, new_n29844_,
    new_n29845_, new_n29846_, new_n29847_, new_n29848_, new_n29849_,
    new_n29850_, new_n29851_, new_n29852_, new_n29853_, new_n29854_,
    new_n29855_, new_n29856_, new_n29857_, new_n29858_, new_n29859_,
    new_n29860_, new_n29861_, new_n29862_, new_n29863_, new_n29864_,
    new_n29865_, new_n29866_, new_n29867_, new_n29868_, new_n29869_,
    new_n29870_, new_n29871_, new_n29872_, new_n29873_, new_n29874_,
    new_n29875_, new_n29876_, new_n29877_, new_n29878_, new_n29879_,
    new_n29880_, new_n29881_, new_n29882_, new_n29883_, new_n29884_,
    new_n29885_, new_n29886_, new_n29887_, new_n29888_, new_n29889_,
    new_n29890_, new_n29891_, new_n29892_, new_n29893_, new_n29894_,
    new_n29895_, new_n29896_, new_n29897_, new_n29898_, new_n29899_,
    new_n29900_, new_n29901_, new_n29902_, new_n29903_, new_n29904_,
    new_n29905_, new_n29906_, new_n29907_, new_n29908_, new_n29909_,
    new_n29910_, new_n29911_, new_n29912_, new_n29913_, new_n29914_,
    new_n29915_, new_n29916_, new_n29917_, new_n29918_, new_n29919_,
    new_n29920_, new_n29921_, new_n29922_, new_n29923_, new_n29924_,
    new_n29925_, new_n29926_, new_n29927_, new_n29928_, new_n29929_,
    new_n29930_, new_n29931_, new_n29932_, new_n29933_, new_n29934_,
    new_n29935_, new_n29936_, new_n29937_, new_n29938_, new_n29939_,
    new_n29940_, new_n29941_, new_n29942_, new_n29943_, new_n29944_,
    new_n29945_, new_n29946_, new_n29947_, new_n29948_, new_n29949_,
    new_n29950_, new_n29951_, new_n29952_, new_n29953_, new_n29954_,
    new_n29955_, new_n29956_, new_n29957_, new_n29958_, new_n29959_,
    new_n29960_, new_n29961_, new_n29962_, new_n29963_, new_n29964_,
    new_n29965_, new_n29966_, new_n29967_, new_n29968_, new_n29969_,
    new_n29970_, new_n29971_, new_n29972_, new_n29973_, new_n29974_,
    new_n29975_, new_n29976_, new_n29977_, new_n29978_, new_n29979_,
    new_n29980_, new_n29981_, new_n29982_, new_n29983_, new_n29984_,
    new_n29985_, new_n29986_, new_n29987_, new_n29988_, new_n29989_,
    new_n29990_, new_n29991_, new_n29992_, new_n29993_, new_n29994_,
    new_n29995_, new_n29996_, new_n29997_, new_n29998_, new_n29999_,
    new_n30000_, new_n30001_, new_n30002_, new_n30003_, new_n30004_,
    new_n30005_, new_n30006_, new_n30007_, new_n30008_, new_n30009_,
    new_n30010_, new_n30011_, new_n30012_, new_n30013_, new_n30014_,
    new_n30015_, new_n30016_, new_n30017_, new_n30018_, new_n30019_,
    new_n30020_, new_n30021_, new_n30022_, new_n30023_, new_n30024_,
    new_n30025_, new_n30026_, new_n30027_, new_n30028_, new_n30029_,
    new_n30030_, new_n30031_, new_n30032_, new_n30033_, new_n30034_,
    new_n30035_, new_n30036_, new_n30037_, new_n30038_, new_n30039_,
    new_n30040_, new_n30041_, new_n30042_, new_n30043_, new_n30044_,
    new_n30045_, new_n30046_, new_n30047_, new_n30048_, new_n30049_,
    new_n30050_, new_n30051_, new_n30052_, new_n30053_, new_n30054_,
    new_n30055_, new_n30056_, new_n30057_, new_n30058_, new_n30059_,
    new_n30060_, new_n30061_, new_n30062_, new_n30063_, new_n30064_,
    new_n30065_, new_n30066_, new_n30067_, new_n30068_, new_n30069_,
    new_n30070_, new_n30071_, new_n30072_, new_n30073_, new_n30074_,
    new_n30075_, new_n30076_, new_n30077_, new_n30078_, new_n30079_,
    new_n30080_, new_n30081_, new_n30082_, new_n30083_, new_n30084_,
    new_n30085_, new_n30086_, new_n30087_, new_n30088_, new_n30089_,
    new_n30090_, new_n30091_, new_n30092_, new_n30093_, new_n30094_,
    new_n30095_, new_n30096_, new_n30097_, new_n30098_, new_n30099_,
    new_n30100_, new_n30101_, new_n30102_, new_n30103_, new_n30104_,
    new_n30105_, new_n30106_, new_n30107_, new_n30108_, new_n30109_,
    new_n30110_, new_n30111_, new_n30112_, new_n30113_, new_n30114_,
    new_n30115_, new_n30116_, new_n30117_, new_n30118_, new_n30119_,
    new_n30120_, new_n30121_, new_n30122_, new_n30123_, new_n30124_,
    new_n30125_, new_n30126_, new_n30127_, new_n30128_, new_n30129_,
    new_n30130_, new_n30131_, new_n30132_, new_n30133_, new_n30134_,
    new_n30135_, new_n30136_, new_n30137_, new_n30138_, new_n30139_,
    new_n30140_, new_n30141_, new_n30142_, new_n30143_, new_n30144_,
    new_n30145_, new_n30146_, new_n30147_, new_n30148_, new_n30149_,
    new_n30150_, new_n30151_, new_n30152_, new_n30153_, new_n30154_,
    new_n30155_, new_n30156_, new_n30157_, new_n30158_, new_n30159_,
    new_n30160_, new_n30161_, new_n30162_, new_n30163_, new_n30164_,
    new_n30165_, new_n30166_, new_n30167_, new_n30168_, new_n30169_,
    new_n30170_, new_n30171_, new_n30172_, new_n30173_, new_n30174_,
    new_n30175_, new_n30176_, new_n30177_, new_n30178_, new_n30179_,
    new_n30180_, new_n30181_, new_n30182_, new_n30183_, new_n30184_,
    new_n30185_, new_n30186_, new_n30187_, new_n30188_, new_n30189_,
    new_n30190_, new_n30191_, new_n30192_, new_n30193_, new_n30194_,
    new_n30195_, new_n30196_, new_n30197_, new_n30198_, new_n30199_,
    new_n30200_, new_n30201_, new_n30202_, new_n30203_, new_n30204_,
    new_n30205_, new_n30206_, new_n30207_, new_n30208_, new_n30209_,
    new_n30210_, new_n30211_, new_n30212_, new_n30213_, new_n30214_,
    new_n30215_, new_n30216_, new_n30217_, new_n30218_, new_n30219_,
    new_n30220_, new_n30221_, new_n30222_, new_n30223_, new_n30224_,
    new_n30225_, new_n30226_, new_n30227_, new_n30228_, new_n30229_,
    new_n30230_, new_n30231_, new_n30232_, new_n30233_, new_n30234_,
    new_n30235_, new_n30236_, new_n30237_, new_n30238_, new_n30239_,
    new_n30241_, new_n30242_, new_n30243_, new_n30245_, new_n30246_,
    new_n30247_, new_n30248_, new_n30249_, new_n30250_, new_n30252_,
    new_n30253_, new_n30254_, new_n30256_, new_n30257_, new_n30259_,
    new_n30260_, new_n30261_, new_n30263_, new_n30264_, new_n30266_,
    new_n30267_, new_n30269_, new_n30270_, new_n30272_, new_n30273_,
    new_n30274_, new_n30275_, new_n30277_, new_n30278_, new_n30279_,
    new_n30280_, new_n30282_, new_n30283_, new_n30284_, new_n30285_,
    new_n30286_, new_n30288_, new_n30289_, new_n30290_, new_n30292_,
    new_n30294_, new_n30296_, new_n30297_, new_n30299_, new_n30301_,
    new_n30303_, new_n30304_, new_n30306_, new_n30307_, new_n30309_,
    new_n30311_, new_n30312_, new_n30314_, new_n30315_, new_n30316_,
    new_n30318_, new_n30319_, new_n30321_, new_n30322_, new_n30323_,
    new_n30325_, new_n30327_, new_n30329_, new_n30331_, new_n30332_,
    new_n30334_, new_n30336_, new_n30338_, new_n30340_, new_n30341_,
    new_n30342_, new_n30344_, new_n30345_, new_n30347_, new_n30348_,
    new_n30349_, new_n30351_, new_n30353_, new_n30355_, new_n30357_,
    new_n30359_, new_n30361_, new_n30362_, new_n30363_, new_n30365_,
    new_n30366_, new_n30367_, new_n30369_, new_n30371_, new_n30373_,
    new_n30374_, new_n30375_, new_n30377_, new_n30378_, new_n30380_,
    new_n30382_, new_n30384_, new_n30386_, new_n30387_, new_n30389_,
    new_n30391_, new_n30393_, new_n30395_, new_n30397_, new_n30398_,
    new_n30400_, new_n30401_, new_n30402_, new_n30404_, new_n30406_,
    new_n30408_, new_n30409_, new_n30410_, new_n30412_, new_n30413_,
    new_n30414_, new_n30416_, new_n30417_, new_n30419_, new_n30420_,
    new_n30422_, new_n30423_, new_n30425_, new_n30426_, new_n30427_,
    new_n30429_, new_n30430_, new_n30431_, new_n30433_, new_n30434_,
    new_n30436_, new_n30437_, new_n30438_, new_n30440_, new_n30441_,
    new_n30443_, new_n30444_, new_n30445_, new_n30446_, new_n30447_,
    new_n30448_, new_n30449_, new_n30450_, new_n30451_, new_n30452_,
    new_n30453_, new_n30455_, new_n30457_, new_n30459_, new_n30461_,
    new_n30462_, new_n30463_, new_n30464_, new_n30465_, new_n30466_,
    new_n30467_, new_n30468_, new_n30469_, new_n30470_, new_n30471_,
    new_n30472_, new_n30473_, new_n30474_, new_n30475_, new_n30476_,
    new_n30477_, new_n30478_, new_n30479_, new_n30480_, new_n30481_,
    new_n30482_, new_n30483_, new_n30484_, new_n30485_, new_n30486_,
    new_n30487_, new_n30488_, new_n30489_, new_n30490_, new_n30492_,
    new_n30493_, new_n30494_, new_n30495_, new_n30496_, new_n30497_,
    new_n30498_, new_n30499_, new_n30500_, new_n30501_, new_n30502_,
    new_n30503_, new_n30504_, new_n30505_, new_n30506_, new_n30507_,
    new_n30508_, new_n30509_, new_n30510_, new_n30511_, new_n30512_,
    new_n30513_, new_n30514_, new_n30515_, new_n30516_, new_n30517_,
    new_n30519_, new_n30521_, new_n30522_, new_n30523_, new_n30524_,
    new_n30525_, new_n30526_, new_n30527_, new_n30528_, new_n30529_,
    new_n30530_, new_n30531_, new_n30532_, new_n30533_, new_n30534_,
    new_n30535_, new_n30536_, new_n30537_, new_n30539_, new_n30540_,
    new_n30541_, new_n30542_, new_n30543_, new_n30544_, new_n30545_,
    new_n30546_, new_n30547_, new_n30548_, new_n30549_, new_n30550_,
    new_n30551_, new_n30552_, new_n30553_, new_n30554_, new_n30555_,
    new_n30556_, new_n30558_, new_n30559_, new_n30560_, new_n30561_,
    new_n30562_, new_n30563_, new_n30564_, new_n30565_, new_n30566_,
    new_n30567_, new_n30568_, new_n30569_, new_n30570_, new_n30571_,
    new_n30572_, new_n30573_, new_n30574_, new_n30575_, new_n30576_,
    new_n30578_, new_n30579_, new_n30580_, new_n30582_, new_n30583_,
    new_n30584_, new_n30585_, new_n30586_, new_n30587_, new_n30588_,
    new_n30589_, new_n30590_, new_n30591_, new_n30592_, new_n30593_,
    new_n30594_, new_n30595_, new_n30596_, new_n30597_, new_n30598_,
    new_n30599_, new_n30601_, new_n30602_, new_n30603_, new_n30604_,
    new_n30605_, new_n30606_, new_n30607_, new_n30608_, new_n30609_,
    new_n30610_, new_n30611_, new_n30612_, new_n30613_, new_n30614_,
    new_n30615_, new_n30616_, new_n30617_, new_n30619_, new_n30620_,
    new_n30621_, new_n30622_, new_n30623_, new_n30624_, new_n30625_,
    new_n30626_, new_n30627_, new_n30628_, new_n30629_, new_n30630_,
    new_n30631_, new_n30632_, new_n30633_, new_n30634_, new_n30635_,
    new_n30636_, new_n30637_, new_n30639_, new_n30640_, new_n30641_,
    new_n30642_, new_n30643_, new_n30644_, new_n30645_, new_n30646_,
    new_n30647_, new_n30648_, new_n30649_, new_n30650_, new_n30651_,
    new_n30652_, new_n30653_, new_n30654_, new_n30655_, new_n30657_,
    new_n30658_, new_n30659_, new_n30660_, new_n30661_, new_n30662_,
    new_n30663_, new_n30664_, new_n30665_, new_n30666_, new_n30667_,
    new_n30668_, new_n30669_, new_n30670_, new_n30671_, new_n30672_,
    new_n30673_, new_n30674_, new_n30675_, new_n30676_, new_n30678_,
    new_n30679_, new_n30680_, new_n30681_, new_n30682_, new_n30683_,
    new_n30684_, new_n30685_, new_n30686_, new_n30687_, new_n30688_,
    new_n30689_, new_n30690_, new_n30691_, new_n30692_, new_n30693_,
    new_n30694_, new_n30695_, new_n30696_, new_n30697_, new_n30699_,
    new_n30700_, new_n30701_, new_n30702_, new_n30703_, new_n30704_,
    new_n30705_, new_n30706_, new_n30707_, new_n30708_, new_n30709_,
    new_n30710_, new_n30711_, new_n30712_, new_n30713_, new_n30714_,
    new_n30715_, new_n30716_, new_n30718_, new_n30719_, new_n30720_,
    new_n30721_, new_n30722_, new_n30723_, new_n30724_, new_n30725_,
    new_n30726_, new_n30727_, new_n30728_, new_n30729_, new_n30730_,
    new_n30731_, new_n30732_, new_n30733_, new_n30734_, new_n30736_,
    new_n30737_, new_n30738_, new_n30739_, new_n30740_, new_n30741_,
    new_n30742_, new_n30743_, new_n30744_, new_n30745_, new_n30746_,
    new_n30747_, new_n30748_, new_n30749_, new_n30750_, new_n30751_,
    new_n30752_, new_n30754_, new_n30755_, new_n30756_, new_n30757_,
    new_n30758_, new_n30759_, new_n30760_, new_n30761_, new_n30762_,
    new_n30763_, new_n30764_, new_n30765_, new_n30766_, new_n30767_,
    new_n30768_, new_n30769_, new_n30770_, new_n30771_, new_n30772_,
    new_n30774_, new_n30776_, new_n30778_, new_n30779_, new_n30780_,
    new_n30781_, new_n30782_, new_n30783_, new_n30784_, new_n30785_,
    new_n30786_, new_n30787_, new_n30788_, new_n30789_, new_n30790_,
    new_n30791_, new_n30792_, new_n30793_, new_n30794_, new_n30796_,
    new_n30798_, new_n30799_, new_n30801_, new_n30802_, new_n30803_,
    new_n30804_, new_n30805_, new_n30806_, new_n30807_, new_n30808_,
    new_n30809_, new_n30810_, new_n30811_, new_n30812_, new_n30813_,
    new_n30814_, new_n30815_, new_n30816_, new_n30817_, new_n30818_,
    new_n30819_, new_n30820_, new_n30822_, new_n30824_, new_n30825_,
    new_n30827_, new_n30829_, new_n30830_, new_n30831_, new_n30832_,
    new_n30833_, new_n30834_, new_n30835_, new_n30836_, new_n30837_,
    new_n30838_, new_n30839_, new_n30840_, new_n30841_, new_n30842_,
    new_n30843_, new_n30845_, new_n30847_, new_n30849_, new_n30850_,
    new_n30851_, new_n30852_, new_n30853_, new_n30854_, new_n30855_,
    new_n30856_, new_n30857_, new_n30858_, new_n30859_, new_n30860_,
    new_n30861_, new_n30862_, new_n30863_, new_n30864_, new_n30865_,
    new_n30866_, new_n30867_, new_n30868_, new_n30869_, new_n30871_,
    new_n30872_, new_n30873_, new_n30875_, new_n30876_, new_n30877_,
    new_n30879_, new_n30880_, new_n30882_, new_n30884_, new_n30885_,
    new_n30887_, new_n30888_, new_n30890_, new_n30892_, new_n30894_,
    new_n30895_, new_n30897_, new_n30898_, new_n30900_, new_n30902_,
    new_n30904_, new_n30906_, new_n30908_, new_n30909_, new_n30910_,
    new_n30911_, new_n30912_, new_n30913_, new_n30914_, new_n30915_,
    new_n30916_, new_n30917_, new_n30918_, new_n30919_, new_n30920_,
    new_n30921_, new_n30922_, new_n30923_, new_n30924_, new_n30925_,
    new_n30926_, new_n30927_, new_n30928_, new_n30929_, new_n30931_,
    new_n30932_, new_n30933_, new_n30934_, new_n30935_, new_n30936_,
    new_n30937_, new_n30938_, new_n30939_, new_n30940_, new_n30941_,
    new_n30942_, new_n30943_, new_n30944_, new_n30945_, new_n30946_,
    new_n30947_, new_n30948_, new_n30949_, new_n30950_, new_n30951_,
    new_n30953_, new_n30954_, new_n30956_, new_n30958_, new_n30959_,
    new_n30960_, new_n30961_, new_n30962_, new_n30963_, new_n30964_,
    new_n30965_, new_n30966_, new_n30967_, new_n30968_, new_n30969_,
    new_n30970_, new_n30971_, new_n30972_, new_n30973_, new_n30975_,
    new_n30976_, new_n30977_, new_n30978_, new_n30979_, new_n30980_,
    new_n30981_, new_n30982_, new_n30983_, new_n30984_, new_n30985_,
    new_n30986_, new_n30987_, new_n30988_, new_n30989_, new_n30990_,
    new_n30991_, new_n30992_, new_n30994_, new_n30995_, new_n30996_,
    new_n30997_, new_n30998_, new_n30999_, new_n31000_, new_n31001_,
    new_n31002_, new_n31003_, new_n31004_, new_n31005_, new_n31006_,
    new_n31007_, new_n31008_, new_n31009_, new_n31011_, new_n31012_,
    new_n31013_, new_n31014_, new_n31015_, new_n31016_, new_n31017_,
    new_n31018_, new_n31019_, new_n31020_, new_n31021_, new_n31022_,
    new_n31023_, new_n31024_, new_n31025_, new_n31026_, new_n31028_,
    new_n31030_, new_n31031_, new_n31032_, new_n31033_, new_n31034_,
    new_n31035_, new_n31036_, new_n31037_, new_n31038_, new_n31039_,
    new_n31040_, new_n31041_, new_n31042_, new_n31043_, new_n31044_,
    new_n31045_, new_n31046_, new_n31047_, new_n31048_, new_n31049_,
    new_n31051_, new_n31052_, new_n31053_, new_n31054_, new_n31055_,
    new_n31056_, new_n31057_, new_n31058_, new_n31059_, new_n31060_,
    new_n31061_, new_n31062_, new_n31063_, new_n31064_, new_n31065_,
    new_n31066_, new_n31067_, new_n31069_, new_n31070_, new_n31071_,
    new_n31072_, new_n31073_, new_n31074_, new_n31075_, new_n31076_,
    new_n31077_, new_n31078_, new_n31079_, new_n31080_, new_n31081_,
    new_n31082_, new_n31083_, new_n31084_, new_n31085_, new_n31086_,
    new_n31087_, new_n31089_, new_n31090_, new_n31091_, new_n31092_,
    new_n31093_, new_n31094_, new_n31095_, new_n31096_, new_n31097_,
    new_n31098_, new_n31099_, new_n31100_, new_n31101_, new_n31102_,
    new_n31103_, new_n31104_, new_n31105_, new_n31107_, new_n31108_,
    new_n31109_, new_n31110_, new_n31111_, new_n31112_, new_n31113_,
    new_n31114_, new_n31115_, new_n31116_, new_n31117_, new_n31118_,
    new_n31119_, new_n31120_, new_n31121_, new_n31122_, new_n31124_,
    new_n31125_, new_n31126_, new_n31127_, new_n31128_, new_n31129_,
    new_n31130_, new_n31131_, new_n31132_, new_n31133_, new_n31134_,
    new_n31135_, new_n31136_, new_n31137_, new_n31138_, new_n31139_,
    new_n31140_, new_n31141_, new_n31142_, new_n31143_, new_n31144_,
    new_n31145_, new_n31146_, new_n31147_, new_n31148_, new_n31149_,
    new_n31150_, new_n31151_, new_n31152_, new_n31153_, new_n31154_,
    new_n31155_, new_n31156_, new_n31157_, new_n31158_, new_n31159_,
    new_n31160_, new_n31161_, new_n31162_, new_n31164_, new_n31165_,
    new_n31166_, new_n31167_, new_n31168_, new_n31169_, new_n31170_,
    new_n31171_, new_n31172_, new_n31173_, new_n31174_, new_n31175_,
    new_n31176_, new_n31177_, new_n31178_, new_n31179_, new_n31180_,
    new_n31181_, new_n31182_, new_n31183_, new_n31185_, new_n31187_,
    new_n31189_, new_n31190_, new_n31192_, new_n31194_, new_n31196_,
    new_n31197_, new_n31199_, new_n31201_, new_n31203_, new_n31204_,
    new_n31205_, new_n31206_, new_n31207_, new_n31208_, new_n31209_,
    new_n31210_, new_n31211_, new_n31212_, new_n31214_, new_n31216_,
    new_n31217_, new_n31218_, new_n31219_, new_n31220_, new_n31221_,
    new_n31222_, new_n31223_, new_n31224_, new_n31225_, new_n31226_,
    new_n31227_, new_n31228_, new_n31229_, new_n31230_, new_n31231_,
    new_n31232_, new_n31233_, new_n31234_, new_n31235_, new_n31237_,
    new_n31238_, new_n31240_, new_n31242_, new_n31244_, new_n31245_,
    new_n31247_, new_n31248_, new_n31250_, new_n31251_, new_n31253_,
    new_n31254_, new_n31256_, new_n31258_, new_n31260_, new_n31261_,
    new_n31263_, new_n31265_, new_n31267_, new_n31268_, new_n31270_,
    new_n31271_, new_n31272_, new_n31273_, new_n31274_, new_n31275_,
    new_n31276_, new_n31278_, new_n31279_, new_n31281_, new_n31282_,
    new_n31284_, new_n31286_, new_n31288_, new_n31290_, new_n31292_,
    new_n31294_, new_n31296_, new_n31298_, new_n31300_, new_n31301_,
    new_n31303_, new_n31304_, new_n31306_, new_n31308_, new_n31310_,
    new_n31312_, new_n31313_, new_n31314_, new_n31316_, new_n31317_,
    new_n31319_, new_n31320_, new_n31322_, new_n31323_, new_n31324_,
    new_n31325_, new_n31326_, new_n31327_, new_n31328_, new_n31329_,
    new_n31330_, new_n31331_, new_n31332_, new_n31333_, new_n31334_,
    new_n31335_, new_n31336_, new_n31337_, new_n31338_, new_n31339_,
    new_n31340_, new_n31341_, new_n31342_, new_n31344_, new_n31345_,
    new_n31347_, new_n31349_, new_n31351_, new_n31352_, new_n31353_,
    new_n31354_, new_n31355_, new_n31356_, new_n31357_, new_n31358_,
    new_n31359_, new_n31360_, new_n31362_, new_n31364_, new_n31365_,
    new_n31366_, new_n31367_, new_n31368_, new_n31369_, new_n31371_,
    new_n31372_, new_n31374_, new_n31375_, new_n31377_, new_n31378_,
    new_n31379_, new_n31380_, new_n31382_, new_n31384_, new_n31385_,
    new_n31386_, new_n31387_, new_n31388_, new_n31389_, new_n31390_,
    new_n31391_, new_n31392_, new_n31394_, new_n31396_, new_n31398_,
    new_n31399_, new_n31400_, new_n31401_, new_n31403_, new_n31407_,
    new_n31419_, new_n31422_, new_n31423_, new_n31424_, new_n31425_,
    new_n31426_, new_n31429_, new_n31434_, new_n31437_, new_n31441_,
    new_n31445_, new_n31448_, new_n31455_, new_n31458_, new_n31461_,
    new_n31462_, new_n31463_, new_n31464_, new_n31465_, new_n31466_,
    new_n31467_, new_n31468_, new_n31469_, new_n31470_, new_n31471_,
    new_n31472_, new_n31475_, new_n31476_, new_n31477_, new_n31478_,
    new_n31479_, new_n31480_, new_n31481_, new_n31482_, new_n31483_,
    new_n31484_, new_n31485_, new_n31488_, new_n31489_, new_n31490_,
    new_n31491_, new_n31492_, new_n31493_, new_n31494_, new_n31495_,
    new_n31496_, new_n31497_, new_n31498_, new_n31499_, new_n31502_,
    new_n31503_, new_n31504_, new_n31505_, new_n31506_, new_n31507_,
    new_n31508_, new_n31509_, new_n31510_, new_n31511_, new_n31512_,
    new_n31514_, new_n31517_, new_n31521_, new_n31522_, new_n31548_,
    new_n31549_, new_n31550_, new_n31559_, new_n31560_, new_n31561_,
    new_n31568_, new_n31569_, new_n31570_, new_n31573_, new_n31574_,
    new_n31575_, new_n31577_, new_n31578_, new_n31579_, new_n31581_,
    new_n31582_, new_n31583_, new_n31629_, new_n31630_, new_n31631_,
    new_n31632_, new_n31633_, new_n31634_, new_n31663_;
  INVX1    g00000(.A(pi0057), .Y(new_n2436_));
  INVX1    g00001(.A(pi0221), .Y(new_n2437_));
  INVX1    g00002(.A(pi0216), .Y(new_n2438_));
  INVX1    g00003(.A(pi1144), .Y(new_n2439_));
  AOI21X1  g00004(.A0(pi0833), .A1(new_n2438_), .B0(new_n2439_), .Y(new_n2440_));
  INVX1    g00005(.A(new_n2440_), .Y(new_n2441_));
  AND2X1   g00006(.A(pi0833), .B(new_n2438_), .Y(new_n2442_));
  AOI21X1  g00007(.A0(new_n2442_), .A1(pi0929), .B0(pi0332), .Y(new_n2443_));
  AOI21X1  g00008(.A0(new_n2443_), .A1(new_n2441_), .B0(new_n2437_), .Y(new_n2444_));
  INVX1    g00009(.A(pi0332), .Y(new_n2445_));
  AOI21X1  g00010(.A0(new_n2445_), .A1(pi0265), .B0(new_n2438_), .Y(new_n2446_));
  INVX1    g00011(.A(new_n2446_), .Y(new_n2447_));
  INVX1    g00012(.A(pi0105), .Y(new_n2448_));
  AND2X1   g00013(.A(new_n2445_), .B(pi0153), .Y(new_n2449_));
  INVX1    g00014(.A(new_n2449_), .Y(new_n2450_));
  NOR3X1   g00015(.A(pi0166), .B(pi0161), .C(pi0152), .Y(new_n2451_));
  INVX1    g00016(.A(new_n2451_), .Y(new_n2452_));
  INVX1    g00017(.A(pi0137), .Y(new_n2453_));
  INVX1    g00018(.A(pi0479), .Y(new_n2454_));
  AND2X1   g00019(.A(new_n2454_), .B(pi0095), .Y(new_n2455_));
  INVX1    g00020(.A(pi0032), .Y(new_n2456_));
  NOR2X1   g00021(.A(pi0072), .B(pi0040), .Y(new_n2457_));
  INVX1    g00022(.A(new_n2457_), .Y(new_n2458_));
  OR4X1    g00023(.A(pi0098), .B(pi0088), .C(pi0077), .D(pi0050), .Y(new_n2459_));
  NOR2X1   g00024(.A(new_n2459_), .B(pi0102), .Y(new_n2460_));
  INVX1    g00025(.A(new_n2460_), .Y(new_n2461_));
  OR2X1    g00026(.A(pi0071), .B(pi0065), .Y(new_n2462_));
  OR2X1    g00027(.A(pi0103), .B(pi0083), .Y(new_n2463_));
  OR2X1    g00028(.A(pi0069), .B(pi0067), .Y(new_n2464_));
  OR2X1    g00029(.A(pi0073), .B(pi0066), .Y(new_n2465_));
  OR4X1    g00030(.A(pi0106), .B(pi0085), .C(pi0076), .D(pi0061), .Y(new_n2466_));
  OR4X1    g00031(.A(new_n2466_), .B(pi0089), .C(pi0049), .D(pi0048), .Y(new_n2467_));
  OR2X1    g00032(.A(pi0111), .B(pi0082), .Y(new_n2468_));
  OR4X1    g00033(.A(new_n2468_), .B(pi0084), .C(pi0068), .D(pi0036), .Y(new_n2469_));
  OR4X1    g00034(.A(new_n2469_), .B(new_n2467_), .C(pi0104), .D(pi0045), .Y(new_n2470_));
  OR4X1    g00035(.A(new_n2470_), .B(new_n2465_), .C(new_n2464_), .D(new_n2463_), .Y(new_n2471_));
  OR2X1    g00036(.A(pi0107), .B(pi0063), .Y(new_n2472_));
  OR4X1    g00037(.A(new_n2472_), .B(new_n2471_), .C(new_n2462_), .D(pi0064), .Y(new_n2473_));
  INVX1    g00038(.A(pi0086), .Y(new_n2474_));
  NOR2X1   g00039(.A(pi0060), .B(pi0053), .Y(new_n2475_));
  NAND2X1  g00040(.A(new_n2475_), .B(new_n2474_), .Y(new_n2476_));
  OR2X1    g00041(.A(pi0108), .B(pi0097), .Y(new_n2477_));
  OR4X1    g00042(.A(new_n2477_), .B(new_n2476_), .C(pi0094), .D(pi0046), .Y(new_n2478_));
  NOR4X1   g00043(.A(new_n2478_), .B(new_n2473_), .C(new_n2461_), .D(pi0081), .Y(new_n2479_));
  INVX1    g00044(.A(new_n2479_), .Y(new_n2480_));
  INVX1    g00045(.A(pi0109), .Y(new_n2481_));
  INVX1    g00046(.A(pi0110), .Y(new_n2482_));
  NOR3X1   g00047(.A(pi0091), .B(pi0058), .C(pi0047), .Y(new_n2483_));
  NAND3X1  g00048(.A(new_n2483_), .B(new_n2482_), .C(new_n2481_), .Y(new_n2484_));
  OR4X1    g00049(.A(pi0096), .B(pi0070), .C(pi0051), .D(pi0035), .Y(new_n2485_));
  NOR3X1   g00050(.A(new_n2485_), .B(pi0093), .C(pi0090), .Y(new_n2486_));
  INVX1    g00051(.A(new_n2486_), .Y(new_n2487_));
  NOR4X1   g00052(.A(new_n2487_), .B(new_n2484_), .C(new_n2480_), .D(new_n2458_), .Y(new_n2488_));
  AOI21X1  g00053(.A0(new_n2488_), .A1(pi0225), .B0(new_n2456_), .Y(new_n2489_));
  NOR2X1   g00054(.A(new_n2489_), .B(pi0095), .Y(new_n2490_));
  NOR2X1   g00055(.A(pi0093), .B(pi0090), .Y(new_n2491_));
  INVX1    g00056(.A(new_n2491_), .Y(new_n2492_));
  INVX1    g00057(.A(pi0053), .Y(new_n2493_));
  INVX1    g00058(.A(pi0060), .Y(new_n2494_));
  OR4X1    g00059(.A(new_n2473_), .B(new_n2461_), .C(pi0081), .D(new_n2494_), .Y(new_n2495_));
  AND2X1   g00060(.A(new_n2495_), .B(new_n2493_), .Y(new_n2496_));
  NOR2X1   g00061(.A(pi0094), .B(pi0086), .Y(new_n2497_));
  INVX1    g00062(.A(new_n2497_), .Y(new_n2498_));
  OR4X1    g00063(.A(new_n2473_), .B(new_n2461_), .C(pi0081), .D(pi0060), .Y(new_n2499_));
  AOI21X1  g00064(.A0(new_n2499_), .A1(pi0053), .B0(new_n2498_), .Y(new_n2500_));
  INVX1    g00065(.A(new_n2500_), .Y(new_n2501_));
  INVX1    g00066(.A(pi0058), .Y(new_n2502_));
  NOR3X1   g00067(.A(pi0110), .B(pi0109), .C(pi0046), .Y(new_n2503_));
  INVX1    g00068(.A(new_n2503_), .Y(new_n2504_));
  NOR4X1   g00069(.A(new_n2504_), .B(new_n2477_), .C(pi0091), .D(pi0047), .Y(new_n2505_));
  NAND2X1  g00070(.A(new_n2505_), .B(new_n2502_), .Y(new_n2506_));
  NOR4X1   g00071(.A(new_n2506_), .B(new_n2501_), .C(new_n2496_), .D(new_n2492_), .Y(new_n2507_));
  NOR2X1   g00072(.A(new_n2507_), .B(pi0035), .Y(new_n2508_));
  INVX1    g00073(.A(pi0081), .Y(new_n2509_));
  NOR4X1   g00074(.A(new_n2472_), .B(new_n2471_), .C(new_n2462_), .D(pi0064), .Y(new_n2510_));
  OR2X1    g00075(.A(pi0110), .B(pi0109), .Y(new_n2511_));
  NOR4X1   g00076(.A(new_n2511_), .B(new_n2478_), .C(pi0091), .D(pi0047), .Y(new_n2512_));
  NAND4X1  g00077(.A(new_n2512_), .B(new_n2510_), .C(new_n2460_), .D(new_n2509_), .Y(new_n2513_));
  OR4X1    g00078(.A(new_n2513_), .B(pi0093), .C(pi0090), .D(pi0058), .Y(new_n2514_));
  AND2X1   g00079(.A(new_n2514_), .B(pi0035), .Y(new_n2515_));
  INVX1    g00080(.A(pi0051), .Y(new_n2516_));
  INVX1    g00081(.A(pi0225), .Y(new_n2517_));
  INVX1    g00082(.A(pi0035), .Y(new_n2518_));
  NOR2X1   g00083(.A(pi0090), .B(pi0058), .Y(new_n2519_));
  INVX1    g00084(.A(new_n2519_), .Y(new_n2520_));
  NOR4X1   g00085(.A(new_n2513_), .B(new_n2520_), .C(pi0093), .D(new_n2518_), .Y(new_n2521_));
  AOI21X1  g00086(.A0(new_n2521_), .A1(new_n2517_), .B0(pi0070), .Y(new_n2522_));
  NAND2X1  g00087(.A(new_n2522_), .B(new_n2516_), .Y(new_n2523_));
  NOR3X1   g00088(.A(new_n2523_), .B(new_n2515_), .C(new_n2508_), .Y(new_n2524_));
  NOR2X1   g00089(.A(new_n2524_), .B(pi0096), .Y(new_n2525_));
  INVX1    g00090(.A(pi0096), .Y(new_n2526_));
  OR2X1    g00091(.A(new_n2473_), .B(pi0081), .Y(new_n2527_));
  NOR3X1   g00092(.A(new_n2511_), .B(new_n2478_), .C(pi0047), .Y(new_n2528_));
  INVX1    g00093(.A(new_n2528_), .Y(new_n2529_));
  INVX1    g00094(.A(pi0091), .Y(new_n2530_));
  INVX1    g00095(.A(pi0093), .Y(new_n2531_));
  NOR3X1   g00096(.A(pi0070), .B(pi0051), .C(pi0035), .Y(new_n2532_));
  NAND4X1  g00097(.A(new_n2532_), .B(new_n2519_), .C(new_n2531_), .D(new_n2530_), .Y(new_n2533_));
  NOR4X1   g00098(.A(new_n2533_), .B(new_n2529_), .C(new_n2527_), .D(new_n2461_), .Y(new_n2534_));
  OR2X1    g00099(.A(new_n2534_), .B(new_n2526_), .Y(new_n2535_));
  AND2X1   g00100(.A(new_n2535_), .B(new_n2457_), .Y(new_n2536_));
  INVX1    g00101(.A(new_n2536_), .Y(new_n2537_));
  OAI21X1  g00102(.A0(new_n2537_), .A1(new_n2525_), .B0(new_n2456_), .Y(new_n2538_));
  AOI21X1  g00103(.A0(new_n2538_), .A1(new_n2490_), .B0(new_n2455_), .Y(new_n2539_));
  INVX1    g00104(.A(pi0095), .Y(new_n2540_));
  NOR2X1   g00105(.A(pi0093), .B(pi0035), .Y(new_n2541_));
  INVX1    g00106(.A(new_n2541_), .Y(new_n2542_));
  NOR4X1   g00107(.A(pi0096), .B(pi0072), .C(pi0070), .D(pi0051), .Y(new_n2543_));
  INVX1    g00108(.A(new_n2543_), .Y(new_n2544_));
  NOR4X1   g00109(.A(new_n2544_), .B(new_n2542_), .C(new_n2513_), .D(new_n2520_), .Y(new_n2545_));
  AOI21X1  g00110(.A0(new_n2545_), .A1(pi0040), .B0(pi0032), .Y(new_n2546_));
  INVX1    g00111(.A(new_n2546_), .Y(new_n2547_));
  INVX1    g00112(.A(pi0072), .Y(new_n2548_));
  INVX1    g00113(.A(pi0040), .Y(new_n2549_));
  NOR4X1   g00114(.A(new_n2484_), .B(new_n2478_), .C(new_n2527_), .D(new_n2461_), .Y(new_n2550_));
  AND2X1   g00115(.A(new_n2486_), .B(new_n2550_), .Y(new_n2551_));
  OR2X1    g00116(.A(new_n2551_), .B(new_n2548_), .Y(new_n2552_));
  AND2X1   g00117(.A(new_n2552_), .B(new_n2549_), .Y(new_n2553_));
  INVX1    g00118(.A(new_n2553_), .Y(new_n2554_));
  OR4X1    g00119(.A(new_n2542_), .B(new_n2513_), .C(new_n2520_), .D(pi0070), .Y(new_n2555_));
  AOI21X1  g00120(.A0(new_n2555_), .A1(pi0051), .B0(pi0096), .Y(new_n2556_));
  INVX1    g00121(.A(new_n2556_), .Y(new_n2557_));
  AOI21X1  g00122(.A0(pi0070), .A1(new_n2516_), .B0(new_n2557_), .Y(new_n2558_));
  OAI21X1  g00123(.A0(new_n2514_), .A1(new_n2517_), .B0(pi0035), .Y(new_n2559_));
  INVX1    g00124(.A(new_n2559_), .Y(new_n2560_));
  OR4X1    g00125(.A(new_n2513_), .B(new_n2531_), .C(pi0090), .D(pi0058), .Y(new_n2561_));
  AND2X1   g00126(.A(new_n2561_), .B(new_n2518_), .Y(new_n2562_));
  NOR4X1   g00127(.A(new_n2529_), .B(new_n2473_), .C(new_n2461_), .D(pi0081), .Y(new_n2563_));
  AOI21X1  g00128(.A0(new_n2563_), .A1(pi0091), .B0(new_n2520_), .Y(new_n2564_));
  INVX1    g00129(.A(new_n2564_), .Y(new_n2565_));
  AOI21X1  g00130(.A0(new_n2479_), .A1(new_n2481_), .B0(new_n2482_), .Y(new_n2566_));
  INVX1    g00131(.A(pi0047), .Y(new_n2567_));
  NOR3X1   g00132(.A(new_n2473_), .B(new_n2461_), .C(pi0081), .Y(new_n2568_));
  NOR2X1   g00133(.A(new_n2511_), .B(new_n2478_), .Y(new_n2569_));
  AOI21X1  g00134(.A0(new_n2569_), .A1(new_n2568_), .B0(new_n2567_), .Y(new_n2570_));
  NOR3X1   g00135(.A(new_n2570_), .B(new_n2566_), .C(pi0091), .Y(new_n2571_));
  INVX1    g00136(.A(new_n2571_), .Y(new_n2572_));
  NOR2X1   g00137(.A(pi0110), .B(pi0047), .Y(new_n2573_));
  NOR2X1   g00138(.A(new_n2479_), .B(new_n2481_), .Y(new_n2574_));
  INVX1    g00139(.A(new_n2574_), .Y(new_n2575_));
  INVX1    g00140(.A(pi0108), .Y(new_n2576_));
  OR2X1    g00141(.A(pi0098), .B(pi0088), .Y(new_n2577_));
  INVX1    g00142(.A(pi0102), .Y(new_n2578_));
  NAND3X1  g00143(.A(new_n2510_), .B(new_n2578_), .C(new_n2509_), .Y(new_n2579_));
  INVX1    g00144(.A(pi0050), .Y(new_n2580_));
  INVX1    g00145(.A(pi0077), .Y(new_n2581_));
  NAND4X1  g00146(.A(new_n2497_), .B(new_n2475_), .C(new_n2581_), .D(new_n2580_), .Y(new_n2582_));
  OR4X1    g00147(.A(new_n2582_), .B(new_n2579_), .C(new_n2577_), .D(pi0097), .Y(new_n2583_));
  AOI21X1  g00148(.A0(new_n2583_), .A1(pi0108), .B0(pi0046), .Y(new_n2584_));
  INVX1    g00149(.A(new_n2584_), .Y(new_n2585_));
  OR4X1    g00150(.A(new_n2473_), .B(new_n2577_), .C(pi0102), .D(pi0081), .Y(new_n2586_));
  OR2X1    g00151(.A(new_n2582_), .B(new_n2586_), .Y(new_n2587_));
  AND2X1   g00152(.A(new_n2587_), .B(pi0097), .Y(new_n2588_));
  INVX1    g00153(.A(new_n2588_), .Y(new_n2589_));
  INVX1    g00154(.A(pi0094), .Y(new_n2590_));
  NAND2X1  g00155(.A(new_n2475_), .B(new_n2580_), .Y(new_n2591_));
  NOR3X1   g00156(.A(new_n2579_), .B(new_n2577_), .C(pi0077), .Y(new_n2592_));
  INVX1    g00157(.A(new_n2592_), .Y(new_n2593_));
  NOR4X1   g00158(.A(new_n2593_), .B(new_n2591_), .C(new_n2590_), .D(pi0086), .Y(new_n2594_));
  NOR2X1   g00159(.A(new_n2594_), .B(pi0097), .Y(new_n2595_));
  INVX1    g00160(.A(new_n2595_), .Y(new_n2596_));
  NOR4X1   g00161(.A(new_n2591_), .B(new_n2579_), .C(new_n2577_), .D(pi0077), .Y(new_n2597_));
  OAI21X1  g00162(.A0(new_n2597_), .A1(new_n2474_), .B0(new_n2590_), .Y(new_n2598_));
  AND2X1   g00163(.A(new_n2499_), .B(pi0053), .Y(new_n2599_));
  NOR2X1   g00164(.A(new_n2586_), .B(new_n2581_), .Y(new_n2600_));
  NOR2X1   g00165(.A(new_n2600_), .B(pi0050), .Y(new_n2601_));
  INVX1    g00166(.A(new_n2601_), .Y(new_n2602_));
  AOI21X1  g00167(.A0(new_n2510_), .A1(new_n2509_), .B0(new_n2578_), .Y(new_n2603_));
  AOI21X1  g00168(.A0(new_n2473_), .A1(pi0081), .B0(new_n2603_), .Y(new_n2604_));
  INVX1    g00169(.A(pi0064), .Y(new_n2605_));
  NOR2X1   g00170(.A(new_n2471_), .B(new_n2462_), .Y(new_n2606_));
  INVX1    g00171(.A(new_n2472_), .Y(new_n2607_));
  AOI21X1  g00172(.A0(new_n2607_), .A1(new_n2606_), .B0(new_n2605_), .Y(new_n2608_));
  INVX1    g00173(.A(pi0107), .Y(new_n2609_));
  AND2X1   g00174(.A(new_n2471_), .B(pi0071), .Y(new_n2610_));
  OR2X1    g00175(.A(new_n2610_), .B(pi0065), .Y(new_n2611_));
  NOR3X1   g00176(.A(new_n2470_), .B(new_n2465_), .C(pi0067), .Y(new_n2612_));
  INVX1    g00177(.A(new_n2612_), .Y(new_n2613_));
  INVX1    g00178(.A(pi0083), .Y(new_n2614_));
  INVX1    g00179(.A(pi0103), .Y(new_n2615_));
  NOR3X1   g00180(.A(new_n2470_), .B(new_n2465_), .C(new_n2464_), .Y(new_n2616_));
  OAI21X1  g00181(.A0(new_n2616_), .A1(new_n2614_), .B0(new_n2615_), .Y(new_n2617_));
  AOI21X1  g00182(.A0(new_n2613_), .A1(pi0069), .B0(new_n2617_), .Y(new_n2618_));
  NOR2X1   g00183(.A(pi0083), .B(pi0069), .Y(new_n2619_));
  NOR2X1   g00184(.A(pi0111), .B(pi0068), .Y(new_n2620_));
  OR4X1    g00185(.A(new_n2467_), .B(new_n2465_), .C(pi0104), .D(pi0045), .Y(new_n2621_));
  AND2X1   g00186(.A(new_n2621_), .B(pi0084), .Y(new_n2622_));
  INVX1    g00187(.A(new_n2465_), .Y(new_n2623_));
  NOR3X1   g00188(.A(new_n2467_), .B(pi0104), .C(pi0045), .Y(new_n2624_));
  NOR2X1   g00189(.A(new_n2467_), .B(pi0104), .Y(new_n2625_));
  OR2X1    g00190(.A(pi0076), .B(pi0061), .Y(new_n2626_));
  OR2X1    g00191(.A(pi0106), .B(pi0085), .Y(new_n2627_));
  OR4X1    g00192(.A(new_n2627_), .B(new_n2626_), .C(pi0089), .D(pi0048), .Y(new_n2628_));
  INVX1    g00193(.A(pi0048), .Y(new_n2629_));
  INVX1    g00194(.A(new_n2466_), .Y(new_n2630_));
  AND2X1   g00195(.A(pi0106), .B(pi0085), .Y(new_n2631_));
  AND2X1   g00196(.A(pi0076), .B(pi0061), .Y(new_n2632_));
  OAI22X1  g00197(.A0(new_n2632_), .A1(new_n2627_), .B0(new_n2631_), .B1(new_n2626_), .Y(new_n2633_));
  AOI21X1  g00198(.A0(new_n2633_), .A1(new_n2629_), .B0(new_n2630_), .Y(new_n2634_));
  INVX1    g00199(.A(pi0089), .Y(new_n2635_));
  AOI21X1  g00200(.A0(new_n2630_), .A1(new_n2629_), .B0(new_n2635_), .Y(new_n2636_));
  OR2X1    g00201(.A(new_n2636_), .B(pi0049), .Y(new_n2637_));
  OAI21X1  g00202(.A0(new_n2637_), .A1(new_n2634_), .B0(new_n2628_), .Y(new_n2638_));
  AOI21X1  g00203(.A0(new_n2467_), .A1(pi0104), .B0(pi0045), .Y(new_n2639_));
  AOI21X1  g00204(.A0(new_n2639_), .A1(new_n2638_), .B0(new_n2625_), .Y(new_n2640_));
  OAI21X1  g00205(.A0(new_n2640_), .A1(new_n2624_), .B0(new_n2623_), .Y(new_n2641_));
  INVX1    g00206(.A(new_n2624_), .Y(new_n2642_));
  AND2X1   g00207(.A(pi0073), .B(pi0066), .Y(new_n2643_));
  AOI21X1  g00208(.A0(new_n2642_), .A1(new_n2465_), .B0(new_n2643_), .Y(new_n2644_));
  AOI21X1  g00209(.A0(new_n2644_), .A1(new_n2641_), .B0(pi0084), .Y(new_n2645_));
  OAI21X1  g00210(.A0(new_n2645_), .A1(new_n2622_), .B0(new_n2620_), .Y(new_n2646_));
  OR2X1    g00211(.A(new_n2621_), .B(pi0084), .Y(new_n2647_));
  INVX1    g00212(.A(pi0082), .Y(new_n2648_));
  INVX1    g00213(.A(pi0111), .Y(new_n2649_));
  NOR3X1   g00214(.A(new_n2621_), .B(pi0084), .C(pi0068), .Y(new_n2650_));
  OAI21X1  g00215(.A0(new_n2650_), .A1(new_n2649_), .B0(new_n2648_), .Y(new_n2651_));
  AOI21X1  g00216(.A0(new_n2647_), .A1(pi0068), .B0(new_n2651_), .Y(new_n2652_));
  NOR2X1   g00217(.A(pi0067), .B(pi0036), .Y(new_n2653_));
  INVX1    g00218(.A(new_n2620_), .Y(new_n2654_));
  OR4X1    g00219(.A(new_n2621_), .B(new_n2654_), .C(pi0084), .D(new_n2648_), .Y(new_n2655_));
  NAND2X1  g00220(.A(new_n2655_), .B(new_n2653_), .Y(new_n2656_));
  AOI21X1  g00221(.A0(new_n2652_), .A1(new_n2646_), .B0(new_n2656_), .Y(new_n2657_));
  INVX1    g00222(.A(pi0036), .Y(new_n2658_));
  OAI21X1  g00223(.A0(new_n2470_), .A1(new_n2465_), .B0(pi0067), .Y(new_n2659_));
  NOR4X1   g00224(.A(new_n2621_), .B(new_n2468_), .C(pi0084), .D(pi0068), .Y(new_n2660_));
  OAI21X1  g00225(.A0(new_n2660_), .A1(new_n2658_), .B0(new_n2659_), .Y(new_n2661_));
  OAI21X1  g00226(.A0(new_n2661_), .A1(new_n2657_), .B0(new_n2619_), .Y(new_n2662_));
  INVX1    g00227(.A(pi0071), .Y(new_n2663_));
  NAND3X1  g00228(.A(new_n2619_), .B(new_n2612_), .C(pi0103), .Y(new_n2664_));
  NAND2X1  g00229(.A(new_n2664_), .B(new_n2663_), .Y(new_n2665_));
  AOI21X1  g00230(.A0(new_n2662_), .A1(new_n2618_), .B0(new_n2665_), .Y(new_n2666_));
  OAI21X1  g00231(.A0(new_n2666_), .A1(new_n2611_), .B0(new_n2609_), .Y(new_n2667_));
  INVX1    g00232(.A(pi0065), .Y(new_n2668_));
  NOR3X1   g00233(.A(new_n2471_), .B(pi0071), .C(new_n2668_), .Y(new_n2669_));
  INVX1    g00234(.A(new_n2606_), .Y(new_n2670_));
  AOI21X1  g00235(.A0(new_n2670_), .A1(pi0107), .B0(pi0063), .Y(new_n2671_));
  OAI21X1  g00236(.A0(new_n2669_), .A1(new_n2667_), .B0(new_n2671_), .Y(new_n2672_));
  AOI21X1  g00237(.A0(new_n2672_), .A1(new_n2605_), .B0(new_n2608_), .Y(new_n2673_));
  INVX1    g00238(.A(pi0063), .Y(new_n2674_));
  OR2X1    g00239(.A(pi0107), .B(new_n2674_), .Y(new_n2675_));
  OAI21X1  g00240(.A0(new_n2675_), .A1(new_n2670_), .B0(new_n2605_), .Y(new_n2676_));
  AOI21X1  g00241(.A0(new_n2671_), .A1(new_n2667_), .B0(new_n2676_), .Y(new_n2677_));
  NOR2X1   g00242(.A(new_n2677_), .B(new_n2608_), .Y(new_n2678_));
  OR4X1    g00243(.A(new_n2678_), .B(new_n2673_), .C(pi0102), .D(pi0081), .Y(new_n2679_));
  AOI21X1  g00244(.A0(new_n2679_), .A1(new_n2604_), .B0(new_n2577_), .Y(new_n2680_));
  INVX1    g00245(.A(pi0088), .Y(new_n2681_));
  OR4X1    g00246(.A(new_n2473_), .B(pi0102), .C(pi0098), .D(pi0081), .Y(new_n2682_));
  INVX1    g00247(.A(new_n2682_), .Y(new_n2683_));
  AOI21X1  g00248(.A0(new_n2579_), .A1(pi0098), .B0(pi0077), .Y(new_n2684_));
  OAI21X1  g00249(.A0(new_n2683_), .A1(new_n2681_), .B0(new_n2684_), .Y(new_n2685_));
  NOR2X1   g00250(.A(new_n2685_), .B(new_n2680_), .Y(new_n2686_));
  AOI21X1  g00251(.A0(new_n2593_), .A1(pi0050), .B0(pi0060), .Y(new_n2687_));
  OAI21X1  g00252(.A0(new_n2686_), .A1(new_n2602_), .B0(new_n2687_), .Y(new_n2688_));
  AND2X1   g00253(.A(new_n2688_), .B(new_n2496_), .Y(new_n2689_));
  OR2X1    g00254(.A(new_n2689_), .B(new_n2599_), .Y(new_n2690_));
  AOI21X1  g00255(.A0(new_n2690_), .A1(new_n2474_), .B0(new_n2598_), .Y(new_n2691_));
  OAI21X1  g00256(.A0(new_n2691_), .A1(new_n2596_), .B0(new_n2589_), .Y(new_n2692_));
  AOI21X1  g00257(.A0(new_n2692_), .A1(new_n2576_), .B0(new_n2585_), .Y(new_n2693_));
  INVX1    g00258(.A(pi0046), .Y(new_n2694_));
  NOR4X1   g00259(.A(new_n2582_), .B(new_n2586_), .C(new_n2477_), .D(new_n2694_), .Y(new_n2695_));
  NOR2X1   g00260(.A(new_n2695_), .B(pi0109), .Y(new_n2696_));
  INVX1    g00261(.A(new_n2696_), .Y(new_n2697_));
  OAI21X1  g00262(.A0(new_n2697_), .A1(new_n2693_), .B0(new_n2575_), .Y(new_n2698_));
  AOI21X1  g00263(.A0(new_n2698_), .A1(new_n2573_), .B0(new_n2572_), .Y(new_n2699_));
  AND2X1   g00264(.A(new_n2513_), .B(pi0058), .Y(new_n2700_));
  INVX1    g00265(.A(pi0090), .Y(new_n2701_));
  NOR2X1   g00266(.A(new_n2550_), .B(new_n2701_), .Y(new_n2702_));
  NOR3X1   g00267(.A(new_n2702_), .B(new_n2700_), .C(pi0093), .Y(new_n2703_));
  OAI21X1  g00268(.A0(new_n2699_), .A1(new_n2565_), .B0(new_n2703_), .Y(new_n2704_));
  AOI21X1  g00269(.A0(new_n2704_), .A1(new_n2562_), .B0(new_n2560_), .Y(new_n2705_));
  OAI21X1  g00270(.A0(new_n2705_), .A1(pi0051), .B0(new_n2558_), .Y(new_n2706_));
  AOI21X1  g00271(.A0(new_n2706_), .A1(new_n2548_), .B0(new_n2554_), .Y(new_n2707_));
  NOR2X1   g00272(.A(new_n2707_), .B(new_n2547_), .Y(new_n2708_));
  OR4X1    g00273(.A(new_n2542_), .B(new_n2513_), .C(pi0090), .D(pi0058), .Y(new_n2709_));
  OR2X1    g00274(.A(pi0072), .B(pi0051), .Y(new_n2710_));
  NOR3X1   g00275(.A(new_n2710_), .B(new_n2709_), .C(pi0040), .Y(new_n2711_));
  NAND3X1  g00276(.A(new_n2711_), .B(new_n2534_), .C(pi0096), .Y(new_n2712_));
  AND2X1   g00277(.A(new_n2712_), .B(new_n2708_), .Y(new_n2713_));
  OAI21X1  g00278(.A0(new_n2713_), .A1(new_n2489_), .B0(new_n2540_), .Y(new_n2714_));
  NOR2X1   g00279(.A(pi0040), .B(pi0032), .Y(new_n2715_));
  AOI21X1  g00280(.A0(new_n2715_), .A1(new_n2545_), .B0(new_n2540_), .Y(new_n2716_));
  AND2X1   g00281(.A(new_n2716_), .B(pi0479), .Y(new_n2717_));
  INVX1    g00282(.A(new_n2717_), .Y(new_n2718_));
  AOI21X1  g00283(.A0(new_n2718_), .A1(new_n2714_), .B0(new_n2453_), .Y(new_n2719_));
  AOI21X1  g00284(.A0(new_n2539_), .A1(new_n2453_), .B0(new_n2719_), .Y(new_n2720_));
  INVX1    g00285(.A(pi0833), .Y(new_n2721_));
  INVX1    g00286(.A(pi1091), .Y(new_n2722_));
  AOI21X1  g00287(.A0(pi0957), .A1(new_n2721_), .B0(new_n2722_), .Y(new_n2723_));
  INVX1    g00288(.A(new_n2723_), .Y(new_n2724_));
  OR2X1    g00289(.A(pi0096), .B(pi0070), .Y(new_n2725_));
  INVX1    g00290(.A(pi0841), .Y(new_n2726_));
  OR4X1    g00291(.A(new_n2513_), .B(new_n2520_), .C(new_n2726_), .D(pi0093), .Y(new_n2727_));
  NAND3X1  g00292(.A(pi0225), .B(new_n2549_), .C(new_n2518_), .Y(new_n2728_));
  NOR4X1   g00293(.A(new_n2728_), .B(new_n2727_), .C(new_n2710_), .D(new_n2725_), .Y(new_n2729_));
  NOR2X1   g00294(.A(new_n2729_), .B(new_n2456_), .Y(new_n2730_));
  OAI21X1  g00295(.A0(new_n2730_), .A1(new_n2713_), .B0(new_n2540_), .Y(new_n2731_));
  AOI21X1  g00296(.A0(new_n2731_), .A1(new_n2718_), .B0(new_n2453_), .Y(new_n2732_));
  INVX1    g00297(.A(new_n2730_), .Y(new_n2733_));
  AND2X1   g00298(.A(new_n2733_), .B(new_n2538_), .Y(new_n2734_));
  MX2X1    g00299(.A(new_n2734_), .B(new_n2454_), .S0(pi0095), .Y(new_n2735_));
  NOR2X1   g00300(.A(new_n2735_), .B(pi0137), .Y(new_n2736_));
  NOR2X1   g00301(.A(new_n2736_), .B(new_n2732_), .Y(new_n2737_));
  NAND2X1  g00302(.A(pi0950), .B(pi0829), .Y(new_n2738_));
  AND2X1   g00303(.A(pi1093), .B(pi1092), .Y(new_n2739_));
  INVX1    g00304(.A(new_n2739_), .Y(new_n2740_));
  OAI21X1  g00305(.A0(new_n2740_), .A1(new_n2738_), .B0(new_n2735_), .Y(new_n2741_));
  NOR2X1   g00306(.A(new_n2523_), .B(new_n2515_), .Y(new_n2742_));
  NOR3X1   g00307(.A(new_n2588_), .B(pi0110), .C(pi0108), .Y(new_n2743_));
  NAND2X1  g00308(.A(new_n2519_), .B(new_n2531_), .Y(new_n2744_));
  INVX1    g00309(.A(new_n2496_), .Y(new_n2745_));
  AOI21X1  g00310(.A0(new_n2500_), .A1(new_n2745_), .B0(pi0097), .Y(new_n2746_));
  NOR4X1   g00311(.A(pi0109), .B(pi0091), .C(pi0047), .D(pi0046), .Y(new_n2747_));
  INVX1    g00312(.A(new_n2747_), .Y(new_n2748_));
  NOR3X1   g00313(.A(new_n2748_), .B(new_n2746_), .C(new_n2744_), .Y(new_n2749_));
  AOI21X1  g00314(.A0(new_n2749_), .A1(new_n2743_), .B0(pi0035), .Y(new_n2750_));
  INVX1    g00315(.A(new_n2750_), .Y(new_n2751_));
  AOI21X1  g00316(.A0(new_n2751_), .A1(new_n2742_), .B0(pi0096), .Y(new_n2752_));
  OAI21X1  g00317(.A0(new_n2752_), .A1(new_n2537_), .B0(new_n2456_), .Y(new_n2753_));
  AOI21X1  g00318(.A0(new_n2753_), .A1(new_n2733_), .B0(pi0095), .Y(new_n2754_));
  INVX1    g00319(.A(pi1092), .Y(new_n2755_));
  INVX1    g00320(.A(pi1093), .Y(new_n2756_));
  NOR3X1   g00321(.A(new_n2738_), .B(new_n2756_), .C(new_n2755_), .Y(new_n2757_));
  OAI21X1  g00322(.A0(new_n2454_), .A1(new_n2540_), .B0(new_n2757_), .Y(new_n2758_));
  OR2X1    g00323(.A(new_n2758_), .B(new_n2754_), .Y(new_n2759_));
  AND2X1   g00324(.A(new_n2759_), .B(new_n2453_), .Y(new_n2760_));
  AND2X1   g00325(.A(new_n2760_), .B(new_n2741_), .Y(new_n2761_));
  NOR3X1   g00326(.A(new_n2761_), .B(new_n2732_), .C(new_n2724_), .Y(new_n2762_));
  AOI21X1  g00327(.A0(new_n2737_), .A1(new_n2724_), .B0(new_n2762_), .Y(new_n2763_));
  INVX1    g00328(.A(new_n2763_), .Y(new_n2764_));
  MX2X1    g00329(.A(new_n2764_), .B(new_n2720_), .S0(pi0210), .Y(new_n2765_));
  INVX1    g00330(.A(pi0210), .Y(new_n2766_));
  NOR3X1   g00331(.A(pi0096), .B(pi0072), .C(pi0040), .Y(new_n2767_));
  INVX1    g00332(.A(new_n2767_), .Y(new_n2768_));
  NOR4X1   g00333(.A(new_n2768_), .B(new_n2523_), .C(new_n2515_), .D(new_n2508_), .Y(new_n2769_));
  OAI21X1  g00334(.A0(new_n2769_), .A1(pi0032), .B0(new_n2490_), .Y(new_n2770_));
  AND2X1   g00335(.A(new_n2770_), .B(new_n2453_), .Y(new_n2771_));
  NOR2X1   g00336(.A(new_n2716_), .B(new_n2455_), .Y(new_n2772_));
  NOR2X1   g00337(.A(new_n2708_), .B(new_n2489_), .Y(new_n2773_));
  OAI21X1  g00338(.A0(new_n2773_), .A1(pi0095), .B0(new_n2772_), .Y(new_n2774_));
  AOI21X1  g00339(.A0(new_n2774_), .A1(pi0137), .B0(new_n2771_), .Y(new_n2775_));
  NOR2X1   g00340(.A(new_n2730_), .B(pi0095), .Y(new_n2776_));
  INVX1    g00341(.A(new_n2776_), .Y(new_n2777_));
  AND2X1   g00342(.A(new_n2757_), .B(new_n2723_), .Y(new_n2778_));
  NOR2X1   g00343(.A(new_n2778_), .B(new_n2508_), .Y(new_n2779_));
  INVX1    g00344(.A(pi0957), .Y(new_n2780_));
  AND2X1   g00345(.A(pi1093), .B(pi1091), .Y(new_n2781_));
  OAI21X1  g00346(.A0(new_n2780_), .A1(pi0833), .B0(new_n2781_), .Y(new_n2782_));
  AND2X1   g00347(.A(pi1092), .B(pi0950), .Y(new_n2783_));
  AND2X1   g00348(.A(new_n2783_), .B(pi0829), .Y(new_n2784_));
  INVX1    g00349(.A(new_n2784_), .Y(new_n2785_));
  NOR3X1   g00350(.A(new_n2785_), .B(new_n2782_), .C(new_n2750_), .Y(new_n2786_));
  NOR3X1   g00351(.A(new_n2768_), .B(new_n2523_), .C(new_n2515_), .Y(new_n2787_));
  OAI21X1  g00352(.A0(new_n2786_), .A1(new_n2779_), .B0(new_n2787_), .Y(new_n2788_));
  AND2X1   g00353(.A(new_n2788_), .B(new_n2456_), .Y(new_n2789_));
  OAI21X1  g00354(.A0(new_n2789_), .A1(new_n2777_), .B0(new_n2453_), .Y(new_n2790_));
  INVX1    g00355(.A(new_n2790_), .Y(new_n2791_));
  OAI21X1  g00356(.A0(new_n2730_), .A1(new_n2708_), .B0(new_n2540_), .Y(new_n2792_));
  AOI21X1  g00357(.A0(new_n2792_), .A1(new_n2772_), .B0(new_n2453_), .Y(new_n2793_));
  OAI21X1  g00358(.A0(new_n2793_), .A1(new_n2791_), .B0(new_n2766_), .Y(new_n2794_));
  OAI21X1  g00359(.A0(new_n2775_), .A1(new_n2766_), .B0(new_n2794_), .Y(new_n2795_));
  OAI21X1  g00360(.A0(new_n2795_), .A1(pi0234), .B0(new_n2445_), .Y(new_n2796_));
  AOI21X1  g00361(.A0(new_n2765_), .A1(pi0234), .B0(new_n2796_), .Y(new_n2797_));
  AND2X1   g00362(.A(new_n2445_), .B(pi0234), .Y(new_n2798_));
  NOR2X1   g00363(.A(new_n2737_), .B(pi0210), .Y(new_n2799_));
  INVX1    g00364(.A(pi0146), .Y(new_n2800_));
  OAI21X1  g00365(.A0(new_n2720_), .A1(new_n2766_), .B0(new_n2800_), .Y(new_n2801_));
  OAI21X1  g00366(.A0(new_n2801_), .A1(new_n2799_), .B0(new_n2798_), .Y(new_n2802_));
  AOI21X1  g00367(.A0(new_n2765_), .A1(pi0146), .B0(new_n2802_), .Y(new_n2803_));
  NOR2X1   g00368(.A(new_n2795_), .B(new_n2800_), .Y(new_n2804_));
  OAI21X1  g00369(.A0(new_n2769_), .A1(pi0032), .B0(new_n2776_), .Y(new_n2805_));
  AND2X1   g00370(.A(new_n2805_), .B(new_n2453_), .Y(new_n2806_));
  OR2X1    g00371(.A(new_n2806_), .B(new_n2793_), .Y(new_n2807_));
  AND2X1   g00372(.A(new_n2807_), .B(new_n2766_), .Y(new_n2808_));
  OAI21X1  g00373(.A0(new_n2775_), .A1(new_n2766_), .B0(new_n2800_), .Y(new_n2809_));
  NOR2X1   g00374(.A(pi0332), .B(pi0234), .Y(new_n2810_));
  OAI21X1  g00375(.A0(new_n2809_), .A1(new_n2808_), .B0(new_n2810_), .Y(new_n2811_));
  OAI21X1  g00376(.A0(new_n2811_), .A1(new_n2804_), .B0(new_n2452_), .Y(new_n2812_));
  OAI22X1  g00377(.A0(new_n2812_), .A1(new_n2803_), .B0(new_n2797_), .B1(new_n2452_), .Y(new_n2813_));
  MX2X1    g00378(.A(new_n2813_), .B(new_n2450_), .S0(new_n2448_), .Y(new_n2814_));
  INVX1    g00379(.A(new_n2716_), .Y(new_n2815_));
  INVX1    g00380(.A(new_n2558_), .Y(new_n2816_));
  INVX1    g00381(.A(new_n2703_), .Y(new_n2817_));
  INVX1    g00382(.A(new_n2573_), .Y(new_n2818_));
  MX2X1    g00383(.A(new_n2693_), .B(new_n2479_), .S0(pi0109), .Y(new_n2819_));
  OAI21X1  g00384(.A0(new_n2819_), .A1(new_n2818_), .B0(new_n2571_), .Y(new_n2820_));
  AND2X1   g00385(.A(new_n2820_), .B(new_n2564_), .Y(new_n2821_));
  OAI21X1  g00386(.A0(new_n2821_), .A1(new_n2817_), .B0(new_n2562_), .Y(new_n2822_));
  AOI21X1  g00387(.A0(new_n2822_), .A1(new_n2559_), .B0(pi0051), .Y(new_n2823_));
  OAI21X1  g00388(.A0(new_n2823_), .A1(new_n2816_), .B0(new_n2548_), .Y(new_n2824_));
  AOI21X1  g00389(.A0(new_n2824_), .A1(new_n2553_), .B0(new_n2547_), .Y(new_n2825_));
  AND2X1   g00390(.A(new_n2825_), .B(new_n2712_), .Y(new_n2826_));
  OAI21X1  g00391(.A0(new_n2826_), .A1(new_n2730_), .B0(new_n2540_), .Y(new_n2827_));
  AOI21X1  g00392(.A0(new_n2827_), .A1(new_n2815_), .B0(new_n2453_), .Y(new_n2828_));
  AND2X1   g00393(.A(pi0957), .B(new_n2721_), .Y(new_n2829_));
  NOR2X1   g00394(.A(new_n2451_), .B(pi0146), .Y(new_n2830_));
  NOR3X1   g00395(.A(new_n2830_), .B(new_n2829_), .C(new_n2722_), .Y(new_n2831_));
  NAND2X1  g00396(.A(new_n2735_), .B(new_n2815_), .Y(new_n2832_));
  AOI21X1  g00397(.A0(new_n2831_), .A1(new_n2741_), .B0(new_n2832_), .Y(new_n2833_));
  NOR4X1   g00398(.A(new_n2830_), .B(new_n2759_), .C(new_n2724_), .D(new_n2716_), .Y(new_n2834_));
  NOR3X1   g00399(.A(new_n2834_), .B(new_n2833_), .C(pi0137), .Y(new_n2835_));
  OAI21X1  g00400(.A0(new_n2835_), .A1(new_n2828_), .B0(new_n2766_), .Y(new_n2836_));
  OAI21X1  g00401(.A0(new_n2825_), .A1(new_n2730_), .B0(new_n2540_), .Y(new_n2837_));
  AOI21X1  g00402(.A0(new_n2837_), .A1(new_n2772_), .B0(new_n2453_), .Y(new_n2838_));
  OR2X1    g00403(.A(pi0234), .B(pi0210), .Y(new_n2839_));
  AOI21X1  g00404(.A0(new_n2830_), .A1(new_n2806_), .B0(new_n2839_), .Y(new_n2840_));
  OAI21X1  g00405(.A0(new_n2830_), .A1(new_n2790_), .B0(new_n2840_), .Y(new_n2841_));
  OAI21X1  g00406(.A0(new_n2825_), .A1(new_n2489_), .B0(new_n2540_), .Y(new_n2842_));
  AOI21X1  g00407(.A0(new_n2842_), .A1(new_n2772_), .B0(new_n2453_), .Y(new_n2843_));
  OR2X1    g00408(.A(new_n2771_), .B(new_n2766_), .Y(new_n2844_));
  OAI22X1  g00409(.A0(new_n2844_), .A1(new_n2843_), .B0(new_n2841_), .B1(new_n2838_), .Y(new_n2845_));
  AOI21X1  g00410(.A0(new_n2836_), .A1(pi0234), .B0(new_n2845_), .Y(new_n2846_));
  OAI21X1  g00411(.A0(new_n2826_), .A1(new_n2489_), .B0(new_n2540_), .Y(new_n2847_));
  NOR2X1   g00412(.A(new_n2716_), .B(new_n2453_), .Y(new_n2848_));
  NOR2X1   g00413(.A(new_n2716_), .B(pi0137), .Y(new_n2849_));
  INVX1    g00414(.A(new_n2849_), .Y(new_n2850_));
  AND2X1   g00415(.A(pi0234), .B(pi0210), .Y(new_n2851_));
  OAI21X1  g00416(.A0(new_n2850_), .A1(new_n2539_), .B0(new_n2851_), .Y(new_n2852_));
  AOI21X1  g00417(.A0(new_n2848_), .A1(new_n2847_), .B0(new_n2852_), .Y(new_n2853_));
  OAI21X1  g00418(.A0(new_n2853_), .A1(new_n2846_), .B0(new_n2449_), .Y(new_n2854_));
  OAI21X1  g00419(.A0(new_n2513_), .A1(new_n2520_), .B0(pi0093), .Y(new_n2855_));
  AND2X1   g00420(.A(new_n2855_), .B(new_n2518_), .Y(new_n2856_));
  NOR2X1   g00421(.A(new_n2702_), .B(new_n2700_), .Y(new_n2857_));
  INVX1    g00422(.A(new_n2857_), .Y(new_n2858_));
  OR2X1    g00423(.A(new_n2688_), .B(pi0053), .Y(new_n2859_));
  AOI21X1  g00424(.A0(new_n2859_), .A1(new_n2474_), .B0(new_n2598_), .Y(new_n2860_));
  NOR2X1   g00425(.A(new_n2860_), .B(new_n2596_), .Y(new_n2861_));
  OAI21X1  g00426(.A0(new_n2861_), .A1(new_n2588_), .B0(new_n2576_), .Y(new_n2862_));
  NAND2X1  g00427(.A(new_n2862_), .B(new_n2584_), .Y(new_n2863_));
  AOI21X1  g00428(.A0(new_n2863_), .A1(new_n2481_), .B0(new_n2574_), .Y(new_n2864_));
  OAI21X1  g00429(.A0(new_n2864_), .A1(new_n2818_), .B0(new_n2571_), .Y(new_n2865_));
  AOI21X1  g00430(.A0(new_n2865_), .A1(new_n2564_), .B0(new_n2858_), .Y(new_n2866_));
  OAI21X1  g00431(.A0(new_n2866_), .A1(pi0093), .B0(new_n2856_), .Y(new_n2867_));
  INVX1    g00432(.A(new_n2867_), .Y(new_n2868_));
  AND2X1   g00433(.A(new_n2555_), .B(pi0051), .Y(new_n2869_));
  AND2X1   g00434(.A(new_n2709_), .B(pi0070), .Y(new_n2870_));
  NOR3X1   g00435(.A(new_n2870_), .B(new_n2869_), .C(pi0096), .Y(new_n2871_));
  OAI21X1  g00436(.A0(new_n2868_), .A1(new_n2523_), .B0(new_n2871_), .Y(new_n2872_));
  AOI21X1  g00437(.A0(new_n2534_), .A1(pi0096), .B0(pi0072), .Y(new_n2873_));
  AOI21X1  g00438(.A0(new_n2873_), .A1(new_n2872_), .B0(new_n2554_), .Y(new_n2874_));
  NOR3X1   g00439(.A(new_n2874_), .B(new_n2778_), .C(new_n2547_), .Y(new_n2875_));
  OAI21X1  g00440(.A0(new_n2726_), .A1(new_n2517_), .B0(new_n2488_), .Y(new_n2876_));
  NAND2X1  g00441(.A(new_n2876_), .B(pi0032), .Y(new_n2877_));
  NAND2X1  g00442(.A(new_n2778_), .B(new_n2546_), .Y(new_n2878_));
  INVX1    g00443(.A(new_n2856_), .Y(new_n2879_));
  INVX1    g00444(.A(pi0097), .Y(new_n2880_));
  OAI21X1  g00445(.A0(new_n2860_), .A1(new_n2594_), .B0(new_n2880_), .Y(new_n2881_));
  AOI21X1  g00446(.A0(new_n2881_), .A1(new_n2576_), .B0(new_n2585_), .Y(new_n2882_));
  OAI21X1  g00447(.A0(new_n2882_), .A1(pi0109), .B0(new_n2575_), .Y(new_n2883_));
  AOI21X1  g00448(.A0(new_n2883_), .A1(new_n2573_), .B0(new_n2572_), .Y(new_n2884_));
  OAI21X1  g00449(.A0(new_n2884_), .A1(new_n2565_), .B0(new_n2857_), .Y(new_n2885_));
  AOI21X1  g00450(.A0(new_n2885_), .A1(new_n2531_), .B0(new_n2879_), .Y(new_n2886_));
  OAI21X1  g00451(.A0(new_n2886_), .A1(new_n2523_), .B0(new_n2871_), .Y(new_n2887_));
  AOI21X1  g00452(.A0(new_n2887_), .A1(new_n2873_), .B0(new_n2554_), .Y(new_n2888_));
  OAI21X1  g00453(.A0(new_n2888_), .A1(new_n2878_), .B0(new_n2877_), .Y(new_n2889_));
  OAI21X1  g00454(.A0(new_n2889_), .A1(new_n2875_), .B0(new_n2540_), .Y(new_n2890_));
  AOI21X1  g00455(.A0(new_n2890_), .A1(new_n2815_), .B0(pi0137), .Y(new_n2891_));
  AOI21X1  g00456(.A0(new_n2876_), .A1(pi0032), .B0(pi0095), .Y(new_n2892_));
  INVX1    g00457(.A(new_n2892_), .Y(new_n2893_));
  OR2X1    g00458(.A(pi0096), .B(pi0051), .Y(new_n2894_));
  NOR4X1   g00459(.A(new_n2894_), .B(new_n2870_), .C(new_n2522_), .D(new_n2458_), .Y(new_n2895_));
  NOR2X1   g00460(.A(new_n2895_), .B(pi0032), .Y(new_n2896_));
  NAND4X1  g00461(.A(new_n2715_), .B(new_n2534_), .C(pi0096), .D(new_n2548_), .Y(new_n2897_));
  AND2X1   g00462(.A(new_n2897_), .B(new_n2896_), .Y(new_n2898_));
  INVX1    g00463(.A(new_n2455_), .Y(new_n2899_));
  INVX1    g00464(.A(new_n2715_), .Y(new_n2900_));
  NOR4X1   g00465(.A(new_n2900_), .B(new_n2544_), .C(new_n2709_), .D(new_n2899_), .Y(new_n2901_));
  NOR2X1   g00466(.A(new_n2901_), .B(new_n2453_), .Y(new_n2902_));
  OAI21X1  g00467(.A0(new_n2898_), .A1(new_n2893_), .B0(new_n2902_), .Y(new_n2903_));
  INVX1    g00468(.A(new_n2903_), .Y(new_n2904_));
  OAI21X1  g00469(.A0(new_n2904_), .A1(new_n2891_), .B0(new_n2766_), .Y(new_n2905_));
  AOI21X1  g00470(.A0(new_n2488_), .A1(new_n2517_), .B0(new_n2456_), .Y(new_n2906_));
  INVX1    g00471(.A(new_n2906_), .Y(new_n2907_));
  OAI21X1  g00472(.A0(new_n2874_), .A1(new_n2547_), .B0(new_n2907_), .Y(new_n2908_));
  AOI21X1  g00473(.A0(new_n2908_), .A1(new_n2540_), .B0(new_n2850_), .Y(new_n2909_));
  NOR3X1   g00474(.A(new_n2906_), .B(new_n2898_), .C(pi0095), .Y(new_n2910_));
  OAI21X1  g00475(.A0(new_n2910_), .A1(new_n2901_), .B0(pi0137), .Y(new_n2911_));
  NAND2X1  g00476(.A(new_n2911_), .B(pi0210), .Y(new_n2912_));
  OAI21X1  g00477(.A0(new_n2912_), .A1(new_n2909_), .B0(new_n2810_), .Y(new_n2913_));
  NOR2X1   g00478(.A(pi0210), .B(pi0146), .Y(new_n2914_));
  OAI21X1  g00479(.A0(new_n2874_), .A1(new_n2547_), .B0(new_n2877_), .Y(new_n2915_));
  AOI21X1  g00480(.A0(new_n2915_), .A1(new_n2540_), .B0(new_n2716_), .Y(new_n2916_));
  OAI21X1  g00481(.A0(new_n2916_), .A1(pi0137), .B0(new_n2903_), .Y(new_n2917_));
  AOI21X1  g00482(.A0(new_n2917_), .A1(new_n2914_), .B0(new_n2913_), .Y(new_n2918_));
  OAI21X1  g00483(.A0(new_n2905_), .A1(new_n2800_), .B0(new_n2918_), .Y(new_n2919_));
  INVX1    g00484(.A(new_n2896_), .Y(new_n2920_));
  AOI21X1  g00485(.A0(new_n2920_), .A1(new_n2892_), .B0(new_n2453_), .Y(new_n2921_));
  AOI21X1  g00486(.A0(new_n2872_), .A1(new_n2548_), .B0(new_n2554_), .Y(new_n2922_));
  NOR3X1   g00487(.A(new_n2922_), .B(new_n2778_), .C(new_n2547_), .Y(new_n2923_));
  AOI21X1  g00488(.A0(new_n2887_), .A1(new_n2548_), .B0(new_n2554_), .Y(new_n2924_));
  OAI21X1  g00489(.A0(new_n2924_), .A1(new_n2878_), .B0(new_n2877_), .Y(new_n2925_));
  OAI21X1  g00490(.A0(new_n2925_), .A1(new_n2923_), .B0(new_n2540_), .Y(new_n2926_));
  AOI21X1  g00491(.A0(new_n2926_), .A1(new_n2772_), .B0(pi0137), .Y(new_n2927_));
  OAI21X1  g00492(.A0(new_n2927_), .A1(new_n2921_), .B0(new_n2766_), .Y(new_n2928_));
  INVX1    g00493(.A(new_n2772_), .Y(new_n2929_));
  OAI21X1  g00494(.A0(new_n2922_), .A1(new_n2547_), .B0(new_n2907_), .Y(new_n2930_));
  AND2X1   g00495(.A(new_n2930_), .B(new_n2540_), .Y(new_n2931_));
  NOR3X1   g00496(.A(new_n2931_), .B(new_n2929_), .C(pi0137), .Y(new_n2932_));
  OR4X1    g00497(.A(new_n2906_), .B(new_n2896_), .C(new_n2453_), .D(pi0095), .Y(new_n2933_));
  AND2X1   g00498(.A(new_n2933_), .B(pi0210), .Y(new_n2934_));
  INVX1    g00499(.A(new_n2934_), .Y(new_n2935_));
  OAI21X1  g00500(.A0(new_n2935_), .A1(new_n2932_), .B0(new_n2798_), .Y(new_n2936_));
  INVX1    g00501(.A(new_n2921_), .Y(new_n2937_));
  OAI21X1  g00502(.A0(new_n2922_), .A1(new_n2547_), .B0(new_n2877_), .Y(new_n2938_));
  AOI21X1  g00503(.A0(new_n2938_), .A1(new_n2540_), .B0(new_n2929_), .Y(new_n2939_));
  OAI21X1  g00504(.A0(new_n2939_), .A1(pi0137), .B0(new_n2937_), .Y(new_n2940_));
  AOI21X1  g00505(.A0(new_n2940_), .A1(new_n2914_), .B0(new_n2936_), .Y(new_n2941_));
  OAI21X1  g00506(.A0(new_n2928_), .A1(new_n2800_), .B0(new_n2941_), .Y(new_n2942_));
  NAND3X1  g00507(.A(new_n2942_), .B(new_n2919_), .C(new_n2452_), .Y(new_n2943_));
  OR2X1    g00508(.A(new_n2935_), .B(new_n2932_), .Y(new_n2944_));
  NAND3X1  g00509(.A(new_n2944_), .B(new_n2928_), .C(new_n2798_), .Y(new_n2945_));
  INVX1    g00510(.A(new_n2913_), .Y(new_n2946_));
  AOI21X1  g00511(.A0(new_n2946_), .A1(new_n2905_), .B0(new_n2452_), .Y(new_n2947_));
  AOI21X1  g00512(.A0(new_n2947_), .A1(new_n2945_), .B0(pi0153), .Y(new_n2948_));
  AOI21X1  g00513(.A0(new_n2948_), .A1(new_n2943_), .B0(pi0228), .Y(new_n2949_));
  AOI22X1  g00514(.A0(new_n2949_), .A1(new_n2854_), .B0(new_n2814_), .B1(pi0228), .Y(new_n2950_));
  OAI21X1  g00515(.A0(new_n2950_), .A1(pi0216), .B0(new_n2447_), .Y(new_n2951_));
  AOI21X1  g00516(.A0(new_n2951_), .A1(new_n2437_), .B0(new_n2444_), .Y(new_n2952_));
  INVX1    g00517(.A(pi0299), .Y(new_n2953_));
  INVX1    g00518(.A(pi0215), .Y(new_n2954_));
  NOR2X1   g00519(.A(pi1144), .B(pi0332), .Y(new_n2955_));
  NOR2X1   g00520(.A(new_n2955_), .B(new_n2954_), .Y(new_n2956_));
  NOR2X1   g00521(.A(new_n2956_), .B(new_n2953_), .Y(new_n2957_));
  OAI21X1  g00522(.A0(new_n2952_), .A1(pi0215), .B0(new_n2957_), .Y(new_n2958_));
  INVX1    g00523(.A(pi0039), .Y(new_n2959_));
  INVX1    g00524(.A(pi0222), .Y(new_n2960_));
  INVX1    g00525(.A(pi0224), .Y(new_n2961_));
  AOI21X1  g00526(.A0(pi0833), .A1(new_n2961_), .B0(new_n2960_), .Y(new_n2962_));
  OAI21X1  g00527(.A0(new_n2962_), .A1(pi0223), .B0(new_n2955_), .Y(new_n2963_));
  INVX1    g00528(.A(pi0223), .Y(new_n2964_));
  AOI21X1  g00529(.A0(new_n2445_), .A1(pi0265), .B0(new_n2961_), .Y(new_n2965_));
  NOR2X1   g00530(.A(new_n2965_), .B(pi0222), .Y(new_n2966_));
  NOR4X1   g00531(.A(pi0929), .B(new_n2721_), .C(pi0332), .D(pi0224), .Y(new_n2967_));
  OAI21X1  g00532(.A0(new_n2967_), .A1(new_n2966_), .B0(new_n2964_), .Y(new_n2968_));
  AOI21X1  g00533(.A0(new_n2968_), .A1(new_n2963_), .B0(pi0299), .Y(new_n2969_));
  NOR2X1   g00534(.A(pi0224), .B(pi0222), .Y(new_n2970_));
  INVX1    g00535(.A(new_n2970_), .Y(new_n2971_));
  INVX1    g00536(.A(pi0142), .Y(new_n2972_));
  INVX1    g00537(.A(pi0198), .Y(new_n2973_));
  OR2X1    g00538(.A(new_n2720_), .B(new_n2973_), .Y(new_n2974_));
  OAI21X1  g00539(.A0(new_n2764_), .A1(pi0198), .B0(new_n2974_), .Y(new_n2975_));
  OAI21X1  g00540(.A0(new_n2736_), .A1(new_n2732_), .B0(new_n2973_), .Y(new_n2976_));
  NAND3X1  g00541(.A(new_n2976_), .B(new_n2974_), .C(new_n2972_), .Y(new_n2977_));
  AND2X1   g00542(.A(new_n2977_), .B(new_n2798_), .Y(new_n2978_));
  OAI21X1  g00543(.A0(new_n2975_), .A1(new_n2972_), .B0(new_n2978_), .Y(new_n2979_));
  NOR3X1   g00544(.A(pi0189), .B(pi0174), .C(pi0144), .Y(new_n2980_));
  OR2X1    g00545(.A(new_n2980_), .B(pi0223), .Y(new_n2981_));
  NOR2X1   g00546(.A(new_n2793_), .B(new_n2791_), .Y(new_n2982_));
  MX2X1    g00547(.A(new_n2982_), .B(new_n2775_), .S0(pi0198), .Y(new_n2983_));
  NAND2X1  g00548(.A(new_n2983_), .B(pi0142), .Y(new_n2984_));
  AOI21X1  g00549(.A0(new_n2807_), .A1(new_n2973_), .B0(pi0142), .Y(new_n2985_));
  OAI21X1  g00550(.A0(new_n2775_), .A1(new_n2973_), .B0(new_n2985_), .Y(new_n2986_));
  AND2X1   g00551(.A(new_n2986_), .B(new_n2810_), .Y(new_n2987_));
  AOI21X1  g00552(.A0(new_n2987_), .A1(new_n2984_), .B0(new_n2981_), .Y(new_n2988_));
  NOR4X1   g00553(.A(pi0223), .B(pi0189), .C(pi0174), .D(pi0144), .Y(new_n2989_));
  INVX1    g00554(.A(pi0234), .Y(new_n2990_));
  AOI21X1  g00555(.A0(new_n2983_), .A1(new_n2990_), .B0(pi0332), .Y(new_n2991_));
  OAI21X1  g00556(.A0(new_n2975_), .A1(new_n2990_), .B0(new_n2991_), .Y(new_n2992_));
  AOI22X1  g00557(.A0(new_n2992_), .A1(new_n2989_), .B0(new_n2988_), .B1(new_n2979_), .Y(new_n2993_));
  OAI21X1  g00558(.A0(new_n2993_), .A1(new_n2971_), .B0(new_n2969_), .Y(new_n2994_));
  AND2X1   g00559(.A(new_n2994_), .B(new_n2959_), .Y(new_n2995_));
  INVX1    g00560(.A(pi0038), .Y(new_n2996_));
  AND2X1   g00561(.A(new_n2968_), .B(new_n2963_), .Y(new_n2997_));
  AOI21X1  g00562(.A0(new_n2455_), .A1(pi0234), .B0(pi0332), .Y(new_n2998_));
  INVX1    g00563(.A(new_n2998_), .Y(new_n2999_));
  NOR4X1   g00564(.A(new_n2900_), .B(new_n2544_), .C(new_n2709_), .D(pi0095), .Y(new_n3000_));
  OAI21X1  g00565(.A0(new_n3000_), .A1(new_n2455_), .B0(pi0234), .Y(new_n3001_));
  NOR4X1   g00566(.A(pi0095), .B(pi0072), .C(pi0040), .D(pi0032), .Y(new_n3002_));
  NAND3X1  g00567(.A(new_n3002_), .B(new_n2526_), .C(new_n2516_), .Y(new_n3003_));
  OR4X1    g00568(.A(new_n3003_), .B(new_n2709_), .C(pi0234), .D(pi0070), .Y(new_n3004_));
  AND2X1   g00569(.A(new_n3004_), .B(new_n3001_), .Y(new_n3005_));
  INVX1    g00570(.A(new_n3005_), .Y(new_n3006_));
  AOI21X1  g00571(.A0(new_n3006_), .A1(pi0137), .B0(new_n2999_), .Y(new_n3007_));
  NOR3X1   g00572(.A(pi0224), .B(pi0223), .C(pi0222), .Y(new_n3008_));
  INVX1    g00573(.A(new_n3008_), .Y(new_n3009_));
  NOR2X1   g00574(.A(new_n3009_), .B(new_n3007_), .Y(new_n3010_));
  NOR2X1   g00575(.A(new_n3010_), .B(new_n2997_), .Y(new_n3011_));
  INVX1    g00576(.A(new_n2444_), .Y(new_n3012_));
  INVX1    g00577(.A(pi0228), .Y(new_n3013_));
  MX2X1    g00578(.A(new_n3007_), .B(new_n2449_), .S0(new_n2448_), .Y(new_n3014_));
  INVX1    g00579(.A(new_n3000_), .Y(new_n3015_));
  NOR4X1   g00580(.A(new_n3015_), .B(pi0332), .C(pi0153), .D(pi0137), .Y(new_n3016_));
  NOR3X1   g00581(.A(new_n3003_), .B(new_n2555_), .C(new_n2453_), .Y(new_n3017_));
  OAI21X1  g00582(.A0(new_n3017_), .A1(new_n2450_), .B0(new_n3013_), .Y(new_n3018_));
  OAI22X1  g00583(.A0(new_n3018_), .A1(new_n3016_), .B0(new_n3014_), .B1(new_n3013_), .Y(new_n3019_));
  AOI21X1  g00584(.A0(new_n3019_), .A1(new_n2438_), .B0(new_n2446_), .Y(new_n3020_));
  OAI21X1  g00585(.A0(new_n3020_), .A1(pi0221), .B0(new_n3012_), .Y(new_n3021_));
  AOI21X1  g00586(.A0(new_n3021_), .A1(new_n2954_), .B0(new_n2956_), .Y(new_n3022_));
  MX2X1    g00587(.A(new_n3022_), .B(new_n3011_), .S0(new_n2953_), .Y(new_n3023_));
  OAI21X1  g00588(.A0(new_n3023_), .A1(new_n2959_), .B0(new_n2996_), .Y(new_n3024_));
  AOI21X1  g00589(.A0(new_n2995_), .A1(new_n2958_), .B0(new_n3024_), .Y(new_n3025_));
  INVX1    g00590(.A(pi0100), .Y(new_n3026_));
  OAI21X1  g00591(.A0(new_n3010_), .A1(new_n2997_), .B0(new_n2953_), .Y(new_n3027_));
  AND2X1   g00592(.A(pi0228), .B(pi0105), .Y(new_n3028_));
  AND2X1   g00593(.A(new_n3028_), .B(new_n2998_), .Y(new_n3029_));
  INVX1    g00594(.A(new_n3028_), .Y(new_n3030_));
  AOI21X1  g00595(.A0(new_n3030_), .A1(new_n2449_), .B0(pi0216), .Y(new_n3031_));
  INVX1    g00596(.A(new_n3031_), .Y(new_n3032_));
  OAI21X1  g00597(.A0(new_n3032_), .A1(new_n3029_), .B0(new_n2447_), .Y(new_n3033_));
  AOI21X1  g00598(.A0(new_n3033_), .A1(new_n2437_), .B0(new_n2444_), .Y(new_n3034_));
  MX2X1    g00599(.A(new_n3034_), .B(new_n2955_), .S0(pi0215), .Y(new_n3035_));
  INVX1    g00600(.A(new_n3035_), .Y(new_n3036_));
  OR2X1    g00601(.A(pi0221), .B(pi0215), .Y(new_n3037_));
  NOR3X1   g00602(.A(new_n3037_), .B(new_n3032_), .C(new_n3007_), .Y(new_n3038_));
  OAI21X1  g00603(.A0(new_n3038_), .A1(new_n3036_), .B0(pi0299), .Y(new_n3039_));
  AOI21X1  g00604(.A0(new_n3039_), .A1(new_n3027_), .B0(pi0039), .Y(new_n3040_));
  NOR2X1   g00605(.A(new_n3009_), .B(new_n2998_), .Y(new_n3041_));
  INVX1    g00606(.A(new_n3041_), .Y(new_n3042_));
  AOI22X1  g00607(.A0(new_n3042_), .A1(new_n2969_), .B0(new_n3035_), .B1(pi0299), .Y(new_n3043_));
  INVX1    g00608(.A(new_n3043_), .Y(new_n3044_));
  OAI21X1  g00609(.A0(new_n3044_), .A1(new_n2959_), .B0(pi0038), .Y(new_n3045_));
  OAI21X1  g00610(.A0(new_n3045_), .A1(new_n3040_), .B0(new_n3026_), .Y(new_n3046_));
  AOI21X1  g00611(.A0(new_n2450_), .A1(new_n2448_), .B0(new_n3013_), .Y(new_n3047_));
  AOI21X1  g00612(.A0(pi0234), .A1(pi0095), .B0(pi0137), .Y(new_n3048_));
  OAI21X1  g00613(.A0(new_n2830_), .A1(pi0210), .B0(new_n3048_), .Y(new_n3049_));
  AOI21X1  g00614(.A0(new_n3049_), .A1(new_n3006_), .B0(pi0332), .Y(new_n3050_));
  OAI21X1  g00615(.A0(new_n3050_), .A1(new_n2448_), .B0(new_n3047_), .Y(new_n3051_));
  INVX1    g00616(.A(new_n3016_), .Y(new_n3052_));
  INVX1    g00617(.A(pi0252), .Y(new_n3053_));
  OAI21X1  g00618(.A0(new_n2766_), .A1(pi0137), .B0(new_n3053_), .Y(new_n3054_));
  NOR4X1   g00619(.A(new_n3054_), .B(new_n3015_), .C(new_n2830_), .D(pi0332), .Y(new_n3055_));
  INVX1    g00620(.A(new_n2830_), .Y(new_n3056_));
  NOR4X1   g00621(.A(new_n3003_), .B(new_n3056_), .C(new_n2555_), .D(new_n2453_), .Y(new_n3057_));
  OR2X1    g00622(.A(new_n3057_), .B(new_n2450_), .Y(new_n3058_));
  AOI21X1  g00623(.A0(new_n3053_), .A1(pi0210), .B0(new_n2830_), .Y(new_n3059_));
  OAI22X1  g00624(.A0(new_n3059_), .A1(new_n3052_), .B0(new_n3058_), .B1(new_n3055_), .Y(new_n3060_));
  AOI21X1  g00625(.A0(new_n3060_), .A1(new_n3013_), .B0(pi0216), .Y(new_n3061_));
  AOI21X1  g00626(.A0(new_n3061_), .A1(new_n3051_), .B0(new_n2446_), .Y(new_n3062_));
  OAI21X1  g00627(.A0(new_n3062_), .A1(pi0221), .B0(new_n3012_), .Y(new_n3063_));
  AOI21X1  g00628(.A0(new_n3063_), .A1(new_n2954_), .B0(new_n2956_), .Y(new_n3064_));
  NOR2X1   g00629(.A(pi0039), .B(pi0038), .Y(new_n3065_));
  INVX1    g00630(.A(new_n3065_), .Y(new_n3066_));
  INVX1    g00631(.A(new_n2997_), .Y(new_n3067_));
  AOI21X1  g00632(.A0(new_n2973_), .A1(pi0142), .B0(pi0137), .Y(new_n3068_));
  OR2X1    g00633(.A(new_n3068_), .B(new_n3005_), .Y(new_n3069_));
  AOI21X1  g00634(.A0(new_n3069_), .A1(new_n2998_), .B0(new_n2981_), .Y(new_n3070_));
  NAND3X1  g00635(.A(pi0198), .B(new_n2453_), .C(new_n2540_), .Y(new_n3071_));
  OAI21X1  g00636(.A0(new_n3000_), .A1(new_n2455_), .B0(new_n3071_), .Y(new_n3072_));
  INVX1    g00637(.A(new_n2810_), .Y(new_n3073_));
  OR2X1    g00638(.A(new_n3003_), .B(new_n2555_), .Y(new_n3074_));
  AOI21X1  g00639(.A0(pi0198), .A1(new_n2453_), .B0(new_n3074_), .Y(new_n3075_));
  OAI21X1  g00640(.A0(new_n3075_), .A1(new_n3073_), .B0(new_n2989_), .Y(new_n3076_));
  AOI21X1  g00641(.A0(new_n3072_), .A1(new_n2798_), .B0(new_n3076_), .Y(new_n3077_));
  OAI21X1  g00642(.A0(new_n3077_), .A1(new_n3070_), .B0(new_n2970_), .Y(new_n3078_));
  AOI21X1  g00643(.A0(new_n3078_), .A1(new_n3067_), .B0(pi0299), .Y(new_n3079_));
  NOR2X1   g00644(.A(new_n3079_), .B(new_n3066_), .Y(new_n3080_));
  OAI21X1  g00645(.A0(new_n3064_), .A1(new_n2953_), .B0(new_n3080_), .Y(new_n3081_));
  AOI21X1  g00646(.A0(new_n3066_), .A1(new_n3044_), .B0(new_n3026_), .Y(new_n3082_));
  AOI21X1  g00647(.A0(new_n3082_), .A1(new_n3081_), .B0(pi0087), .Y(new_n3083_));
  OAI21X1  g00648(.A0(new_n3046_), .A1(new_n3025_), .B0(new_n3083_), .Y(new_n3084_));
  NOR3X1   g00649(.A(pi0100), .B(pi0039), .C(pi0038), .Y(new_n3085_));
  MX2X1    g00650(.A(new_n3044_), .B(new_n3023_), .S0(new_n3085_), .Y(new_n3086_));
  AOI21X1  g00651(.A0(new_n3086_), .A1(pi0087), .B0(pi0075), .Y(new_n3087_));
  AOI21X1  g00652(.A0(new_n3051_), .A1(new_n3031_), .B0(new_n2446_), .Y(new_n3088_));
  OAI21X1  g00653(.A0(new_n3088_), .A1(pi0221), .B0(new_n3012_), .Y(new_n3089_));
  AOI21X1  g00654(.A0(new_n3089_), .A1(new_n2954_), .B0(new_n2956_), .Y(new_n3090_));
  NOR4X1   g00655(.A(pi0100), .B(pi0087), .C(pi0039), .D(pi0038), .Y(new_n3091_));
  INVX1    g00656(.A(new_n3091_), .Y(new_n3092_));
  NOR2X1   g00657(.A(new_n3092_), .B(new_n3079_), .Y(new_n3093_));
  OAI21X1  g00658(.A0(new_n3090_), .A1(new_n2953_), .B0(new_n3093_), .Y(new_n3094_));
  INVX1    g00659(.A(pi0075), .Y(new_n3095_));
  AOI21X1  g00660(.A0(new_n3092_), .A1(new_n3044_), .B0(new_n3095_), .Y(new_n3096_));
  AOI22X1  g00661(.A0(new_n3096_), .A1(new_n3094_), .B0(new_n3087_), .B1(new_n3084_), .Y(new_n3097_));
  NOR2X1   g00662(.A(pi0087), .B(pi0075), .Y(new_n3098_));
  NAND2X1  g00663(.A(new_n3098_), .B(new_n3086_), .Y(new_n3099_));
  INVX1    g00664(.A(pi0092), .Y(new_n3100_));
  INVX1    g00665(.A(new_n3098_), .Y(new_n3101_));
  AOI21X1  g00666(.A0(new_n3101_), .A1(new_n3044_), .B0(new_n3100_), .Y(new_n3102_));
  AOI21X1  g00667(.A0(new_n3102_), .A1(new_n3099_), .B0(pi0054), .Y(new_n3103_));
  OAI21X1  g00668(.A0(new_n3097_), .A1(pi0092), .B0(new_n3103_), .Y(new_n3104_));
  NOR2X1   g00669(.A(pi0092), .B(pi0075), .Y(new_n3105_));
  AND2X1   g00670(.A(new_n3105_), .B(new_n3091_), .Y(new_n3106_));
  INVX1    g00671(.A(new_n3106_), .Y(new_n3107_));
  NOR3X1   g00672(.A(pi0100), .B(pi0087), .C(pi0038), .Y(new_n3108_));
  AND2X1   g00673(.A(new_n3108_), .B(new_n3105_), .Y(new_n3109_));
  AOI22X1  g00674(.A0(new_n3109_), .A1(new_n3040_), .B0(new_n3107_), .B1(new_n3043_), .Y(new_n3110_));
  AOI21X1  g00675(.A0(new_n3110_), .A1(pi0054), .B0(pi0074), .Y(new_n3111_));
  INVX1    g00676(.A(pi0054), .Y(new_n3112_));
  OAI21X1  g00677(.A0(new_n3043_), .A1(new_n3112_), .B0(pi0074), .Y(new_n3113_));
  AOI21X1  g00678(.A0(new_n3110_), .A1(new_n3112_), .B0(new_n3113_), .Y(new_n3114_));
  AOI21X1  g00679(.A0(new_n3111_), .A1(new_n3104_), .B0(new_n3114_), .Y(new_n3115_));
  INVX1    g00680(.A(new_n3047_), .Y(new_n3116_));
  NAND3X1  g00681(.A(new_n3004_), .B(new_n3001_), .C(new_n2445_), .Y(new_n3117_));
  AOI21X1  g00682(.A0(new_n3117_), .A1(pi0105), .B0(new_n3116_), .Y(new_n3118_));
  NAND3X1  g00683(.A(new_n3074_), .B(new_n2449_), .C(new_n3013_), .Y(new_n3119_));
  NAND2X1  g00684(.A(new_n3119_), .B(new_n2438_), .Y(new_n3120_));
  OAI21X1  g00685(.A0(new_n3120_), .A1(new_n3118_), .B0(new_n2447_), .Y(new_n3121_));
  AOI21X1  g00686(.A0(new_n3121_), .A1(new_n2437_), .B0(new_n2444_), .Y(new_n3122_));
  NOR2X1   g00687(.A(pi0100), .B(pi0087), .Y(new_n3123_));
  INVX1    g00688(.A(new_n3123_), .Y(new_n3124_));
  OR4X1    g00689(.A(pi0092), .B(pi0075), .C(pi0074), .D(pi0054), .Y(new_n3125_));
  NOR4X1   g00690(.A(new_n3125_), .B(new_n3124_), .C(new_n3066_), .D(new_n2956_), .Y(new_n3126_));
  OAI21X1  g00691(.A0(new_n3122_), .A1(pi0215), .B0(new_n3126_), .Y(new_n3127_));
  INVX1    g00692(.A(pi0055), .Y(new_n3128_));
  NOR3X1   g00693(.A(new_n3125_), .B(pi0100), .C(pi0087), .Y(new_n3129_));
  AND2X1   g00694(.A(new_n3129_), .B(new_n3065_), .Y(new_n3130_));
  INVX1    g00695(.A(new_n3130_), .Y(new_n3131_));
  AOI21X1  g00696(.A0(new_n3131_), .A1(new_n3035_), .B0(new_n3128_), .Y(new_n3132_));
  AOI21X1  g00697(.A0(new_n3132_), .A1(new_n3127_), .B0(pi0056), .Y(new_n3133_));
  OAI21X1  g00698(.A0(new_n3115_), .A1(pi0055), .B0(new_n3133_), .Y(new_n3134_));
  NOR2X1   g00699(.A(pi0074), .B(pi0054), .Y(new_n3135_));
  INVX1    g00700(.A(new_n3135_), .Y(new_n3136_));
  NOR3X1   g00701(.A(pi0100), .B(pi0039), .C(pi0038), .Y(new_n3137_));
  INVX1    g00702(.A(new_n3137_), .Y(new_n3138_));
  NAND2X1  g00703(.A(new_n3098_), .B(new_n3100_), .Y(new_n3139_));
  NOR4X1   g00704(.A(new_n3139_), .B(new_n3138_), .C(new_n3136_), .D(pi0055), .Y(new_n3140_));
  MX2X1    g00705(.A(new_n3035_), .B(new_n3022_), .S0(new_n3140_), .Y(new_n3141_));
  AOI21X1  g00706(.A0(new_n3141_), .A1(pi0056), .B0(pi0062), .Y(new_n3142_));
  INVX1    g00707(.A(pi0056), .Y(new_n3143_));
  OAI21X1  g00708(.A0(new_n3036_), .A1(new_n3143_), .B0(pi0062), .Y(new_n3144_));
  AOI21X1  g00709(.A0(new_n3141_), .A1(new_n3143_), .B0(new_n3144_), .Y(new_n3145_));
  OR2X1    g00710(.A(new_n3145_), .B(pi0059), .Y(new_n3146_));
  AOI21X1  g00711(.A0(new_n3142_), .A1(new_n3134_), .B0(new_n3146_), .Y(new_n3147_));
  NOR2X1   g00712(.A(pi0062), .B(pi0056), .Y(new_n3148_));
  NAND2X1  g00713(.A(new_n3148_), .B(new_n3140_), .Y(new_n3149_));
  NOR4X1   g00714(.A(new_n3149_), .B(new_n3037_), .C(new_n3032_), .D(new_n3007_), .Y(new_n3150_));
  NAND2X1  g00715(.A(new_n3035_), .B(pi0059), .Y(new_n3151_));
  OAI21X1  g00716(.A0(new_n3151_), .A1(new_n3150_), .B0(new_n2436_), .Y(new_n3152_));
  INVX1    g00717(.A(pi0059), .Y(new_n3153_));
  AOI21X1  g00718(.A0(new_n3150_), .A1(new_n3153_), .B0(new_n3036_), .Y(new_n3154_));
  OAI22X1  g00719(.A0(new_n3154_), .A1(new_n2436_), .B0(new_n3152_), .B1(new_n3147_), .Y(po0153));
  INVX1    g00720(.A(pi0087), .Y(new_n3156_));
  INVX1    g00721(.A(new_n3085_), .Y(new_n3157_));
  INVX1    g00722(.A(pi0154), .Y(new_n3158_));
  AND2X1   g00723(.A(pi0833), .B(new_n2961_), .Y(new_n3159_));
  INVX1    g00724(.A(pi0939), .Y(new_n3160_));
  AOI21X1  g00725(.A0(new_n3159_), .A1(new_n3160_), .B0(new_n2960_), .Y(new_n3161_));
  OAI21X1  g00726(.A0(new_n3159_), .A1(pi1146), .B0(new_n3161_), .Y(new_n3162_));
  AND2X1   g00727(.A(pi0224), .B(new_n2960_), .Y(new_n3163_));
  AOI21X1  g00728(.A0(new_n3163_), .A1(pi0276), .B0(pi0223), .Y(new_n3164_));
  INVX1    g00729(.A(pi1146), .Y(new_n3165_));
  AOI21X1  g00730(.A0(new_n3165_), .A1(pi0223), .B0(pi0299), .Y(new_n3166_));
  INVX1    g00731(.A(new_n3166_), .Y(new_n3167_));
  AOI21X1  g00732(.A0(new_n3164_), .A1(new_n3162_), .B0(new_n3167_), .Y(new_n3168_));
  INVX1    g00733(.A(new_n3168_), .Y(new_n3169_));
  AOI21X1  g00734(.A0(new_n2442_), .A1(new_n3160_), .B0(new_n2437_), .Y(new_n3170_));
  OAI21X1  g00735(.A0(new_n2442_), .A1(pi1146), .B0(new_n3170_), .Y(new_n3171_));
  OAI21X1  g00736(.A0(new_n3165_), .A1(new_n2954_), .B0(new_n3171_), .Y(new_n3172_));
  NOR4X1   g00737(.A(new_n3172_), .B(new_n3074_), .C(pi0228), .D(pi0216), .Y(new_n3173_));
  AND2X1   g00738(.A(pi1146), .B(pi0215), .Y(new_n3174_));
  INVX1    g00739(.A(pi0276), .Y(new_n3175_));
  NOR3X1   g00740(.A(new_n3175_), .B(pi0221), .C(new_n2438_), .Y(new_n3176_));
  AOI21X1  g00741(.A0(new_n3030_), .A1(new_n2438_), .B0(new_n3176_), .Y(new_n3177_));
  OAI21X1  g00742(.A0(new_n3177_), .A1(pi0221), .B0(new_n3171_), .Y(new_n3178_));
  AOI21X1  g00743(.A0(new_n3178_), .A1(new_n2954_), .B0(new_n3174_), .Y(new_n3179_));
  OR2X1    g00744(.A(new_n3179_), .B(new_n2953_), .Y(new_n3180_));
  OAI21X1  g00745(.A0(new_n3180_), .A1(new_n3173_), .B0(new_n3169_), .Y(new_n3181_));
  INVX1    g00746(.A(new_n3176_), .Y(new_n3182_));
  AOI21X1  g00747(.A0(new_n3182_), .A1(new_n3171_), .B0(pi0215), .Y(new_n3183_));
  NOR2X1   g00748(.A(new_n3183_), .B(new_n3174_), .Y(new_n3184_));
  OAI21X1  g00749(.A0(new_n3184_), .A1(new_n2953_), .B0(new_n3169_), .Y(new_n3185_));
  AND2X1   g00750(.A(new_n3185_), .B(pi0154), .Y(new_n3186_));
  OR2X1    g00751(.A(new_n3186_), .B(new_n3157_), .Y(new_n3187_));
  AOI21X1  g00752(.A0(new_n3181_), .A1(new_n3158_), .B0(new_n3187_), .Y(new_n3188_));
  MX2X1    g00753(.A(new_n3184_), .B(new_n3179_), .S0(new_n3158_), .Y(new_n3189_));
  INVX1    g00754(.A(new_n3189_), .Y(new_n3190_));
  AOI21X1  g00755(.A0(new_n3190_), .A1(pi0299), .B0(new_n3168_), .Y(new_n3191_));
  AOI21X1  g00756(.A0(new_n3191_), .A1(new_n3157_), .B0(new_n3188_), .Y(new_n3192_));
  AND2X1   g00757(.A(new_n3074_), .B(pi0039), .Y(new_n3193_));
  INVX1    g00758(.A(new_n2873_), .Y(new_n3194_));
  AOI22X1  g00759(.A0(new_n2709_), .A1(pi0070), .B0(new_n2514_), .B1(pi0035), .Y(new_n3195_));
  OAI21X1  g00760(.A0(new_n2822_), .A1(pi0070), .B0(new_n3195_), .Y(new_n3196_));
  AOI21X1  g00761(.A0(new_n3196_), .A1(new_n2516_), .B0(new_n2557_), .Y(new_n3197_));
  OAI21X1  g00762(.A0(new_n3197_), .A1(new_n3194_), .B0(new_n2552_), .Y(new_n3198_));
  NOR2X1   g00763(.A(new_n2545_), .B(new_n2549_), .Y(new_n3199_));
  NOR2X1   g00764(.A(new_n2488_), .B(new_n2456_), .Y(new_n3200_));
  NOR2X1   g00765(.A(new_n3200_), .B(new_n3199_), .Y(new_n3201_));
  INVX1    g00766(.A(new_n3201_), .Y(new_n3202_));
  AOI21X1  g00767(.A0(new_n3198_), .A1(new_n2715_), .B0(new_n3202_), .Y(new_n3203_));
  OAI21X1  g00768(.A0(new_n3203_), .A1(pi0095), .B0(new_n2815_), .Y(new_n3204_));
  AOI21X1  g00769(.A0(new_n3204_), .A1(new_n2959_), .B0(new_n3193_), .Y(new_n3205_));
  NOR3X1   g00770(.A(new_n3172_), .B(pi0228), .C(pi0216), .Y(new_n3206_));
  AOI21X1  g00771(.A0(new_n3206_), .A1(new_n3205_), .B0(new_n3180_), .Y(new_n3207_));
  OAI21X1  g00772(.A0(new_n3207_), .A1(new_n3168_), .B0(new_n3158_), .Y(new_n3208_));
  AOI21X1  g00773(.A0(new_n3185_), .A1(pi0154), .B0(pi0038), .Y(new_n3209_));
  INVX1    g00774(.A(new_n3191_), .Y(new_n3210_));
  OAI21X1  g00775(.A0(new_n3210_), .A1(new_n2996_), .B0(new_n3026_), .Y(new_n3211_));
  AOI21X1  g00776(.A0(new_n3209_), .A1(new_n3208_), .B0(new_n3211_), .Y(new_n3212_));
  AOI21X1  g00777(.A0(pi0252), .A1(pi0146), .B0(new_n3074_), .Y(new_n3213_));
  INVX1    g00778(.A(new_n3213_), .Y(new_n3214_));
  NOR2X1   g00779(.A(pi0166), .B(pi0161), .Y(new_n3215_));
  NOR3X1   g00780(.A(new_n3003_), .B(new_n2555_), .C(pi0252), .Y(new_n3216_));
  AOI21X1  g00781(.A0(new_n3215_), .A1(new_n3216_), .B0(pi0152), .Y(new_n3217_));
  OAI21X1  g00782(.A0(new_n3215_), .A1(new_n3214_), .B0(new_n3217_), .Y(new_n3218_));
  INVX1    g00783(.A(new_n3218_), .Y(new_n3219_));
  AOI21X1  g00784(.A0(new_n3214_), .A1(pi0152), .B0(new_n3219_), .Y(new_n3220_));
  INVX1    g00785(.A(new_n3220_), .Y(new_n3221_));
  NOR3X1   g00786(.A(pi0228), .B(pi0216), .C(pi0038), .Y(new_n3222_));
  NAND4X1  g00787(.A(new_n3222_), .B(pi0299), .C(new_n3158_), .D(new_n2959_), .Y(new_n3223_));
  NOR3X1   g00788(.A(new_n3223_), .B(new_n3221_), .C(new_n3172_), .Y(new_n3224_));
  OR2X1    g00789(.A(new_n3191_), .B(new_n3026_), .Y(new_n3225_));
  OAI21X1  g00790(.A0(new_n3225_), .A1(new_n3224_), .B0(new_n3156_), .Y(new_n3226_));
  OAI22X1  g00791(.A0(new_n3226_), .A1(new_n3212_), .B0(new_n3192_), .B1(new_n3156_), .Y(new_n3227_));
  OAI21X1  g00792(.A0(new_n3210_), .A1(new_n3095_), .B0(new_n3100_), .Y(new_n3228_));
  AOI21X1  g00793(.A0(new_n3227_), .A1(new_n3095_), .B0(new_n3228_), .Y(new_n3229_));
  AND2X1   g00794(.A(new_n3137_), .B(new_n3098_), .Y(new_n3230_));
  OAI21X1  g00795(.A0(new_n3230_), .A1(new_n3210_), .B0(pi0092), .Y(new_n3231_));
  AOI21X1  g00796(.A0(new_n3188_), .A1(new_n3098_), .B0(new_n3231_), .Y(new_n3232_));
  NOR3X1   g00797(.A(new_n3232_), .B(new_n3229_), .C(new_n3136_), .Y(new_n3233_));
  OAI21X1  g00798(.A0(new_n3210_), .A1(new_n3135_), .B0(new_n3128_), .Y(new_n3234_));
  OAI21X1  g00799(.A0(new_n3184_), .A1(new_n3158_), .B0(new_n3173_), .Y(new_n3235_));
  NOR2X1   g00800(.A(new_n3189_), .B(new_n3128_), .Y(new_n3236_));
  OAI21X1  g00801(.A0(new_n3235_), .A1(new_n3131_), .B0(new_n3236_), .Y(new_n3237_));
  AND2X1   g00802(.A(new_n3237_), .B(new_n3143_), .Y(new_n3238_));
  OAI21X1  g00803(.A0(new_n3234_), .A1(new_n3233_), .B0(new_n3238_), .Y(new_n3239_));
  NOR3X1   g00804(.A(new_n3189_), .B(new_n3131_), .C(pi0055), .Y(new_n3240_));
  NAND2X1  g00805(.A(new_n3240_), .B(new_n3235_), .Y(new_n3241_));
  INVX1    g00806(.A(new_n3140_), .Y(new_n3242_));
  AOI21X1  g00807(.A0(new_n3190_), .A1(new_n3242_), .B0(new_n3143_), .Y(new_n3243_));
  AOI21X1  g00808(.A0(new_n3243_), .A1(new_n3241_), .B0(pi0062), .Y(new_n3244_));
  INVX1    g00809(.A(pi0062), .Y(new_n3245_));
  NOR2X1   g00810(.A(pi0059), .B(pi0057), .Y(new_n3246_));
  NOR4X1   g00811(.A(new_n3139_), .B(new_n3136_), .C(pi0056), .D(pi0055), .Y(new_n3247_));
  AND2X1   g00812(.A(new_n3247_), .B(new_n3137_), .Y(new_n3248_));
  INVX1    g00813(.A(new_n3248_), .Y(new_n3249_));
  AOI22X1  g00814(.A0(new_n3249_), .A1(new_n3190_), .B0(new_n3240_), .B1(new_n3235_), .Y(new_n3250_));
  OAI21X1  g00815(.A0(new_n3250_), .A1(new_n3245_), .B0(new_n3246_), .Y(new_n3251_));
  AOI21X1  g00816(.A0(new_n3244_), .A1(new_n3239_), .B0(new_n3251_), .Y(new_n3252_));
  INVX1    g00817(.A(pi0239), .Y(new_n3253_));
  OAI21X1  g00818(.A0(new_n3246_), .A1(new_n3190_), .B0(new_n3253_), .Y(new_n3254_));
  INVX1    g00819(.A(new_n2563_), .Y(new_n3255_));
  INVX1    g00820(.A(new_n3002_), .Y(new_n3256_));
  NOR4X1   g00821(.A(new_n3256_), .B(new_n2533_), .C(new_n3255_), .D(new_n2526_), .Y(new_n3257_));
  NOR2X1   g00822(.A(new_n3257_), .B(new_n2455_), .Y(new_n3258_));
  INVX1    g00823(.A(new_n3258_), .Y(new_n3259_));
  AOI21X1  g00824(.A0(new_n3175_), .A1(pi0224), .B0(pi0222), .Y(new_n3260_));
  OAI21X1  g00825(.A0(new_n3259_), .A1(pi0224), .B0(new_n3260_), .Y(new_n3261_));
  AND2X1   g00826(.A(new_n3162_), .B(new_n2964_), .Y(new_n3262_));
  AOI22X1  g00827(.A0(new_n3262_), .A1(new_n3261_), .B0(new_n3165_), .B1(pi0223), .Y(new_n3263_));
  MX2X1    g00828(.A(new_n3197_), .B(new_n2551_), .S0(pi0072), .Y(new_n3264_));
  OAI21X1  g00829(.A0(new_n3264_), .A1(new_n2900_), .B0(new_n3201_), .Y(new_n3265_));
  AOI21X1  g00830(.A0(new_n3265_), .A1(new_n2540_), .B0(new_n2929_), .Y(new_n3266_));
  AOI22X1  g00831(.A0(new_n3266_), .A1(new_n3013_), .B0(new_n3258_), .B1(new_n3028_), .Y(new_n3267_));
  INVX1    g00832(.A(new_n3267_), .Y(new_n3268_));
  NOR3X1   g00833(.A(pi0221), .B(pi0216), .C(pi0215), .Y(new_n3269_));
  NOR2X1   g00834(.A(new_n3258_), .B(new_n2448_), .Y(new_n3270_));
  NOR2X1   g00835(.A(new_n3258_), .B(new_n2716_), .Y(new_n3271_));
  MX2X1    g00836(.A(new_n3271_), .B(new_n3270_), .S0(pi0228), .Y(new_n3272_));
  OAI21X1  g00837(.A0(new_n3272_), .A1(new_n3158_), .B0(new_n3269_), .Y(new_n3273_));
  AOI21X1  g00838(.A0(new_n3268_), .A1(new_n3158_), .B0(new_n3273_), .Y(new_n3274_));
  NAND2X1  g00839(.A(new_n3184_), .B(pi0299), .Y(new_n3275_));
  OAI22X1  g00840(.A0(new_n3275_), .A1(new_n3274_), .B0(new_n3263_), .B1(pi0299), .Y(new_n3276_));
  NOR2X1   g00841(.A(pi0100), .B(pi0038), .Y(new_n3277_));
  OR2X1    g00842(.A(new_n3179_), .B(pi0154), .Y(new_n3278_));
  INVX1    g00843(.A(new_n3184_), .Y(new_n3279_));
  NOR4X1   g00844(.A(pi0479), .B(new_n3013_), .C(new_n2448_), .D(new_n2540_), .Y(new_n3280_));
  AND2X1   g00845(.A(new_n3280_), .B(new_n3269_), .Y(new_n3281_));
  OAI21X1  g00846(.A0(new_n3281_), .A1(new_n3279_), .B0(new_n2954_), .Y(new_n3282_));
  OAI21X1  g00847(.A0(new_n3281_), .A1(new_n3279_), .B0(pi0154), .Y(new_n3283_));
  NAND3X1  g00848(.A(new_n3283_), .B(new_n3282_), .C(new_n3278_), .Y(new_n3284_));
  OR4X1    g00849(.A(pi0299), .B(pi0224), .C(pi0223), .D(pi0222), .Y(new_n3285_));
  NOR3X1   g00850(.A(new_n3285_), .B(pi0479), .C(new_n2540_), .Y(new_n3286_));
  OR2X1    g00851(.A(new_n3286_), .B(new_n3168_), .Y(new_n3287_));
  AOI21X1  g00852(.A0(new_n3284_), .A1(pi0299), .B0(new_n3287_), .Y(new_n3288_));
  NAND2X1  g00853(.A(new_n3283_), .B(new_n3173_), .Y(new_n3289_));
  AOI21X1  g00854(.A0(new_n3289_), .A1(new_n3284_), .B0(new_n2953_), .Y(new_n3290_));
  OAI21X1  g00855(.A0(new_n3290_), .A1(new_n3288_), .B0(pi0039), .Y(new_n3291_));
  NAND2X1  g00856(.A(new_n3291_), .B(new_n3277_), .Y(new_n3292_));
  AOI21X1  g00857(.A0(new_n3276_), .A1(new_n2959_), .B0(new_n3292_), .Y(new_n3293_));
  NOR4X1   g00858(.A(new_n3223_), .B(new_n3221_), .C(new_n3172_), .D(new_n3026_), .Y(new_n3294_));
  NOR3X1   g00859(.A(new_n3294_), .B(new_n3288_), .C(new_n3277_), .Y(new_n3295_));
  OAI21X1  g00860(.A0(new_n3295_), .A1(new_n3293_), .B0(new_n3156_), .Y(new_n3296_));
  OR2X1    g00861(.A(new_n3288_), .B(new_n3156_), .Y(new_n3297_));
  AOI21X1  g00862(.A0(new_n3290_), .A1(new_n3085_), .B0(new_n3297_), .Y(new_n3298_));
  NOR2X1   g00863(.A(new_n3298_), .B(pi0075), .Y(new_n3299_));
  AND2X1   g00864(.A(new_n3288_), .B(pi0075), .Y(new_n3300_));
  OR2X1    g00865(.A(new_n3300_), .B(pi0092), .Y(new_n3301_));
  AOI21X1  g00866(.A0(new_n3299_), .A1(new_n3296_), .B0(new_n3301_), .Y(new_n3302_));
  OR2X1    g00867(.A(new_n3288_), .B(new_n3100_), .Y(new_n3303_));
  AOI21X1  g00868(.A0(new_n3290_), .A1(new_n3230_), .B0(new_n3303_), .Y(new_n3304_));
  OR2X1    g00869(.A(new_n3304_), .B(new_n3136_), .Y(new_n3305_));
  AOI21X1  g00870(.A0(new_n3288_), .A1(new_n3136_), .B0(pi0055), .Y(new_n3306_));
  OAI21X1  g00871(.A0(new_n3305_), .A1(new_n3302_), .B0(new_n3306_), .Y(new_n3307_));
  NAND3X1  g00872(.A(new_n3283_), .B(new_n3173_), .C(new_n3130_), .Y(new_n3308_));
  NAND3X1  g00873(.A(new_n3308_), .B(new_n3284_), .C(pi0055), .Y(new_n3309_));
  NAND3X1  g00874(.A(new_n3309_), .B(new_n3307_), .C(new_n3143_), .Y(new_n3310_));
  NAND4X1  g00875(.A(new_n3289_), .B(new_n3284_), .C(new_n3130_), .D(new_n3128_), .Y(new_n3311_));
  AOI21X1  g00876(.A0(new_n3284_), .A1(new_n3242_), .B0(new_n3143_), .Y(new_n3312_));
  AOI21X1  g00877(.A0(new_n3312_), .A1(new_n3311_), .B0(pi0062), .Y(new_n3313_));
  NOR2X1   g00878(.A(new_n3311_), .B(pi0056), .Y(new_n3314_));
  AOI21X1  g00879(.A0(new_n3284_), .A1(new_n3249_), .B0(new_n3314_), .Y(new_n3315_));
  OAI21X1  g00880(.A0(new_n3315_), .A1(new_n3245_), .B0(new_n3246_), .Y(new_n3316_));
  AOI21X1  g00881(.A0(new_n3313_), .A1(new_n3310_), .B0(new_n3316_), .Y(new_n3317_));
  OAI21X1  g00882(.A0(new_n3284_), .A1(new_n3246_), .B0(pi0239), .Y(new_n3318_));
  OAI22X1  g00883(.A0(new_n3318_), .A1(new_n3317_), .B0(new_n3254_), .B1(new_n3252_), .Y(po0154));
  INVX1    g00884(.A(pi0927), .Y(new_n3320_));
  AOI21X1  g00885(.A0(new_n2442_), .A1(new_n3320_), .B0(new_n2437_), .Y(new_n3321_));
  OAI21X1  g00886(.A0(new_n2442_), .A1(pi1145), .B0(new_n3321_), .Y(new_n3322_));
  AOI21X1  g00887(.A0(pi0274), .A1(pi0216), .B0(pi0221), .Y(new_n3323_));
  INVX1    g00888(.A(new_n3323_), .Y(new_n3324_));
  INVX1    g00889(.A(pi0151), .Y(new_n3325_));
  INVX1    g00890(.A(new_n3272_), .Y(new_n3326_));
  OAI21X1  g00891(.A0(new_n3326_), .A1(new_n3325_), .B0(new_n2438_), .Y(new_n3327_));
  AOI21X1  g00892(.A0(new_n3267_), .A1(new_n3325_), .B0(new_n3327_), .Y(new_n3328_));
  OAI21X1  g00893(.A0(new_n3328_), .A1(new_n3324_), .B0(new_n3322_), .Y(new_n3329_));
  AND2X1   g00894(.A(pi1145), .B(pi0215), .Y(new_n3330_));
  OR2X1    g00895(.A(new_n3330_), .B(new_n2953_), .Y(new_n3331_));
  AOI21X1  g00896(.A0(new_n3329_), .A1(new_n2954_), .B0(new_n3331_), .Y(new_n3332_));
  AOI21X1  g00897(.A0(new_n3159_), .A1(new_n3320_), .B0(new_n2960_), .Y(new_n3333_));
  OAI21X1  g00898(.A0(new_n3159_), .A1(pi1145), .B0(new_n3333_), .Y(new_n3334_));
  AOI21X1  g00899(.A0(pi0274), .A1(pi0224), .B0(pi0222), .Y(new_n3335_));
  OAI21X1  g00900(.A0(new_n3259_), .A1(pi0224), .B0(new_n3335_), .Y(new_n3336_));
  AOI21X1  g00901(.A0(new_n3336_), .A1(new_n3334_), .B0(pi0223), .Y(new_n3337_));
  NAND2X1  g00902(.A(pi1145), .B(pi0223), .Y(new_n3338_));
  NAND2X1  g00903(.A(new_n3338_), .B(new_n2953_), .Y(new_n3339_));
  OAI21X1  g00904(.A0(new_n3339_), .A1(new_n3337_), .B0(new_n2959_), .Y(new_n3340_));
  INVX1    g00905(.A(new_n3334_), .Y(new_n3341_));
  NOR3X1   g00906(.A(pi0274), .B(new_n2961_), .C(pi0222), .Y(new_n3342_));
  OAI21X1  g00907(.A0(new_n3342_), .A1(new_n3341_), .B0(new_n2964_), .Y(new_n3343_));
  AOI21X1  g00908(.A0(new_n3343_), .A1(new_n3338_), .B0(pi0299), .Y(new_n3344_));
  NOR2X1   g00909(.A(new_n3344_), .B(new_n3286_), .Y(new_n3345_));
  INVX1    g00910(.A(pi1145), .Y(new_n3346_));
  INVX1    g00911(.A(new_n3322_), .Y(new_n3347_));
  AOI21X1  g00912(.A0(pi0228), .A1(pi0105), .B0(pi0151), .Y(new_n3348_));
  NOR2X1   g00913(.A(new_n3348_), .B(new_n3280_), .Y(new_n3349_));
  NOR4X1   g00914(.A(new_n3003_), .B(new_n2555_), .C(pi0228), .D(pi0151), .Y(new_n3350_));
  OAI21X1  g00915(.A0(new_n3350_), .A1(new_n3349_), .B0(new_n2438_), .Y(new_n3351_));
  AOI21X1  g00916(.A0(new_n3351_), .A1(new_n3323_), .B0(new_n3347_), .Y(new_n3352_));
  MX2X1    g00917(.A(new_n3352_), .B(new_n3346_), .S0(pi0215), .Y(new_n3353_));
  OAI21X1  g00918(.A0(new_n3353_), .A1(new_n2953_), .B0(new_n3345_), .Y(new_n3354_));
  AOI21X1  g00919(.A0(new_n3354_), .A1(pi0039), .B0(pi0038), .Y(new_n3355_));
  OAI21X1  g00920(.A0(new_n3340_), .A1(new_n3332_), .B0(new_n3355_), .Y(new_n3356_));
  OAI21X1  g00921(.A0(new_n3348_), .A1(pi0216), .B0(new_n3323_), .Y(new_n3357_));
  AOI21X1  g00922(.A0(new_n3357_), .A1(new_n3322_), .B0(pi0215), .Y(new_n3358_));
  NOR2X1   g00923(.A(new_n3358_), .B(new_n3330_), .Y(new_n3359_));
  INVX1    g00924(.A(pi0274), .Y(new_n3360_));
  NOR4X1   g00925(.A(new_n3037_), .B(new_n3030_), .C(pi0479), .D(new_n2540_), .Y(new_n3361_));
  OAI21X1  g00926(.A0(new_n3360_), .A1(new_n2438_), .B0(new_n3361_), .Y(new_n3362_));
  AND2X1   g00927(.A(new_n3362_), .B(new_n3359_), .Y(new_n3363_));
  OAI21X1  g00928(.A0(new_n3363_), .A1(new_n2953_), .B0(new_n3345_), .Y(new_n3364_));
  INVX1    g00929(.A(new_n3364_), .Y(new_n3365_));
  AOI21X1  g00930(.A0(new_n3365_), .A1(pi0038), .B0(pi0100), .Y(new_n3366_));
  AOI22X1  g00931(.A0(new_n3220_), .A1(new_n3013_), .B0(new_n3028_), .B1(new_n2899_), .Y(new_n3367_));
  AOI21X1  g00932(.A0(new_n3367_), .A1(new_n3325_), .B0(new_n3351_), .Y(new_n3368_));
  OAI21X1  g00933(.A0(new_n3368_), .A1(new_n3324_), .B0(new_n3322_), .Y(new_n3369_));
  AOI21X1  g00934(.A0(new_n3369_), .A1(new_n2954_), .B0(new_n3330_), .Y(new_n3370_));
  NOR3X1   g00935(.A(new_n3344_), .B(new_n3286_), .C(new_n3066_), .Y(new_n3371_));
  OAI21X1  g00936(.A0(new_n3370_), .A1(new_n2953_), .B0(new_n3371_), .Y(new_n3372_));
  AOI21X1  g00937(.A0(new_n3365_), .A1(new_n3066_), .B0(new_n3026_), .Y(new_n3373_));
  AOI22X1  g00938(.A0(new_n3373_), .A1(new_n3372_), .B0(new_n3366_), .B1(new_n3356_), .Y(new_n3374_));
  MX2X1    g00939(.A(new_n3364_), .B(new_n3354_), .S0(new_n3085_), .Y(new_n3375_));
  AOI21X1  g00940(.A0(new_n3375_), .A1(pi0087), .B0(pi0075), .Y(new_n3376_));
  OAI21X1  g00941(.A0(new_n3374_), .A1(pi0087), .B0(new_n3376_), .Y(new_n3377_));
  AOI21X1  g00942(.A0(new_n3365_), .A1(pi0075), .B0(pi0092), .Y(new_n3378_));
  NOR2X1   g00943(.A(new_n3375_), .B(new_n3101_), .Y(new_n3379_));
  OAI21X1  g00944(.A0(new_n3364_), .A1(new_n3098_), .B0(pi0092), .Y(new_n3380_));
  OAI21X1  g00945(.A0(new_n3380_), .A1(new_n3379_), .B0(new_n3135_), .Y(new_n3381_));
  AOI21X1  g00946(.A0(new_n3378_), .A1(new_n3377_), .B0(new_n3381_), .Y(new_n3382_));
  OAI21X1  g00947(.A0(new_n3364_), .A1(new_n3135_), .B0(new_n3128_), .Y(new_n3383_));
  NAND2X1  g00948(.A(new_n3353_), .B(new_n3130_), .Y(new_n3384_));
  AOI21X1  g00949(.A0(new_n3363_), .A1(new_n3131_), .B0(new_n3128_), .Y(new_n3385_));
  AOI21X1  g00950(.A0(new_n3385_), .A1(new_n3384_), .B0(pi0056), .Y(new_n3386_));
  OAI21X1  g00951(.A0(new_n3383_), .A1(new_n3382_), .B0(new_n3386_), .Y(new_n3387_));
  INVX1    g00952(.A(new_n3363_), .Y(new_n3388_));
  AOI21X1  g00953(.A0(new_n3388_), .A1(new_n3242_), .B0(new_n3143_), .Y(new_n3389_));
  OAI21X1  g00954(.A0(new_n3353_), .A1(new_n3242_), .B0(new_n3389_), .Y(new_n3390_));
  NAND3X1  g00955(.A(new_n3390_), .B(new_n3387_), .C(new_n3245_), .Y(new_n3391_));
  INVX1    g00956(.A(pi0235), .Y(new_n3392_));
  INVX1    g00957(.A(new_n3246_), .Y(new_n3393_));
  OAI21X1  g00958(.A0(new_n3388_), .A1(new_n3248_), .B0(pi0062), .Y(new_n3394_));
  AOI21X1  g00959(.A0(new_n3353_), .A1(new_n3248_), .B0(new_n3394_), .Y(new_n3395_));
  NOR3X1   g00960(.A(new_n3395_), .B(new_n3393_), .C(new_n3392_), .Y(new_n3396_));
  INVX1    g00961(.A(new_n3359_), .Y(new_n3397_));
  OAI21X1  g00962(.A0(new_n3346_), .A1(new_n2954_), .B0(new_n3322_), .Y(new_n3398_));
  NOR4X1   g00963(.A(new_n3398_), .B(new_n3074_), .C(pi0228), .D(pi0216), .Y(new_n3399_));
  INVX1    g00964(.A(new_n3399_), .Y(new_n3400_));
  NOR2X1   g00965(.A(new_n3359_), .B(new_n2953_), .Y(new_n3401_));
  OR2X1    g00966(.A(new_n3344_), .B(new_n3138_), .Y(new_n3402_));
  AOI21X1  g00967(.A0(new_n3401_), .A1(new_n3400_), .B0(new_n3402_), .Y(new_n3403_));
  NOR3X1   g00968(.A(new_n3401_), .B(new_n3344_), .C(new_n3085_), .Y(new_n3404_));
  OAI21X1  g00969(.A0(new_n3404_), .A1(new_n3403_), .B0(pi0087), .Y(new_n3405_));
  INVX1    g00970(.A(new_n3401_), .Y(new_n3406_));
  INVX1    g00971(.A(new_n3205_), .Y(new_n3407_));
  OR2X1    g00972(.A(new_n3026_), .B(pi0039), .Y(new_n3408_));
  OAI22X1  g00973(.A0(new_n3408_), .A1(new_n3221_), .B0(new_n3407_), .B1(pi0100), .Y(new_n3409_));
  NOR4X1   g00974(.A(new_n3398_), .B(pi0228), .C(pi0216), .D(pi0038), .Y(new_n3410_));
  AOI21X1  g00975(.A0(new_n3410_), .A1(new_n3409_), .B0(new_n3406_), .Y(new_n3411_));
  OR2X1    g00976(.A(new_n3344_), .B(pi0087), .Y(new_n3412_));
  OAI21X1  g00977(.A0(new_n3412_), .A1(new_n3411_), .B0(new_n3405_), .Y(new_n3413_));
  NOR2X1   g00978(.A(new_n3401_), .B(new_n3344_), .Y(new_n3414_));
  INVX1    g00979(.A(new_n3414_), .Y(new_n3415_));
  OAI21X1  g00980(.A0(new_n3415_), .A1(new_n3095_), .B0(new_n3100_), .Y(new_n3416_));
  AOI21X1  g00981(.A0(new_n3413_), .A1(new_n3095_), .B0(new_n3416_), .Y(new_n3417_));
  OAI21X1  g00982(.A0(new_n3415_), .A1(new_n3230_), .B0(pi0092), .Y(new_n3418_));
  AOI21X1  g00983(.A0(new_n3403_), .A1(new_n3098_), .B0(new_n3418_), .Y(new_n3419_));
  OR2X1    g00984(.A(new_n3419_), .B(new_n3136_), .Y(new_n3420_));
  AOI21X1  g00985(.A0(new_n3414_), .A1(new_n3136_), .B0(pi0055), .Y(new_n3421_));
  OAI21X1  g00986(.A0(new_n3420_), .A1(new_n3417_), .B0(new_n3421_), .Y(new_n3422_));
  NAND2X1  g00987(.A(new_n3399_), .B(new_n3130_), .Y(new_n3423_));
  NOR2X1   g00988(.A(new_n3359_), .B(new_n3128_), .Y(new_n3424_));
  AOI21X1  g00989(.A0(new_n3424_), .A1(new_n3423_), .B0(pi0056), .Y(new_n3425_));
  AOI21X1  g00990(.A0(new_n3399_), .A1(new_n3140_), .B0(new_n3359_), .Y(new_n3426_));
  OAI21X1  g00991(.A0(new_n3426_), .A1(new_n3143_), .B0(new_n3245_), .Y(new_n3427_));
  AOI21X1  g00992(.A0(new_n3425_), .A1(new_n3422_), .B0(new_n3427_), .Y(new_n3428_));
  NOR3X1   g00993(.A(new_n3400_), .B(new_n3242_), .C(pi0056), .Y(new_n3429_));
  OAI21X1  g00994(.A0(new_n3358_), .A1(new_n3330_), .B0(pi0062), .Y(new_n3430_));
  NOR3X1   g00995(.A(pi0235), .B(pi0059), .C(pi0057), .Y(new_n3431_));
  OAI21X1  g00996(.A0(new_n3430_), .A1(new_n3429_), .B0(new_n3431_), .Y(new_n3432_));
  OAI21X1  g00997(.A0(new_n3362_), .A1(new_n3392_), .B0(new_n3393_), .Y(new_n3433_));
  OAI22X1  g00998(.A0(new_n3433_), .A1(new_n3397_), .B0(new_n3432_), .B1(new_n3428_), .Y(new_n3434_));
  AOI21X1  g00999(.A0(new_n3396_), .A1(new_n3391_), .B0(new_n3434_), .Y(po0155));
  AND2X1   g01000(.A(pi1143), .B(pi0215), .Y(new_n3436_));
  OR2X1    g01001(.A(new_n3436_), .B(new_n2953_), .Y(new_n3437_));
  INVX1    g01002(.A(pi0944), .Y(new_n3438_));
  AOI21X1  g01003(.A0(new_n2442_), .A1(new_n3438_), .B0(new_n2437_), .Y(new_n3439_));
  OAI21X1  g01004(.A0(new_n2442_), .A1(pi1143), .B0(new_n3439_), .Y(new_n3440_));
  AOI21X1  g01005(.A0(pi0264), .A1(pi0216), .B0(pi0221), .Y(new_n3441_));
  INVX1    g01006(.A(new_n3441_), .Y(new_n3442_));
  NOR2X1   g01007(.A(new_n3266_), .B(pi0146), .Y(new_n3443_));
  AOI21X1  g01008(.A0(new_n3271_), .A1(pi0146), .B0(pi0284), .Y(new_n3444_));
  AND2X1   g01009(.A(pi0284), .B(pi0146), .Y(new_n3445_));
  AOI21X1  g01010(.A0(new_n3445_), .A1(new_n3204_), .B0(new_n3444_), .Y(new_n3446_));
  OAI21X1  g01011(.A0(new_n3446_), .A1(new_n3443_), .B0(new_n3013_), .Y(new_n3447_));
  INVX1    g01012(.A(pi0284), .Y(new_n3448_));
  AOI21X1  g01013(.A0(new_n2454_), .A1(pi0095), .B0(new_n3448_), .Y(new_n3449_));
  AOI21X1  g01014(.A0(pi0146), .A1(new_n2448_), .B0(new_n3013_), .Y(new_n3450_));
  OAI21X1  g01015(.A0(new_n3449_), .A1(new_n2448_), .B0(new_n3450_), .Y(new_n3451_));
  INVX1    g01016(.A(new_n3451_), .Y(new_n3452_));
  AOI21X1  g01017(.A0(new_n3259_), .A1(new_n3028_), .B0(new_n3452_), .Y(new_n3453_));
  AOI21X1  g01018(.A0(new_n3453_), .A1(new_n3447_), .B0(pi0216), .Y(new_n3454_));
  OAI21X1  g01019(.A0(new_n3454_), .A1(new_n3442_), .B0(new_n3440_), .Y(new_n3455_));
  AOI21X1  g01020(.A0(new_n3455_), .A1(new_n2954_), .B0(new_n3437_), .Y(new_n3456_));
  AOI21X1  g01021(.A0(pi1143), .A1(pi0223), .B0(pi0299), .Y(new_n3457_));
  INVX1    g01022(.A(new_n3457_), .Y(new_n3458_));
  AOI21X1  g01023(.A0(new_n3159_), .A1(new_n3438_), .B0(new_n2960_), .Y(new_n3459_));
  OAI21X1  g01024(.A0(new_n3159_), .A1(pi1143), .B0(new_n3459_), .Y(new_n3460_));
  AOI21X1  g01025(.A0(pi0264), .A1(pi0224), .B0(pi0222), .Y(new_n3461_));
  INVX1    g01026(.A(new_n3461_), .Y(new_n3462_));
  AOI21X1  g01027(.A0(new_n3258_), .A1(new_n3448_), .B0(pi0224), .Y(new_n3463_));
  OAI21X1  g01028(.A0(new_n3463_), .A1(new_n3462_), .B0(new_n3460_), .Y(new_n3464_));
  AOI21X1  g01029(.A0(new_n3461_), .A1(new_n3259_), .B0(new_n3464_), .Y(new_n3465_));
  OAI21X1  g01030(.A0(new_n3465_), .A1(pi0223), .B0(new_n3457_), .Y(new_n3466_));
  AND2X1   g01031(.A(new_n3466_), .B(new_n2959_), .Y(new_n3467_));
  OAI21X1  g01032(.A0(new_n3464_), .A1(new_n3458_), .B0(new_n3467_), .Y(new_n3468_));
  AND2X1   g01033(.A(pi1143), .B(pi0223), .Y(new_n3469_));
  AOI21X1  g01034(.A0(new_n3449_), .A1(new_n2961_), .B0(new_n3462_), .Y(new_n3470_));
  INVX1    g01035(.A(new_n3470_), .Y(new_n3471_));
  AOI21X1  g01036(.A0(new_n3471_), .A1(new_n3460_), .B0(pi0223), .Y(new_n3472_));
  OAI21X1  g01037(.A0(new_n3472_), .A1(new_n3469_), .B0(new_n2953_), .Y(new_n3473_));
  AOI21X1  g01038(.A0(new_n3008_), .A1(new_n2455_), .B0(new_n3473_), .Y(new_n3474_));
  INVX1    g01039(.A(new_n3474_), .Y(new_n3475_));
  MX2X1    g01040(.A(new_n3448_), .B(pi0146), .S0(new_n3074_), .Y(new_n3476_));
  NOR2X1   g01041(.A(new_n3476_), .B(pi0228), .Y(new_n3477_));
  INVX1    g01042(.A(new_n3477_), .Y(new_n3478_));
  INVX1    g01043(.A(new_n3280_), .Y(new_n3479_));
  AND2X1   g01044(.A(new_n3451_), .B(new_n3479_), .Y(new_n3480_));
  AOI21X1  g01045(.A0(new_n3480_), .A1(new_n3478_), .B0(pi0216), .Y(new_n3481_));
  OAI21X1  g01046(.A0(new_n3481_), .A1(new_n3442_), .B0(new_n3440_), .Y(new_n3482_));
  AOI21X1  g01047(.A0(new_n3482_), .A1(new_n2954_), .B0(new_n3436_), .Y(new_n3483_));
  OAI21X1  g01048(.A0(new_n3483_), .A1(new_n2953_), .B0(new_n3475_), .Y(new_n3484_));
  AOI21X1  g01049(.A0(new_n3484_), .A1(pi0039), .B0(pi0038), .Y(new_n3485_));
  OAI21X1  g01050(.A0(new_n3468_), .A1(new_n3456_), .B0(new_n3485_), .Y(new_n3486_));
  INVX1    g01051(.A(new_n3480_), .Y(new_n3487_));
  AOI21X1  g01052(.A0(new_n3013_), .A1(new_n2800_), .B0(new_n3487_), .Y(new_n3488_));
  OAI21X1  g01053(.A0(new_n3488_), .A1(pi0216), .B0(new_n3441_), .Y(new_n3489_));
  AOI21X1  g01054(.A0(new_n3489_), .A1(new_n3440_), .B0(pi0215), .Y(new_n3490_));
  NOR2X1   g01055(.A(new_n3490_), .B(new_n3436_), .Y(new_n3491_));
  INVX1    g01056(.A(new_n3491_), .Y(new_n3492_));
  AOI21X1  g01057(.A0(new_n3492_), .A1(pi0299), .B0(new_n3474_), .Y(new_n3493_));
  AOI21X1  g01058(.A0(new_n3493_), .A1(pi0038), .B0(pi0100), .Y(new_n3494_));
  INVX1    g01059(.A(pi1143), .Y(new_n3495_));
  INVX1    g01060(.A(new_n3440_), .Y(new_n3496_));
  INVX1    g01061(.A(new_n3216_), .Y(new_n3497_));
  OAI21X1  g01062(.A0(new_n2452_), .A1(new_n3053_), .B0(new_n3448_), .Y(new_n3498_));
  OAI21X1  g01063(.A0(new_n3498_), .A1(new_n3074_), .B0(new_n3013_), .Y(new_n3499_));
  AOI21X1  g01064(.A0(new_n3497_), .A1(pi0146), .B0(new_n3499_), .Y(new_n3500_));
  OAI21X1  g01065(.A0(new_n3500_), .A1(new_n3487_), .B0(new_n2438_), .Y(new_n3501_));
  AOI21X1  g01066(.A0(new_n3501_), .A1(new_n3441_), .B0(new_n3496_), .Y(new_n3502_));
  MX2X1    g01067(.A(new_n3502_), .B(new_n3495_), .S0(pi0215), .Y(new_n3503_));
  NOR2X1   g01068(.A(new_n3474_), .B(new_n3066_), .Y(new_n3504_));
  OAI21X1  g01069(.A0(new_n3503_), .A1(new_n2953_), .B0(new_n3504_), .Y(new_n3505_));
  AOI21X1  g01070(.A0(new_n3493_), .A1(new_n3066_), .B0(new_n3026_), .Y(new_n3506_));
  AOI22X1  g01071(.A0(new_n3506_), .A1(new_n3505_), .B0(new_n3494_), .B1(new_n3486_), .Y(new_n3507_));
  INVX1    g01072(.A(new_n3493_), .Y(new_n3508_));
  MX2X1    g01073(.A(new_n3508_), .B(new_n3484_), .S0(new_n3085_), .Y(new_n3509_));
  AOI21X1  g01074(.A0(new_n3509_), .A1(pi0087), .B0(pi0075), .Y(new_n3510_));
  OAI21X1  g01075(.A0(new_n3507_), .A1(pi0087), .B0(new_n3510_), .Y(new_n3511_));
  AOI21X1  g01076(.A0(new_n3493_), .A1(pi0075), .B0(pi0092), .Y(new_n3512_));
  NOR2X1   g01077(.A(new_n3509_), .B(new_n3101_), .Y(new_n3513_));
  OAI21X1  g01078(.A0(new_n3508_), .A1(new_n3098_), .B0(pi0092), .Y(new_n3514_));
  OAI21X1  g01079(.A0(new_n3514_), .A1(new_n3513_), .B0(new_n3135_), .Y(new_n3515_));
  AOI21X1  g01080(.A0(new_n3512_), .A1(new_n3511_), .B0(new_n3515_), .Y(new_n3516_));
  OAI21X1  g01081(.A0(new_n3508_), .A1(new_n3135_), .B0(new_n3128_), .Y(new_n3517_));
  NAND2X1  g01082(.A(new_n3483_), .B(new_n3130_), .Y(new_n3518_));
  AOI21X1  g01083(.A0(new_n3491_), .A1(new_n3131_), .B0(new_n3128_), .Y(new_n3519_));
  AOI21X1  g01084(.A0(new_n3519_), .A1(new_n3518_), .B0(pi0056), .Y(new_n3520_));
  OAI21X1  g01085(.A0(new_n3517_), .A1(new_n3516_), .B0(new_n3520_), .Y(new_n3521_));
  AOI21X1  g01086(.A0(new_n3492_), .A1(new_n3242_), .B0(new_n3143_), .Y(new_n3522_));
  OAI21X1  g01087(.A0(new_n3483_), .A1(new_n3242_), .B0(new_n3522_), .Y(new_n3523_));
  AND2X1   g01088(.A(new_n3523_), .B(new_n3245_), .Y(new_n3524_));
  OAI21X1  g01089(.A0(new_n3492_), .A1(new_n3248_), .B0(pi0062), .Y(new_n3525_));
  AOI21X1  g01090(.A0(new_n3483_), .A1(new_n3248_), .B0(new_n3525_), .Y(new_n3526_));
  OR4X1    g01091(.A(new_n3526_), .B(pi0238), .C(pi0059), .D(pi0057), .Y(new_n3527_));
  AOI21X1  g01092(.A0(new_n3524_), .A1(new_n3521_), .B0(new_n3527_), .Y(new_n3528_));
  INVX1    g01093(.A(new_n3467_), .Y(new_n3529_));
  OAI21X1  g01094(.A0(new_n3258_), .A1(new_n2448_), .B0(new_n3452_), .Y(new_n3530_));
  INVX1    g01095(.A(new_n3266_), .Y(new_n3531_));
  INVX1    g01096(.A(new_n3271_), .Y(new_n3532_));
  OAI21X1  g01097(.A0(new_n3532_), .A1(pi0146), .B0(pi0284), .Y(new_n3533_));
  AOI21X1  g01098(.A0(new_n3531_), .A1(pi0146), .B0(new_n3533_), .Y(new_n3534_));
  INVX1    g01099(.A(new_n3204_), .Y(new_n3535_));
  NOR3X1   g01100(.A(new_n3535_), .B(pi0284), .C(pi0146), .Y(new_n3536_));
  OAI21X1  g01101(.A0(new_n3536_), .A1(new_n3534_), .B0(new_n3013_), .Y(new_n3537_));
  AOI21X1  g01102(.A0(new_n3537_), .A1(new_n3530_), .B0(pi0216), .Y(new_n3538_));
  OAI21X1  g01103(.A0(new_n3538_), .A1(new_n3442_), .B0(new_n3440_), .Y(new_n3539_));
  AOI21X1  g01104(.A0(new_n3539_), .A1(new_n2954_), .B0(new_n3437_), .Y(new_n3540_));
  AOI21X1  g01105(.A0(new_n3478_), .A1(new_n3451_), .B0(pi0216), .Y(new_n3541_));
  OAI21X1  g01106(.A0(new_n3541_), .A1(new_n3442_), .B0(new_n3440_), .Y(new_n3542_));
  AOI21X1  g01107(.A0(new_n3542_), .A1(new_n2954_), .B0(new_n3436_), .Y(new_n3543_));
  OAI21X1  g01108(.A0(new_n3543_), .A1(new_n2953_), .B0(new_n3473_), .Y(new_n3544_));
  AOI21X1  g01109(.A0(new_n3544_), .A1(pi0039), .B0(pi0038), .Y(new_n3545_));
  OAI21X1  g01110(.A0(new_n3540_), .A1(new_n3529_), .B0(new_n3545_), .Y(new_n3546_));
  INVX1    g01111(.A(new_n3473_), .Y(new_n3547_));
  INVX1    g01112(.A(new_n3361_), .Y(new_n3548_));
  AOI21X1  g01113(.A0(pi0264), .A1(pi0216), .B0(new_n3548_), .Y(new_n3549_));
  NOR3X1   g01114(.A(new_n3549_), .B(new_n3490_), .C(new_n3436_), .Y(new_n3550_));
  INVX1    g01115(.A(new_n3550_), .Y(new_n3551_));
  AOI21X1  g01116(.A0(new_n3551_), .A1(pi0299), .B0(new_n3547_), .Y(new_n3552_));
  AOI21X1  g01117(.A0(new_n3552_), .A1(pi0038), .B0(pi0100), .Y(new_n3553_));
  OAI21X1  g01118(.A0(new_n3500_), .A1(new_n3452_), .B0(new_n2438_), .Y(new_n3554_));
  AOI21X1  g01119(.A0(new_n3554_), .A1(new_n3441_), .B0(new_n3496_), .Y(new_n3555_));
  MX2X1    g01120(.A(new_n3555_), .B(new_n3495_), .S0(pi0215), .Y(new_n3556_));
  AND2X1   g01121(.A(new_n3473_), .B(new_n3065_), .Y(new_n3557_));
  OAI21X1  g01122(.A0(new_n3556_), .A1(new_n2953_), .B0(new_n3557_), .Y(new_n3558_));
  AOI21X1  g01123(.A0(new_n3552_), .A1(new_n3066_), .B0(new_n3026_), .Y(new_n3559_));
  AOI22X1  g01124(.A0(new_n3559_), .A1(new_n3558_), .B0(new_n3553_), .B1(new_n3546_), .Y(new_n3560_));
  INVX1    g01125(.A(new_n3552_), .Y(new_n3561_));
  MX2X1    g01126(.A(new_n3561_), .B(new_n3544_), .S0(new_n3085_), .Y(new_n3562_));
  AOI21X1  g01127(.A0(new_n3562_), .A1(pi0087), .B0(pi0075), .Y(new_n3563_));
  OAI21X1  g01128(.A0(new_n3560_), .A1(pi0087), .B0(new_n3563_), .Y(new_n3564_));
  AOI21X1  g01129(.A0(new_n3552_), .A1(pi0075), .B0(pi0092), .Y(new_n3565_));
  NOR2X1   g01130(.A(new_n3562_), .B(new_n3101_), .Y(new_n3566_));
  OAI21X1  g01131(.A0(new_n3561_), .A1(new_n3098_), .B0(pi0092), .Y(new_n3567_));
  OAI21X1  g01132(.A0(new_n3567_), .A1(new_n3566_), .B0(new_n3135_), .Y(new_n3568_));
  AOI21X1  g01133(.A0(new_n3565_), .A1(new_n3564_), .B0(new_n3568_), .Y(new_n3569_));
  OAI21X1  g01134(.A0(new_n3561_), .A1(new_n3135_), .B0(new_n3128_), .Y(new_n3570_));
  NAND2X1  g01135(.A(new_n3543_), .B(new_n3130_), .Y(new_n3571_));
  AOI21X1  g01136(.A0(new_n3550_), .A1(new_n3131_), .B0(new_n3128_), .Y(new_n3572_));
  AOI21X1  g01137(.A0(new_n3572_), .A1(new_n3571_), .B0(pi0056), .Y(new_n3573_));
  OAI21X1  g01138(.A0(new_n3570_), .A1(new_n3569_), .B0(new_n3573_), .Y(new_n3574_));
  AOI21X1  g01139(.A0(new_n3551_), .A1(new_n3242_), .B0(new_n3143_), .Y(new_n3575_));
  OAI21X1  g01140(.A0(new_n3543_), .A1(new_n3242_), .B0(new_n3575_), .Y(new_n3576_));
  AND2X1   g01141(.A(new_n3576_), .B(new_n3245_), .Y(new_n3577_));
  INVX1    g01142(.A(pi0238), .Y(new_n3578_));
  OAI21X1  g01143(.A0(new_n3551_), .A1(new_n3248_), .B0(pi0062), .Y(new_n3579_));
  AOI21X1  g01144(.A0(new_n3543_), .A1(new_n3248_), .B0(new_n3579_), .Y(new_n3580_));
  OR4X1    g01145(.A(new_n3580_), .B(new_n3578_), .C(pi0059), .D(pi0057), .Y(new_n3581_));
  AOI21X1  g01146(.A0(new_n3577_), .A1(new_n3574_), .B0(new_n3581_), .Y(new_n3582_));
  AND2X1   g01147(.A(new_n3549_), .B(pi0238), .Y(new_n3583_));
  NOR4X1   g01148(.A(new_n3583_), .B(new_n3490_), .C(new_n3436_), .D(new_n3246_), .Y(new_n3584_));
  NOR3X1   g01149(.A(new_n3584_), .B(new_n3582_), .C(new_n3528_), .Y(po0156));
  AND2X1   g01150(.A(pi1142), .B(pi0215), .Y(new_n3586_));
  NOR2X1   g01151(.A(new_n3586_), .B(new_n2953_), .Y(new_n3587_));
  INVX1    g01152(.A(pi0932), .Y(new_n3588_));
  AOI21X1  g01153(.A0(new_n2442_), .A1(new_n3588_), .B0(new_n2437_), .Y(new_n3589_));
  OAI21X1  g01154(.A0(new_n2442_), .A1(pi1142), .B0(new_n3589_), .Y(new_n3590_));
  INVX1    g01155(.A(new_n3590_), .Y(new_n3591_));
  AOI21X1  g01156(.A0(pi0277), .A1(pi0216), .B0(pi0221), .Y(new_n3592_));
  INVX1    g01157(.A(pi0262), .Y(new_n3593_));
  AOI21X1  g01158(.A0(new_n3271_), .A1(new_n3593_), .B0(pi0172), .Y(new_n3594_));
  AND2X1   g01159(.A(new_n3593_), .B(pi0172), .Y(new_n3595_));
  AOI21X1  g01160(.A0(new_n3595_), .A1(new_n3266_), .B0(new_n3594_), .Y(new_n3596_));
  OAI21X1  g01161(.A0(new_n3204_), .A1(new_n3593_), .B0(new_n3013_), .Y(new_n3597_));
  INVX1    g01162(.A(new_n3257_), .Y(new_n3598_));
  AOI21X1  g01163(.A0(new_n2454_), .A1(pi0095), .B0(new_n3593_), .Y(new_n3599_));
  AND2X1   g01164(.A(new_n3599_), .B(pi0105), .Y(new_n3600_));
  INVX1    g01165(.A(pi0172), .Y(new_n3601_));
  OAI21X1  g01166(.A0(new_n3601_), .A1(pi0105), .B0(pi0228), .Y(new_n3602_));
  AOI21X1  g01167(.A0(new_n3600_), .A1(new_n3598_), .B0(new_n3602_), .Y(new_n3603_));
  OAI21X1  g01168(.A0(new_n3258_), .A1(new_n2448_), .B0(new_n3603_), .Y(new_n3604_));
  AND2X1   g01169(.A(new_n3604_), .B(new_n2438_), .Y(new_n3605_));
  OAI21X1  g01170(.A0(new_n3597_), .A1(new_n3596_), .B0(new_n3605_), .Y(new_n3606_));
  AOI21X1  g01171(.A0(new_n3606_), .A1(new_n3592_), .B0(new_n3591_), .Y(new_n3607_));
  OAI21X1  g01172(.A0(new_n3607_), .A1(pi0215), .B0(new_n3587_), .Y(new_n3608_));
  AOI21X1  g01173(.A0(pi1142), .A1(pi0223), .B0(pi0299), .Y(new_n3609_));
  INVX1    g01174(.A(new_n3609_), .Y(new_n3610_));
  AOI21X1  g01175(.A0(new_n3159_), .A1(new_n3588_), .B0(new_n2960_), .Y(new_n3611_));
  OAI21X1  g01176(.A0(new_n3159_), .A1(pi1142), .B0(new_n3611_), .Y(new_n3612_));
  AOI21X1  g01177(.A0(pi0277), .A1(pi0224), .B0(pi0222), .Y(new_n3613_));
  INVX1    g01178(.A(new_n3613_), .Y(new_n3614_));
  AOI21X1  g01179(.A0(new_n3258_), .A1(new_n3593_), .B0(pi0224), .Y(new_n3615_));
  OAI21X1  g01180(.A0(new_n3615_), .A1(new_n3614_), .B0(new_n3612_), .Y(new_n3616_));
  OR2X1    g01181(.A(new_n3616_), .B(new_n3610_), .Y(new_n3617_));
  NOR2X1   g01182(.A(new_n3614_), .B(new_n3258_), .Y(new_n3618_));
  OAI21X1  g01183(.A0(new_n3618_), .A1(new_n3616_), .B0(new_n2964_), .Y(new_n3619_));
  AOI21X1  g01184(.A0(new_n3619_), .A1(new_n3609_), .B0(pi0039), .Y(new_n3620_));
  NAND3X1  g01185(.A(new_n3620_), .B(new_n3617_), .C(new_n3608_), .Y(new_n3621_));
  AND2X1   g01186(.A(pi1142), .B(pi0223), .Y(new_n3622_));
  AOI21X1  g01187(.A0(new_n3599_), .A1(new_n2961_), .B0(new_n3614_), .Y(new_n3623_));
  INVX1    g01188(.A(new_n3623_), .Y(new_n3624_));
  AOI21X1  g01189(.A0(new_n3624_), .A1(new_n3612_), .B0(pi0223), .Y(new_n3625_));
  OAI21X1  g01190(.A0(new_n3625_), .A1(new_n3622_), .B0(new_n2953_), .Y(new_n3626_));
  AOI21X1  g01191(.A0(new_n3008_), .A1(new_n2455_), .B0(new_n3626_), .Y(new_n3627_));
  INVX1    g01192(.A(new_n3627_), .Y(new_n3628_));
  INVX1    g01193(.A(new_n3592_), .Y(new_n3629_));
  INVX1    g01194(.A(new_n3074_), .Y(new_n3630_));
  NOR3X1   g01195(.A(new_n3003_), .B(new_n2555_), .C(pi0228), .Y(new_n3631_));
  INVX1    g01196(.A(new_n3631_), .Y(new_n3632_));
  AND2X1   g01197(.A(new_n3013_), .B(pi0172), .Y(new_n3633_));
  INVX1    g01198(.A(new_n3633_), .Y(new_n3634_));
  AOI22X1  g01199(.A0(new_n3634_), .A1(new_n3632_), .B0(new_n3630_), .B1(new_n3593_), .Y(new_n3635_));
  INVX1    g01200(.A(new_n3635_), .Y(new_n3636_));
  AND2X1   g01201(.A(pi0172), .B(new_n2448_), .Y(new_n3637_));
  OAI21X1  g01202(.A0(new_n3637_), .A1(new_n3600_), .B0(pi0228), .Y(new_n3638_));
  AND2X1   g01203(.A(new_n3638_), .B(new_n3479_), .Y(new_n3639_));
  AOI21X1  g01204(.A0(new_n3639_), .A1(new_n3636_), .B0(pi0216), .Y(new_n3640_));
  OAI21X1  g01205(.A0(new_n3640_), .A1(new_n3629_), .B0(new_n3590_), .Y(new_n3641_));
  AOI21X1  g01206(.A0(new_n3641_), .A1(new_n2954_), .B0(new_n3586_), .Y(new_n3642_));
  OAI21X1  g01207(.A0(new_n3642_), .A1(new_n2953_), .B0(new_n3628_), .Y(new_n3643_));
  AOI21X1  g01208(.A0(new_n3643_), .A1(pi0039), .B0(pi0038), .Y(new_n3644_));
  AOI21X1  g01209(.A0(new_n3638_), .A1(new_n3634_), .B0(pi0216), .Y(new_n3645_));
  OAI21X1  g01210(.A0(new_n3645_), .A1(new_n3629_), .B0(new_n3590_), .Y(new_n3646_));
  AOI21X1  g01211(.A0(new_n3646_), .A1(new_n2954_), .B0(new_n3586_), .Y(new_n3647_));
  NOR2X1   g01212(.A(new_n3647_), .B(new_n3281_), .Y(new_n3648_));
  AOI21X1  g01213(.A0(new_n3648_), .A1(pi0299), .B0(new_n3627_), .Y(new_n3649_));
  INVX1    g01214(.A(new_n3649_), .Y(new_n3650_));
  OAI21X1  g01215(.A0(new_n3650_), .A1(new_n2996_), .B0(new_n3026_), .Y(new_n3651_));
  AOI21X1  g01216(.A0(new_n3644_), .A1(new_n3621_), .B0(new_n3651_), .Y(new_n3652_));
  INVX1    g01217(.A(new_n3638_), .Y(new_n3653_));
  AND2X1   g01218(.A(new_n3220_), .B(new_n3013_), .Y(new_n3654_));
  INVX1    g01219(.A(new_n3654_), .Y(new_n3655_));
  AOI22X1  g01220(.A0(new_n3634_), .A1(new_n3655_), .B0(new_n3220_), .B1(new_n3593_), .Y(new_n3656_));
  NOR3X1   g01221(.A(new_n3656_), .B(new_n3653_), .C(new_n3280_), .Y(new_n3657_));
  OAI21X1  g01222(.A0(new_n3657_), .A1(pi0216), .B0(new_n3592_), .Y(new_n3658_));
  AOI21X1  g01223(.A0(new_n3658_), .A1(new_n3590_), .B0(pi0215), .Y(new_n3659_));
  OAI21X1  g01224(.A0(new_n3659_), .A1(new_n3586_), .B0(pi0299), .Y(new_n3660_));
  NOR2X1   g01225(.A(new_n3627_), .B(new_n3066_), .Y(new_n3661_));
  OAI21X1  g01226(.A0(new_n3650_), .A1(new_n3065_), .B0(pi0100), .Y(new_n3662_));
  AOI21X1  g01227(.A0(new_n3661_), .A1(new_n3660_), .B0(new_n3662_), .Y(new_n3663_));
  OAI21X1  g01228(.A0(new_n3663_), .A1(new_n3652_), .B0(new_n3156_), .Y(new_n3664_));
  MX2X1    g01229(.A(new_n3650_), .B(new_n3643_), .S0(new_n3085_), .Y(new_n3665_));
  AOI21X1  g01230(.A0(new_n3665_), .A1(pi0087), .B0(pi0075), .Y(new_n3666_));
  OAI21X1  g01231(.A0(new_n3650_), .A1(new_n3095_), .B0(new_n3100_), .Y(new_n3667_));
  AOI21X1  g01232(.A0(new_n3666_), .A1(new_n3664_), .B0(new_n3667_), .Y(new_n3668_));
  NOR2X1   g01233(.A(new_n3665_), .B(new_n3101_), .Y(new_n3669_));
  OAI21X1  g01234(.A0(new_n3650_), .A1(new_n3098_), .B0(pi0092), .Y(new_n3670_));
  OAI21X1  g01235(.A0(new_n3670_), .A1(new_n3669_), .B0(new_n3135_), .Y(new_n3671_));
  AOI21X1  g01236(.A0(new_n3649_), .A1(new_n3136_), .B0(pi0055), .Y(new_n3672_));
  OAI21X1  g01237(.A0(new_n3671_), .A1(new_n3668_), .B0(new_n3672_), .Y(new_n3673_));
  NAND2X1  g01238(.A(new_n3642_), .B(new_n3130_), .Y(new_n3674_));
  INVX1    g01239(.A(new_n3648_), .Y(new_n3675_));
  AOI21X1  g01240(.A0(new_n3675_), .A1(new_n3131_), .B0(new_n3128_), .Y(new_n3676_));
  AOI21X1  g01241(.A0(new_n3676_), .A1(new_n3674_), .B0(pi0056), .Y(new_n3677_));
  AOI21X1  g01242(.A0(new_n3648_), .A1(new_n3242_), .B0(new_n3143_), .Y(new_n3678_));
  OAI21X1  g01243(.A0(new_n3642_), .A1(new_n3242_), .B0(new_n3678_), .Y(new_n3679_));
  NAND2X1  g01244(.A(new_n3679_), .B(new_n3245_), .Y(new_n3680_));
  AOI21X1  g01245(.A0(new_n3677_), .A1(new_n3673_), .B0(new_n3680_), .Y(new_n3681_));
  OAI21X1  g01246(.A0(new_n3648_), .A1(new_n3248_), .B0(pi0062), .Y(new_n3682_));
  AOI21X1  g01247(.A0(new_n3642_), .A1(new_n3248_), .B0(new_n3682_), .Y(new_n3683_));
  OR2X1    g01248(.A(new_n3683_), .B(new_n3393_), .Y(new_n3684_));
  AOI21X1  g01249(.A0(new_n3675_), .A1(new_n3393_), .B0(pi0249), .Y(new_n3685_));
  OAI21X1  g01250(.A0(new_n3684_), .A1(new_n3681_), .B0(new_n3685_), .Y(new_n3686_));
  INVX1    g01251(.A(new_n3620_), .Y(new_n3687_));
  INVX1    g01252(.A(new_n3587_), .Y(new_n3688_));
  OAI21X1  g01253(.A0(new_n3531_), .A1(new_n3593_), .B0(new_n3601_), .Y(new_n3689_));
  AOI21X1  g01254(.A0(new_n3532_), .A1(pi0262), .B0(new_n3601_), .Y(new_n3690_));
  OAI21X1  g01255(.A0(new_n3535_), .A1(pi0262), .B0(new_n3690_), .Y(new_n3691_));
  AOI21X1  g01256(.A0(new_n3691_), .A1(new_n3689_), .B0(pi0228), .Y(new_n3692_));
  NOR3X1   g01257(.A(new_n3692_), .B(new_n3603_), .C(pi0216), .Y(new_n3693_));
  OAI21X1  g01258(.A0(new_n3693_), .A1(new_n3629_), .B0(new_n3590_), .Y(new_n3694_));
  AOI21X1  g01259(.A0(new_n3694_), .A1(new_n2954_), .B0(new_n3688_), .Y(new_n3695_));
  AOI21X1  g01260(.A0(new_n3638_), .A1(new_n3636_), .B0(pi0216), .Y(new_n3696_));
  OAI21X1  g01261(.A0(new_n3696_), .A1(new_n3629_), .B0(new_n3590_), .Y(new_n3697_));
  AOI21X1  g01262(.A0(new_n3697_), .A1(new_n2954_), .B0(new_n3586_), .Y(new_n3698_));
  OAI21X1  g01263(.A0(new_n3698_), .A1(new_n2953_), .B0(new_n3626_), .Y(new_n3699_));
  AOI21X1  g01264(.A0(new_n3699_), .A1(pi0039), .B0(pi0038), .Y(new_n3700_));
  OAI21X1  g01265(.A0(new_n3695_), .A1(new_n3687_), .B0(new_n3700_), .Y(new_n3701_));
  INVX1    g01266(.A(new_n3626_), .Y(new_n3702_));
  INVX1    g01267(.A(new_n3647_), .Y(new_n3703_));
  AOI21X1  g01268(.A0(new_n3703_), .A1(pi0299), .B0(new_n3702_), .Y(new_n3704_));
  AOI21X1  g01269(.A0(new_n3704_), .A1(pi0038), .B0(pi0100), .Y(new_n3705_));
  INVX1    g01270(.A(pi1142), .Y(new_n3706_));
  OAI21X1  g01271(.A0(new_n3656_), .A1(new_n3653_), .B0(new_n2438_), .Y(new_n3707_));
  AOI21X1  g01272(.A0(new_n3707_), .A1(new_n3592_), .B0(new_n3591_), .Y(new_n3708_));
  MX2X1    g01273(.A(new_n3708_), .B(new_n3706_), .S0(pi0215), .Y(new_n3709_));
  AND2X1   g01274(.A(new_n3626_), .B(new_n3065_), .Y(new_n3710_));
  OAI21X1  g01275(.A0(new_n3709_), .A1(new_n2953_), .B0(new_n3710_), .Y(new_n3711_));
  AOI21X1  g01276(.A0(new_n3704_), .A1(new_n3066_), .B0(new_n3026_), .Y(new_n3712_));
  AOI22X1  g01277(.A0(new_n3712_), .A1(new_n3711_), .B0(new_n3705_), .B1(new_n3701_), .Y(new_n3713_));
  INVX1    g01278(.A(new_n3704_), .Y(new_n3714_));
  MX2X1    g01279(.A(new_n3714_), .B(new_n3699_), .S0(new_n3085_), .Y(new_n3715_));
  AOI21X1  g01280(.A0(new_n3715_), .A1(pi0087), .B0(pi0075), .Y(new_n3716_));
  OAI21X1  g01281(.A0(new_n3713_), .A1(pi0087), .B0(new_n3716_), .Y(new_n3717_));
  AOI21X1  g01282(.A0(new_n3704_), .A1(pi0075), .B0(pi0092), .Y(new_n3718_));
  NOR2X1   g01283(.A(new_n3715_), .B(new_n3101_), .Y(new_n3719_));
  OAI21X1  g01284(.A0(new_n3714_), .A1(new_n3098_), .B0(pi0092), .Y(new_n3720_));
  OAI21X1  g01285(.A0(new_n3720_), .A1(new_n3719_), .B0(new_n3135_), .Y(new_n3721_));
  AOI21X1  g01286(.A0(new_n3718_), .A1(new_n3717_), .B0(new_n3721_), .Y(new_n3722_));
  OAI21X1  g01287(.A0(new_n3714_), .A1(new_n3135_), .B0(new_n3128_), .Y(new_n3723_));
  NAND2X1  g01288(.A(new_n3698_), .B(new_n3130_), .Y(new_n3724_));
  AOI21X1  g01289(.A0(new_n3647_), .A1(new_n3131_), .B0(new_n3128_), .Y(new_n3725_));
  AOI21X1  g01290(.A0(new_n3725_), .A1(new_n3724_), .B0(pi0056), .Y(new_n3726_));
  OAI21X1  g01291(.A0(new_n3723_), .A1(new_n3722_), .B0(new_n3726_), .Y(new_n3727_));
  AOI21X1  g01292(.A0(new_n3703_), .A1(new_n3242_), .B0(new_n3143_), .Y(new_n3728_));
  OAI21X1  g01293(.A0(new_n3698_), .A1(new_n3242_), .B0(new_n3728_), .Y(new_n3729_));
  AND2X1   g01294(.A(new_n3729_), .B(new_n3245_), .Y(new_n3730_));
  OAI21X1  g01295(.A0(new_n3703_), .A1(new_n3248_), .B0(pi0062), .Y(new_n3731_));
  AOI21X1  g01296(.A0(new_n3698_), .A1(new_n3248_), .B0(new_n3731_), .Y(new_n3732_));
  OR2X1    g01297(.A(new_n3732_), .B(new_n3393_), .Y(new_n3733_));
  AOI21X1  g01298(.A0(new_n3730_), .A1(new_n3727_), .B0(new_n3733_), .Y(new_n3734_));
  OAI21X1  g01299(.A0(new_n3703_), .A1(new_n3246_), .B0(pi0249), .Y(new_n3735_));
  OAI21X1  g01300(.A0(new_n3735_), .A1(new_n3734_), .B0(new_n3686_), .Y(po0157));
  AND2X1   g01301(.A(pi1141), .B(pi0215), .Y(new_n3737_));
  OR2X1    g01302(.A(new_n3737_), .B(new_n2953_), .Y(new_n3738_));
  INVX1    g01303(.A(pi0935), .Y(new_n3739_));
  AOI21X1  g01304(.A0(new_n2442_), .A1(new_n3739_), .B0(new_n2437_), .Y(new_n3740_));
  OAI21X1  g01305(.A0(new_n2442_), .A1(pi1141), .B0(new_n3740_), .Y(new_n3741_));
  AOI21X1  g01306(.A0(pi0270), .A1(pi0216), .B0(pi0221), .Y(new_n3742_));
  INVX1    g01307(.A(new_n3742_), .Y(new_n3743_));
  INVX1    g01308(.A(pi0861), .Y(new_n3744_));
  AOI21X1  g01309(.A0(new_n3271_), .A1(pi0861), .B0(pi0171), .Y(new_n3745_));
  AOI21X1  g01310(.A0(new_n3266_), .A1(pi0171), .B0(new_n3745_), .Y(new_n3746_));
  NAND2X1  g01311(.A(new_n3745_), .B(new_n3204_), .Y(new_n3747_));
  OAI21X1  g01312(.A0(new_n3746_), .A1(new_n3744_), .B0(new_n3747_), .Y(new_n3748_));
  AOI21X1  g01313(.A0(new_n2454_), .A1(pi0095), .B0(new_n3744_), .Y(new_n3749_));
  AOI21X1  g01314(.A0(pi0171), .A1(new_n2448_), .B0(new_n3013_), .Y(new_n3750_));
  OAI21X1  g01315(.A0(new_n3749_), .A1(new_n2448_), .B0(new_n3750_), .Y(new_n3751_));
  OAI21X1  g01316(.A0(new_n3751_), .A1(new_n3270_), .B0(new_n2438_), .Y(new_n3752_));
  AOI21X1  g01317(.A0(new_n3748_), .A1(new_n3013_), .B0(new_n3752_), .Y(new_n3753_));
  OAI21X1  g01318(.A0(new_n3753_), .A1(new_n3743_), .B0(new_n3741_), .Y(new_n3754_));
  AOI21X1  g01319(.A0(new_n3754_), .A1(new_n2954_), .B0(new_n3738_), .Y(new_n3755_));
  AOI21X1  g01320(.A0(pi1141), .A1(pi0223), .B0(pi0299), .Y(new_n3756_));
  INVX1    g01321(.A(new_n3756_), .Y(new_n3757_));
  AOI21X1  g01322(.A0(new_n3159_), .A1(new_n3739_), .B0(new_n2960_), .Y(new_n3758_));
  OAI21X1  g01323(.A0(new_n3159_), .A1(pi1141), .B0(new_n3758_), .Y(new_n3759_));
  AOI21X1  g01324(.A0(pi0270), .A1(pi0224), .B0(pi0222), .Y(new_n3760_));
  INVX1    g01325(.A(new_n3760_), .Y(new_n3761_));
  AOI21X1  g01326(.A0(new_n3258_), .A1(pi0861), .B0(pi0224), .Y(new_n3762_));
  OAI21X1  g01327(.A0(new_n3762_), .A1(new_n3761_), .B0(new_n3759_), .Y(new_n3763_));
  NOR2X1   g01328(.A(new_n3761_), .B(new_n3258_), .Y(new_n3764_));
  OAI21X1  g01329(.A0(new_n3764_), .A1(new_n3763_), .B0(new_n2964_), .Y(new_n3765_));
  AOI21X1  g01330(.A0(new_n3765_), .A1(new_n3756_), .B0(pi0039), .Y(new_n3766_));
  OAI21X1  g01331(.A0(new_n3763_), .A1(new_n3757_), .B0(new_n3766_), .Y(new_n3767_));
  AND2X1   g01332(.A(pi1141), .B(pi0223), .Y(new_n3768_));
  OAI21X1  g01333(.A0(new_n3749_), .A1(pi0224), .B0(new_n3760_), .Y(new_n3769_));
  AOI21X1  g01334(.A0(new_n3769_), .A1(new_n3759_), .B0(pi0223), .Y(new_n3770_));
  OAI21X1  g01335(.A0(new_n3770_), .A1(new_n3768_), .B0(new_n2953_), .Y(new_n3771_));
  AND2X1   g01336(.A(new_n3751_), .B(new_n2438_), .Y(new_n3772_));
  INVX1    g01337(.A(new_n3772_), .Y(new_n3773_));
  INVX1    g01338(.A(pi0171), .Y(new_n3774_));
  OAI21X1  g01339(.A0(new_n3630_), .A1(new_n3774_), .B0(new_n3013_), .Y(new_n3775_));
  AOI21X1  g01340(.A0(new_n3630_), .A1(new_n3744_), .B0(new_n3775_), .Y(new_n3776_));
  OAI21X1  g01341(.A0(new_n3776_), .A1(new_n3773_), .B0(new_n3742_), .Y(new_n3777_));
  AOI21X1  g01342(.A0(new_n3777_), .A1(new_n3741_), .B0(pi0215), .Y(new_n3778_));
  OAI21X1  g01343(.A0(new_n3778_), .A1(new_n3737_), .B0(pi0299), .Y(new_n3779_));
  NAND2X1  g01344(.A(new_n3779_), .B(new_n3771_), .Y(new_n3780_));
  AOI21X1  g01345(.A0(new_n3780_), .A1(pi0039), .B0(pi0038), .Y(new_n3781_));
  OAI21X1  g01346(.A0(new_n3767_), .A1(new_n3755_), .B0(new_n3781_), .Y(new_n3782_));
  INVX1    g01347(.A(new_n3771_), .Y(new_n3783_));
  AOI21X1  g01348(.A0(new_n3013_), .A1(new_n3774_), .B0(new_n3773_), .Y(new_n3784_));
  OAI21X1  g01349(.A0(new_n3784_), .A1(new_n3743_), .B0(new_n3741_), .Y(new_n3785_));
  AOI21X1  g01350(.A0(new_n3785_), .A1(new_n2954_), .B0(new_n3737_), .Y(new_n3786_));
  INVX1    g01351(.A(new_n3786_), .Y(new_n3787_));
  AOI21X1  g01352(.A0(new_n3787_), .A1(pi0299), .B0(new_n3783_), .Y(new_n3788_));
  AOI21X1  g01353(.A0(new_n3788_), .A1(pi0038), .B0(pi0100), .Y(new_n3789_));
  INVX1    g01354(.A(new_n3737_), .Y(new_n3790_));
  INVX1    g01355(.A(new_n3741_), .Y(new_n3791_));
  AOI21X1  g01356(.A0(new_n3221_), .A1(pi0171), .B0(pi0228), .Y(new_n3792_));
  OAI21X1  g01357(.A0(new_n3221_), .A1(pi0861), .B0(new_n3792_), .Y(new_n3793_));
  AOI21X1  g01358(.A0(new_n3793_), .A1(new_n3772_), .B0(new_n3743_), .Y(new_n3794_));
  OAI21X1  g01359(.A0(new_n3794_), .A1(new_n3791_), .B0(new_n2954_), .Y(new_n3795_));
  AOI21X1  g01360(.A0(new_n3795_), .A1(new_n3790_), .B0(new_n2953_), .Y(new_n3796_));
  OR4X1    g01361(.A(new_n3796_), .B(new_n3783_), .C(pi0039), .D(pi0038), .Y(new_n3797_));
  AOI21X1  g01362(.A0(new_n3788_), .A1(new_n3066_), .B0(new_n3026_), .Y(new_n3798_));
  AOI22X1  g01363(.A0(new_n3798_), .A1(new_n3797_), .B0(new_n3789_), .B1(new_n3782_), .Y(new_n3799_));
  INVX1    g01364(.A(new_n3788_), .Y(new_n3800_));
  MX2X1    g01365(.A(new_n3800_), .B(new_n3780_), .S0(new_n3085_), .Y(new_n3801_));
  AOI21X1  g01366(.A0(new_n3801_), .A1(pi0087), .B0(pi0075), .Y(new_n3802_));
  OAI21X1  g01367(.A0(new_n3799_), .A1(pi0087), .B0(new_n3802_), .Y(new_n3803_));
  AOI21X1  g01368(.A0(new_n3788_), .A1(pi0075), .B0(pi0092), .Y(new_n3804_));
  NOR2X1   g01369(.A(new_n3801_), .B(new_n3101_), .Y(new_n3805_));
  OAI21X1  g01370(.A0(new_n3800_), .A1(new_n3098_), .B0(pi0092), .Y(new_n3806_));
  OAI21X1  g01371(.A0(new_n3806_), .A1(new_n3805_), .B0(new_n3135_), .Y(new_n3807_));
  AOI21X1  g01372(.A0(new_n3804_), .A1(new_n3803_), .B0(new_n3807_), .Y(new_n3808_));
  OAI21X1  g01373(.A0(new_n3800_), .A1(new_n3135_), .B0(new_n3128_), .Y(new_n3809_));
  INVX1    g01374(.A(new_n3129_), .Y(new_n3810_));
  OR4X1    g01375(.A(new_n3778_), .B(new_n3737_), .C(new_n3810_), .D(new_n3066_), .Y(new_n3811_));
  AOI21X1  g01376(.A0(new_n3786_), .A1(new_n3131_), .B0(new_n3128_), .Y(new_n3812_));
  AOI21X1  g01377(.A0(new_n3812_), .A1(new_n3811_), .B0(pi0056), .Y(new_n3813_));
  OAI21X1  g01378(.A0(new_n3809_), .A1(new_n3808_), .B0(new_n3813_), .Y(new_n3814_));
  OAI21X1  g01379(.A0(new_n3778_), .A1(new_n3737_), .B0(new_n3140_), .Y(new_n3815_));
  AOI21X1  g01380(.A0(new_n3787_), .A1(new_n3242_), .B0(new_n3143_), .Y(new_n3816_));
  AOI21X1  g01381(.A0(new_n3816_), .A1(new_n3815_), .B0(pi0062), .Y(new_n3817_));
  NOR3X1   g01382(.A(new_n3778_), .B(new_n3737_), .C(new_n3249_), .Y(new_n3818_));
  OAI21X1  g01383(.A0(new_n3787_), .A1(new_n3248_), .B0(pi0062), .Y(new_n3819_));
  NOR3X1   g01384(.A(pi0241), .B(pi0059), .C(pi0057), .Y(new_n3820_));
  OAI21X1  g01385(.A0(new_n3819_), .A1(new_n3818_), .B0(new_n3820_), .Y(new_n3821_));
  AOI21X1  g01386(.A0(new_n3817_), .A1(new_n3814_), .B0(new_n3821_), .Y(new_n3822_));
  OAI21X1  g01387(.A0(new_n3531_), .A1(pi0861), .B0(new_n3774_), .Y(new_n3823_));
  AOI21X1  g01388(.A0(new_n3532_), .A1(new_n3744_), .B0(new_n3774_), .Y(new_n3824_));
  OAI21X1  g01389(.A0(new_n3535_), .A1(new_n3744_), .B0(new_n3824_), .Y(new_n3825_));
  AOI21X1  g01390(.A0(new_n3825_), .A1(new_n3823_), .B0(pi0228), .Y(new_n3826_));
  OAI21X1  g01391(.A0(new_n3258_), .A1(new_n3030_), .B0(new_n3772_), .Y(new_n3827_));
  OAI21X1  g01392(.A0(new_n3827_), .A1(new_n3826_), .B0(new_n3742_), .Y(new_n3828_));
  AOI21X1  g01393(.A0(new_n3828_), .A1(new_n3741_), .B0(pi0215), .Y(new_n3829_));
  OAI21X1  g01394(.A0(new_n3829_), .A1(new_n3738_), .B0(new_n3766_), .Y(new_n3830_));
  INVX1    g01395(.A(new_n3286_), .Y(new_n3831_));
  AND2X1   g01396(.A(new_n3771_), .B(new_n3831_), .Y(new_n3832_));
  NAND3X1  g01397(.A(new_n3751_), .B(new_n3479_), .C(new_n2438_), .Y(new_n3833_));
  OAI21X1  g01398(.A0(new_n3833_), .A1(new_n3776_), .B0(new_n3742_), .Y(new_n3834_));
  AOI21X1  g01399(.A0(new_n3834_), .A1(new_n3741_), .B0(pi0215), .Y(new_n3835_));
  OAI21X1  g01400(.A0(new_n3835_), .A1(new_n3737_), .B0(pi0299), .Y(new_n3836_));
  NAND2X1  g01401(.A(new_n3836_), .B(new_n3832_), .Y(new_n3837_));
  AOI21X1  g01402(.A0(new_n3837_), .A1(pi0039), .B0(pi0038), .Y(new_n3838_));
  INVX1    g01403(.A(new_n3832_), .Y(new_n3839_));
  AOI21X1  g01404(.A0(pi0270), .A1(pi0216), .B0(new_n3548_), .Y(new_n3840_));
  NOR2X1   g01405(.A(new_n3840_), .B(new_n3787_), .Y(new_n3841_));
  INVX1    g01406(.A(new_n3841_), .Y(new_n3842_));
  AOI21X1  g01407(.A0(new_n3842_), .A1(pi0299), .B0(new_n3839_), .Y(new_n3843_));
  INVX1    g01408(.A(new_n3843_), .Y(new_n3844_));
  OAI21X1  g01409(.A0(new_n3844_), .A1(new_n2996_), .B0(new_n3026_), .Y(new_n3845_));
  AOI21X1  g01410(.A0(new_n3838_), .A1(new_n3830_), .B0(new_n3845_), .Y(new_n3846_));
  INVX1    g01411(.A(pi1141), .Y(new_n3847_));
  NAND3X1  g01412(.A(new_n3793_), .B(new_n3772_), .C(new_n3479_), .Y(new_n3848_));
  AOI21X1  g01413(.A0(new_n3848_), .A1(new_n3742_), .B0(new_n3791_), .Y(new_n3849_));
  MX2X1    g01414(.A(new_n3849_), .B(new_n3847_), .S0(pi0215), .Y(new_n3850_));
  AND2X1   g01415(.A(new_n3832_), .B(new_n3065_), .Y(new_n3851_));
  OAI21X1  g01416(.A0(new_n3850_), .A1(new_n2953_), .B0(new_n3851_), .Y(new_n3852_));
  AOI21X1  g01417(.A0(new_n3843_), .A1(new_n3066_), .B0(new_n3026_), .Y(new_n3853_));
  AND2X1   g01418(.A(new_n3853_), .B(new_n3852_), .Y(new_n3854_));
  OAI21X1  g01419(.A0(new_n3854_), .A1(new_n3846_), .B0(new_n3156_), .Y(new_n3855_));
  MX2X1    g01420(.A(new_n3844_), .B(new_n3837_), .S0(new_n3085_), .Y(new_n3856_));
  AOI21X1  g01421(.A0(new_n3856_), .A1(pi0087), .B0(pi0075), .Y(new_n3857_));
  OAI21X1  g01422(.A0(new_n3844_), .A1(new_n3095_), .B0(new_n3100_), .Y(new_n3858_));
  AOI21X1  g01423(.A0(new_n3857_), .A1(new_n3855_), .B0(new_n3858_), .Y(new_n3859_));
  OR2X1    g01424(.A(new_n3856_), .B(new_n3101_), .Y(new_n3860_));
  AOI21X1  g01425(.A0(new_n3843_), .A1(new_n3101_), .B0(new_n3100_), .Y(new_n3861_));
  AND2X1   g01426(.A(new_n3861_), .B(new_n3860_), .Y(new_n3862_));
  NOR3X1   g01427(.A(new_n3862_), .B(new_n3859_), .C(new_n3136_), .Y(new_n3863_));
  OAI21X1  g01428(.A0(new_n3844_), .A1(new_n3135_), .B0(new_n3128_), .Y(new_n3864_));
  OR4X1    g01429(.A(new_n3835_), .B(new_n3737_), .C(new_n3810_), .D(new_n3066_), .Y(new_n3865_));
  AOI21X1  g01430(.A0(new_n3841_), .A1(new_n3131_), .B0(new_n3128_), .Y(new_n3866_));
  AOI21X1  g01431(.A0(new_n3866_), .A1(new_n3865_), .B0(pi0056), .Y(new_n3867_));
  OAI21X1  g01432(.A0(new_n3864_), .A1(new_n3863_), .B0(new_n3867_), .Y(new_n3868_));
  OAI21X1  g01433(.A0(new_n3835_), .A1(new_n3737_), .B0(new_n3140_), .Y(new_n3869_));
  AOI21X1  g01434(.A0(new_n3842_), .A1(new_n3242_), .B0(new_n3143_), .Y(new_n3870_));
  AOI21X1  g01435(.A0(new_n3870_), .A1(new_n3869_), .B0(pi0062), .Y(new_n3871_));
  NOR3X1   g01436(.A(new_n3835_), .B(new_n3737_), .C(new_n3249_), .Y(new_n3872_));
  OAI21X1  g01437(.A0(new_n3842_), .A1(new_n3248_), .B0(pi0062), .Y(new_n3873_));
  AND2X1   g01438(.A(new_n3246_), .B(pi0241), .Y(new_n3874_));
  OAI21X1  g01439(.A0(new_n3873_), .A1(new_n3872_), .B0(new_n3874_), .Y(new_n3875_));
  AOI21X1  g01440(.A0(new_n3871_), .A1(new_n3868_), .B0(new_n3875_), .Y(new_n3876_));
  AOI21X1  g01441(.A0(new_n3840_), .A1(pi0241), .B0(new_n3246_), .Y(new_n3877_));
  AND2X1   g01442(.A(new_n3877_), .B(new_n3786_), .Y(new_n3878_));
  NOR3X1   g01443(.A(new_n3878_), .B(new_n3876_), .C(new_n3822_), .Y(po0158));
  AND2X1   g01444(.A(pi1140), .B(pi0215), .Y(new_n3880_));
  OR2X1    g01445(.A(new_n3880_), .B(new_n2953_), .Y(new_n3881_));
  INVX1    g01446(.A(pi0921), .Y(new_n3882_));
  AOI21X1  g01447(.A0(new_n2442_), .A1(new_n3882_), .B0(new_n2437_), .Y(new_n3883_));
  OAI21X1  g01448(.A0(new_n2442_), .A1(pi1140), .B0(new_n3883_), .Y(new_n3884_));
  AOI21X1  g01449(.A0(pi0282), .A1(pi0216), .B0(pi0221), .Y(new_n3885_));
  INVX1    g01450(.A(new_n3885_), .Y(new_n3886_));
  INVX1    g01451(.A(pi0869), .Y(new_n3887_));
  AOI21X1  g01452(.A0(new_n3271_), .A1(pi0869), .B0(pi0170), .Y(new_n3888_));
  AOI21X1  g01453(.A0(new_n3266_), .A1(pi0170), .B0(new_n3888_), .Y(new_n3889_));
  NAND2X1  g01454(.A(new_n3888_), .B(new_n3204_), .Y(new_n3890_));
  OAI21X1  g01455(.A0(new_n3889_), .A1(new_n3887_), .B0(new_n3890_), .Y(new_n3891_));
  AOI21X1  g01456(.A0(new_n2454_), .A1(pi0095), .B0(new_n3887_), .Y(new_n3892_));
  AOI21X1  g01457(.A0(pi0170), .A1(new_n2448_), .B0(new_n3013_), .Y(new_n3893_));
  OAI21X1  g01458(.A0(new_n3892_), .A1(new_n2448_), .B0(new_n3893_), .Y(new_n3894_));
  OAI21X1  g01459(.A0(new_n3894_), .A1(new_n3270_), .B0(new_n2438_), .Y(new_n3895_));
  AOI21X1  g01460(.A0(new_n3891_), .A1(new_n3013_), .B0(new_n3895_), .Y(new_n3896_));
  OAI21X1  g01461(.A0(new_n3896_), .A1(new_n3886_), .B0(new_n3884_), .Y(new_n3897_));
  AOI21X1  g01462(.A0(new_n3897_), .A1(new_n2954_), .B0(new_n3881_), .Y(new_n3898_));
  AOI21X1  g01463(.A0(pi1140), .A1(pi0223), .B0(pi0299), .Y(new_n3899_));
  INVX1    g01464(.A(new_n3899_), .Y(new_n3900_));
  AOI21X1  g01465(.A0(new_n3159_), .A1(new_n3882_), .B0(new_n2960_), .Y(new_n3901_));
  OAI21X1  g01466(.A0(new_n3159_), .A1(pi1140), .B0(new_n3901_), .Y(new_n3902_));
  AOI21X1  g01467(.A0(pi0282), .A1(pi0224), .B0(pi0222), .Y(new_n3903_));
  INVX1    g01468(.A(new_n3903_), .Y(new_n3904_));
  AOI21X1  g01469(.A0(new_n3258_), .A1(pi0869), .B0(pi0224), .Y(new_n3905_));
  OAI21X1  g01470(.A0(new_n3905_), .A1(new_n3904_), .B0(new_n3902_), .Y(new_n3906_));
  NOR2X1   g01471(.A(new_n3904_), .B(new_n3258_), .Y(new_n3907_));
  OAI21X1  g01472(.A0(new_n3907_), .A1(new_n3906_), .B0(new_n2964_), .Y(new_n3908_));
  AOI21X1  g01473(.A0(new_n3908_), .A1(new_n3899_), .B0(pi0039), .Y(new_n3909_));
  OAI21X1  g01474(.A0(new_n3906_), .A1(new_n3900_), .B0(new_n3909_), .Y(new_n3910_));
  AND2X1   g01475(.A(pi1140), .B(pi0223), .Y(new_n3911_));
  OAI21X1  g01476(.A0(new_n3892_), .A1(pi0224), .B0(new_n3903_), .Y(new_n3912_));
  AOI21X1  g01477(.A0(new_n3912_), .A1(new_n3902_), .B0(pi0223), .Y(new_n3913_));
  OAI21X1  g01478(.A0(new_n3913_), .A1(new_n3911_), .B0(new_n2953_), .Y(new_n3914_));
  AND2X1   g01479(.A(new_n3894_), .B(new_n2438_), .Y(new_n3915_));
  INVX1    g01480(.A(new_n3915_), .Y(new_n3916_));
  INVX1    g01481(.A(pi0170), .Y(new_n3917_));
  OAI21X1  g01482(.A0(new_n3630_), .A1(new_n3917_), .B0(new_n3013_), .Y(new_n3918_));
  AOI21X1  g01483(.A0(new_n3630_), .A1(new_n3887_), .B0(new_n3918_), .Y(new_n3919_));
  OAI21X1  g01484(.A0(new_n3919_), .A1(new_n3916_), .B0(new_n3885_), .Y(new_n3920_));
  AOI21X1  g01485(.A0(new_n3920_), .A1(new_n3884_), .B0(pi0215), .Y(new_n3921_));
  OAI21X1  g01486(.A0(new_n3921_), .A1(new_n3880_), .B0(pi0299), .Y(new_n3922_));
  NAND2X1  g01487(.A(new_n3922_), .B(new_n3914_), .Y(new_n3923_));
  AOI21X1  g01488(.A0(new_n3923_), .A1(pi0039), .B0(pi0038), .Y(new_n3924_));
  OAI21X1  g01489(.A0(new_n3910_), .A1(new_n3898_), .B0(new_n3924_), .Y(new_n3925_));
  INVX1    g01490(.A(new_n3914_), .Y(new_n3926_));
  AOI21X1  g01491(.A0(new_n3013_), .A1(new_n3917_), .B0(new_n3916_), .Y(new_n3927_));
  OAI21X1  g01492(.A0(new_n3927_), .A1(new_n3886_), .B0(new_n3884_), .Y(new_n3928_));
  AOI21X1  g01493(.A0(new_n3928_), .A1(new_n2954_), .B0(new_n3880_), .Y(new_n3929_));
  INVX1    g01494(.A(new_n3929_), .Y(new_n3930_));
  AOI21X1  g01495(.A0(new_n3930_), .A1(pi0299), .B0(new_n3926_), .Y(new_n3931_));
  AOI21X1  g01496(.A0(new_n3931_), .A1(pi0038), .B0(pi0100), .Y(new_n3932_));
  INVX1    g01497(.A(new_n3880_), .Y(new_n3933_));
  INVX1    g01498(.A(new_n3884_), .Y(new_n3934_));
  AOI21X1  g01499(.A0(new_n3221_), .A1(pi0170), .B0(pi0228), .Y(new_n3935_));
  OAI21X1  g01500(.A0(new_n3221_), .A1(pi0869), .B0(new_n3935_), .Y(new_n3936_));
  AOI21X1  g01501(.A0(new_n3936_), .A1(new_n3915_), .B0(new_n3886_), .Y(new_n3937_));
  OAI21X1  g01502(.A0(new_n3937_), .A1(new_n3934_), .B0(new_n2954_), .Y(new_n3938_));
  AOI21X1  g01503(.A0(new_n3938_), .A1(new_n3933_), .B0(new_n2953_), .Y(new_n3939_));
  OR4X1    g01504(.A(new_n3939_), .B(new_n3926_), .C(pi0039), .D(pi0038), .Y(new_n3940_));
  AOI21X1  g01505(.A0(new_n3931_), .A1(new_n3066_), .B0(new_n3026_), .Y(new_n3941_));
  AOI22X1  g01506(.A0(new_n3941_), .A1(new_n3940_), .B0(new_n3932_), .B1(new_n3925_), .Y(new_n3942_));
  INVX1    g01507(.A(new_n3931_), .Y(new_n3943_));
  MX2X1    g01508(.A(new_n3943_), .B(new_n3923_), .S0(new_n3085_), .Y(new_n3944_));
  AOI21X1  g01509(.A0(new_n3944_), .A1(pi0087), .B0(pi0075), .Y(new_n3945_));
  OAI21X1  g01510(.A0(new_n3942_), .A1(pi0087), .B0(new_n3945_), .Y(new_n3946_));
  AOI21X1  g01511(.A0(new_n3931_), .A1(pi0075), .B0(pi0092), .Y(new_n3947_));
  NOR2X1   g01512(.A(new_n3944_), .B(new_n3101_), .Y(new_n3948_));
  OAI21X1  g01513(.A0(new_n3943_), .A1(new_n3098_), .B0(pi0092), .Y(new_n3949_));
  OAI21X1  g01514(.A0(new_n3949_), .A1(new_n3948_), .B0(new_n3135_), .Y(new_n3950_));
  AOI21X1  g01515(.A0(new_n3947_), .A1(new_n3946_), .B0(new_n3950_), .Y(new_n3951_));
  OAI21X1  g01516(.A0(new_n3943_), .A1(new_n3135_), .B0(new_n3128_), .Y(new_n3952_));
  OR4X1    g01517(.A(new_n3921_), .B(new_n3880_), .C(new_n3810_), .D(new_n3066_), .Y(new_n3953_));
  AOI21X1  g01518(.A0(new_n3929_), .A1(new_n3131_), .B0(new_n3128_), .Y(new_n3954_));
  AOI21X1  g01519(.A0(new_n3954_), .A1(new_n3953_), .B0(pi0056), .Y(new_n3955_));
  OAI21X1  g01520(.A0(new_n3952_), .A1(new_n3951_), .B0(new_n3955_), .Y(new_n3956_));
  OAI21X1  g01521(.A0(new_n3921_), .A1(new_n3880_), .B0(new_n3140_), .Y(new_n3957_));
  AOI21X1  g01522(.A0(new_n3930_), .A1(new_n3242_), .B0(new_n3143_), .Y(new_n3958_));
  AOI21X1  g01523(.A0(new_n3958_), .A1(new_n3957_), .B0(pi0062), .Y(new_n3959_));
  NOR3X1   g01524(.A(new_n3921_), .B(new_n3880_), .C(new_n3249_), .Y(new_n3960_));
  OAI21X1  g01525(.A0(new_n3930_), .A1(new_n3248_), .B0(pi0062), .Y(new_n3961_));
  NOR3X1   g01526(.A(pi0248), .B(pi0059), .C(pi0057), .Y(new_n3962_));
  OAI21X1  g01527(.A0(new_n3961_), .A1(new_n3960_), .B0(new_n3962_), .Y(new_n3963_));
  AOI21X1  g01528(.A0(new_n3959_), .A1(new_n3956_), .B0(new_n3963_), .Y(new_n3964_));
  OAI21X1  g01529(.A0(new_n3531_), .A1(pi0869), .B0(new_n3917_), .Y(new_n3965_));
  AOI21X1  g01530(.A0(new_n3532_), .A1(new_n3887_), .B0(new_n3917_), .Y(new_n3966_));
  OAI21X1  g01531(.A0(new_n3535_), .A1(new_n3887_), .B0(new_n3966_), .Y(new_n3967_));
  AOI21X1  g01532(.A0(new_n3967_), .A1(new_n3965_), .B0(pi0228), .Y(new_n3968_));
  OAI21X1  g01533(.A0(new_n3258_), .A1(new_n3030_), .B0(new_n3915_), .Y(new_n3969_));
  OAI21X1  g01534(.A0(new_n3969_), .A1(new_n3968_), .B0(new_n3885_), .Y(new_n3970_));
  AOI21X1  g01535(.A0(new_n3970_), .A1(new_n3884_), .B0(pi0215), .Y(new_n3971_));
  OAI21X1  g01536(.A0(new_n3971_), .A1(new_n3881_), .B0(new_n3909_), .Y(new_n3972_));
  AND2X1   g01537(.A(new_n3914_), .B(new_n3831_), .Y(new_n3973_));
  NAND3X1  g01538(.A(new_n3894_), .B(new_n3479_), .C(new_n2438_), .Y(new_n3974_));
  OAI21X1  g01539(.A0(new_n3974_), .A1(new_n3919_), .B0(new_n3885_), .Y(new_n3975_));
  AOI21X1  g01540(.A0(new_n3975_), .A1(new_n3884_), .B0(pi0215), .Y(new_n3976_));
  OAI21X1  g01541(.A0(new_n3976_), .A1(new_n3880_), .B0(pi0299), .Y(new_n3977_));
  NAND2X1  g01542(.A(new_n3977_), .B(new_n3973_), .Y(new_n3978_));
  AOI21X1  g01543(.A0(new_n3978_), .A1(pi0039), .B0(pi0038), .Y(new_n3979_));
  INVX1    g01544(.A(new_n3973_), .Y(new_n3980_));
  AOI21X1  g01545(.A0(pi0282), .A1(pi0216), .B0(new_n3548_), .Y(new_n3981_));
  NOR2X1   g01546(.A(new_n3981_), .B(new_n3930_), .Y(new_n3982_));
  INVX1    g01547(.A(new_n3982_), .Y(new_n3983_));
  AOI21X1  g01548(.A0(new_n3983_), .A1(pi0299), .B0(new_n3980_), .Y(new_n3984_));
  INVX1    g01549(.A(new_n3984_), .Y(new_n3985_));
  OAI21X1  g01550(.A0(new_n3985_), .A1(new_n2996_), .B0(new_n3026_), .Y(new_n3986_));
  AOI21X1  g01551(.A0(new_n3979_), .A1(new_n3972_), .B0(new_n3986_), .Y(new_n3987_));
  INVX1    g01552(.A(pi1140), .Y(new_n3988_));
  NAND3X1  g01553(.A(new_n3936_), .B(new_n3915_), .C(new_n3479_), .Y(new_n3989_));
  AOI21X1  g01554(.A0(new_n3989_), .A1(new_n3885_), .B0(new_n3934_), .Y(new_n3990_));
  MX2X1    g01555(.A(new_n3990_), .B(new_n3988_), .S0(pi0215), .Y(new_n3991_));
  AND2X1   g01556(.A(new_n3973_), .B(new_n3065_), .Y(new_n3992_));
  OAI21X1  g01557(.A0(new_n3991_), .A1(new_n2953_), .B0(new_n3992_), .Y(new_n3993_));
  AOI21X1  g01558(.A0(new_n3984_), .A1(new_n3066_), .B0(new_n3026_), .Y(new_n3994_));
  AND2X1   g01559(.A(new_n3994_), .B(new_n3993_), .Y(new_n3995_));
  OAI21X1  g01560(.A0(new_n3995_), .A1(new_n3987_), .B0(new_n3156_), .Y(new_n3996_));
  MX2X1    g01561(.A(new_n3985_), .B(new_n3978_), .S0(new_n3085_), .Y(new_n3997_));
  AOI21X1  g01562(.A0(new_n3997_), .A1(pi0087), .B0(pi0075), .Y(new_n3998_));
  OAI21X1  g01563(.A0(new_n3985_), .A1(new_n3095_), .B0(new_n3100_), .Y(new_n3999_));
  AOI21X1  g01564(.A0(new_n3998_), .A1(new_n3996_), .B0(new_n3999_), .Y(new_n4000_));
  OR2X1    g01565(.A(new_n3997_), .B(new_n3101_), .Y(new_n4001_));
  AOI21X1  g01566(.A0(new_n3984_), .A1(new_n3101_), .B0(new_n3100_), .Y(new_n4002_));
  AND2X1   g01567(.A(new_n4002_), .B(new_n4001_), .Y(new_n4003_));
  NOR3X1   g01568(.A(new_n4003_), .B(new_n4000_), .C(new_n3136_), .Y(new_n4004_));
  OAI21X1  g01569(.A0(new_n3985_), .A1(new_n3135_), .B0(new_n3128_), .Y(new_n4005_));
  OR4X1    g01570(.A(new_n3976_), .B(new_n3880_), .C(new_n3810_), .D(new_n3066_), .Y(new_n4006_));
  AOI21X1  g01571(.A0(new_n3982_), .A1(new_n3131_), .B0(new_n3128_), .Y(new_n4007_));
  AOI21X1  g01572(.A0(new_n4007_), .A1(new_n4006_), .B0(pi0056), .Y(new_n4008_));
  OAI21X1  g01573(.A0(new_n4005_), .A1(new_n4004_), .B0(new_n4008_), .Y(new_n4009_));
  OAI21X1  g01574(.A0(new_n3976_), .A1(new_n3880_), .B0(new_n3140_), .Y(new_n4010_));
  AOI21X1  g01575(.A0(new_n3983_), .A1(new_n3242_), .B0(new_n3143_), .Y(new_n4011_));
  AOI21X1  g01576(.A0(new_n4011_), .A1(new_n4010_), .B0(pi0062), .Y(new_n4012_));
  NOR3X1   g01577(.A(new_n3976_), .B(new_n3880_), .C(new_n3249_), .Y(new_n4013_));
  OAI21X1  g01578(.A0(new_n3983_), .A1(new_n3248_), .B0(pi0062), .Y(new_n4014_));
  AND2X1   g01579(.A(new_n3246_), .B(pi0248), .Y(new_n4015_));
  OAI21X1  g01580(.A0(new_n4014_), .A1(new_n4013_), .B0(new_n4015_), .Y(new_n4016_));
  AOI21X1  g01581(.A0(new_n4012_), .A1(new_n4009_), .B0(new_n4016_), .Y(new_n4017_));
  AOI21X1  g01582(.A0(new_n3981_), .A1(pi0248), .B0(new_n3246_), .Y(new_n4018_));
  AND2X1   g01583(.A(new_n4018_), .B(new_n3929_), .Y(new_n4019_));
  NOR3X1   g01584(.A(new_n4019_), .B(new_n4017_), .C(new_n3964_), .Y(po0159));
  NOR2X1   g01585(.A(pi0215), .B(pi0148), .Y(new_n4021_));
  INVX1    g01586(.A(new_n4021_), .Y(new_n4022_));
  AND2X1   g01587(.A(pi0920), .B(pi0833), .Y(new_n4023_));
  INVX1    g01588(.A(new_n4023_), .Y(new_n4024_));
  AOI21X1  g01589(.A0(pi1139), .A1(new_n2721_), .B0(pi0216), .Y(new_n4025_));
  AOI21X1  g01590(.A0(new_n4025_), .A1(new_n4024_), .B0(new_n2437_), .Y(new_n4026_));
  OAI21X1  g01591(.A0(pi1139), .A1(new_n2438_), .B0(new_n4026_), .Y(new_n4027_));
  INVX1    g01592(.A(new_n4027_), .Y(new_n4028_));
  AOI21X1  g01593(.A0(pi0281), .A1(pi0216), .B0(pi0221), .Y(new_n4029_));
  AOI21X1  g01594(.A0(new_n3479_), .A1(pi0862), .B0(pi0216), .Y(new_n4030_));
  OAI21X1  g01595(.A0(new_n3631_), .A1(new_n3028_), .B0(new_n4030_), .Y(new_n4031_));
  AOI21X1  g01596(.A0(new_n4031_), .A1(new_n4029_), .B0(new_n4028_), .Y(new_n4032_));
  NAND3X1  g01597(.A(new_n4029_), .B(new_n3655_), .C(new_n3030_), .Y(new_n4033_));
  AOI21X1  g01598(.A0(new_n4033_), .A1(new_n4032_), .B0(new_n4022_), .Y(new_n4034_));
  INVX1    g01599(.A(pi1139), .Y(new_n4035_));
  INVX1    g01600(.A(pi0148), .Y(new_n4036_));
  INVX1    g01601(.A(new_n4029_), .Y(new_n4037_));
  AOI21X1  g01602(.A0(new_n3028_), .A1(new_n2899_), .B0(new_n3631_), .Y(new_n4038_));
  NOR3X1   g01603(.A(new_n4038_), .B(pi0862), .C(pi0216), .Y(new_n4039_));
  OAI21X1  g01604(.A0(new_n4039_), .A1(new_n4037_), .B0(new_n4027_), .Y(new_n4040_));
  AOI21X1  g01605(.A0(new_n4029_), .A1(new_n3367_), .B0(new_n4040_), .Y(new_n4041_));
  NOR2X1   g01606(.A(new_n4026_), .B(pi0216), .Y(new_n4042_));
  AND2X1   g01607(.A(new_n4042_), .B(new_n3367_), .Y(new_n4043_));
  OR4X1    g01608(.A(new_n4043_), .B(new_n4041_), .C(pi0215), .D(new_n4036_), .Y(new_n4044_));
  OAI21X1  g01609(.A0(new_n4035_), .A1(new_n2954_), .B0(new_n4044_), .Y(new_n4045_));
  OAI21X1  g01610(.A0(new_n4045_), .A1(new_n4034_), .B0(pi0299), .Y(new_n4046_));
  AOI21X1  g01611(.A0(pi0833), .A1(new_n2961_), .B0(pi1139), .Y(new_n4047_));
  NOR3X1   g01612(.A(pi0920), .B(new_n2721_), .C(pi0224), .Y(new_n4048_));
  NOR3X1   g01613(.A(new_n4048_), .B(new_n4047_), .C(new_n2960_), .Y(new_n4049_));
  AND2X1   g01614(.A(pi1139), .B(pi0223), .Y(new_n4050_));
  NOR4X1   g01615(.A(new_n4050_), .B(new_n4049_), .C(new_n2899_), .D(pi0224), .Y(new_n4051_));
  NOR4X1   g01616(.A(new_n4050_), .B(new_n4049_), .C(pi0862), .D(pi0224), .Y(new_n4052_));
  AOI21X1  g01617(.A0(pi0281), .A1(pi0224), .B0(pi0222), .Y(new_n4053_));
  NOR2X1   g01618(.A(new_n4053_), .B(new_n4049_), .Y(new_n4054_));
  MX2X1    g01619(.A(new_n4054_), .B(new_n4035_), .S0(pi0223), .Y(new_n4055_));
  NOR4X1   g01620(.A(new_n4055_), .B(new_n4052_), .C(new_n4051_), .D(pi0299), .Y(new_n4056_));
  NOR2X1   g01621(.A(new_n4056_), .B(new_n3066_), .Y(new_n4057_));
  NOR4X1   g01622(.A(new_n3030_), .B(new_n2455_), .C(pi0862), .D(pi0216), .Y(new_n4058_));
  OAI21X1  g01623(.A0(new_n4058_), .A1(new_n4037_), .B0(new_n4027_), .Y(new_n4059_));
  NOR4X1   g01624(.A(new_n4026_), .B(new_n3028_), .C(pi0216), .D(new_n4036_), .Y(new_n4060_));
  NOR2X1   g01625(.A(new_n4060_), .B(pi0215), .Y(new_n4061_));
  AOI22X1  g01626(.A0(new_n4061_), .A1(new_n4059_), .B0(pi1139), .B1(pi0215), .Y(new_n4062_));
  NOR2X1   g01627(.A(new_n4062_), .B(new_n3281_), .Y(new_n4063_));
  AOI21X1  g01628(.A0(new_n4063_), .A1(pi0299), .B0(new_n4056_), .Y(new_n4064_));
  INVX1    g01629(.A(new_n4064_), .Y(new_n4065_));
  OAI21X1  g01630(.A0(new_n4065_), .A1(new_n3065_), .B0(pi0100), .Y(new_n4066_));
  AOI21X1  g01631(.A0(new_n4057_), .A1(new_n4046_), .B0(new_n4066_), .Y(new_n4067_));
  OAI21X1  g01632(.A0(new_n3204_), .A1(pi0228), .B0(new_n3030_), .Y(new_n4068_));
  AOI21X1  g01633(.A0(new_n3326_), .A1(pi0862), .B0(pi0216), .Y(new_n4069_));
  OAI21X1  g01634(.A0(new_n4068_), .A1(pi0862), .B0(new_n4069_), .Y(new_n4070_));
  AOI21X1  g01635(.A0(new_n4070_), .A1(new_n4029_), .B0(new_n4028_), .Y(new_n4071_));
  NOR2X1   g01636(.A(new_n4071_), .B(new_n4022_), .Y(new_n4072_));
  NOR3X1   g01637(.A(new_n3267_), .B(pi0862), .C(pi0216), .Y(new_n4073_));
  OAI21X1  g01638(.A0(new_n4073_), .A1(new_n4037_), .B0(new_n4027_), .Y(new_n4074_));
  INVX1    g01639(.A(new_n4074_), .Y(new_n4075_));
  AND2X1   g01640(.A(new_n2954_), .B(pi0148), .Y(new_n4076_));
  INVX1    g01641(.A(new_n4076_), .Y(new_n4077_));
  AND2X1   g01642(.A(new_n4042_), .B(new_n3267_), .Y(new_n4078_));
  OR2X1    g01643(.A(new_n4078_), .B(new_n4077_), .Y(new_n4079_));
  AOI21X1  g01644(.A0(pi1139), .A1(pi0215), .B0(new_n2953_), .Y(new_n4080_));
  OAI21X1  g01645(.A0(new_n4079_), .A1(new_n4075_), .B0(new_n4080_), .Y(new_n4081_));
  NOR4X1   g01646(.A(new_n4050_), .B(new_n4049_), .C(new_n3258_), .D(pi0224), .Y(new_n4082_));
  OR2X1    g01647(.A(new_n4055_), .B(new_n4052_), .Y(new_n4083_));
  OAI21X1  g01648(.A0(new_n4083_), .A1(new_n4082_), .B0(new_n2953_), .Y(new_n4084_));
  AND2X1   g01649(.A(new_n4084_), .B(new_n2959_), .Y(new_n4085_));
  OAI21X1  g01650(.A0(new_n4081_), .A1(new_n4072_), .B0(new_n4085_), .Y(new_n4086_));
  AOI21X1  g01651(.A0(new_n4042_), .A1(new_n4038_), .B0(new_n4077_), .Y(new_n4087_));
  AOI22X1  g01652(.A0(new_n4087_), .A1(new_n4040_), .B0(pi1139), .B1(pi0215), .Y(new_n4088_));
  OAI21X1  g01653(.A0(new_n4032_), .A1(new_n4022_), .B0(new_n4088_), .Y(new_n4089_));
  AOI21X1  g01654(.A0(new_n4089_), .A1(pi0299), .B0(new_n4056_), .Y(new_n4090_));
  INVX1    g01655(.A(new_n4090_), .Y(new_n4091_));
  AOI21X1  g01656(.A0(new_n4091_), .A1(pi0039), .B0(pi0038), .Y(new_n4092_));
  OAI21X1  g01657(.A0(new_n4065_), .A1(new_n2996_), .B0(new_n3026_), .Y(new_n4093_));
  AOI21X1  g01658(.A0(new_n4092_), .A1(new_n4086_), .B0(new_n4093_), .Y(new_n4094_));
  OAI21X1  g01659(.A0(new_n4094_), .A1(new_n4067_), .B0(new_n3156_), .Y(new_n4095_));
  MX2X1    g01660(.A(new_n4065_), .B(new_n4091_), .S0(new_n3085_), .Y(new_n4096_));
  AOI21X1  g01661(.A0(new_n4096_), .A1(pi0087), .B0(pi0075), .Y(new_n4097_));
  OAI21X1  g01662(.A0(new_n4065_), .A1(new_n3095_), .B0(new_n3100_), .Y(new_n4098_));
  AOI21X1  g01663(.A0(new_n4097_), .A1(new_n4095_), .B0(new_n4098_), .Y(new_n4099_));
  OR2X1    g01664(.A(new_n4096_), .B(new_n3101_), .Y(new_n4100_));
  AOI21X1  g01665(.A0(new_n4064_), .A1(new_n3101_), .B0(new_n3100_), .Y(new_n4101_));
  AND2X1   g01666(.A(new_n4101_), .B(new_n4100_), .Y(new_n4102_));
  NOR3X1   g01667(.A(new_n4102_), .B(new_n4099_), .C(new_n3136_), .Y(new_n4103_));
  OAI21X1  g01668(.A0(new_n4065_), .A1(new_n3135_), .B0(new_n3128_), .Y(new_n4104_));
  OAI21X1  g01669(.A0(new_n4062_), .A1(new_n3281_), .B0(new_n3131_), .Y(new_n4105_));
  AND2X1   g01670(.A(new_n4105_), .B(pi0055), .Y(new_n4106_));
  OAI21X1  g01671(.A0(new_n4089_), .A1(new_n3131_), .B0(new_n4106_), .Y(new_n4107_));
  AND2X1   g01672(.A(new_n4107_), .B(new_n3143_), .Y(new_n4108_));
  OAI21X1  g01673(.A0(new_n4104_), .A1(new_n4103_), .B0(new_n4108_), .Y(new_n4109_));
  NAND2X1  g01674(.A(new_n4089_), .B(new_n3140_), .Y(new_n4110_));
  AOI21X1  g01675(.A0(new_n4063_), .A1(new_n3242_), .B0(new_n3143_), .Y(new_n4111_));
  AOI21X1  g01676(.A0(new_n4111_), .A1(new_n4110_), .B0(pi0062), .Y(new_n4112_));
  NOR2X1   g01677(.A(new_n4089_), .B(new_n3249_), .Y(new_n4113_));
  OAI21X1  g01678(.A0(new_n4063_), .A1(new_n3248_), .B0(pi0062), .Y(new_n4114_));
  OAI21X1  g01679(.A0(new_n4114_), .A1(new_n4113_), .B0(new_n3246_), .Y(new_n4115_));
  AOI21X1  g01680(.A0(new_n4112_), .A1(new_n4109_), .B0(new_n4115_), .Y(new_n4116_));
  INVX1    g01681(.A(pi0247), .Y(new_n4117_));
  OAI21X1  g01682(.A0(new_n4063_), .A1(new_n3246_), .B0(new_n4117_), .Y(new_n4118_));
  NOR2X1   g01683(.A(new_n4041_), .B(new_n4022_), .Y(new_n4119_));
  NOR4X1   g01684(.A(new_n4028_), .B(new_n3654_), .C(new_n3028_), .D(pi0216), .Y(new_n4120_));
  NAND2X1  g01685(.A(new_n4076_), .B(new_n4040_), .Y(new_n4121_));
  OAI22X1  g01686(.A0(new_n4121_), .A1(new_n4120_), .B0(new_n4035_), .B1(new_n2954_), .Y(new_n4122_));
  OAI21X1  g01687(.A0(new_n4122_), .A1(new_n4119_), .B0(pi0299), .Y(new_n4123_));
  NOR3X1   g01688(.A(new_n4055_), .B(new_n4052_), .C(pi0299), .Y(new_n4124_));
  NOR3X1   g01689(.A(new_n4124_), .B(new_n3286_), .C(new_n3066_), .Y(new_n4125_));
  INVX1    g01690(.A(new_n4062_), .Y(new_n4126_));
  NOR2X1   g01691(.A(new_n4124_), .B(new_n3286_), .Y(new_n4127_));
  INVX1    g01692(.A(new_n4127_), .Y(new_n4128_));
  AOI21X1  g01693(.A0(new_n4126_), .A1(pi0299), .B0(new_n4128_), .Y(new_n4129_));
  INVX1    g01694(.A(new_n4129_), .Y(new_n4130_));
  OAI21X1  g01695(.A0(new_n4130_), .A1(new_n3065_), .B0(pi0100), .Y(new_n4131_));
  AOI21X1  g01696(.A0(new_n4125_), .A1(new_n4123_), .B0(new_n4131_), .Y(new_n4132_));
  OR2X1    g01697(.A(new_n4055_), .B(pi0299), .Y(new_n4133_));
  AOI21X1  g01698(.A0(new_n4052_), .A1(new_n3258_), .B0(new_n4133_), .Y(new_n4134_));
  OAI21X1  g01699(.A0(new_n3326_), .A1(pi0862), .B0(new_n2438_), .Y(new_n4135_));
  AOI21X1  g01700(.A0(new_n4068_), .A1(pi0862), .B0(new_n4135_), .Y(new_n4136_));
  OAI21X1  g01701(.A0(new_n4136_), .A1(new_n4037_), .B0(new_n4027_), .Y(new_n4137_));
  NAND2X1  g01702(.A(new_n4137_), .B(new_n4076_), .Y(new_n4138_));
  AOI22X1  g01703(.A0(new_n4074_), .A1(new_n4021_), .B0(pi1139), .B1(pi0215), .Y(new_n4139_));
  AOI21X1  g01704(.A0(new_n4139_), .A1(new_n4138_), .B0(new_n2953_), .Y(new_n4140_));
  OAI21X1  g01705(.A0(new_n4140_), .A1(new_n4134_), .B0(new_n2959_), .Y(new_n4141_));
  NAND2X1  g01706(.A(new_n4061_), .B(new_n4040_), .Y(new_n4142_));
  AOI21X1  g01707(.A0(new_n4142_), .A1(new_n4088_), .B0(new_n2953_), .Y(new_n4143_));
  NOR2X1   g01708(.A(new_n4143_), .B(new_n4128_), .Y(new_n4144_));
  INVX1    g01709(.A(new_n4144_), .Y(new_n4145_));
  AOI21X1  g01710(.A0(new_n4145_), .A1(pi0039), .B0(pi0038), .Y(new_n4146_));
  OAI21X1  g01711(.A0(new_n4130_), .A1(new_n2996_), .B0(new_n3026_), .Y(new_n4147_));
  AOI21X1  g01712(.A0(new_n4146_), .A1(new_n4141_), .B0(new_n4147_), .Y(new_n4148_));
  OAI21X1  g01713(.A0(new_n4148_), .A1(new_n4132_), .B0(new_n3156_), .Y(new_n4149_));
  MX2X1    g01714(.A(new_n4130_), .B(new_n4145_), .S0(new_n3085_), .Y(new_n4150_));
  AOI21X1  g01715(.A0(new_n4150_), .A1(pi0087), .B0(pi0075), .Y(new_n4151_));
  OAI21X1  g01716(.A0(new_n4130_), .A1(new_n3095_), .B0(new_n3100_), .Y(new_n4152_));
  AOI21X1  g01717(.A0(new_n4151_), .A1(new_n4149_), .B0(new_n4152_), .Y(new_n4153_));
  OR2X1    g01718(.A(new_n4150_), .B(new_n3101_), .Y(new_n4154_));
  AOI21X1  g01719(.A0(new_n4129_), .A1(new_n3101_), .B0(new_n3100_), .Y(new_n4155_));
  AND2X1   g01720(.A(new_n4155_), .B(new_n4154_), .Y(new_n4156_));
  NOR3X1   g01721(.A(new_n4156_), .B(new_n4153_), .C(new_n3136_), .Y(new_n4157_));
  OAI21X1  g01722(.A0(new_n4130_), .A1(new_n3135_), .B0(new_n3128_), .Y(new_n4158_));
  NAND3X1  g01723(.A(new_n4142_), .B(new_n4088_), .C(new_n3130_), .Y(new_n4159_));
  AOI21X1  g01724(.A0(new_n4062_), .A1(new_n3131_), .B0(new_n3128_), .Y(new_n4160_));
  AOI21X1  g01725(.A0(new_n4160_), .A1(new_n4159_), .B0(pi0056), .Y(new_n4161_));
  OAI21X1  g01726(.A0(new_n4158_), .A1(new_n4157_), .B0(new_n4161_), .Y(new_n4162_));
  AND2X1   g01727(.A(new_n4142_), .B(new_n4088_), .Y(new_n4163_));
  AOI21X1  g01728(.A0(new_n4126_), .A1(new_n3242_), .B0(new_n3143_), .Y(new_n4164_));
  OAI21X1  g01729(.A0(new_n4163_), .A1(new_n3242_), .B0(new_n4164_), .Y(new_n4165_));
  AND2X1   g01730(.A(new_n4165_), .B(new_n3245_), .Y(new_n4166_));
  OAI21X1  g01731(.A0(new_n4126_), .A1(new_n3248_), .B0(pi0062), .Y(new_n4167_));
  AOI21X1  g01732(.A0(new_n4163_), .A1(new_n3248_), .B0(new_n4167_), .Y(new_n4168_));
  OR2X1    g01733(.A(new_n4168_), .B(new_n3393_), .Y(new_n4169_));
  AOI21X1  g01734(.A0(new_n4166_), .A1(new_n4162_), .B0(new_n4169_), .Y(new_n4170_));
  OAI21X1  g01735(.A0(new_n4126_), .A1(new_n3246_), .B0(pi0247), .Y(new_n4171_));
  OAI22X1  g01736(.A0(new_n4171_), .A1(new_n4170_), .B0(new_n4118_), .B1(new_n4116_), .Y(po0160));
  AND2X1   g01737(.A(pi1138), .B(pi0215), .Y(new_n4173_));
  OR2X1    g01738(.A(new_n4173_), .B(new_n2953_), .Y(new_n4174_));
  INVX1    g01739(.A(pi0940), .Y(new_n4175_));
  AOI21X1  g01740(.A0(new_n2442_), .A1(new_n4175_), .B0(new_n2437_), .Y(new_n4176_));
  OAI21X1  g01741(.A0(new_n2442_), .A1(pi1138), .B0(new_n4176_), .Y(new_n4177_));
  AOI21X1  g01742(.A0(pi0269), .A1(pi0216), .B0(pi0221), .Y(new_n4178_));
  INVX1    g01743(.A(new_n4178_), .Y(new_n4179_));
  INVX1    g01744(.A(pi0877), .Y(new_n4180_));
  AOI21X1  g01745(.A0(new_n3271_), .A1(pi0877), .B0(pi0169), .Y(new_n4181_));
  AOI21X1  g01746(.A0(new_n3266_), .A1(pi0169), .B0(new_n4181_), .Y(new_n4182_));
  NAND2X1  g01747(.A(new_n4181_), .B(new_n3204_), .Y(new_n4183_));
  OAI21X1  g01748(.A0(new_n4182_), .A1(new_n4180_), .B0(new_n4183_), .Y(new_n4184_));
  AOI21X1  g01749(.A0(new_n2454_), .A1(pi0095), .B0(new_n4180_), .Y(new_n4185_));
  AOI21X1  g01750(.A0(pi0169), .A1(new_n2448_), .B0(new_n3013_), .Y(new_n4186_));
  OAI21X1  g01751(.A0(new_n4185_), .A1(new_n2448_), .B0(new_n4186_), .Y(new_n4187_));
  OAI21X1  g01752(.A0(new_n4187_), .A1(new_n3270_), .B0(new_n2438_), .Y(new_n4188_));
  AOI21X1  g01753(.A0(new_n4184_), .A1(new_n3013_), .B0(new_n4188_), .Y(new_n4189_));
  OAI21X1  g01754(.A0(new_n4189_), .A1(new_n4179_), .B0(new_n4177_), .Y(new_n4190_));
  AOI21X1  g01755(.A0(new_n4190_), .A1(new_n2954_), .B0(new_n4174_), .Y(new_n4191_));
  AOI21X1  g01756(.A0(pi1138), .A1(pi0223), .B0(pi0299), .Y(new_n4192_));
  INVX1    g01757(.A(new_n4192_), .Y(new_n4193_));
  AOI21X1  g01758(.A0(new_n3159_), .A1(new_n4175_), .B0(new_n2960_), .Y(new_n4194_));
  OAI21X1  g01759(.A0(new_n3159_), .A1(pi1138), .B0(new_n4194_), .Y(new_n4195_));
  AOI21X1  g01760(.A0(pi0269), .A1(pi0224), .B0(pi0222), .Y(new_n4196_));
  INVX1    g01761(.A(new_n4196_), .Y(new_n4197_));
  AOI21X1  g01762(.A0(new_n3258_), .A1(pi0877), .B0(pi0224), .Y(new_n4198_));
  OAI21X1  g01763(.A0(new_n4198_), .A1(new_n4197_), .B0(new_n4195_), .Y(new_n4199_));
  NOR2X1   g01764(.A(new_n4197_), .B(new_n3258_), .Y(new_n4200_));
  OAI21X1  g01765(.A0(new_n4200_), .A1(new_n4199_), .B0(new_n2964_), .Y(new_n4201_));
  AOI21X1  g01766(.A0(new_n4201_), .A1(new_n4192_), .B0(pi0039), .Y(new_n4202_));
  OAI21X1  g01767(.A0(new_n4199_), .A1(new_n4193_), .B0(new_n4202_), .Y(new_n4203_));
  AND2X1   g01768(.A(pi1138), .B(pi0223), .Y(new_n4204_));
  OAI21X1  g01769(.A0(new_n4185_), .A1(pi0224), .B0(new_n4196_), .Y(new_n4205_));
  AOI21X1  g01770(.A0(new_n4205_), .A1(new_n4195_), .B0(pi0223), .Y(new_n4206_));
  OAI21X1  g01771(.A0(new_n4206_), .A1(new_n4204_), .B0(new_n2953_), .Y(new_n4207_));
  AND2X1   g01772(.A(new_n4187_), .B(new_n2438_), .Y(new_n4208_));
  INVX1    g01773(.A(new_n4208_), .Y(new_n4209_));
  INVX1    g01774(.A(pi0169), .Y(new_n4210_));
  OAI21X1  g01775(.A0(new_n3630_), .A1(new_n4210_), .B0(new_n3013_), .Y(new_n4211_));
  AOI21X1  g01776(.A0(new_n3630_), .A1(new_n4180_), .B0(new_n4211_), .Y(new_n4212_));
  OAI21X1  g01777(.A0(new_n4212_), .A1(new_n4209_), .B0(new_n4178_), .Y(new_n4213_));
  AOI21X1  g01778(.A0(new_n4213_), .A1(new_n4177_), .B0(pi0215), .Y(new_n4214_));
  OAI21X1  g01779(.A0(new_n4214_), .A1(new_n4173_), .B0(pi0299), .Y(new_n4215_));
  NAND2X1  g01780(.A(new_n4215_), .B(new_n4207_), .Y(new_n4216_));
  AOI21X1  g01781(.A0(new_n4216_), .A1(pi0039), .B0(pi0038), .Y(new_n4217_));
  OAI21X1  g01782(.A0(new_n4203_), .A1(new_n4191_), .B0(new_n4217_), .Y(new_n4218_));
  INVX1    g01783(.A(new_n4207_), .Y(new_n4219_));
  AOI21X1  g01784(.A0(new_n3013_), .A1(new_n4210_), .B0(new_n4209_), .Y(new_n4220_));
  OAI21X1  g01785(.A0(new_n4220_), .A1(new_n4179_), .B0(new_n4177_), .Y(new_n4221_));
  AOI21X1  g01786(.A0(new_n4221_), .A1(new_n2954_), .B0(new_n4173_), .Y(new_n4222_));
  INVX1    g01787(.A(new_n4222_), .Y(new_n4223_));
  AOI21X1  g01788(.A0(new_n4223_), .A1(pi0299), .B0(new_n4219_), .Y(new_n4224_));
  AOI21X1  g01789(.A0(new_n4224_), .A1(pi0038), .B0(pi0100), .Y(new_n4225_));
  INVX1    g01790(.A(new_n4173_), .Y(new_n4226_));
  INVX1    g01791(.A(new_n4177_), .Y(new_n4227_));
  AOI21X1  g01792(.A0(new_n3221_), .A1(pi0169), .B0(pi0228), .Y(new_n4228_));
  OAI21X1  g01793(.A0(new_n3221_), .A1(pi0877), .B0(new_n4228_), .Y(new_n4229_));
  AOI21X1  g01794(.A0(new_n4229_), .A1(new_n4208_), .B0(new_n4179_), .Y(new_n4230_));
  OAI21X1  g01795(.A0(new_n4230_), .A1(new_n4227_), .B0(new_n2954_), .Y(new_n4231_));
  AOI21X1  g01796(.A0(new_n4231_), .A1(new_n4226_), .B0(new_n2953_), .Y(new_n4232_));
  OR4X1    g01797(.A(new_n4232_), .B(new_n4219_), .C(pi0039), .D(pi0038), .Y(new_n4233_));
  AOI21X1  g01798(.A0(new_n4224_), .A1(new_n3066_), .B0(new_n3026_), .Y(new_n4234_));
  AOI22X1  g01799(.A0(new_n4234_), .A1(new_n4233_), .B0(new_n4225_), .B1(new_n4218_), .Y(new_n4235_));
  INVX1    g01800(.A(new_n4224_), .Y(new_n4236_));
  MX2X1    g01801(.A(new_n4236_), .B(new_n4216_), .S0(new_n3085_), .Y(new_n4237_));
  AOI21X1  g01802(.A0(new_n4237_), .A1(pi0087), .B0(pi0075), .Y(new_n4238_));
  OAI21X1  g01803(.A0(new_n4235_), .A1(pi0087), .B0(new_n4238_), .Y(new_n4239_));
  AOI21X1  g01804(.A0(new_n4224_), .A1(pi0075), .B0(pi0092), .Y(new_n4240_));
  NOR2X1   g01805(.A(new_n4237_), .B(new_n3101_), .Y(new_n4241_));
  OAI21X1  g01806(.A0(new_n4236_), .A1(new_n3098_), .B0(pi0092), .Y(new_n4242_));
  OAI21X1  g01807(.A0(new_n4242_), .A1(new_n4241_), .B0(new_n3135_), .Y(new_n4243_));
  AOI21X1  g01808(.A0(new_n4240_), .A1(new_n4239_), .B0(new_n4243_), .Y(new_n4244_));
  OAI21X1  g01809(.A0(new_n4236_), .A1(new_n3135_), .B0(new_n3128_), .Y(new_n4245_));
  OR4X1    g01810(.A(new_n4214_), .B(new_n4173_), .C(new_n3810_), .D(new_n3066_), .Y(new_n4246_));
  AOI21X1  g01811(.A0(new_n4222_), .A1(new_n3131_), .B0(new_n3128_), .Y(new_n4247_));
  AOI21X1  g01812(.A0(new_n4247_), .A1(new_n4246_), .B0(pi0056), .Y(new_n4248_));
  OAI21X1  g01813(.A0(new_n4245_), .A1(new_n4244_), .B0(new_n4248_), .Y(new_n4249_));
  OAI21X1  g01814(.A0(new_n4214_), .A1(new_n4173_), .B0(new_n3140_), .Y(new_n4250_));
  AOI21X1  g01815(.A0(new_n4223_), .A1(new_n3242_), .B0(new_n3143_), .Y(new_n4251_));
  AOI21X1  g01816(.A0(new_n4251_), .A1(new_n4250_), .B0(pi0062), .Y(new_n4252_));
  NOR3X1   g01817(.A(new_n4214_), .B(new_n4173_), .C(new_n3249_), .Y(new_n4253_));
  OAI21X1  g01818(.A0(new_n4223_), .A1(new_n3248_), .B0(pi0062), .Y(new_n4254_));
  NOR3X1   g01819(.A(pi0246), .B(pi0059), .C(pi0057), .Y(new_n4255_));
  OAI21X1  g01820(.A0(new_n4254_), .A1(new_n4253_), .B0(new_n4255_), .Y(new_n4256_));
  AOI21X1  g01821(.A0(new_n4252_), .A1(new_n4249_), .B0(new_n4256_), .Y(new_n4257_));
  OAI21X1  g01822(.A0(new_n3531_), .A1(pi0877), .B0(new_n4210_), .Y(new_n4258_));
  AOI21X1  g01823(.A0(new_n3532_), .A1(new_n4180_), .B0(new_n4210_), .Y(new_n4259_));
  OAI21X1  g01824(.A0(new_n3535_), .A1(new_n4180_), .B0(new_n4259_), .Y(new_n4260_));
  AOI21X1  g01825(.A0(new_n4260_), .A1(new_n4258_), .B0(pi0228), .Y(new_n4261_));
  OAI21X1  g01826(.A0(new_n3258_), .A1(new_n3030_), .B0(new_n4208_), .Y(new_n4262_));
  OAI21X1  g01827(.A0(new_n4262_), .A1(new_n4261_), .B0(new_n4178_), .Y(new_n4263_));
  AOI21X1  g01828(.A0(new_n4263_), .A1(new_n4177_), .B0(pi0215), .Y(new_n4264_));
  OAI21X1  g01829(.A0(new_n4264_), .A1(new_n4174_), .B0(new_n4202_), .Y(new_n4265_));
  AND2X1   g01830(.A(new_n4207_), .B(new_n3831_), .Y(new_n4266_));
  NAND3X1  g01831(.A(new_n4187_), .B(new_n3479_), .C(new_n2438_), .Y(new_n4267_));
  OAI21X1  g01832(.A0(new_n4267_), .A1(new_n4212_), .B0(new_n4178_), .Y(new_n4268_));
  AOI21X1  g01833(.A0(new_n4268_), .A1(new_n4177_), .B0(pi0215), .Y(new_n4269_));
  OAI21X1  g01834(.A0(new_n4269_), .A1(new_n4173_), .B0(pi0299), .Y(new_n4270_));
  NAND2X1  g01835(.A(new_n4270_), .B(new_n4266_), .Y(new_n4271_));
  AOI21X1  g01836(.A0(new_n4271_), .A1(pi0039), .B0(pi0038), .Y(new_n4272_));
  INVX1    g01837(.A(new_n4266_), .Y(new_n4273_));
  AOI21X1  g01838(.A0(pi0269), .A1(pi0216), .B0(new_n3548_), .Y(new_n4274_));
  NOR2X1   g01839(.A(new_n4274_), .B(new_n4223_), .Y(new_n4275_));
  INVX1    g01840(.A(new_n4275_), .Y(new_n4276_));
  AOI21X1  g01841(.A0(new_n4276_), .A1(pi0299), .B0(new_n4273_), .Y(new_n4277_));
  INVX1    g01842(.A(new_n4277_), .Y(new_n4278_));
  OAI21X1  g01843(.A0(new_n4278_), .A1(new_n2996_), .B0(new_n3026_), .Y(new_n4279_));
  AOI21X1  g01844(.A0(new_n4272_), .A1(new_n4265_), .B0(new_n4279_), .Y(new_n4280_));
  INVX1    g01845(.A(pi1138), .Y(new_n4281_));
  NAND3X1  g01846(.A(new_n4229_), .B(new_n4208_), .C(new_n3479_), .Y(new_n4282_));
  AOI21X1  g01847(.A0(new_n4282_), .A1(new_n4178_), .B0(new_n4227_), .Y(new_n4283_));
  MX2X1    g01848(.A(new_n4283_), .B(new_n4281_), .S0(pi0215), .Y(new_n4284_));
  AND2X1   g01849(.A(new_n4266_), .B(new_n3065_), .Y(new_n4285_));
  OAI21X1  g01850(.A0(new_n4284_), .A1(new_n2953_), .B0(new_n4285_), .Y(new_n4286_));
  AOI21X1  g01851(.A0(new_n4277_), .A1(new_n3066_), .B0(new_n3026_), .Y(new_n4287_));
  AND2X1   g01852(.A(new_n4287_), .B(new_n4286_), .Y(new_n4288_));
  OAI21X1  g01853(.A0(new_n4288_), .A1(new_n4280_), .B0(new_n3156_), .Y(new_n4289_));
  MX2X1    g01854(.A(new_n4278_), .B(new_n4271_), .S0(new_n3085_), .Y(new_n4290_));
  AOI21X1  g01855(.A0(new_n4290_), .A1(pi0087), .B0(pi0075), .Y(new_n4291_));
  OAI21X1  g01856(.A0(new_n4278_), .A1(new_n3095_), .B0(new_n3100_), .Y(new_n4292_));
  AOI21X1  g01857(.A0(new_n4291_), .A1(new_n4289_), .B0(new_n4292_), .Y(new_n4293_));
  OR2X1    g01858(.A(new_n4290_), .B(new_n3101_), .Y(new_n4294_));
  AOI21X1  g01859(.A0(new_n4277_), .A1(new_n3101_), .B0(new_n3100_), .Y(new_n4295_));
  AND2X1   g01860(.A(new_n4295_), .B(new_n4294_), .Y(new_n4296_));
  NOR3X1   g01861(.A(new_n4296_), .B(new_n4293_), .C(new_n3136_), .Y(new_n4297_));
  OAI21X1  g01862(.A0(new_n4278_), .A1(new_n3135_), .B0(new_n3128_), .Y(new_n4298_));
  OR4X1    g01863(.A(new_n4269_), .B(new_n4173_), .C(new_n3810_), .D(new_n3066_), .Y(new_n4299_));
  AOI21X1  g01864(.A0(new_n4275_), .A1(new_n3131_), .B0(new_n3128_), .Y(new_n4300_));
  AOI21X1  g01865(.A0(new_n4300_), .A1(new_n4299_), .B0(pi0056), .Y(new_n4301_));
  OAI21X1  g01866(.A0(new_n4298_), .A1(new_n4297_), .B0(new_n4301_), .Y(new_n4302_));
  OAI21X1  g01867(.A0(new_n4269_), .A1(new_n4173_), .B0(new_n3140_), .Y(new_n4303_));
  AOI21X1  g01868(.A0(new_n4276_), .A1(new_n3242_), .B0(new_n3143_), .Y(new_n4304_));
  AOI21X1  g01869(.A0(new_n4304_), .A1(new_n4303_), .B0(pi0062), .Y(new_n4305_));
  NOR3X1   g01870(.A(new_n4269_), .B(new_n4173_), .C(new_n3249_), .Y(new_n4306_));
  OAI21X1  g01871(.A0(new_n4276_), .A1(new_n3248_), .B0(pi0062), .Y(new_n4307_));
  AND2X1   g01872(.A(new_n3246_), .B(pi0246), .Y(new_n4308_));
  OAI21X1  g01873(.A0(new_n4307_), .A1(new_n4306_), .B0(new_n4308_), .Y(new_n4309_));
  AOI21X1  g01874(.A0(new_n4305_), .A1(new_n4302_), .B0(new_n4309_), .Y(new_n4310_));
  AOI21X1  g01875(.A0(new_n4274_), .A1(pi0246), .B0(new_n3246_), .Y(new_n4311_));
  AND2X1   g01876(.A(new_n4311_), .B(new_n4222_), .Y(new_n4312_));
  NOR3X1   g01877(.A(new_n4312_), .B(new_n4310_), .C(new_n4257_), .Y(po0161));
  AND2X1   g01878(.A(pi1137), .B(pi0215), .Y(new_n4314_));
  OR2X1    g01879(.A(new_n4314_), .B(new_n2953_), .Y(new_n4315_));
  INVX1    g01880(.A(pi0933), .Y(new_n4316_));
  AOI21X1  g01881(.A0(new_n2442_), .A1(new_n4316_), .B0(new_n2437_), .Y(new_n4317_));
  OAI21X1  g01882(.A0(new_n2442_), .A1(pi1137), .B0(new_n4317_), .Y(new_n4318_));
  AOI21X1  g01883(.A0(pi0280), .A1(pi0216), .B0(pi0221), .Y(new_n4319_));
  INVX1    g01884(.A(new_n4319_), .Y(new_n4320_));
  INVX1    g01885(.A(pi0878), .Y(new_n4321_));
  AOI21X1  g01886(.A0(new_n3271_), .A1(pi0878), .B0(pi0168), .Y(new_n4322_));
  AOI21X1  g01887(.A0(new_n3266_), .A1(pi0168), .B0(new_n4322_), .Y(new_n4323_));
  NAND2X1  g01888(.A(new_n4322_), .B(new_n3204_), .Y(new_n4324_));
  OAI21X1  g01889(.A0(new_n4323_), .A1(new_n4321_), .B0(new_n4324_), .Y(new_n4325_));
  AOI21X1  g01890(.A0(new_n2454_), .A1(pi0095), .B0(new_n4321_), .Y(new_n4326_));
  AOI21X1  g01891(.A0(pi0168), .A1(new_n2448_), .B0(new_n3013_), .Y(new_n4327_));
  OAI21X1  g01892(.A0(new_n4326_), .A1(new_n2448_), .B0(new_n4327_), .Y(new_n4328_));
  OAI21X1  g01893(.A0(new_n4328_), .A1(new_n3270_), .B0(new_n2438_), .Y(new_n4329_));
  AOI21X1  g01894(.A0(new_n4325_), .A1(new_n3013_), .B0(new_n4329_), .Y(new_n4330_));
  OAI21X1  g01895(.A0(new_n4330_), .A1(new_n4320_), .B0(new_n4318_), .Y(new_n4331_));
  AOI21X1  g01896(.A0(new_n4331_), .A1(new_n2954_), .B0(new_n4315_), .Y(new_n4332_));
  AOI21X1  g01897(.A0(pi1137), .A1(pi0223), .B0(pi0299), .Y(new_n4333_));
  INVX1    g01898(.A(new_n4333_), .Y(new_n4334_));
  AOI21X1  g01899(.A0(new_n3159_), .A1(new_n4316_), .B0(new_n2960_), .Y(new_n4335_));
  OAI21X1  g01900(.A0(new_n3159_), .A1(pi1137), .B0(new_n4335_), .Y(new_n4336_));
  AOI21X1  g01901(.A0(pi0280), .A1(pi0224), .B0(pi0222), .Y(new_n4337_));
  INVX1    g01902(.A(new_n4337_), .Y(new_n4338_));
  AOI21X1  g01903(.A0(new_n3258_), .A1(pi0878), .B0(pi0224), .Y(new_n4339_));
  OAI21X1  g01904(.A0(new_n4339_), .A1(new_n4338_), .B0(new_n4336_), .Y(new_n4340_));
  NOR2X1   g01905(.A(new_n4338_), .B(new_n3258_), .Y(new_n4341_));
  OAI21X1  g01906(.A0(new_n4341_), .A1(new_n4340_), .B0(new_n2964_), .Y(new_n4342_));
  AOI21X1  g01907(.A0(new_n4342_), .A1(new_n4333_), .B0(pi0039), .Y(new_n4343_));
  OAI21X1  g01908(.A0(new_n4340_), .A1(new_n4334_), .B0(new_n4343_), .Y(new_n4344_));
  AND2X1   g01909(.A(pi1137), .B(pi0223), .Y(new_n4345_));
  OAI21X1  g01910(.A0(new_n4326_), .A1(pi0224), .B0(new_n4337_), .Y(new_n4346_));
  AOI21X1  g01911(.A0(new_n4346_), .A1(new_n4336_), .B0(pi0223), .Y(new_n4347_));
  OAI21X1  g01912(.A0(new_n4347_), .A1(new_n4345_), .B0(new_n2953_), .Y(new_n4348_));
  AND2X1   g01913(.A(new_n4328_), .B(new_n2438_), .Y(new_n4349_));
  INVX1    g01914(.A(new_n4349_), .Y(new_n4350_));
  INVX1    g01915(.A(pi0168), .Y(new_n4351_));
  OAI21X1  g01916(.A0(new_n3630_), .A1(new_n4351_), .B0(new_n3013_), .Y(new_n4352_));
  AOI21X1  g01917(.A0(new_n3630_), .A1(new_n4321_), .B0(new_n4352_), .Y(new_n4353_));
  OAI21X1  g01918(.A0(new_n4353_), .A1(new_n4350_), .B0(new_n4319_), .Y(new_n4354_));
  AOI21X1  g01919(.A0(new_n4354_), .A1(new_n4318_), .B0(pi0215), .Y(new_n4355_));
  OAI21X1  g01920(.A0(new_n4355_), .A1(new_n4314_), .B0(pi0299), .Y(new_n4356_));
  NAND2X1  g01921(.A(new_n4356_), .B(new_n4348_), .Y(new_n4357_));
  AOI21X1  g01922(.A0(new_n4357_), .A1(pi0039), .B0(pi0038), .Y(new_n4358_));
  OAI21X1  g01923(.A0(new_n4344_), .A1(new_n4332_), .B0(new_n4358_), .Y(new_n4359_));
  INVX1    g01924(.A(new_n4348_), .Y(new_n4360_));
  AOI21X1  g01925(.A0(new_n3013_), .A1(new_n4351_), .B0(new_n4350_), .Y(new_n4361_));
  OAI21X1  g01926(.A0(new_n4361_), .A1(new_n4320_), .B0(new_n4318_), .Y(new_n4362_));
  AOI21X1  g01927(.A0(new_n4362_), .A1(new_n2954_), .B0(new_n4314_), .Y(new_n4363_));
  INVX1    g01928(.A(new_n4363_), .Y(new_n4364_));
  AOI21X1  g01929(.A0(new_n4364_), .A1(pi0299), .B0(new_n4360_), .Y(new_n4365_));
  AOI21X1  g01930(.A0(new_n4365_), .A1(pi0038), .B0(pi0100), .Y(new_n4366_));
  INVX1    g01931(.A(new_n4314_), .Y(new_n4367_));
  INVX1    g01932(.A(new_n4318_), .Y(new_n4368_));
  AOI21X1  g01933(.A0(new_n3221_), .A1(pi0168), .B0(pi0228), .Y(new_n4369_));
  OAI21X1  g01934(.A0(new_n3221_), .A1(pi0878), .B0(new_n4369_), .Y(new_n4370_));
  AOI21X1  g01935(.A0(new_n4370_), .A1(new_n4349_), .B0(new_n4320_), .Y(new_n4371_));
  OAI21X1  g01936(.A0(new_n4371_), .A1(new_n4368_), .B0(new_n2954_), .Y(new_n4372_));
  AOI21X1  g01937(.A0(new_n4372_), .A1(new_n4367_), .B0(new_n2953_), .Y(new_n4373_));
  OR4X1    g01938(.A(new_n4373_), .B(new_n4360_), .C(pi0039), .D(pi0038), .Y(new_n4374_));
  AOI21X1  g01939(.A0(new_n4365_), .A1(new_n3066_), .B0(new_n3026_), .Y(new_n4375_));
  AOI22X1  g01940(.A0(new_n4375_), .A1(new_n4374_), .B0(new_n4366_), .B1(new_n4359_), .Y(new_n4376_));
  INVX1    g01941(.A(new_n4365_), .Y(new_n4377_));
  MX2X1    g01942(.A(new_n4377_), .B(new_n4357_), .S0(new_n3085_), .Y(new_n4378_));
  AOI21X1  g01943(.A0(new_n4378_), .A1(pi0087), .B0(pi0075), .Y(new_n4379_));
  OAI21X1  g01944(.A0(new_n4376_), .A1(pi0087), .B0(new_n4379_), .Y(new_n4380_));
  AOI21X1  g01945(.A0(new_n4365_), .A1(pi0075), .B0(pi0092), .Y(new_n4381_));
  NOR2X1   g01946(.A(new_n4378_), .B(new_n3101_), .Y(new_n4382_));
  OAI21X1  g01947(.A0(new_n4377_), .A1(new_n3098_), .B0(pi0092), .Y(new_n4383_));
  OAI21X1  g01948(.A0(new_n4383_), .A1(new_n4382_), .B0(new_n3135_), .Y(new_n4384_));
  AOI21X1  g01949(.A0(new_n4381_), .A1(new_n4380_), .B0(new_n4384_), .Y(new_n4385_));
  OAI21X1  g01950(.A0(new_n4377_), .A1(new_n3135_), .B0(new_n3128_), .Y(new_n4386_));
  OR4X1    g01951(.A(new_n4355_), .B(new_n4314_), .C(new_n3810_), .D(new_n3066_), .Y(new_n4387_));
  AOI21X1  g01952(.A0(new_n4363_), .A1(new_n3131_), .B0(new_n3128_), .Y(new_n4388_));
  AOI21X1  g01953(.A0(new_n4388_), .A1(new_n4387_), .B0(pi0056), .Y(new_n4389_));
  OAI21X1  g01954(.A0(new_n4386_), .A1(new_n4385_), .B0(new_n4389_), .Y(new_n4390_));
  OAI21X1  g01955(.A0(new_n4355_), .A1(new_n4314_), .B0(new_n3140_), .Y(new_n4391_));
  AOI21X1  g01956(.A0(new_n4364_), .A1(new_n3242_), .B0(new_n3143_), .Y(new_n4392_));
  AOI21X1  g01957(.A0(new_n4392_), .A1(new_n4391_), .B0(pi0062), .Y(new_n4393_));
  NOR3X1   g01958(.A(new_n4355_), .B(new_n4314_), .C(new_n3249_), .Y(new_n4394_));
  OAI21X1  g01959(.A0(new_n4364_), .A1(new_n3248_), .B0(pi0062), .Y(new_n4395_));
  NOR3X1   g01960(.A(pi0240), .B(pi0059), .C(pi0057), .Y(new_n4396_));
  OAI21X1  g01961(.A0(new_n4395_), .A1(new_n4394_), .B0(new_n4396_), .Y(new_n4397_));
  AOI21X1  g01962(.A0(new_n4393_), .A1(new_n4390_), .B0(new_n4397_), .Y(new_n4398_));
  OAI21X1  g01963(.A0(new_n3531_), .A1(pi0878), .B0(new_n4351_), .Y(new_n4399_));
  AOI21X1  g01964(.A0(new_n3532_), .A1(new_n4321_), .B0(new_n4351_), .Y(new_n4400_));
  OAI21X1  g01965(.A0(new_n3535_), .A1(new_n4321_), .B0(new_n4400_), .Y(new_n4401_));
  AOI21X1  g01966(.A0(new_n4401_), .A1(new_n4399_), .B0(pi0228), .Y(new_n4402_));
  OAI21X1  g01967(.A0(new_n3258_), .A1(new_n3030_), .B0(new_n4349_), .Y(new_n4403_));
  OAI21X1  g01968(.A0(new_n4403_), .A1(new_n4402_), .B0(new_n4319_), .Y(new_n4404_));
  AOI21X1  g01969(.A0(new_n4404_), .A1(new_n4318_), .B0(pi0215), .Y(new_n4405_));
  OAI21X1  g01970(.A0(new_n4405_), .A1(new_n4315_), .B0(new_n4343_), .Y(new_n4406_));
  AND2X1   g01971(.A(new_n4348_), .B(new_n3831_), .Y(new_n4407_));
  NAND3X1  g01972(.A(new_n4328_), .B(new_n3479_), .C(new_n2438_), .Y(new_n4408_));
  OAI21X1  g01973(.A0(new_n4408_), .A1(new_n4353_), .B0(new_n4319_), .Y(new_n4409_));
  AOI21X1  g01974(.A0(new_n4409_), .A1(new_n4318_), .B0(pi0215), .Y(new_n4410_));
  OAI21X1  g01975(.A0(new_n4410_), .A1(new_n4314_), .B0(pi0299), .Y(new_n4411_));
  NAND2X1  g01976(.A(new_n4411_), .B(new_n4407_), .Y(new_n4412_));
  AOI21X1  g01977(.A0(new_n4412_), .A1(pi0039), .B0(pi0038), .Y(new_n4413_));
  INVX1    g01978(.A(new_n4407_), .Y(new_n4414_));
  AOI21X1  g01979(.A0(pi0280), .A1(pi0216), .B0(new_n3548_), .Y(new_n4415_));
  NOR2X1   g01980(.A(new_n4415_), .B(new_n4364_), .Y(new_n4416_));
  INVX1    g01981(.A(new_n4416_), .Y(new_n4417_));
  AOI21X1  g01982(.A0(new_n4417_), .A1(pi0299), .B0(new_n4414_), .Y(new_n4418_));
  INVX1    g01983(.A(new_n4418_), .Y(new_n4419_));
  OAI21X1  g01984(.A0(new_n4419_), .A1(new_n2996_), .B0(new_n3026_), .Y(new_n4420_));
  AOI21X1  g01985(.A0(new_n4413_), .A1(new_n4406_), .B0(new_n4420_), .Y(new_n4421_));
  INVX1    g01986(.A(pi1137), .Y(new_n4422_));
  NAND3X1  g01987(.A(new_n4370_), .B(new_n4349_), .C(new_n3479_), .Y(new_n4423_));
  AOI21X1  g01988(.A0(new_n4423_), .A1(new_n4319_), .B0(new_n4368_), .Y(new_n4424_));
  MX2X1    g01989(.A(new_n4424_), .B(new_n4422_), .S0(pi0215), .Y(new_n4425_));
  AND2X1   g01990(.A(new_n4407_), .B(new_n3065_), .Y(new_n4426_));
  OAI21X1  g01991(.A0(new_n4425_), .A1(new_n2953_), .B0(new_n4426_), .Y(new_n4427_));
  AOI21X1  g01992(.A0(new_n4418_), .A1(new_n3066_), .B0(new_n3026_), .Y(new_n4428_));
  AND2X1   g01993(.A(new_n4428_), .B(new_n4427_), .Y(new_n4429_));
  OAI21X1  g01994(.A0(new_n4429_), .A1(new_n4421_), .B0(new_n3156_), .Y(new_n4430_));
  MX2X1    g01995(.A(new_n4419_), .B(new_n4412_), .S0(new_n3085_), .Y(new_n4431_));
  AOI21X1  g01996(.A0(new_n4431_), .A1(pi0087), .B0(pi0075), .Y(new_n4432_));
  OAI21X1  g01997(.A0(new_n4419_), .A1(new_n3095_), .B0(new_n3100_), .Y(new_n4433_));
  AOI21X1  g01998(.A0(new_n4432_), .A1(new_n4430_), .B0(new_n4433_), .Y(new_n4434_));
  OR2X1    g01999(.A(new_n4431_), .B(new_n3101_), .Y(new_n4435_));
  AOI21X1  g02000(.A0(new_n4418_), .A1(new_n3101_), .B0(new_n3100_), .Y(new_n4436_));
  AND2X1   g02001(.A(new_n4436_), .B(new_n4435_), .Y(new_n4437_));
  NOR3X1   g02002(.A(new_n4437_), .B(new_n4434_), .C(new_n3136_), .Y(new_n4438_));
  OAI21X1  g02003(.A0(new_n4419_), .A1(new_n3135_), .B0(new_n3128_), .Y(new_n4439_));
  OR4X1    g02004(.A(new_n4410_), .B(new_n4314_), .C(new_n3810_), .D(new_n3066_), .Y(new_n4440_));
  AOI21X1  g02005(.A0(new_n4416_), .A1(new_n3131_), .B0(new_n3128_), .Y(new_n4441_));
  AOI21X1  g02006(.A0(new_n4441_), .A1(new_n4440_), .B0(pi0056), .Y(new_n4442_));
  OAI21X1  g02007(.A0(new_n4439_), .A1(new_n4438_), .B0(new_n4442_), .Y(new_n4443_));
  OAI21X1  g02008(.A0(new_n4410_), .A1(new_n4314_), .B0(new_n3140_), .Y(new_n4444_));
  AOI21X1  g02009(.A0(new_n4417_), .A1(new_n3242_), .B0(new_n3143_), .Y(new_n4445_));
  AOI21X1  g02010(.A0(new_n4445_), .A1(new_n4444_), .B0(pi0062), .Y(new_n4446_));
  NOR3X1   g02011(.A(new_n4410_), .B(new_n4314_), .C(new_n3249_), .Y(new_n4447_));
  OAI21X1  g02012(.A0(new_n4417_), .A1(new_n3248_), .B0(pi0062), .Y(new_n4448_));
  AND2X1   g02013(.A(new_n3246_), .B(pi0240), .Y(new_n4449_));
  OAI21X1  g02014(.A0(new_n4448_), .A1(new_n4447_), .B0(new_n4449_), .Y(new_n4450_));
  AOI21X1  g02015(.A0(new_n4446_), .A1(new_n4443_), .B0(new_n4450_), .Y(new_n4451_));
  AOI21X1  g02016(.A0(new_n4415_), .A1(pi0240), .B0(new_n3246_), .Y(new_n4452_));
  AND2X1   g02017(.A(new_n4452_), .B(new_n4363_), .Y(new_n4453_));
  NOR3X1   g02018(.A(new_n4453_), .B(new_n4451_), .C(new_n4398_), .Y(po0162));
  INVX1    g02019(.A(pi0928), .Y(new_n4455_));
  AOI21X1  g02020(.A0(new_n2442_), .A1(new_n4455_), .B0(new_n2437_), .Y(new_n4456_));
  OAI21X1  g02021(.A0(new_n2442_), .A1(pi1136), .B0(new_n4456_), .Y(new_n4457_));
  AND2X1   g02022(.A(pi0266), .B(pi0216), .Y(new_n4458_));
  OAI21X1  g02023(.A0(new_n3258_), .A1(new_n2448_), .B0(pi0228), .Y(new_n4459_));
  INVX1    g02024(.A(pi0875), .Y(new_n4460_));
  AOI21X1  g02025(.A0(new_n2454_), .A1(pi0095), .B0(new_n4460_), .Y(new_n4461_));
  MX2X1    g02026(.A(new_n4461_), .B(pi0166), .S0(new_n2448_), .Y(new_n4462_));
  OAI21X1  g02027(.A0(new_n4462_), .A1(new_n4459_), .B0(new_n2438_), .Y(new_n4463_));
  INVX1    g02028(.A(pi0166), .Y(new_n4464_));
  OAI21X1  g02029(.A0(new_n3532_), .A1(new_n4464_), .B0(pi0875), .Y(new_n4465_));
  AOI21X1  g02030(.A0(new_n3531_), .A1(new_n4464_), .B0(new_n4465_), .Y(new_n4466_));
  NOR3X1   g02031(.A(new_n3535_), .B(pi0875), .C(new_n4464_), .Y(new_n4467_));
  OAI21X1  g02032(.A0(new_n4467_), .A1(new_n4466_), .B0(new_n3013_), .Y(new_n4468_));
  AOI21X1  g02033(.A0(new_n4468_), .A1(new_n4459_), .B0(new_n4463_), .Y(new_n4469_));
  OAI21X1  g02034(.A0(new_n4469_), .A1(new_n4458_), .B0(new_n2437_), .Y(new_n4470_));
  AOI21X1  g02035(.A0(new_n4470_), .A1(new_n4457_), .B0(pi0215), .Y(new_n4471_));
  AND2X1   g02036(.A(pi1136), .B(pi0215), .Y(new_n4472_));
  NOR2X1   g02037(.A(new_n4472_), .B(new_n2953_), .Y(new_n4473_));
  INVX1    g02038(.A(new_n4473_), .Y(new_n4474_));
  NOR3X1   g02039(.A(new_n2455_), .B(pi0875), .C(pi0224), .Y(new_n4475_));
  OAI21X1  g02040(.A0(pi0266), .A1(new_n2961_), .B0(new_n2960_), .Y(new_n4476_));
  OR2X1    g02041(.A(new_n4476_), .B(new_n4475_), .Y(new_n4477_));
  NOR2X1   g02042(.A(new_n3258_), .B(new_n2971_), .Y(new_n4478_));
  AOI21X1  g02043(.A0(new_n3159_), .A1(new_n4455_), .B0(new_n2960_), .Y(new_n4479_));
  OAI21X1  g02044(.A0(new_n3159_), .A1(pi1136), .B0(new_n4479_), .Y(new_n4480_));
  AOI21X1  g02045(.A0(pi1136), .A1(pi0223), .B0(pi0299), .Y(new_n4481_));
  AND2X1   g02046(.A(new_n4481_), .B(new_n4480_), .Y(new_n4482_));
  OAI21X1  g02047(.A0(new_n4478_), .A1(new_n4477_), .B0(new_n4482_), .Y(new_n4483_));
  NAND2X1  g02048(.A(new_n4480_), .B(new_n4477_), .Y(new_n4484_));
  NOR2X1   g02049(.A(new_n4484_), .B(new_n4478_), .Y(new_n4485_));
  OAI21X1  g02050(.A0(new_n4485_), .A1(pi0223), .B0(new_n4481_), .Y(new_n4486_));
  AND2X1   g02051(.A(new_n4486_), .B(new_n2959_), .Y(new_n4487_));
  AND2X1   g02052(.A(new_n4487_), .B(new_n4483_), .Y(new_n4488_));
  OAI21X1  g02053(.A0(new_n4474_), .A1(new_n4471_), .B0(new_n4488_), .Y(new_n4489_));
  AND2X1   g02054(.A(pi1136), .B(pi0223), .Y(new_n4490_));
  AOI21X1  g02055(.A0(new_n4480_), .A1(new_n4477_), .B0(pi0223), .Y(new_n4491_));
  OAI21X1  g02056(.A0(new_n4491_), .A1(new_n4490_), .B0(new_n2953_), .Y(new_n4492_));
  INVX1    g02057(.A(new_n4492_), .Y(new_n4493_));
  OAI21X1  g02058(.A0(new_n4461_), .A1(new_n3009_), .B0(new_n4493_), .Y(new_n4494_));
  AND2X1   g02059(.A(new_n4462_), .B(pi0228), .Y(new_n4495_));
  INVX1    g02060(.A(new_n4495_), .Y(new_n4496_));
  AOI21X1  g02061(.A0(new_n3630_), .A1(new_n4460_), .B0(pi0228), .Y(new_n4497_));
  OAI21X1  g02062(.A0(new_n3630_), .A1(pi0166), .B0(new_n4497_), .Y(new_n4498_));
  AOI21X1  g02063(.A0(new_n4498_), .A1(new_n4496_), .B0(pi0216), .Y(new_n4499_));
  OAI21X1  g02064(.A0(new_n4499_), .A1(new_n4458_), .B0(new_n2437_), .Y(new_n4500_));
  AOI21X1  g02065(.A0(new_n4500_), .A1(new_n4457_), .B0(pi0215), .Y(new_n4501_));
  OAI21X1  g02066(.A0(new_n4501_), .A1(new_n4472_), .B0(pi0299), .Y(new_n4502_));
  NAND2X1  g02067(.A(new_n4502_), .B(new_n4494_), .Y(new_n4503_));
  AOI21X1  g02068(.A0(new_n4503_), .A1(pi0039), .B0(pi0038), .Y(new_n4504_));
  INVX1    g02069(.A(pi0266), .Y(new_n4505_));
  AOI21X1  g02070(.A0(new_n3013_), .A1(pi0166), .B0(new_n4495_), .Y(new_n4506_));
  MX2X1    g02071(.A(new_n4506_), .B(new_n4505_), .S0(pi0216), .Y(new_n4507_));
  OAI21X1  g02072(.A0(new_n4507_), .A1(pi0221), .B0(new_n4457_), .Y(new_n4508_));
  AOI21X1  g02073(.A0(new_n4508_), .A1(new_n2954_), .B0(new_n4472_), .Y(new_n4509_));
  OAI21X1  g02074(.A0(new_n4509_), .A1(new_n2953_), .B0(new_n4494_), .Y(new_n4510_));
  OAI21X1  g02075(.A0(new_n4510_), .A1(new_n2996_), .B0(new_n3026_), .Y(new_n4511_));
  AOI21X1  g02076(.A0(new_n4504_), .A1(new_n4489_), .B0(new_n4511_), .Y(new_n4512_));
  AOI21X1  g02077(.A0(new_n3213_), .A1(new_n4460_), .B0(new_n4464_), .Y(new_n4513_));
  INVX1    g02078(.A(new_n4513_), .Y(new_n4514_));
  NOR2X1   g02079(.A(pi0161), .B(pi0152), .Y(new_n4515_));
  AOI21X1  g02080(.A0(new_n3497_), .A1(new_n4515_), .B0(new_n4460_), .Y(new_n4516_));
  OAI21X1  g02081(.A0(new_n3213_), .A1(new_n4515_), .B0(new_n4516_), .Y(new_n4517_));
  AOI21X1  g02082(.A0(new_n4517_), .A1(new_n4514_), .B0(pi0228), .Y(new_n4518_));
  OR2X1    g02083(.A(new_n4518_), .B(new_n4495_), .Y(new_n4519_));
  AOI21X1  g02084(.A0(new_n4519_), .A1(new_n2438_), .B0(new_n4458_), .Y(new_n4520_));
  OAI21X1  g02085(.A0(new_n4520_), .A1(pi0221), .B0(new_n4457_), .Y(new_n4521_));
  AOI21X1  g02086(.A0(new_n4521_), .A1(new_n2954_), .B0(new_n4472_), .Y(new_n4522_));
  AND2X1   g02087(.A(new_n4494_), .B(new_n3065_), .Y(new_n4523_));
  OAI21X1  g02088(.A0(new_n4522_), .A1(new_n2953_), .B0(new_n4523_), .Y(new_n4524_));
  INVX1    g02089(.A(new_n4510_), .Y(new_n4525_));
  AOI21X1  g02090(.A0(new_n4525_), .A1(new_n3066_), .B0(new_n3026_), .Y(new_n4526_));
  AND2X1   g02091(.A(new_n4526_), .B(new_n4524_), .Y(new_n4527_));
  OAI21X1  g02092(.A0(new_n4527_), .A1(new_n4512_), .B0(new_n3156_), .Y(new_n4528_));
  MX2X1    g02093(.A(new_n4510_), .B(new_n4503_), .S0(new_n3085_), .Y(new_n4529_));
  AOI21X1  g02094(.A0(new_n4529_), .A1(pi0087), .B0(pi0075), .Y(new_n4530_));
  OAI21X1  g02095(.A0(new_n4510_), .A1(new_n3095_), .B0(new_n3100_), .Y(new_n4531_));
  AOI21X1  g02096(.A0(new_n4530_), .A1(new_n4528_), .B0(new_n4531_), .Y(new_n4532_));
  OR2X1    g02097(.A(new_n4529_), .B(new_n3101_), .Y(new_n4533_));
  AOI21X1  g02098(.A0(new_n4525_), .A1(new_n3101_), .B0(new_n3100_), .Y(new_n4534_));
  AND2X1   g02099(.A(new_n4534_), .B(new_n4533_), .Y(new_n4535_));
  NOR3X1   g02100(.A(new_n4535_), .B(new_n4532_), .C(new_n3136_), .Y(new_n4536_));
  OAI21X1  g02101(.A0(new_n4510_), .A1(new_n3135_), .B0(new_n3128_), .Y(new_n4537_));
  OR4X1    g02102(.A(new_n4501_), .B(new_n4472_), .C(new_n3810_), .D(new_n3066_), .Y(new_n4538_));
  AOI21X1  g02103(.A0(new_n4509_), .A1(new_n3131_), .B0(new_n3128_), .Y(new_n4539_));
  AOI21X1  g02104(.A0(new_n4539_), .A1(new_n4538_), .B0(pi0056), .Y(new_n4540_));
  OAI21X1  g02105(.A0(new_n4537_), .A1(new_n4536_), .B0(new_n4540_), .Y(new_n4541_));
  OAI21X1  g02106(.A0(new_n4501_), .A1(new_n4472_), .B0(new_n3140_), .Y(new_n4542_));
  INVX1    g02107(.A(new_n4509_), .Y(new_n4543_));
  AOI21X1  g02108(.A0(new_n4543_), .A1(new_n3242_), .B0(new_n3143_), .Y(new_n4544_));
  AOI21X1  g02109(.A0(new_n4544_), .A1(new_n4542_), .B0(pi0062), .Y(new_n4545_));
  NOR3X1   g02110(.A(new_n4501_), .B(new_n4472_), .C(new_n3249_), .Y(new_n4546_));
  OAI21X1  g02111(.A0(new_n4543_), .A1(new_n3248_), .B0(pi0062), .Y(new_n4547_));
  OAI21X1  g02112(.A0(new_n4547_), .A1(new_n4546_), .B0(new_n3246_), .Y(new_n4548_));
  AOI21X1  g02113(.A0(new_n4545_), .A1(new_n4541_), .B0(new_n4548_), .Y(new_n4549_));
  INVX1    g02114(.A(pi0245), .Y(new_n4550_));
  OAI21X1  g02115(.A0(new_n4543_), .A1(new_n3246_), .B0(new_n4550_), .Y(new_n4551_));
  INVX1    g02116(.A(new_n4457_), .Y(new_n4552_));
  INVX1    g02117(.A(new_n4458_), .Y(new_n4553_));
  OAI21X1  g02118(.A0(new_n3271_), .A1(pi0166), .B0(new_n4460_), .Y(new_n4554_));
  AOI21X1  g02119(.A0(new_n3266_), .A1(pi0166), .B0(new_n4554_), .Y(new_n4555_));
  AOI21X1  g02120(.A0(new_n3204_), .A1(new_n4464_), .B0(new_n4460_), .Y(new_n4556_));
  NOR3X1   g02121(.A(new_n4556_), .B(new_n4555_), .C(pi0228), .Y(new_n4557_));
  OAI21X1  g02122(.A0(new_n4557_), .A1(new_n4463_), .B0(new_n4553_), .Y(new_n4558_));
  AOI21X1  g02123(.A0(new_n4558_), .A1(new_n2437_), .B0(new_n4552_), .Y(new_n4559_));
  OAI21X1  g02124(.A0(new_n4559_), .A1(pi0215), .B0(new_n4473_), .Y(new_n4560_));
  AOI21X1  g02125(.A0(new_n4462_), .A1(pi0228), .B0(new_n3280_), .Y(new_n4561_));
  AOI21X1  g02126(.A0(new_n4561_), .A1(new_n4498_), .B0(pi0216), .Y(new_n4562_));
  OAI21X1  g02127(.A0(new_n4562_), .A1(new_n4458_), .B0(new_n2437_), .Y(new_n4563_));
  AOI21X1  g02128(.A0(new_n4563_), .A1(new_n4457_), .B0(pi0215), .Y(new_n4564_));
  OR2X1    g02129(.A(new_n4564_), .B(new_n4472_), .Y(new_n4565_));
  AOI21X1  g02130(.A0(new_n4565_), .A1(pi0299), .B0(new_n4493_), .Y(new_n4566_));
  OAI21X1  g02131(.A0(new_n4566_), .A1(new_n2959_), .B0(new_n2996_), .Y(new_n4567_));
  AOI21X1  g02132(.A0(new_n4560_), .A1(new_n4487_), .B0(new_n4567_), .Y(new_n4568_));
  NOR2X1   g02133(.A(new_n4543_), .B(new_n3281_), .Y(new_n4569_));
  INVX1    g02134(.A(new_n4569_), .Y(new_n4570_));
  AOI21X1  g02135(.A0(new_n4570_), .A1(pi0299), .B0(new_n4493_), .Y(new_n4571_));
  INVX1    g02136(.A(new_n4571_), .Y(new_n4572_));
  OAI21X1  g02137(.A0(new_n4572_), .A1(new_n2996_), .B0(new_n3026_), .Y(new_n4573_));
  INVX1    g02138(.A(new_n4472_), .Y(new_n4574_));
  INVX1    g02139(.A(new_n4561_), .Y(new_n4575_));
  OAI21X1  g02140(.A0(new_n4575_), .A1(new_n4518_), .B0(new_n2438_), .Y(new_n4576_));
  AOI21X1  g02141(.A0(new_n4576_), .A1(new_n4553_), .B0(pi0221), .Y(new_n4577_));
  OAI21X1  g02142(.A0(new_n4577_), .A1(new_n4552_), .B0(new_n2954_), .Y(new_n4578_));
  AOI21X1  g02143(.A0(new_n4578_), .A1(new_n4574_), .B0(new_n2953_), .Y(new_n4579_));
  NOR3X1   g02144(.A(new_n4579_), .B(new_n4493_), .C(new_n3066_), .Y(new_n4580_));
  OAI21X1  g02145(.A0(new_n4572_), .A1(new_n3065_), .B0(pi0100), .Y(new_n4581_));
  OAI22X1  g02146(.A0(new_n4581_), .A1(new_n4580_), .B0(new_n4573_), .B1(new_n4568_), .Y(new_n4582_));
  MX2X1    g02147(.A(new_n4571_), .B(new_n4566_), .S0(new_n3085_), .Y(new_n4583_));
  OAI21X1  g02148(.A0(new_n4583_), .A1(new_n3156_), .B0(new_n3095_), .Y(new_n4584_));
  AOI21X1  g02149(.A0(new_n4582_), .A1(new_n3156_), .B0(new_n4584_), .Y(new_n4585_));
  OAI21X1  g02150(.A0(new_n4572_), .A1(new_n3095_), .B0(new_n3100_), .Y(new_n4586_));
  NAND2X1  g02151(.A(new_n4583_), .B(new_n3098_), .Y(new_n4587_));
  AOI21X1  g02152(.A0(new_n4571_), .A1(new_n3101_), .B0(new_n3100_), .Y(new_n4588_));
  AOI21X1  g02153(.A0(new_n4588_), .A1(new_n4587_), .B0(new_n3136_), .Y(new_n4589_));
  OAI21X1  g02154(.A0(new_n4586_), .A1(new_n4585_), .B0(new_n4589_), .Y(new_n4590_));
  AOI21X1  g02155(.A0(new_n4571_), .A1(new_n3136_), .B0(pi0055), .Y(new_n4591_));
  NOR3X1   g02156(.A(new_n4564_), .B(new_n4472_), .C(new_n3131_), .Y(new_n4592_));
  OAI21X1  g02157(.A0(new_n4570_), .A1(new_n3130_), .B0(pi0055), .Y(new_n4593_));
  OAI21X1  g02158(.A0(new_n4593_), .A1(new_n4592_), .B0(new_n3143_), .Y(new_n4594_));
  AOI21X1  g02159(.A0(new_n4591_), .A1(new_n4590_), .B0(new_n4594_), .Y(new_n4595_));
  OAI21X1  g02160(.A0(new_n4569_), .A1(new_n3140_), .B0(pi0056), .Y(new_n4596_));
  AOI21X1  g02161(.A0(new_n4565_), .A1(new_n3140_), .B0(new_n4596_), .Y(new_n4597_));
  NOR3X1   g02162(.A(new_n4597_), .B(new_n4595_), .C(pi0062), .Y(new_n4598_));
  NOR3X1   g02163(.A(new_n4564_), .B(new_n4472_), .C(new_n3249_), .Y(new_n4599_));
  OAI21X1  g02164(.A0(new_n4570_), .A1(new_n3248_), .B0(pi0062), .Y(new_n4600_));
  OAI21X1  g02165(.A0(new_n4600_), .A1(new_n4599_), .B0(new_n3246_), .Y(new_n4601_));
  AOI21X1  g02166(.A0(new_n4569_), .A1(new_n3393_), .B0(new_n4550_), .Y(new_n4602_));
  OAI21X1  g02167(.A0(new_n4601_), .A1(new_n4598_), .B0(new_n4602_), .Y(new_n4603_));
  OAI21X1  g02168(.A0(new_n4551_), .A1(new_n4549_), .B0(new_n4603_), .Y(po0163));
  INVX1    g02169(.A(pi0938), .Y(new_n4605_));
  AOI21X1  g02170(.A0(new_n2442_), .A1(new_n4605_), .B0(new_n2437_), .Y(new_n4606_));
  OAI21X1  g02171(.A0(new_n2442_), .A1(pi1135), .B0(new_n4606_), .Y(new_n4607_));
  AND2X1   g02172(.A(pi0279), .B(pi0216), .Y(new_n4608_));
  INVX1    g02173(.A(pi0879), .Y(new_n4609_));
  AOI21X1  g02174(.A0(new_n2454_), .A1(pi0095), .B0(new_n4609_), .Y(new_n4610_));
  MX2X1    g02175(.A(new_n4610_), .B(pi0161), .S0(new_n2448_), .Y(new_n4611_));
  OAI21X1  g02176(.A0(new_n4611_), .A1(new_n4459_), .B0(new_n2438_), .Y(new_n4612_));
  INVX1    g02177(.A(pi0161), .Y(new_n4613_));
  OAI21X1  g02178(.A0(new_n3532_), .A1(new_n4613_), .B0(pi0879), .Y(new_n4614_));
  AOI21X1  g02179(.A0(new_n3531_), .A1(new_n4613_), .B0(new_n4614_), .Y(new_n4615_));
  NOR3X1   g02180(.A(new_n3535_), .B(pi0879), .C(new_n4613_), .Y(new_n4616_));
  OAI21X1  g02181(.A0(new_n4616_), .A1(new_n4615_), .B0(new_n3013_), .Y(new_n4617_));
  AOI21X1  g02182(.A0(new_n4617_), .A1(new_n4459_), .B0(new_n4612_), .Y(new_n4618_));
  OAI21X1  g02183(.A0(new_n4618_), .A1(new_n4608_), .B0(new_n2437_), .Y(new_n4619_));
  AOI21X1  g02184(.A0(new_n4619_), .A1(new_n4607_), .B0(pi0215), .Y(new_n4620_));
  AND2X1   g02185(.A(pi1135), .B(pi0215), .Y(new_n4621_));
  NOR2X1   g02186(.A(new_n4621_), .B(new_n2953_), .Y(new_n4622_));
  INVX1    g02187(.A(new_n4622_), .Y(new_n4623_));
  AOI21X1  g02188(.A0(pi1135), .A1(pi0223), .B0(pi0299), .Y(new_n4624_));
  AOI21X1  g02189(.A0(new_n3159_), .A1(new_n4605_), .B0(new_n2960_), .Y(new_n4625_));
  OAI21X1  g02190(.A0(new_n3159_), .A1(pi1135), .B0(new_n4625_), .Y(new_n4626_));
  NOR3X1   g02191(.A(new_n2455_), .B(pi0879), .C(pi0224), .Y(new_n4627_));
  OAI21X1  g02192(.A0(pi0279), .A1(new_n2961_), .B0(new_n2960_), .Y(new_n4628_));
  OAI21X1  g02193(.A0(new_n4628_), .A1(new_n4627_), .B0(new_n4626_), .Y(new_n4629_));
  INVX1    g02194(.A(new_n4626_), .Y(new_n4630_));
  OR4X1    g02195(.A(new_n4630_), .B(new_n3258_), .C(pi0224), .D(pi0222), .Y(new_n4631_));
  NAND3X1  g02196(.A(new_n4631_), .B(new_n4629_), .C(new_n2964_), .Y(new_n4632_));
  AOI21X1  g02197(.A0(new_n4632_), .A1(new_n4624_), .B0(pi0039), .Y(new_n4633_));
  OAI21X1  g02198(.A0(new_n4623_), .A1(new_n4620_), .B0(new_n4633_), .Y(new_n4634_));
  AND2X1   g02199(.A(pi1135), .B(pi0223), .Y(new_n4635_));
  AOI21X1  g02200(.A0(new_n4629_), .A1(new_n2964_), .B0(new_n4635_), .Y(new_n4636_));
  OR2X1    g02201(.A(new_n4636_), .B(pi0299), .Y(new_n4637_));
  INVX1    g02202(.A(new_n4637_), .Y(new_n4638_));
  OAI21X1  g02203(.A0(new_n4610_), .A1(new_n3009_), .B0(new_n4638_), .Y(new_n4639_));
  AND2X1   g02204(.A(new_n4611_), .B(pi0228), .Y(new_n4640_));
  INVX1    g02205(.A(new_n4640_), .Y(new_n4641_));
  AND2X1   g02206(.A(new_n3013_), .B(pi0161), .Y(new_n4642_));
  OAI22X1  g02207(.A0(new_n4642_), .A1(new_n3631_), .B0(new_n3074_), .B1(pi0879), .Y(new_n4643_));
  AOI21X1  g02208(.A0(new_n4643_), .A1(new_n4641_), .B0(pi0216), .Y(new_n4644_));
  OAI21X1  g02209(.A0(new_n4644_), .A1(new_n4608_), .B0(new_n2437_), .Y(new_n4645_));
  AOI21X1  g02210(.A0(new_n4645_), .A1(new_n4607_), .B0(pi0215), .Y(new_n4646_));
  OAI21X1  g02211(.A0(new_n4646_), .A1(new_n4621_), .B0(pi0299), .Y(new_n4647_));
  AND2X1   g02212(.A(new_n4647_), .B(new_n4639_), .Y(new_n4648_));
  INVX1    g02213(.A(new_n4648_), .Y(new_n4649_));
  AOI21X1  g02214(.A0(new_n4649_), .A1(pi0039), .B0(pi0038), .Y(new_n4650_));
  INVX1    g02215(.A(new_n4639_), .Y(new_n4651_));
  INVX1    g02216(.A(pi0279), .Y(new_n4652_));
  AOI21X1  g02217(.A0(new_n4611_), .A1(pi0228), .B0(new_n4642_), .Y(new_n4653_));
  MX2X1    g02218(.A(new_n4653_), .B(new_n4652_), .S0(pi0216), .Y(new_n4654_));
  OAI21X1  g02219(.A0(new_n4654_), .A1(pi0221), .B0(new_n4607_), .Y(new_n4655_));
  AOI21X1  g02220(.A0(new_n4655_), .A1(new_n2954_), .B0(new_n4621_), .Y(new_n4656_));
  INVX1    g02221(.A(new_n4656_), .Y(new_n4657_));
  AOI21X1  g02222(.A0(new_n4657_), .A1(pi0299), .B0(new_n4651_), .Y(new_n4658_));
  INVX1    g02223(.A(new_n4658_), .Y(new_n4659_));
  OAI21X1  g02224(.A0(new_n4659_), .A1(new_n2996_), .B0(new_n3026_), .Y(new_n4660_));
  AOI21X1  g02225(.A0(new_n4650_), .A1(new_n4634_), .B0(new_n4660_), .Y(new_n4661_));
  AOI21X1  g02226(.A0(new_n3213_), .A1(new_n4609_), .B0(new_n4613_), .Y(new_n4662_));
  INVX1    g02227(.A(new_n4662_), .Y(new_n4663_));
  NOR2X1   g02228(.A(pi0166), .B(pi0152), .Y(new_n4664_));
  AOI21X1  g02229(.A0(new_n4664_), .A1(new_n3497_), .B0(new_n4609_), .Y(new_n4665_));
  OAI21X1  g02230(.A0(new_n4664_), .A1(new_n3213_), .B0(new_n4665_), .Y(new_n4666_));
  AOI21X1  g02231(.A0(new_n4666_), .A1(new_n4663_), .B0(pi0228), .Y(new_n4667_));
  OR2X1    g02232(.A(new_n4667_), .B(new_n4640_), .Y(new_n4668_));
  AOI21X1  g02233(.A0(new_n4668_), .A1(new_n2438_), .B0(new_n4608_), .Y(new_n4669_));
  OAI21X1  g02234(.A0(new_n4669_), .A1(pi0221), .B0(new_n4607_), .Y(new_n4670_));
  AOI21X1  g02235(.A0(new_n4670_), .A1(new_n2954_), .B0(new_n4621_), .Y(new_n4671_));
  AND2X1   g02236(.A(new_n4639_), .B(new_n3065_), .Y(new_n4672_));
  OAI21X1  g02237(.A0(new_n4671_), .A1(new_n2953_), .B0(new_n4672_), .Y(new_n4673_));
  AOI21X1  g02238(.A0(new_n4658_), .A1(new_n3066_), .B0(new_n3026_), .Y(new_n4674_));
  AND2X1   g02239(.A(new_n4674_), .B(new_n4673_), .Y(new_n4675_));
  OAI21X1  g02240(.A0(new_n4675_), .A1(new_n4661_), .B0(new_n3156_), .Y(new_n4676_));
  MX2X1    g02241(.A(new_n4659_), .B(new_n4649_), .S0(new_n3085_), .Y(new_n4677_));
  AOI21X1  g02242(.A0(new_n4677_), .A1(pi0087), .B0(pi0075), .Y(new_n4678_));
  OAI21X1  g02243(.A0(new_n4659_), .A1(new_n3095_), .B0(new_n3100_), .Y(new_n4679_));
  AOI21X1  g02244(.A0(new_n4678_), .A1(new_n4676_), .B0(new_n4679_), .Y(new_n4680_));
  OR2X1    g02245(.A(new_n4677_), .B(new_n3101_), .Y(new_n4681_));
  AOI21X1  g02246(.A0(new_n4658_), .A1(new_n3101_), .B0(new_n3100_), .Y(new_n4682_));
  AND2X1   g02247(.A(new_n4682_), .B(new_n4681_), .Y(new_n4683_));
  NOR3X1   g02248(.A(new_n4683_), .B(new_n4680_), .C(new_n3136_), .Y(new_n4684_));
  OAI21X1  g02249(.A0(new_n4659_), .A1(new_n3135_), .B0(new_n3128_), .Y(new_n4685_));
  OR4X1    g02250(.A(new_n4646_), .B(new_n4621_), .C(new_n3810_), .D(new_n3066_), .Y(new_n4686_));
  AOI21X1  g02251(.A0(new_n4656_), .A1(new_n3131_), .B0(new_n3128_), .Y(new_n4687_));
  AOI21X1  g02252(.A0(new_n4687_), .A1(new_n4686_), .B0(pi0056), .Y(new_n4688_));
  OAI21X1  g02253(.A0(new_n4685_), .A1(new_n4684_), .B0(new_n4688_), .Y(new_n4689_));
  OAI21X1  g02254(.A0(new_n4646_), .A1(new_n4621_), .B0(new_n3140_), .Y(new_n4690_));
  AOI21X1  g02255(.A0(new_n4657_), .A1(new_n3242_), .B0(new_n3143_), .Y(new_n4691_));
  AOI21X1  g02256(.A0(new_n4691_), .A1(new_n4690_), .B0(pi0062), .Y(new_n4692_));
  NOR3X1   g02257(.A(new_n4646_), .B(new_n4621_), .C(new_n3249_), .Y(new_n4693_));
  OAI21X1  g02258(.A0(new_n4657_), .A1(new_n3248_), .B0(pi0062), .Y(new_n4694_));
  OAI21X1  g02259(.A0(new_n4694_), .A1(new_n4693_), .B0(new_n3246_), .Y(new_n4695_));
  AOI21X1  g02260(.A0(new_n4692_), .A1(new_n4689_), .B0(new_n4695_), .Y(new_n4696_));
  INVX1    g02261(.A(pi0244), .Y(new_n4697_));
  OAI21X1  g02262(.A0(new_n4657_), .A1(new_n3246_), .B0(new_n4697_), .Y(new_n4698_));
  INVX1    g02263(.A(new_n4607_), .Y(new_n4699_));
  INVX1    g02264(.A(new_n4608_), .Y(new_n4700_));
  OAI21X1  g02265(.A0(new_n3271_), .A1(pi0161), .B0(new_n4609_), .Y(new_n4701_));
  AOI21X1  g02266(.A0(new_n3266_), .A1(pi0161), .B0(new_n4701_), .Y(new_n4702_));
  AOI21X1  g02267(.A0(new_n3204_), .A1(new_n4613_), .B0(new_n4609_), .Y(new_n4703_));
  NOR3X1   g02268(.A(new_n4703_), .B(new_n4702_), .C(pi0228), .Y(new_n4704_));
  OAI21X1  g02269(.A0(new_n4704_), .A1(new_n4612_), .B0(new_n4700_), .Y(new_n4705_));
  AOI21X1  g02270(.A0(new_n4705_), .A1(new_n2437_), .B0(new_n4699_), .Y(new_n4706_));
  OAI21X1  g02271(.A0(new_n4706_), .A1(pi0215), .B0(new_n4622_), .Y(new_n4707_));
  OAI21X1  g02272(.A0(new_n4629_), .A1(new_n4478_), .B0(new_n2964_), .Y(new_n4708_));
  AOI21X1  g02273(.A0(new_n4708_), .A1(new_n4624_), .B0(pi0039), .Y(new_n4709_));
  AOI21X1  g02274(.A0(new_n4611_), .A1(pi0228), .B0(new_n3280_), .Y(new_n4710_));
  AOI21X1  g02275(.A0(new_n4710_), .A1(new_n4643_), .B0(pi0216), .Y(new_n4711_));
  OAI21X1  g02276(.A0(new_n4711_), .A1(new_n4608_), .B0(new_n2437_), .Y(new_n4712_));
  AOI21X1  g02277(.A0(new_n4712_), .A1(new_n4607_), .B0(pi0215), .Y(new_n4713_));
  NOR2X1   g02278(.A(new_n4713_), .B(new_n4621_), .Y(new_n4714_));
  MX2X1    g02279(.A(new_n4714_), .B(new_n4636_), .S0(new_n2953_), .Y(new_n4715_));
  OAI21X1  g02280(.A0(new_n4715_), .A1(new_n2959_), .B0(new_n2996_), .Y(new_n4716_));
  AOI21X1  g02281(.A0(new_n4709_), .A1(new_n4707_), .B0(new_n4716_), .Y(new_n4717_));
  NOR2X1   g02282(.A(new_n4657_), .B(new_n3281_), .Y(new_n4718_));
  MX2X1    g02283(.A(new_n4718_), .B(new_n4636_), .S0(new_n2953_), .Y(new_n4719_));
  INVX1    g02284(.A(new_n4719_), .Y(new_n4720_));
  OAI21X1  g02285(.A0(new_n4720_), .A1(new_n2996_), .B0(new_n3026_), .Y(new_n4721_));
  INVX1    g02286(.A(new_n4621_), .Y(new_n4722_));
  INVX1    g02287(.A(new_n4710_), .Y(new_n4723_));
  OAI21X1  g02288(.A0(new_n4723_), .A1(new_n4667_), .B0(new_n2438_), .Y(new_n4724_));
  AOI21X1  g02289(.A0(new_n4724_), .A1(new_n4700_), .B0(pi0221), .Y(new_n4725_));
  OAI21X1  g02290(.A0(new_n4725_), .A1(new_n4699_), .B0(new_n2954_), .Y(new_n4726_));
  AOI21X1  g02291(.A0(new_n4726_), .A1(new_n4722_), .B0(new_n2953_), .Y(new_n4727_));
  NOR3X1   g02292(.A(new_n4727_), .B(new_n4638_), .C(new_n3066_), .Y(new_n4728_));
  OAI21X1  g02293(.A0(new_n4720_), .A1(new_n3065_), .B0(pi0100), .Y(new_n4729_));
  OAI22X1  g02294(.A0(new_n4729_), .A1(new_n4728_), .B0(new_n4721_), .B1(new_n4717_), .Y(new_n4730_));
  MX2X1    g02295(.A(new_n4719_), .B(new_n4715_), .S0(new_n3085_), .Y(new_n4731_));
  OAI21X1  g02296(.A0(new_n4731_), .A1(new_n3156_), .B0(new_n3095_), .Y(new_n4732_));
  AOI21X1  g02297(.A0(new_n4730_), .A1(new_n3156_), .B0(new_n4732_), .Y(new_n4733_));
  OAI21X1  g02298(.A0(new_n4720_), .A1(new_n3095_), .B0(new_n3100_), .Y(new_n4734_));
  NAND2X1  g02299(.A(new_n4731_), .B(new_n3098_), .Y(new_n4735_));
  AOI21X1  g02300(.A0(new_n4719_), .A1(new_n3101_), .B0(new_n3100_), .Y(new_n4736_));
  AOI21X1  g02301(.A0(new_n4736_), .A1(new_n4735_), .B0(new_n3136_), .Y(new_n4737_));
  OAI21X1  g02302(.A0(new_n4734_), .A1(new_n4733_), .B0(new_n4737_), .Y(new_n4738_));
  AOI21X1  g02303(.A0(new_n4719_), .A1(new_n3136_), .B0(pi0055), .Y(new_n4739_));
  NOR3X1   g02304(.A(new_n4713_), .B(new_n4621_), .C(new_n3131_), .Y(new_n4740_));
  INVX1    g02305(.A(new_n4718_), .Y(new_n4741_));
  OAI21X1  g02306(.A0(new_n4741_), .A1(new_n3130_), .B0(pi0055), .Y(new_n4742_));
  OAI21X1  g02307(.A0(new_n4742_), .A1(new_n4740_), .B0(new_n3143_), .Y(new_n4743_));
  AOI21X1  g02308(.A0(new_n4739_), .A1(new_n4738_), .B0(new_n4743_), .Y(new_n4744_));
  OAI21X1  g02309(.A0(new_n4713_), .A1(new_n4621_), .B0(new_n3140_), .Y(new_n4745_));
  AOI21X1  g02310(.A0(new_n4741_), .A1(new_n3242_), .B0(new_n3143_), .Y(new_n4746_));
  AND2X1   g02311(.A(new_n4746_), .B(new_n4745_), .Y(new_n4747_));
  NOR3X1   g02312(.A(new_n4747_), .B(new_n4744_), .C(pi0062), .Y(new_n4748_));
  NOR3X1   g02313(.A(new_n4713_), .B(new_n4621_), .C(new_n3249_), .Y(new_n4749_));
  OAI21X1  g02314(.A0(new_n4741_), .A1(new_n3248_), .B0(pi0062), .Y(new_n4750_));
  OAI21X1  g02315(.A0(new_n4750_), .A1(new_n4749_), .B0(new_n3246_), .Y(new_n4751_));
  AOI21X1  g02316(.A0(new_n4718_), .A1(new_n3393_), .B0(new_n4697_), .Y(new_n4752_));
  OAI21X1  g02317(.A0(new_n4751_), .A1(new_n4748_), .B0(new_n4752_), .Y(new_n4753_));
  OAI21X1  g02318(.A0(new_n4698_), .A1(new_n4696_), .B0(new_n4753_), .Y(po0164));
  INVX1    g02319(.A(pi1134), .Y(new_n4755_));
  NOR4X1   g02320(.A(pi0930), .B(new_n2721_), .C(new_n2437_), .D(pi0216), .Y(new_n4756_));
  AOI21X1  g02321(.A0(pi0278), .A1(pi0216), .B0(pi0221), .Y(new_n4757_));
  INVX1    g02322(.A(new_n4757_), .Y(new_n4758_));
  AOI21X1  g02323(.A0(pi0152), .A1(new_n2448_), .B0(new_n3013_), .Y(new_n4759_));
  INVX1    g02324(.A(new_n4759_), .Y(new_n4760_));
  INVX1    g02325(.A(pi0846), .Y(new_n4761_));
  AOI21X1  g02326(.A0(new_n3258_), .A1(new_n4761_), .B0(new_n2448_), .Y(new_n4762_));
  OAI21X1  g02327(.A0(new_n4762_), .A1(new_n4760_), .B0(new_n2438_), .Y(new_n4763_));
  INVX1    g02328(.A(new_n4763_), .Y(new_n4764_));
  OAI21X1  g02329(.A0(new_n3532_), .A1(pi0152), .B0(new_n4761_), .Y(new_n4765_));
  AOI21X1  g02330(.A0(new_n3531_), .A1(pi0152), .B0(new_n4765_), .Y(new_n4766_));
  NOR3X1   g02331(.A(new_n3535_), .B(new_n4761_), .C(pi0152), .Y(new_n4767_));
  OAI21X1  g02332(.A0(new_n4767_), .A1(new_n4766_), .B0(new_n3013_), .Y(new_n4768_));
  AOI21X1  g02333(.A0(new_n4768_), .A1(new_n4764_), .B0(new_n4758_), .Y(new_n4769_));
  AOI21X1  g02334(.A0(pi0833), .A1(new_n2438_), .B0(new_n2437_), .Y(new_n4770_));
  NOR3X1   g02335(.A(new_n4770_), .B(new_n2953_), .C(pi0215), .Y(new_n4771_));
  INVX1    g02336(.A(new_n4771_), .Y(new_n4772_));
  NOR3X1   g02337(.A(new_n4772_), .B(new_n4769_), .C(new_n4756_), .Y(new_n4773_));
  NOR4X1   g02338(.A(pi0930), .B(new_n2721_), .C(pi0224), .D(new_n2960_), .Y(new_n4774_));
  INVX1    g02339(.A(new_n4774_), .Y(new_n4775_));
  AOI21X1  g02340(.A0(pi0278), .A1(pi0224), .B0(pi0222), .Y(new_n4776_));
  INVX1    g02341(.A(new_n4776_), .Y(new_n4777_));
  AOI21X1  g02342(.A0(new_n3258_), .A1(new_n4761_), .B0(pi0224), .Y(new_n4778_));
  OAI21X1  g02343(.A0(new_n4778_), .A1(new_n4777_), .B0(new_n4775_), .Y(new_n4779_));
  NOR2X1   g02344(.A(pi0299), .B(pi0223), .Y(new_n4780_));
  INVX1    g02345(.A(new_n4780_), .Y(new_n4781_));
  NOR2X1   g02346(.A(new_n4781_), .B(new_n2962_), .Y(new_n4782_));
  INVX1    g02347(.A(new_n4782_), .Y(new_n4783_));
  OAI21X1  g02348(.A0(new_n4783_), .A1(new_n4779_), .B0(new_n2959_), .Y(new_n4784_));
  AOI21X1  g02349(.A0(new_n2454_), .A1(pi0095), .B0(new_n4761_), .Y(new_n4785_));
  AOI21X1  g02350(.A0(new_n4785_), .A1(new_n2961_), .B0(new_n4777_), .Y(new_n4786_));
  NOR4X1   g02351(.A(new_n4786_), .B(new_n4774_), .C(new_n2962_), .D(pi0223), .Y(new_n4787_));
  NOR2X1   g02352(.A(new_n4787_), .B(pi0299), .Y(new_n4788_));
  INVX1    g02353(.A(new_n4788_), .Y(new_n4789_));
  AOI21X1  g02354(.A0(new_n3008_), .A1(new_n2455_), .B0(new_n4789_), .Y(new_n4790_));
  INVX1    g02355(.A(new_n4790_), .Y(new_n4791_));
  NOR3X1   g02356(.A(new_n4770_), .B(new_n4756_), .C(pi0215), .Y(new_n4792_));
  INVX1    g02357(.A(new_n4792_), .Y(new_n4793_));
  MX2X1    g02358(.A(new_n4785_), .B(pi0152), .S0(new_n2448_), .Y(new_n4794_));
  AOI21X1  g02359(.A0(new_n4794_), .A1(pi0228), .B0(new_n3280_), .Y(new_n4795_));
  AOI21X1  g02360(.A0(new_n3630_), .A1(new_n4761_), .B0(pi0228), .Y(new_n4796_));
  OAI21X1  g02361(.A0(new_n3630_), .A1(pi0152), .B0(new_n4796_), .Y(new_n4797_));
  AOI21X1  g02362(.A0(new_n4797_), .A1(new_n4795_), .B0(pi0216), .Y(new_n4798_));
  NOR2X1   g02363(.A(new_n4798_), .B(new_n4758_), .Y(new_n4799_));
  NOR2X1   g02364(.A(new_n4799_), .B(new_n4793_), .Y(new_n4800_));
  OAI21X1  g02365(.A0(new_n4800_), .A1(new_n2953_), .B0(new_n4791_), .Y(new_n4801_));
  AOI21X1  g02366(.A0(new_n4801_), .A1(pi0039), .B0(pi0038), .Y(new_n4802_));
  OAI21X1  g02367(.A0(new_n4784_), .A1(new_n4773_), .B0(new_n4802_), .Y(new_n4803_));
  AND2X1   g02368(.A(new_n4794_), .B(pi0228), .Y(new_n4804_));
  AOI21X1  g02369(.A0(new_n3013_), .A1(pi0152), .B0(new_n4804_), .Y(new_n4805_));
  OAI21X1  g02370(.A0(new_n4805_), .A1(pi0216), .B0(new_n4757_), .Y(new_n4806_));
  AOI21X1  g02371(.A0(new_n4806_), .A1(new_n4792_), .B0(new_n3281_), .Y(new_n4807_));
  AOI21X1  g02372(.A0(new_n4807_), .A1(pi0299), .B0(new_n4790_), .Y(new_n4808_));
  AOI21X1  g02373(.A0(new_n4808_), .A1(pi0038), .B0(pi0100), .Y(new_n4809_));
  AOI22X1  g02374(.A0(new_n3218_), .A1(pi0846), .B0(new_n3214_), .B1(pi0152), .Y(new_n4810_));
  OAI21X1  g02375(.A0(new_n4810_), .A1(pi0228), .B0(new_n4795_), .Y(new_n4811_));
  AOI21X1  g02376(.A0(new_n4811_), .A1(new_n2438_), .B0(new_n4758_), .Y(new_n4812_));
  OAI21X1  g02377(.A0(new_n4812_), .A1(new_n4793_), .B0(pi0299), .Y(new_n4813_));
  NAND3X1  g02378(.A(new_n4813_), .B(new_n4791_), .C(new_n3065_), .Y(new_n4814_));
  AOI21X1  g02379(.A0(new_n4808_), .A1(new_n3066_), .B0(new_n3026_), .Y(new_n4815_));
  AOI22X1  g02380(.A0(new_n4815_), .A1(new_n4814_), .B0(new_n4809_), .B1(new_n4803_), .Y(new_n4816_));
  INVX1    g02381(.A(new_n4808_), .Y(new_n4817_));
  MX2X1    g02382(.A(new_n4817_), .B(new_n4801_), .S0(new_n3085_), .Y(new_n4818_));
  AOI21X1  g02383(.A0(new_n4818_), .A1(pi0087), .B0(pi0075), .Y(new_n4819_));
  OAI21X1  g02384(.A0(new_n4816_), .A1(pi0087), .B0(new_n4819_), .Y(new_n4820_));
  AOI21X1  g02385(.A0(new_n4808_), .A1(pi0075), .B0(pi0092), .Y(new_n4821_));
  NOR2X1   g02386(.A(new_n4818_), .B(new_n3101_), .Y(new_n4822_));
  OAI21X1  g02387(.A0(new_n4817_), .A1(new_n3098_), .B0(pi0092), .Y(new_n4823_));
  OAI21X1  g02388(.A0(new_n4823_), .A1(new_n4822_), .B0(new_n3135_), .Y(new_n4824_));
  AOI21X1  g02389(.A0(new_n4821_), .A1(new_n4820_), .B0(new_n4824_), .Y(new_n4825_));
  OAI21X1  g02390(.A0(new_n4817_), .A1(new_n3135_), .B0(new_n3128_), .Y(new_n4826_));
  NOR2X1   g02391(.A(new_n4770_), .B(pi0215), .Y(new_n4827_));
  INVX1    g02392(.A(new_n4827_), .Y(new_n4828_));
  OR4X1    g02393(.A(new_n4799_), .B(new_n4828_), .C(new_n4756_), .D(new_n3131_), .Y(new_n4829_));
  OR2X1    g02394(.A(new_n4807_), .B(new_n3130_), .Y(new_n4830_));
  AND2X1   g02395(.A(new_n4830_), .B(pi0055), .Y(new_n4831_));
  AOI21X1  g02396(.A0(new_n4831_), .A1(new_n4829_), .B0(pi0056), .Y(new_n4832_));
  OAI21X1  g02397(.A0(new_n4826_), .A1(new_n4825_), .B0(new_n4832_), .Y(new_n4833_));
  OAI21X1  g02398(.A0(new_n4799_), .A1(new_n4793_), .B0(new_n3140_), .Y(new_n4834_));
  AOI21X1  g02399(.A0(new_n4807_), .A1(new_n3242_), .B0(new_n3143_), .Y(new_n4835_));
  AOI21X1  g02400(.A0(new_n4835_), .A1(new_n4834_), .B0(pi0062), .Y(new_n4836_));
  NOR3X1   g02401(.A(new_n4799_), .B(new_n4793_), .C(new_n3249_), .Y(new_n4837_));
  OAI21X1  g02402(.A0(new_n4807_), .A1(new_n3248_), .B0(pi0062), .Y(new_n4838_));
  OAI21X1  g02403(.A0(new_n4838_), .A1(new_n4837_), .B0(new_n3246_), .Y(new_n4839_));
  AOI21X1  g02404(.A0(new_n4836_), .A1(new_n4833_), .B0(new_n4839_), .Y(new_n4840_));
  OAI21X1  g02405(.A0(new_n4807_), .A1(new_n3246_), .B0(pi0242), .Y(new_n4841_));
  INVX1    g02406(.A(new_n4756_), .Y(new_n4842_));
  AOI21X1  g02407(.A0(new_n3271_), .A1(pi0152), .B0(new_n4761_), .Y(new_n4843_));
  OAI21X1  g02408(.A0(new_n3266_), .A1(pi0152), .B0(new_n4843_), .Y(new_n4844_));
  AND2X1   g02409(.A(new_n4761_), .B(pi0152), .Y(new_n4845_));
  AOI21X1  g02410(.A0(new_n4845_), .A1(new_n3204_), .B0(pi0228), .Y(new_n4846_));
  AOI21X1  g02411(.A0(new_n4759_), .A1(new_n3259_), .B0(new_n4763_), .Y(new_n4847_));
  INVX1    g02412(.A(new_n4847_), .Y(new_n4848_));
  AOI21X1  g02413(.A0(new_n4846_), .A1(new_n4844_), .B0(new_n4848_), .Y(new_n4849_));
  OAI21X1  g02414(.A0(new_n4849_), .A1(new_n4758_), .B0(new_n4842_), .Y(new_n4850_));
  OR4X1    g02415(.A(new_n3257_), .B(new_n2455_), .C(new_n4761_), .D(pi0224), .Y(new_n4851_));
  AND2X1   g02416(.A(new_n4851_), .B(new_n4776_), .Y(new_n4852_));
  OR4X1    g02417(.A(new_n4852_), .B(new_n4774_), .C(new_n4781_), .D(new_n2962_), .Y(new_n4853_));
  AND2X1   g02418(.A(new_n4853_), .B(new_n2959_), .Y(new_n4854_));
  OAI21X1  g02419(.A0(new_n4850_), .A1(new_n4772_), .B0(new_n4854_), .Y(new_n4855_));
  INVX1    g02420(.A(new_n4804_), .Y(new_n4856_));
  AOI21X1  g02421(.A0(new_n4797_), .A1(new_n4856_), .B0(pi0216), .Y(new_n4857_));
  NOR2X1   g02422(.A(new_n4857_), .B(new_n4758_), .Y(new_n4858_));
  OAI21X1  g02423(.A0(new_n4858_), .A1(new_n4793_), .B0(pi0299), .Y(new_n4859_));
  NAND2X1  g02424(.A(new_n4859_), .B(new_n4789_), .Y(new_n4860_));
  AOI21X1  g02425(.A0(new_n4860_), .A1(pi0039), .B0(pi0038), .Y(new_n4861_));
  AND2X1   g02426(.A(new_n4806_), .B(new_n4792_), .Y(new_n4862_));
  MX2X1    g02427(.A(new_n4862_), .B(new_n4787_), .S0(new_n2953_), .Y(new_n4863_));
  INVX1    g02428(.A(new_n4863_), .Y(new_n4864_));
  OAI21X1  g02429(.A0(new_n4864_), .A1(new_n2996_), .B0(new_n3026_), .Y(new_n4865_));
  AOI21X1  g02430(.A0(new_n4861_), .A1(new_n4855_), .B0(new_n4865_), .Y(new_n4866_));
  OAI21X1  g02431(.A0(new_n4810_), .A1(pi0228), .B0(new_n4856_), .Y(new_n4867_));
  AOI21X1  g02432(.A0(new_n4867_), .A1(new_n2438_), .B0(new_n4758_), .Y(new_n4868_));
  OAI21X1  g02433(.A0(new_n4868_), .A1(new_n4793_), .B0(pi0299), .Y(new_n4869_));
  NAND3X1  g02434(.A(new_n4869_), .B(new_n4789_), .C(new_n3065_), .Y(new_n4870_));
  AOI21X1  g02435(.A0(new_n4863_), .A1(new_n3066_), .B0(new_n3026_), .Y(new_n4871_));
  AOI21X1  g02436(.A0(new_n4871_), .A1(new_n4870_), .B0(new_n4866_), .Y(new_n4872_));
  MX2X1    g02437(.A(new_n4864_), .B(new_n4860_), .S0(new_n3085_), .Y(new_n4873_));
  AOI21X1  g02438(.A0(new_n4873_), .A1(pi0087), .B0(pi0075), .Y(new_n4874_));
  OAI21X1  g02439(.A0(new_n4872_), .A1(pi0087), .B0(new_n4874_), .Y(new_n4875_));
  AOI21X1  g02440(.A0(new_n4863_), .A1(pi0075), .B0(pi0092), .Y(new_n4876_));
  NOR2X1   g02441(.A(new_n4873_), .B(new_n3101_), .Y(new_n4877_));
  OAI21X1  g02442(.A0(new_n4864_), .A1(new_n3098_), .B0(pi0092), .Y(new_n4878_));
  OAI21X1  g02443(.A0(new_n4878_), .A1(new_n4877_), .B0(new_n3135_), .Y(new_n4879_));
  AOI21X1  g02444(.A0(new_n4876_), .A1(new_n4875_), .B0(new_n4879_), .Y(new_n4880_));
  OAI21X1  g02445(.A0(new_n4864_), .A1(new_n3135_), .B0(new_n3128_), .Y(new_n4881_));
  OR4X1    g02446(.A(new_n4858_), .B(new_n4828_), .C(new_n4756_), .D(new_n3131_), .Y(new_n4882_));
  AOI21X1  g02447(.A0(new_n4862_), .A1(new_n3131_), .B0(new_n3128_), .Y(new_n4883_));
  AOI21X1  g02448(.A0(new_n4883_), .A1(new_n4882_), .B0(pi0056), .Y(new_n4884_));
  OAI21X1  g02449(.A0(new_n4881_), .A1(new_n4880_), .B0(new_n4884_), .Y(new_n4885_));
  OAI21X1  g02450(.A0(new_n4858_), .A1(new_n4793_), .B0(new_n3140_), .Y(new_n4886_));
  INVX1    g02451(.A(new_n4862_), .Y(new_n4887_));
  AOI21X1  g02452(.A0(new_n4887_), .A1(new_n3242_), .B0(new_n3143_), .Y(new_n4888_));
  AOI21X1  g02453(.A0(new_n4888_), .A1(new_n4886_), .B0(pi0062), .Y(new_n4889_));
  NOR3X1   g02454(.A(new_n4858_), .B(new_n4793_), .C(new_n3249_), .Y(new_n4890_));
  OAI21X1  g02455(.A0(new_n4887_), .A1(new_n3248_), .B0(pi0062), .Y(new_n4891_));
  OAI21X1  g02456(.A0(new_n4891_), .A1(new_n4890_), .B0(new_n3246_), .Y(new_n4892_));
  AOI21X1  g02457(.A0(new_n4889_), .A1(new_n4885_), .B0(new_n4892_), .Y(new_n4893_));
  INVX1    g02458(.A(pi0242), .Y(new_n4894_));
  OAI21X1  g02459(.A0(new_n4887_), .A1(new_n3246_), .B0(new_n4894_), .Y(new_n4895_));
  OAI22X1  g02460(.A0(new_n4895_), .A1(new_n4893_), .B0(new_n4841_), .B1(new_n4840_), .Y(new_n4896_));
  AOI21X1  g02461(.A0(new_n4779_), .A1(new_n4780_), .B0(pi0039), .Y(new_n4897_));
  AND2X1   g02462(.A(pi0299), .B(new_n2954_), .Y(new_n4898_));
  OAI21X1  g02463(.A0(new_n4769_), .A1(new_n4756_), .B0(new_n4898_), .Y(new_n4899_));
  NOR2X1   g02464(.A(new_n2962_), .B(pi0223), .Y(new_n4900_));
  AOI21X1  g02465(.A0(new_n4790_), .A1(new_n4900_), .B0(pi0299), .Y(new_n4901_));
  OAI21X1  g02466(.A0(new_n4799_), .A1(new_n4756_), .B0(new_n2954_), .Y(new_n4902_));
  AOI21X1  g02467(.A0(new_n4902_), .A1(pi0299), .B0(new_n4901_), .Y(new_n4903_));
  OAI21X1  g02468(.A0(new_n4903_), .A1(new_n2959_), .B0(new_n2996_), .Y(new_n4904_));
  AOI21X1  g02469(.A0(new_n4899_), .A1(new_n4897_), .B0(new_n4904_), .Y(new_n4905_));
  AOI21X1  g02470(.A0(new_n4806_), .A1(new_n4842_), .B0(pi0215), .Y(new_n4906_));
  INVX1    g02471(.A(new_n4906_), .Y(new_n4907_));
  NOR2X1   g02472(.A(new_n4907_), .B(new_n3281_), .Y(new_n4908_));
  INVX1    g02473(.A(new_n4908_), .Y(new_n4909_));
  AOI21X1  g02474(.A0(new_n4909_), .A1(pi0299), .B0(new_n4901_), .Y(new_n4910_));
  INVX1    g02475(.A(new_n4910_), .Y(new_n4911_));
  OAI21X1  g02476(.A0(new_n4911_), .A1(new_n2996_), .B0(new_n3026_), .Y(new_n4912_));
  OAI21X1  g02477(.A0(new_n4812_), .A1(new_n4756_), .B0(new_n2954_), .Y(new_n4913_));
  OR2X1    g02478(.A(new_n4901_), .B(new_n3066_), .Y(new_n4914_));
  AOI21X1  g02479(.A0(new_n4913_), .A1(pi0299), .B0(new_n4914_), .Y(new_n4915_));
  OAI21X1  g02480(.A0(new_n4911_), .A1(new_n3065_), .B0(pi0100), .Y(new_n4916_));
  OAI22X1  g02481(.A0(new_n4916_), .A1(new_n4915_), .B0(new_n4912_), .B1(new_n4905_), .Y(new_n4917_));
  MX2X1    g02482(.A(new_n4910_), .B(new_n4903_), .S0(new_n3085_), .Y(new_n4918_));
  OAI21X1  g02483(.A0(new_n4918_), .A1(new_n3156_), .B0(new_n3095_), .Y(new_n4919_));
  AOI21X1  g02484(.A0(new_n4917_), .A1(new_n3156_), .B0(new_n4919_), .Y(new_n4920_));
  OAI21X1  g02485(.A0(new_n4911_), .A1(new_n3095_), .B0(new_n3100_), .Y(new_n4921_));
  NAND2X1  g02486(.A(new_n4918_), .B(new_n3098_), .Y(new_n4922_));
  AOI21X1  g02487(.A0(new_n4910_), .A1(new_n3101_), .B0(new_n3100_), .Y(new_n4923_));
  AOI21X1  g02488(.A0(new_n4923_), .A1(new_n4922_), .B0(new_n3136_), .Y(new_n4924_));
  OAI21X1  g02489(.A0(new_n4921_), .A1(new_n4920_), .B0(new_n4924_), .Y(new_n4925_));
  AOI21X1  g02490(.A0(new_n4910_), .A1(new_n3136_), .B0(pi0055), .Y(new_n4926_));
  NOR2X1   g02491(.A(new_n4902_), .B(new_n3131_), .Y(new_n4927_));
  OAI21X1  g02492(.A0(new_n4909_), .A1(new_n3130_), .B0(pi0055), .Y(new_n4928_));
  OAI21X1  g02493(.A0(new_n4928_), .A1(new_n4927_), .B0(new_n3143_), .Y(new_n4929_));
  AOI21X1  g02494(.A0(new_n4926_), .A1(new_n4925_), .B0(new_n4929_), .Y(new_n4930_));
  OAI21X1  g02495(.A0(new_n4908_), .A1(new_n3140_), .B0(pi0056), .Y(new_n4931_));
  AOI21X1  g02496(.A0(new_n4902_), .A1(new_n3140_), .B0(new_n4931_), .Y(new_n4932_));
  NOR3X1   g02497(.A(new_n4932_), .B(new_n4930_), .C(pi0062), .Y(new_n4933_));
  NOR2X1   g02498(.A(new_n4902_), .B(new_n3249_), .Y(new_n4934_));
  OAI21X1  g02499(.A0(new_n4909_), .A1(new_n3248_), .B0(pi0062), .Y(new_n4935_));
  OAI21X1  g02500(.A0(new_n4935_), .A1(new_n4934_), .B0(new_n3246_), .Y(new_n4936_));
  AOI21X1  g02501(.A0(new_n4908_), .A1(new_n3393_), .B0(new_n4894_), .Y(new_n4937_));
  OAI21X1  g02502(.A0(new_n4936_), .A1(new_n4933_), .B0(new_n4937_), .Y(new_n4938_));
  NAND2X1  g02503(.A(new_n4850_), .B(new_n4898_), .Y(new_n4939_));
  NAND3X1  g02504(.A(new_n4851_), .B(new_n4776_), .C(new_n4780_), .Y(new_n4940_));
  NAND3X1  g02505(.A(new_n4940_), .B(new_n4939_), .C(new_n4897_), .Y(new_n4941_));
  NAND2X1  g02506(.A(new_n4786_), .B(new_n2964_), .Y(new_n4942_));
  AND2X1   g02507(.A(new_n4942_), .B(new_n4901_), .Y(new_n4943_));
  OAI21X1  g02508(.A0(new_n4858_), .A1(new_n4756_), .B0(new_n2954_), .Y(new_n4944_));
  AOI21X1  g02509(.A0(new_n4944_), .A1(pi0299), .B0(new_n4943_), .Y(new_n4945_));
  INVX1    g02510(.A(new_n4945_), .Y(new_n4946_));
  AOI21X1  g02511(.A0(new_n4946_), .A1(pi0039), .B0(pi0038), .Y(new_n4947_));
  AOI22X1  g02512(.A0(new_n4942_), .A1(new_n4901_), .B0(new_n4907_), .B1(pi0299), .Y(new_n4948_));
  INVX1    g02513(.A(new_n4948_), .Y(new_n4949_));
  OAI21X1  g02514(.A0(new_n4949_), .A1(new_n2996_), .B0(new_n3026_), .Y(new_n4950_));
  AOI21X1  g02515(.A0(new_n4947_), .A1(new_n4941_), .B0(new_n4950_), .Y(new_n4951_));
  OAI21X1  g02516(.A0(new_n4868_), .A1(new_n4756_), .B0(new_n2954_), .Y(new_n4952_));
  OR2X1    g02517(.A(new_n4943_), .B(new_n3066_), .Y(new_n4953_));
  AOI21X1  g02518(.A0(new_n4952_), .A1(pi0299), .B0(new_n4953_), .Y(new_n4954_));
  AND2X1   g02519(.A(new_n4948_), .B(new_n3066_), .Y(new_n4955_));
  NOR3X1   g02520(.A(new_n4955_), .B(new_n4954_), .C(new_n3026_), .Y(new_n4956_));
  OAI21X1  g02521(.A0(new_n4956_), .A1(new_n4951_), .B0(new_n3156_), .Y(new_n4957_));
  MX2X1    g02522(.A(new_n4949_), .B(new_n4946_), .S0(new_n3085_), .Y(new_n4958_));
  AOI21X1  g02523(.A0(new_n4958_), .A1(pi0087), .B0(pi0075), .Y(new_n4959_));
  OAI21X1  g02524(.A0(new_n4949_), .A1(new_n3095_), .B0(new_n3100_), .Y(new_n4960_));
  AOI21X1  g02525(.A0(new_n4959_), .A1(new_n4957_), .B0(new_n4960_), .Y(new_n4961_));
  AOI21X1  g02526(.A0(new_n4948_), .A1(new_n3101_), .B0(new_n3100_), .Y(new_n4962_));
  OAI21X1  g02527(.A0(new_n4958_), .A1(new_n3101_), .B0(new_n4962_), .Y(new_n4963_));
  NAND2X1  g02528(.A(new_n4963_), .B(new_n3135_), .Y(new_n4964_));
  OR2X1    g02529(.A(new_n4964_), .B(new_n4961_), .Y(new_n4965_));
  AOI21X1  g02530(.A0(new_n4948_), .A1(new_n3136_), .B0(pi0055), .Y(new_n4966_));
  NOR2X1   g02531(.A(new_n4944_), .B(new_n3131_), .Y(new_n4967_));
  OAI21X1  g02532(.A0(new_n4907_), .A1(new_n3130_), .B0(pi0055), .Y(new_n4968_));
  OAI21X1  g02533(.A0(new_n4968_), .A1(new_n4967_), .B0(new_n3143_), .Y(new_n4969_));
  AOI21X1  g02534(.A0(new_n4966_), .A1(new_n4965_), .B0(new_n4969_), .Y(new_n4970_));
  OAI21X1  g02535(.A0(new_n4906_), .A1(new_n3140_), .B0(pi0056), .Y(new_n4971_));
  AOI21X1  g02536(.A0(new_n4944_), .A1(new_n3140_), .B0(new_n4971_), .Y(new_n4972_));
  OR2X1    g02537(.A(new_n4972_), .B(pi0062), .Y(new_n4973_));
  AOI21X1  g02538(.A0(new_n4906_), .A1(new_n3249_), .B0(new_n3245_), .Y(new_n4974_));
  OAI21X1  g02539(.A0(new_n4944_), .A1(new_n3249_), .B0(new_n4974_), .Y(new_n4975_));
  AND2X1   g02540(.A(new_n4975_), .B(new_n3246_), .Y(new_n4976_));
  OAI21X1  g02541(.A0(new_n4973_), .A1(new_n4970_), .B0(new_n4976_), .Y(new_n4977_));
  AOI21X1  g02542(.A0(new_n4906_), .A1(new_n3393_), .B0(pi0242), .Y(new_n4978_));
  AOI21X1  g02543(.A0(new_n4978_), .A1(new_n4977_), .B0(new_n4755_), .Y(new_n4979_));
  AOI22X1  g02544(.A0(new_n4979_), .A1(new_n4938_), .B0(new_n4896_), .B1(new_n4755_), .Y(po0165));
  AND2X1   g02545(.A(pi0059), .B(pi0057), .Y(new_n4982_));
  INVX1    g02546(.A(new_n4982_), .Y(new_n4983_));
  NOR3X1   g02547(.A(new_n3149_), .B(new_n3003_), .C(new_n2555_), .Y(new_n4984_));
  OAI21X1  g02548(.A0(new_n4984_), .A1(new_n3246_), .B0(new_n4983_), .Y(new_n4985_));
  INVX1    g02549(.A(new_n4985_), .Y(new_n4986_));
  NOR3X1   g02550(.A(new_n3139_), .B(new_n3136_), .C(pi0055), .Y(new_n4987_));
  AND2X1   g02551(.A(new_n3085_), .B(new_n3000_), .Y(new_n4988_));
  AOI21X1  g02552(.A0(new_n4988_), .A1(new_n4987_), .B0(new_n3143_), .Y(new_n4989_));
  INVX1    g02553(.A(new_n4989_), .Y(new_n4990_));
  INVX1    g02554(.A(pi0074), .Y(new_n4991_));
  NOR4X1   g02555(.A(pi0092), .B(pi0087), .C(pi0075), .D(pi0054), .Y(new_n4992_));
  AOI21X1  g02556(.A0(new_n4992_), .A1(new_n4988_), .B0(new_n4991_), .Y(new_n4993_));
  OR2X1    g02557(.A(new_n4993_), .B(pi0055), .Y(new_n4994_));
  AND2X1   g02558(.A(new_n3000_), .B(new_n2959_), .Y(new_n4995_));
  INVX1    g02559(.A(new_n4995_), .Y(new_n4996_));
  AOI21X1  g02560(.A0(new_n4996_), .A1(pi0038), .B0(pi0100), .Y(new_n4997_));
  INVX1    g02561(.A(new_n4997_), .Y(new_n4998_));
  NOR2X1   g02562(.A(new_n2513_), .B(new_n2502_), .Y(new_n4999_));
  NOR2X1   g02563(.A(new_n4999_), .B(pi0090), .Y(new_n5000_));
  OR4X1    g02564(.A(new_n2685_), .B(new_n2680_), .C(new_n2591_), .D(new_n2498_), .Y(new_n5001_));
  AOI21X1  g02565(.A0(new_n5001_), .A1(new_n2595_), .B0(new_n2588_), .Y(new_n5002_));
  OAI21X1  g02566(.A0(new_n5002_), .A1(pi0108), .B0(new_n2584_), .Y(new_n5003_));
  NOR3X1   g02567(.A(new_n2695_), .B(pi0110), .C(pi0109), .Y(new_n5004_));
  OR2X1    g02568(.A(new_n2574_), .B(new_n2566_), .Y(new_n5005_));
  AOI21X1  g02569(.A0(new_n5004_), .A1(new_n5003_), .B0(new_n5005_), .Y(new_n5006_));
  OR2X1    g02570(.A(pi0091), .B(pi0058), .Y(new_n5007_));
  NOR2X1   g02571(.A(new_n2570_), .B(new_n5007_), .Y(new_n5008_));
  OAI21X1  g02572(.A0(new_n5006_), .A1(pi0047), .B0(new_n5008_), .Y(new_n5009_));
  AOI21X1  g02573(.A0(new_n5009_), .A1(new_n5000_), .B0(new_n2702_), .Y(new_n5010_));
  NOR2X1   g02574(.A(new_n2513_), .B(new_n2520_), .Y(new_n5011_));
  AOI21X1  g02575(.A0(new_n5011_), .A1(new_n2726_), .B0(new_n2531_), .Y(new_n5012_));
  INVX1    g02576(.A(new_n5012_), .Y(new_n5013_));
  OAI21X1  g02577(.A0(new_n5010_), .A1(pi0093), .B0(new_n5013_), .Y(new_n5014_));
  OR2X1    g02578(.A(new_n2515_), .B(pi0070), .Y(new_n5015_));
  AOI21X1  g02579(.A0(new_n5014_), .A1(new_n2518_), .B0(new_n5015_), .Y(new_n5016_));
  OAI21X1  g02580(.A0(new_n5016_), .A1(pi0051), .B0(new_n2556_), .Y(new_n5017_));
  AOI21X1  g02581(.A0(new_n5017_), .A1(new_n2873_), .B0(new_n2554_), .Y(new_n5018_));
  MX2X1    g02582(.A(pi0198), .B(pi0210), .S0(pi0299), .Y(new_n5019_));
  NAND3X1  g02583(.A(new_n2543_), .B(new_n2549_), .C(new_n2518_), .Y(new_n5020_));
  NOR2X1   g02584(.A(new_n5020_), .B(new_n2727_), .Y(new_n5021_));
  NOR2X1   g02585(.A(new_n5021_), .B(new_n2456_), .Y(new_n5022_));
  MX2X1    g02586(.A(new_n5022_), .B(new_n3200_), .S0(new_n5019_), .Y(new_n5023_));
  INVX1    g02587(.A(new_n5023_), .Y(new_n5024_));
  OAI21X1  g02588(.A0(new_n5018_), .A1(new_n2547_), .B0(new_n5024_), .Y(new_n5025_));
  AOI21X1  g02589(.A0(new_n5025_), .A1(new_n2540_), .B0(new_n2716_), .Y(new_n5026_));
  INVX1    g02590(.A(pi0603), .Y(new_n5027_));
  NOR4X1   g02591(.A(pi0642), .B(pi0616), .C(pi0614), .D(new_n5027_), .Y(new_n5028_));
  INVX1    g02592(.A(pi0680), .Y(new_n5029_));
  NOR4X1   g02593(.A(pi0681), .B(new_n5029_), .C(pi0662), .D(pi0661), .Y(new_n5030_));
  NOR2X1   g02594(.A(new_n5030_), .B(new_n5028_), .Y(new_n5031_));
  INVX1    g02595(.A(new_n5031_), .Y(po1101));
  NOR2X1   g02596(.A(pi0468), .B(pi0332), .Y(new_n5033_));
  AND2X1   g02597(.A(pi0984), .B(pi0835), .Y(new_n5034_));
  INVX1    g02598(.A(pi0979), .Y(new_n5035_));
  OR2X1    g02599(.A(pi1001), .B(pi0252), .Y(new_n5036_));
  NAND2X1  g02600(.A(new_n5036_), .B(new_n5035_), .Y(new_n5037_));
  NAND2X1  g02601(.A(pi0950), .B(pi0835), .Y(new_n5038_));
  NOR4X1   g02602(.A(new_n5038_), .B(new_n5037_), .C(new_n5034_), .D(pi0287), .Y(new_n5039_));
  INVX1    g02603(.A(new_n5039_), .Y(new_n5040_));
  NOR2X1   g02604(.A(pi0829), .B(pi0824), .Y(new_n5041_));
  AND2X1   g02605(.A(new_n2722_), .B(pi0824), .Y(new_n5042_));
  NOR3X1   g02606(.A(new_n5042_), .B(new_n2723_), .C(new_n2756_), .Y(new_n5043_));
  NOR4X1   g02607(.A(new_n5043_), .B(new_n5041_), .C(new_n5040_), .D(new_n2755_), .Y(new_n5044_));
  OAI21X1  g02608(.A0(new_n5044_), .A1(new_n5033_), .B0(po1101), .Y(new_n5045_));
  AND2X1   g02609(.A(new_n5033_), .B(new_n3000_), .Y(new_n5046_));
  AOI22X1  g02610(.A0(new_n5046_), .A1(po1101), .B0(new_n5045_), .B1(new_n3630_), .Y(new_n5047_));
  NOR4X1   g02611(.A(pi0977), .B(pi0974), .C(pi0971), .D(pi0969), .Y(new_n5048_));
  NOR4X1   g02612(.A(pi0967), .B(pi0961), .C(pi0602), .D(pi0587), .Y(new_n5049_));
  AND2X1   g02613(.A(new_n5049_), .B(new_n5048_), .Y(new_n5050_));
  INVX1    g02614(.A(new_n5050_), .Y(new_n5051_));
  NOR3X1   g02615(.A(new_n5033_), .B(new_n5030_), .C(new_n5028_), .Y(new_n5052_));
  INVX1    g02616(.A(new_n5052_), .Y(new_n5053_));
  AOI21X1  g02617(.A0(new_n5053_), .A1(new_n5044_), .B0(new_n3074_), .Y(new_n5054_));
  AOI21X1  g02618(.A0(new_n5054_), .A1(new_n5051_), .B0(new_n2964_), .Y(new_n5055_));
  OAI21X1  g02619(.A0(new_n5051_), .A1(new_n5047_), .B0(new_n5055_), .Y(new_n5056_));
  INVX1    g02620(.A(new_n5033_), .Y(new_n5057_));
  MX2X1    g02621(.A(new_n5050_), .B(new_n5031_), .S0(new_n5057_), .Y(new_n5058_));
  AND2X1   g02622(.A(new_n5039_), .B(new_n2778_), .Y(new_n5059_));
  INVX1    g02623(.A(new_n5059_), .Y(new_n5060_));
  NOR4X1   g02624(.A(new_n5060_), .B(new_n5058_), .C(new_n2961_), .D(new_n2960_), .Y(new_n5061_));
  OAI21X1  g02625(.A0(new_n5061_), .A1(new_n3074_), .B0(new_n2964_), .Y(new_n5062_));
  NAND3X1  g02626(.A(new_n5062_), .B(new_n5056_), .C(new_n2953_), .Y(new_n5063_));
  NOR2X1   g02627(.A(pi0947), .B(pi0907), .Y(new_n5064_));
  INVX1    g02628(.A(new_n5064_), .Y(new_n5065_));
  INVX1    g02629(.A(pi0960), .Y(new_n5066_));
  INVX1    g02630(.A(pi0963), .Y(new_n5067_));
  NOR4X1   g02631(.A(pi0978), .B(pi0975), .C(pi0972), .D(pi0970), .Y(new_n5068_));
  NAND3X1  g02632(.A(new_n5068_), .B(new_n5067_), .C(new_n5066_), .Y(new_n5069_));
  NOR2X1   g02633(.A(new_n5069_), .B(new_n5065_), .Y(new_n5070_));
  INVX1    g02634(.A(new_n5070_), .Y(new_n5071_));
  AOI21X1  g02635(.A0(new_n5071_), .A1(new_n5054_), .B0(new_n2954_), .Y(new_n5072_));
  OAI21X1  g02636(.A0(new_n5071_), .A1(new_n5047_), .B0(new_n5072_), .Y(new_n5073_));
  MX2X1    g02637(.A(new_n5070_), .B(new_n5031_), .S0(new_n5057_), .Y(new_n5074_));
  NOR4X1   g02638(.A(new_n5074_), .B(new_n5060_), .C(new_n2437_), .D(new_n2438_), .Y(new_n5075_));
  OAI21X1  g02639(.A0(new_n5075_), .A1(new_n3074_), .B0(new_n2954_), .Y(new_n5076_));
  NAND3X1  g02640(.A(new_n5076_), .B(new_n5073_), .C(pi0299), .Y(new_n5077_));
  NAND3X1  g02641(.A(new_n5077_), .B(new_n5063_), .C(pi0039), .Y(new_n5078_));
  OAI21X1  g02642(.A0(new_n5026_), .A1(pi0039), .B0(new_n5078_), .Y(new_n5079_));
  AOI21X1  g02643(.A0(new_n5079_), .A1(new_n2996_), .B0(new_n4998_), .Y(new_n5080_));
  NOR2X1   g02644(.A(new_n2980_), .B(pi0142), .Y(new_n5081_));
  INVX1    g02645(.A(new_n5081_), .Y(new_n5082_));
  MX2X1    g02646(.A(new_n5082_), .B(new_n3056_), .S0(pi0299), .Y(new_n5083_));
  INVX1    g02647(.A(new_n5083_), .Y(new_n5084_));
  AND2X1   g02648(.A(pi0100), .B(new_n2996_), .Y(new_n5085_));
  INVX1    g02649(.A(new_n5085_), .Y(new_n5086_));
  NOR4X1   g02650(.A(new_n5086_), .B(new_n3003_), .C(new_n2555_), .D(pi0039), .Y(new_n5087_));
  INVX1    g02651(.A(pi0683), .Y(new_n5088_));
  NOR3X1   g02652(.A(pi0101), .B(pi0099), .C(pi0041), .Y(new_n5089_));
  INVX1    g02653(.A(new_n5089_), .Y(new_n5090_));
  OR4X1    g02654(.A(pi0116), .B(pi0115), .C(pi0114), .D(pi0113), .Y(new_n5091_));
  NOR4X1   g02655(.A(new_n5091_), .B(pi0052), .C(pi0043), .D(pi0042), .Y(new_n5092_));
  INVX1    g02656(.A(new_n5092_), .Y(new_n5093_));
  NOR3X1   g02657(.A(new_n5093_), .B(new_n5090_), .C(pi0044), .Y(new_n5094_));
  INVX1    g02658(.A(pi0129), .Y(new_n5095_));
  INVX1    g02659(.A(pi0950), .Y(new_n5096_));
  NOR4X1   g02660(.A(new_n5041_), .B(pi1093), .C(new_n2755_), .D(new_n5096_), .Y(po0740));
  MX2X1    g02661(.A(po0740), .B(new_n5095_), .S0(pi0250), .Y(new_n5098_));
  OR4X1    g02662(.A(new_n5098_), .B(new_n5094_), .C(new_n5083_), .D(new_n5088_), .Y(new_n5099_));
  AND2X1   g02663(.A(new_n5099_), .B(new_n5087_), .Y(new_n5100_));
  OAI21X1  g02664(.A0(new_n5084_), .A1(new_n3216_), .B0(new_n5100_), .Y(new_n5101_));
  AND2X1   g02665(.A(new_n5101_), .B(new_n3156_), .Y(new_n5102_));
  INVX1    g02666(.A(new_n5102_), .Y(new_n5103_));
  OR2X1    g02667(.A(new_n4988_), .B(new_n3156_), .Y(new_n5104_));
  AND2X1   g02668(.A(new_n5104_), .B(new_n3095_), .Y(new_n5105_));
  INVX1    g02669(.A(new_n5105_), .Y(new_n5106_));
  OR2X1    g02670(.A(pi0092), .B(pi0054), .Y(new_n5107_));
  NOR2X1   g02671(.A(new_n5107_), .B(new_n5106_), .Y(new_n5108_));
  OAI21X1  g02672(.A0(new_n5103_), .A1(new_n5080_), .B0(new_n5108_), .Y(new_n5109_));
  AOI21X1  g02673(.A0(new_n5109_), .A1(new_n4991_), .B0(new_n4994_), .Y(new_n5110_));
  OAI21X1  g02674(.A0(new_n5110_), .A1(pi0056), .B0(new_n4990_), .Y(new_n5111_));
  AOI21X1  g02675(.A0(new_n4988_), .A1(new_n3247_), .B0(new_n3245_), .Y(new_n5112_));
  OR2X1    g02676(.A(new_n5112_), .B(pi0059), .Y(new_n5113_));
  AOI21X1  g02677(.A0(new_n5111_), .A1(new_n3245_), .B0(new_n5113_), .Y(new_n5114_));
  MX2X1    g02678(.A(new_n5114_), .B(new_n4986_), .S0(pi0057), .Y(po0167));
  INVX1    g02679(.A(pi1090), .Y(po0170));
  NOR4X1   g02680(.A(pi0062), .B(pi0059), .C(pi0056), .D(pi0055), .Y(new_n5117_));
  INVX1    g02681(.A(new_n5117_), .Y(new_n5118_));
  AOI21X1  g02682(.A0(new_n5118_), .A1(new_n3013_), .B0(new_n2436_), .Y(new_n5119_));
  MX2X1    g02683(.A(pi0907), .B(new_n5030_), .S0(new_n5057_), .Y(new_n5120_));
  AND2X1   g02684(.A(pi0228), .B(pi0030), .Y(new_n5121_));
  INVX1    g02685(.A(new_n5121_), .Y(new_n5122_));
  AOI22X1  g02686(.A0(new_n5122_), .A1(new_n3632_), .B0(new_n3131_), .B1(new_n3013_), .Y(new_n5123_));
  AND2X1   g02687(.A(new_n5123_), .B(new_n5120_), .Y(new_n5124_));
  AND2X1   g02688(.A(new_n5121_), .B(new_n5120_), .Y(new_n5125_));
  OR2X1    g02689(.A(new_n5125_), .B(new_n2953_), .Y(new_n5126_));
  INVX1    g02690(.A(new_n5120_), .Y(new_n5127_));
  INVX1    g02691(.A(pi0158), .Y(new_n5128_));
  INVX1    g02692(.A(pi0159), .Y(new_n5129_));
  NAND2X1  g02693(.A(pi0197), .B(pi0160), .Y(new_n5130_));
  NOR3X1   g02694(.A(new_n5130_), .B(new_n5129_), .C(new_n5128_), .Y(new_n5131_));
  INVX1    g02695(.A(new_n2901_), .Y(new_n5132_));
  NOR3X1   g02696(.A(new_n2870_), .B(pi0096), .C(pi0051), .Y(new_n5133_));
  INVX1    g02697(.A(pi0070), .Y(new_n5134_));
  INVX1    g02698(.A(new_n2702_), .Y(new_n5135_));
  OR2X1    g02699(.A(pi0314), .B(pi0091), .Y(new_n5136_));
  NOR2X1   g02700(.A(new_n2574_), .B(new_n2818_), .Y(new_n5137_));
  INVX1    g02701(.A(new_n2599_), .Y(new_n5138_));
  INVX1    g02702(.A(new_n2687_), .Y(new_n5139_));
  INVX1    g02703(.A(new_n2618_), .Y(new_n5140_));
  INVX1    g02704(.A(new_n2653_), .Y(new_n5141_));
  INVX1    g02705(.A(new_n2468_), .Y(new_n5142_));
  INVX1    g02706(.A(new_n2655_), .Y(new_n5143_));
  NOR2X1   g02707(.A(pi0084), .B(pi0068), .Y(new_n5144_));
  INVX1    g02708(.A(pi0085), .Y(new_n5145_));
  NOR3X1   g02709(.A(new_n2640_), .B(new_n2624_), .C(new_n5145_), .Y(new_n5146_));
  OAI21X1  g02710(.A0(new_n5146_), .A1(new_n2465_), .B0(new_n2644_), .Y(new_n5147_));
  AOI21X1  g02711(.A0(new_n2647_), .A1(pi0068), .B0(new_n2622_), .Y(new_n5148_));
  INVX1    g02712(.A(new_n5148_), .Y(new_n5149_));
  AOI21X1  g02713(.A0(new_n5147_), .A1(new_n5144_), .B0(new_n5149_), .Y(new_n5150_));
  AOI21X1  g02714(.A0(new_n5150_), .A1(new_n5142_), .B0(new_n5143_), .Y(new_n5151_));
  OR2X1    g02715(.A(new_n5151_), .B(new_n5141_), .Y(new_n5152_));
  INVX1    g02716(.A(pi0067), .Y(new_n5153_));
  NOR3X1   g02717(.A(new_n2470_), .B(new_n2465_), .C(new_n5153_), .Y(new_n5154_));
  NOR3X1   g02718(.A(new_n5154_), .B(pi0083), .C(pi0069), .Y(new_n5155_));
  AOI21X1  g02719(.A0(new_n5155_), .A1(new_n5152_), .B0(new_n5140_), .Y(new_n5156_));
  OR2X1    g02720(.A(new_n2472_), .B(pi0064), .Y(po1049));
  NOR3X1   g02721(.A(po1049), .B(new_n2610_), .C(pi0065), .Y(new_n5158_));
  OAI21X1  g02722(.A0(new_n5156_), .A1(pi0071), .B0(new_n5158_), .Y(new_n5159_));
  NAND2X1  g02723(.A(new_n5159_), .B(new_n2509_), .Y(new_n5160_));
  NOR4X1   g02724(.A(po1049), .B(new_n2664_), .C(new_n2610_), .D(pi0065), .Y(new_n5161_));
  OAI21X1  g02725(.A0(new_n2510_), .A1(new_n2509_), .B0(new_n2578_), .Y(new_n5162_));
  NOR3X1   g02726(.A(new_n5162_), .B(new_n2577_), .C(pi0077), .Y(new_n5163_));
  OAI21X1  g02727(.A0(new_n5161_), .A1(new_n5160_), .B0(new_n5163_), .Y(new_n5164_));
  AOI21X1  g02728(.A0(new_n5164_), .A1(new_n2601_), .B0(new_n5139_), .Y(new_n5165_));
  OAI21X1  g02729(.A0(new_n5165_), .A1(new_n2745_), .B0(new_n5138_), .Y(new_n5166_));
  NOR3X1   g02730(.A(new_n2598_), .B(new_n2477_), .C(pi0046), .Y(new_n5167_));
  INVX1    g02731(.A(new_n5167_), .Y(new_n5168_));
  AOI21X1  g02732(.A0(new_n5166_), .A1(new_n2474_), .B0(new_n5168_), .Y(new_n5169_));
  OR2X1    g02733(.A(new_n5169_), .B(new_n2697_), .Y(new_n5170_));
  AOI21X1  g02734(.A0(new_n5170_), .A1(new_n5137_), .B0(new_n5136_), .Y(new_n5171_));
  AOI21X1  g02735(.A0(new_n3255_), .A1(pi0091), .B0(pi0058), .Y(new_n5172_));
  AND2X1   g02736(.A(pi0314), .B(new_n2530_), .Y(new_n5173_));
  INVX1    g02737(.A(new_n5173_), .Y(new_n5174_));
  INVX1    g02738(.A(new_n5137_), .Y(new_n5175_));
  AOI21X1  g02739(.A0(new_n5163_), .A1(new_n5160_), .B0(new_n2602_), .Y(new_n5176_));
  OAI21X1  g02740(.A0(new_n5176_), .A1(new_n5139_), .B0(new_n2496_), .Y(new_n5177_));
  AOI21X1  g02741(.A0(new_n5177_), .A1(new_n5138_), .B0(pi0086), .Y(new_n5178_));
  NOR2X1   g02742(.A(new_n5178_), .B(new_n5168_), .Y(new_n5179_));
  INVX1    g02743(.A(new_n5179_), .Y(new_n5180_));
  AOI21X1  g02744(.A0(new_n5180_), .A1(new_n2696_), .B0(new_n5175_), .Y(new_n5181_));
  OAI21X1  g02745(.A0(new_n5181_), .A1(new_n5174_), .B0(new_n5172_), .Y(new_n5182_));
  OAI21X1  g02746(.A0(new_n5182_), .A1(new_n5171_), .B0(new_n2701_), .Y(new_n5183_));
  AOI21X1  g02747(.A0(new_n5183_), .A1(new_n5135_), .B0(pi0093), .Y(new_n5184_));
  NOR3X1   g02748(.A(new_n2513_), .B(new_n2520_), .C(new_n2726_), .Y(new_n5185_));
  OAI21X1  g02749(.A0(new_n5185_), .A1(new_n2531_), .B0(new_n2518_), .Y(new_n5186_));
  OAI21X1  g02750(.A0(new_n5186_), .A1(new_n5184_), .B0(new_n5134_), .Y(new_n5187_));
  AOI21X1  g02751(.A0(new_n5187_), .A1(new_n5133_), .B0(pi0072), .Y(new_n5188_));
  NOR3X1   g02752(.A(pi0095), .B(pi0040), .C(pi0032), .Y(new_n5189_));
  AND2X1   g02753(.A(new_n5189_), .B(new_n2552_), .Y(new_n5190_));
  INVX1    g02754(.A(new_n5190_), .Y(new_n5191_));
  OAI21X1  g02755(.A0(new_n5191_), .A1(new_n5188_), .B0(new_n5132_), .Y(new_n5192_));
  INVX1    g02756(.A(new_n2532_), .Y(new_n5193_));
  OR4X1    g02757(.A(new_n2513_), .B(new_n2520_), .C(pi0841), .D(pi0093), .Y(new_n5194_));
  OR4X1    g02758(.A(new_n5194_), .B(new_n2768_), .C(new_n5193_), .D(new_n2456_), .Y(new_n5195_));
  NOR3X1   g02759(.A(new_n5195_), .B(pi0210), .C(pi0095), .Y(new_n5196_));
  NOR2X1   g02760(.A(new_n5196_), .B(new_n5192_), .Y(new_n5197_));
  INVX1    g02761(.A(new_n5197_), .Y(new_n5198_));
  NOR3X1   g02762(.A(pi0110), .B(pi0109), .C(pi0047), .Y(new_n5199_));
  OR2X1    g02763(.A(new_n5169_), .B(new_n2695_), .Y(new_n5200_));
  AOI21X1  g02764(.A0(new_n5200_), .A1(new_n5199_), .B0(new_n5136_), .Y(new_n5201_));
  INVX1    g02765(.A(new_n2695_), .Y(new_n5202_));
  INVX1    g02766(.A(new_n5199_), .Y(new_n5203_));
  AOI21X1  g02767(.A0(new_n5180_), .A1(new_n5202_), .B0(new_n5203_), .Y(new_n5204_));
  OAI21X1  g02768(.A0(new_n5204_), .A1(new_n5174_), .B0(new_n5172_), .Y(new_n5205_));
  OAI21X1  g02769(.A0(new_n5205_), .A1(new_n5201_), .B0(new_n2701_), .Y(new_n5206_));
  AOI21X1  g02770(.A0(new_n5206_), .A1(new_n5135_), .B0(pi0093), .Y(new_n5207_));
  OAI21X1  g02771(.A0(new_n5207_), .A1(new_n5186_), .B0(new_n5134_), .Y(new_n5208_));
  AOI21X1  g02772(.A0(new_n5208_), .A1(new_n5133_), .B0(pi0072), .Y(new_n5209_));
  OAI21X1  g02773(.A0(new_n5209_), .A1(new_n5191_), .B0(new_n5132_), .Y(new_n5210_));
  OAI21X1  g02774(.A0(new_n5210_), .A1(new_n5196_), .B0(new_n5033_), .Y(new_n5211_));
  INVX1    g02775(.A(new_n5211_), .Y(new_n5212_));
  AOI21X1  g02776(.A0(new_n5198_), .A1(new_n5057_), .B0(new_n5212_), .Y(new_n5213_));
  OAI21X1  g02777(.A0(new_n5213_), .A1(new_n5127_), .B0(new_n5131_), .Y(new_n5214_));
  INVX1    g02778(.A(new_n5131_), .Y(new_n5215_));
  OAI21X1  g02779(.A0(new_n5196_), .A1(new_n5192_), .B0(new_n5120_), .Y(new_n5216_));
  AOI21X1  g02780(.A0(new_n5216_), .A1(new_n5215_), .B0(pi0228), .Y(new_n5217_));
  AOI21X1  g02781(.A0(new_n5217_), .A1(new_n5214_), .B0(new_n5126_), .Y(new_n5218_));
  MX2X1    g02782(.A(pi0602), .B(new_n5030_), .S0(new_n5057_), .Y(new_n5219_));
  NOR3X1   g02783(.A(new_n5195_), .B(pi0198), .C(pi0095), .Y(new_n5220_));
  OR2X1    g02784(.A(new_n5220_), .B(new_n5192_), .Y(new_n5221_));
  MX2X1    g02785(.A(new_n5221_), .B(pi0030), .S0(pi0228), .Y(new_n5222_));
  AOI21X1  g02786(.A0(new_n5222_), .A1(new_n5219_), .B0(pi0299), .Y(new_n5223_));
  INVX1    g02787(.A(pi0145), .Y(new_n5224_));
  INVX1    g02788(.A(pi0180), .Y(new_n5225_));
  INVX1    g02789(.A(pi0181), .Y(new_n5226_));
  INVX1    g02790(.A(pi0182), .Y(new_n5227_));
  NOR4X1   g02791(.A(new_n5227_), .B(new_n5226_), .C(new_n5225_), .D(new_n5224_), .Y(new_n5228_));
  AOI21X1  g02792(.A0(new_n5228_), .A1(new_n2953_), .B0(new_n5223_), .Y(new_n5229_));
  INVX1    g02793(.A(new_n5228_), .Y(new_n5230_));
  NAND2X1  g02794(.A(new_n5219_), .B(new_n5121_), .Y(new_n5231_));
  OR2X1    g02795(.A(new_n5220_), .B(new_n5210_), .Y(new_n5232_));
  MX2X1    g02796(.A(new_n5232_), .B(new_n5221_), .S0(new_n5057_), .Y(new_n5233_));
  NAND3X1  g02797(.A(new_n5233_), .B(new_n5219_), .C(new_n3013_), .Y(new_n5234_));
  AOI21X1  g02798(.A0(new_n5234_), .A1(new_n5231_), .B0(new_n5230_), .Y(new_n5235_));
  OAI21X1  g02799(.A0(new_n5235_), .A1(new_n5229_), .B0(pi0232), .Y(new_n5236_));
  INVX1    g02800(.A(pi0232), .Y(new_n5237_));
  NOR2X1   g02801(.A(new_n5216_), .B(pi0228), .Y(new_n5238_));
  OAI21X1  g02802(.A0(new_n5238_), .A1(new_n5126_), .B0(new_n5237_), .Y(new_n5239_));
  OAI22X1  g02803(.A0(new_n5239_), .A1(new_n5223_), .B0(new_n5236_), .B1(new_n5218_), .Y(new_n5240_));
  AND2X1   g02804(.A(pi0221), .B(new_n2954_), .Y(new_n5241_));
  INVX1    g02805(.A(new_n5241_), .Y(new_n5242_));
  OR4X1    g02806(.A(new_n3003_), .B(new_n2709_), .C(pi0287), .D(pi0070), .Y(new_n5243_));
  INVX1    g02807(.A(pi0984), .Y(new_n5244_));
  NAND4X1  g02808(.A(new_n5036_), .B(new_n5244_), .C(new_n5035_), .D(pi0835), .Y(new_n5245_));
  AND2X1   g02809(.A(pi1093), .B(pi0824), .Y(new_n5246_));
  AND2X1   g02810(.A(new_n5246_), .B(new_n2783_), .Y(new_n5247_));
  INVX1    g02811(.A(new_n5247_), .Y(new_n5248_));
  NOR4X1   g02812(.A(new_n5248_), .B(new_n5245_), .C(new_n5243_), .D(pi1091), .Y(new_n5249_));
  INVX1    g02813(.A(new_n2778_), .Y(new_n5250_));
  INVX1    g02814(.A(pi0824), .Y(new_n5251_));
  INVX1    g02815(.A(new_n2783_), .Y(new_n5252_));
  NOR3X1   g02816(.A(new_n2722_), .B(new_n2780_), .C(pi0833), .Y(new_n5253_));
  OR4X1    g02817(.A(new_n5253_), .B(new_n5252_), .C(new_n2756_), .D(new_n5251_), .Y(new_n5254_));
  AND2X1   g02818(.A(new_n5254_), .B(new_n5250_), .Y(new_n5255_));
  NOR4X1   g02819(.A(new_n5255_), .B(new_n5245_), .C(new_n5243_), .D(new_n2722_), .Y(new_n5256_));
  NOR2X1   g02820(.A(new_n5256_), .B(new_n5249_), .Y(new_n5257_));
  INVX1    g02821(.A(pi0829), .Y(new_n5258_));
  OAI21X1  g02822(.A0(new_n2780_), .A1(pi0833), .B0(new_n5258_), .Y(new_n5259_));
  AND2X1   g02823(.A(new_n5259_), .B(pi1091), .Y(new_n5260_));
  NOR4X1   g02824(.A(new_n5260_), .B(new_n5248_), .C(new_n5245_), .D(new_n5243_), .Y(new_n5261_));
  INVX1    g02825(.A(new_n5261_), .Y(new_n5262_));
  MX2X1    g02826(.A(new_n5262_), .B(new_n5257_), .S0(pi0216), .Y(new_n5263_));
  OR2X1    g02827(.A(new_n5263_), .B(pi0228), .Y(new_n5264_));
  OAI21X1  g02828(.A0(new_n5264_), .A1(new_n5242_), .B0(new_n5122_), .Y(new_n5265_));
  AOI21X1  g02829(.A0(new_n5265_), .A1(new_n5120_), .B0(new_n2953_), .Y(new_n5266_));
  NOR3X1   g02830(.A(new_n5256_), .B(new_n5249_), .C(new_n2961_), .Y(new_n5267_));
  NOR2X1   g02831(.A(new_n5261_), .B(pi0224), .Y(new_n5268_));
  OR4X1    g02832(.A(new_n5268_), .B(new_n5267_), .C(pi0223), .D(new_n2960_), .Y(new_n5269_));
  OAI21X1  g02833(.A0(new_n5269_), .A1(pi0228), .B0(new_n5122_), .Y(new_n5270_));
  AOI21X1  g02834(.A0(new_n5270_), .A1(new_n5219_), .B0(pi0299), .Y(new_n5271_));
  OR2X1    g02835(.A(new_n5271_), .B(new_n2959_), .Y(new_n5272_));
  OAI21X1  g02836(.A0(new_n5272_), .A1(new_n5266_), .B0(new_n2996_), .Y(new_n5273_));
  AOI21X1  g02837(.A0(new_n5240_), .A1(new_n2959_), .B0(new_n5273_), .Y(new_n5274_));
  INVX1    g02838(.A(new_n5219_), .Y(new_n5275_));
  MX2X1    g02839(.A(new_n5275_), .B(new_n5127_), .S0(pi0299), .Y(new_n5276_));
  OAI21X1  g02840(.A0(new_n5121_), .A1(new_n3631_), .B0(new_n2959_), .Y(new_n5277_));
  NOR2X1   g02841(.A(new_n5277_), .B(new_n5276_), .Y(new_n5278_));
  NOR2X1   g02842(.A(new_n5276_), .B(new_n5122_), .Y(new_n5279_));
  NOR3X1   g02843(.A(new_n5279_), .B(new_n5278_), .C(new_n2996_), .Y(new_n5280_));
  OAI21X1  g02844(.A0(new_n5280_), .A1(new_n5274_), .B0(new_n3026_), .Y(new_n5281_));
  INVX1    g02845(.A(new_n5030_), .Y(new_n5282_));
  NOR4X1   g02846(.A(new_n5098_), .B(new_n5094_), .C(new_n3074_), .D(new_n5088_), .Y(new_n5283_));
  INVX1    g02847(.A(new_n5283_), .Y(new_n5284_));
  AOI21X1  g02848(.A0(new_n5057_), .A1(new_n5282_), .B0(new_n5284_), .Y(new_n5285_));
  NAND2X1  g02849(.A(new_n5285_), .B(new_n5081_), .Y(new_n5286_));
  NOR2X1   g02850(.A(new_n5081_), .B(new_n3053_), .Y(new_n5287_));
  INVX1    g02851(.A(new_n5287_), .Y(new_n5288_));
  NAND3X1  g02852(.A(new_n5033_), .B(new_n3000_), .C(pi0252), .Y(new_n5289_));
  OR4X1    g02853(.A(new_n3003_), .B(new_n2709_), .C(new_n3053_), .D(pi0070), .Y(new_n5290_));
  MX2X1    g02854(.A(new_n5290_), .B(new_n5289_), .S0(new_n5282_), .Y(new_n5291_));
  OAI21X1  g02855(.A0(new_n5291_), .A1(new_n5288_), .B0(new_n5286_), .Y(new_n5292_));
  INVX1    g02856(.A(pi0602), .Y(new_n5293_));
  AOI21X1  g02857(.A0(new_n5033_), .A1(new_n5293_), .B0(pi0228), .Y(new_n5294_));
  NAND2X1  g02858(.A(new_n5231_), .B(new_n2953_), .Y(new_n5295_));
  AOI21X1  g02859(.A0(new_n5294_), .A1(new_n5292_), .B0(new_n5295_), .Y(new_n5296_));
  INVX1    g02860(.A(pi0907), .Y(new_n5297_));
  AOI21X1  g02861(.A0(new_n5033_), .A1(new_n5297_), .B0(pi0228), .Y(new_n5298_));
  OAI21X1  g02862(.A0(new_n5285_), .A1(new_n3056_), .B0(new_n5298_), .Y(new_n5299_));
  AOI21X1  g02863(.A0(new_n5291_), .A1(new_n3056_), .B0(new_n5299_), .Y(new_n5300_));
  OAI21X1  g02864(.A0(new_n5300_), .A1(new_n5126_), .B0(new_n3065_), .Y(new_n5301_));
  AOI21X1  g02865(.A0(new_n5279_), .A1(new_n3066_), .B0(new_n3026_), .Y(new_n5302_));
  OAI21X1  g02866(.A0(new_n5301_), .A1(new_n5296_), .B0(new_n5302_), .Y(new_n5303_));
  AND2X1   g02867(.A(new_n5303_), .B(new_n3156_), .Y(new_n5304_));
  INVX1    g02868(.A(new_n5279_), .Y(new_n5305_));
  OAI21X1  g02869(.A0(new_n5305_), .A1(new_n3156_), .B0(new_n3095_), .Y(new_n5306_));
  AOI21X1  g02870(.A0(new_n5304_), .A1(new_n5281_), .B0(new_n5306_), .Y(new_n5307_));
  AOI22X1  g02871(.A0(new_n5279_), .A1(new_n3092_), .B0(new_n5278_), .B1(new_n3108_), .Y(new_n5308_));
  INVX1    g02872(.A(new_n5308_), .Y(new_n5309_));
  OAI21X1  g02873(.A0(new_n5309_), .A1(new_n3095_), .B0(new_n3100_), .Y(new_n5310_));
  NAND2X1  g02874(.A(new_n5308_), .B(new_n3095_), .Y(new_n5311_));
  AOI21X1  g02875(.A0(new_n5305_), .A1(pi0075), .B0(new_n3100_), .Y(new_n5312_));
  AOI21X1  g02876(.A0(new_n5312_), .A1(new_n5311_), .B0(pi0054), .Y(new_n5313_));
  OAI21X1  g02877(.A0(new_n5310_), .A1(new_n5307_), .B0(new_n5313_), .Y(new_n5314_));
  INVX1    g02878(.A(new_n3105_), .Y(new_n5315_));
  MX2X1    g02879(.A(new_n5308_), .B(new_n5305_), .S0(new_n5315_), .Y(new_n5316_));
  AOI21X1  g02880(.A0(new_n5316_), .A1(pi0054), .B0(pi0074), .Y(new_n5317_));
  NOR3X1   g02881(.A(new_n5309_), .B(new_n5315_), .C(pi0054), .Y(new_n5318_));
  NOR3X1   g02882(.A(pi0092), .B(pi0075), .C(pi0054), .Y(new_n5319_));
  OAI21X1  g02883(.A0(new_n5319_), .A1(new_n5279_), .B0(pi0074), .Y(new_n5320_));
  OAI21X1  g02884(.A0(new_n5320_), .A1(new_n5318_), .B0(new_n3128_), .Y(new_n5321_));
  AOI21X1  g02885(.A0(new_n5317_), .A1(new_n5314_), .B0(new_n5321_), .Y(new_n5322_));
  OAI21X1  g02886(.A0(new_n5124_), .A1(new_n3128_), .B0(new_n3148_), .Y(new_n5323_));
  INVX1    g02887(.A(new_n3148_), .Y(new_n5324_));
  AOI21X1  g02888(.A0(new_n5125_), .A1(new_n5324_), .B0(pi0059), .Y(new_n5325_));
  OAI21X1  g02889(.A0(new_n5323_), .A1(new_n5322_), .B0(new_n5325_), .Y(new_n5326_));
  NOR3X1   g02890(.A(pi0062), .B(pi0056), .C(pi0055), .Y(new_n5327_));
  OAI21X1  g02891(.A0(new_n5327_), .A1(pi0228), .B0(new_n5124_), .Y(new_n5328_));
  AOI21X1  g02892(.A0(new_n5328_), .A1(pi0059), .B0(pi0057), .Y(new_n5329_));
  AOI22X1  g02893(.A0(new_n5329_), .A1(new_n5326_), .B0(new_n5124_), .B1(new_n5119_), .Y(po0171));
  MX2X1    g02894(.A(new_n5028_), .B(pi0947), .S0(new_n5033_), .Y(new_n5331_));
  AND2X1   g02895(.A(new_n5331_), .B(new_n5123_), .Y(new_n5332_));
  AND2X1   g02896(.A(new_n5331_), .B(new_n5121_), .Y(new_n5333_));
  OR2X1    g02897(.A(new_n5333_), .B(new_n2953_), .Y(new_n5334_));
  INVX1    g02898(.A(new_n5331_), .Y(new_n5335_));
  OAI21X1  g02899(.A0(new_n5335_), .A1(new_n5213_), .B0(new_n5131_), .Y(new_n5336_));
  OAI21X1  g02900(.A0(new_n5196_), .A1(new_n5192_), .B0(new_n5331_), .Y(new_n5337_));
  AOI21X1  g02901(.A0(new_n5337_), .A1(new_n5215_), .B0(pi0228), .Y(new_n5338_));
  AOI21X1  g02902(.A0(new_n5338_), .A1(new_n5336_), .B0(new_n5334_), .Y(new_n5339_));
  MX2X1    g02903(.A(new_n5028_), .B(pi0587), .S0(new_n5033_), .Y(new_n5340_));
  NAND2X1  g02904(.A(new_n5340_), .B(new_n5121_), .Y(new_n5341_));
  NAND3X1  g02905(.A(new_n5340_), .B(new_n5233_), .C(new_n3013_), .Y(new_n5342_));
  AOI21X1  g02906(.A0(new_n5342_), .A1(new_n5341_), .B0(new_n5230_), .Y(new_n5343_));
  NAND3X1  g02907(.A(new_n5340_), .B(new_n5230_), .C(new_n5222_), .Y(new_n5344_));
  NAND2X1  g02908(.A(new_n5344_), .B(new_n2953_), .Y(new_n5345_));
  OAI21X1  g02909(.A0(new_n5345_), .A1(new_n5343_), .B0(pi0232), .Y(new_n5346_));
  AOI21X1  g02910(.A0(new_n5340_), .A1(new_n5222_), .B0(pi0299), .Y(new_n5347_));
  NOR2X1   g02911(.A(new_n5337_), .B(pi0228), .Y(new_n5348_));
  OAI21X1  g02912(.A0(new_n5348_), .A1(new_n5334_), .B0(new_n5237_), .Y(new_n5349_));
  OAI22X1  g02913(.A0(new_n5349_), .A1(new_n5347_), .B0(new_n5346_), .B1(new_n5339_), .Y(new_n5350_));
  AOI21X1  g02914(.A0(new_n5264_), .A1(new_n5122_), .B0(new_n5242_), .Y(new_n5351_));
  NOR3X1   g02915(.A(new_n2953_), .B(new_n2437_), .C(pi0215), .Y(new_n5352_));
  INVX1    g02916(.A(new_n5352_), .Y(new_n5353_));
  AOI22X1  g02917(.A0(new_n5353_), .A1(new_n5334_), .B0(new_n5331_), .B1(new_n5351_), .Y(new_n5354_));
  AOI21X1  g02918(.A0(new_n5340_), .A1(new_n5270_), .B0(pi0299), .Y(new_n5355_));
  OR2X1    g02919(.A(new_n5355_), .B(new_n2959_), .Y(new_n5356_));
  OAI21X1  g02920(.A0(new_n5356_), .A1(new_n5354_), .B0(new_n2996_), .Y(new_n5357_));
  AOI21X1  g02921(.A0(new_n5350_), .A1(new_n2959_), .B0(new_n5357_), .Y(new_n5358_));
  MX2X1    g02922(.A(new_n5340_), .B(new_n5331_), .S0(pi0299), .Y(new_n5359_));
  INVX1    g02923(.A(new_n5359_), .Y(new_n5360_));
  NOR2X1   g02924(.A(new_n5360_), .B(new_n5277_), .Y(new_n5361_));
  AND2X1   g02925(.A(new_n5359_), .B(new_n5121_), .Y(new_n5362_));
  NOR3X1   g02926(.A(new_n5362_), .B(new_n5361_), .C(new_n2996_), .Y(new_n5363_));
  OAI21X1  g02927(.A0(new_n5363_), .A1(new_n5358_), .B0(new_n3026_), .Y(new_n5364_));
  NOR3X1   g02928(.A(pi0587), .B(pi0468), .C(pi0332), .Y(new_n5365_));
  NOR4X1   g02929(.A(pi0228), .B(pi0189), .C(pi0174), .D(pi0144), .Y(new_n5366_));
  INVX1    g02930(.A(new_n5028_), .Y(new_n5367_));
  MX2X1    g02931(.A(new_n5290_), .B(new_n5289_), .S0(new_n5367_), .Y(new_n5368_));
  OAI21X1  g02932(.A0(new_n5368_), .A1(new_n5365_), .B0(new_n5366_), .Y(new_n5369_));
  AND2X1   g02933(.A(new_n5368_), .B(pi0142), .Y(new_n5370_));
  NOR2X1   g02934(.A(new_n5033_), .B(new_n5028_), .Y(new_n5371_));
  OAI21X1  g02935(.A0(new_n5284_), .A1(new_n5371_), .B0(new_n2972_), .Y(new_n5372_));
  AND2X1   g02936(.A(new_n5057_), .B(new_n5028_), .Y(new_n5373_));
  OR2X1    g02937(.A(new_n5373_), .B(pi0587), .Y(new_n5374_));
  NAND3X1  g02938(.A(new_n5374_), .B(new_n5372_), .C(new_n3013_), .Y(new_n5375_));
  AOI21X1  g02939(.A0(new_n5340_), .A1(new_n5121_), .B0(new_n5366_), .Y(new_n5376_));
  OAI21X1  g02940(.A0(new_n5375_), .A1(new_n5370_), .B0(new_n5376_), .Y(new_n5377_));
  AOI21X1  g02941(.A0(new_n5377_), .A1(new_n5369_), .B0(pi0299), .Y(new_n5378_));
  OAI21X1  g02942(.A0(new_n5057_), .A1(pi0947), .B0(new_n2830_), .Y(new_n5379_));
  NOR3X1   g02943(.A(new_n5379_), .B(new_n5284_), .C(new_n5371_), .Y(new_n5380_));
  OAI21X1  g02944(.A0(new_n5373_), .A1(pi0947), .B0(new_n3056_), .Y(new_n5381_));
  NOR2X1   g02945(.A(new_n5381_), .B(new_n5368_), .Y(new_n5382_));
  OR2X1    g02946(.A(new_n5382_), .B(new_n5380_), .Y(new_n5383_));
  AOI21X1  g02947(.A0(new_n5383_), .A1(new_n3013_), .B0(new_n5334_), .Y(new_n5384_));
  OR4X1    g02948(.A(new_n5384_), .B(new_n5378_), .C(pi0039), .D(pi0038), .Y(new_n5385_));
  AOI21X1  g02949(.A0(new_n5362_), .A1(new_n3066_), .B0(new_n3026_), .Y(new_n5386_));
  AOI21X1  g02950(.A0(new_n5386_), .A1(new_n5385_), .B0(pi0087), .Y(new_n5387_));
  INVX1    g02951(.A(new_n5362_), .Y(new_n5388_));
  OAI21X1  g02952(.A0(new_n5388_), .A1(new_n3156_), .B0(new_n3095_), .Y(new_n5389_));
  AOI21X1  g02953(.A0(new_n5387_), .A1(new_n5364_), .B0(new_n5389_), .Y(new_n5390_));
  AOI22X1  g02954(.A0(new_n5362_), .A1(new_n3092_), .B0(new_n5361_), .B1(new_n3108_), .Y(new_n5391_));
  INVX1    g02955(.A(new_n5391_), .Y(new_n5392_));
  OAI21X1  g02956(.A0(new_n5392_), .A1(new_n3095_), .B0(new_n3100_), .Y(new_n5393_));
  NAND2X1  g02957(.A(new_n5391_), .B(new_n3095_), .Y(new_n5394_));
  AOI21X1  g02958(.A0(new_n5388_), .A1(pi0075), .B0(new_n3100_), .Y(new_n5395_));
  AOI21X1  g02959(.A0(new_n5395_), .A1(new_n5394_), .B0(pi0054), .Y(new_n5396_));
  OAI21X1  g02960(.A0(new_n5393_), .A1(new_n5390_), .B0(new_n5396_), .Y(new_n5397_));
  MX2X1    g02961(.A(new_n5391_), .B(new_n5388_), .S0(new_n5315_), .Y(new_n5398_));
  AOI21X1  g02962(.A0(new_n5398_), .A1(pi0054), .B0(pi0074), .Y(new_n5399_));
  NOR3X1   g02963(.A(new_n5392_), .B(new_n5315_), .C(pi0054), .Y(new_n5400_));
  OAI21X1  g02964(.A0(new_n5362_), .A1(new_n5319_), .B0(pi0074), .Y(new_n5401_));
  OAI21X1  g02965(.A0(new_n5401_), .A1(new_n5400_), .B0(new_n3128_), .Y(new_n5402_));
  AOI21X1  g02966(.A0(new_n5399_), .A1(new_n5397_), .B0(new_n5402_), .Y(new_n5403_));
  OAI21X1  g02967(.A0(new_n5332_), .A1(new_n3128_), .B0(new_n3148_), .Y(new_n5404_));
  AOI21X1  g02968(.A0(new_n5333_), .A1(new_n5324_), .B0(pi0059), .Y(new_n5405_));
  OAI21X1  g02969(.A0(new_n5404_), .A1(new_n5403_), .B0(new_n5405_), .Y(new_n5406_));
  OAI21X1  g02970(.A0(new_n5327_), .A1(pi0228), .B0(new_n5332_), .Y(new_n5407_));
  AOI21X1  g02971(.A0(new_n5407_), .A1(pi0059), .B0(pi0057), .Y(new_n5408_));
  AOI22X1  g02972(.A0(new_n5408_), .A1(new_n5406_), .B0(new_n5332_), .B1(new_n5119_), .Y(po0172));
  INVX1    g02973(.A(pi0970), .Y(new_n5410_));
  INVX1    g02974(.A(pi0030), .Y(new_n5411_));
  NOR4X1   g02975(.A(pi0468), .B(pi0332), .C(new_n3013_), .D(new_n5411_), .Y(new_n5412_));
  INVX1    g02976(.A(new_n5412_), .Y(new_n5413_));
  AND2X1   g02977(.A(pi0970), .B(new_n3013_), .Y(new_n5414_));
  NAND4X1  g02978(.A(new_n5414_), .B(new_n5117_), .C(new_n5046_), .D(new_n3130_), .Y(new_n5415_));
  OAI21X1  g02979(.A0(new_n5413_), .A1(new_n5410_), .B0(new_n5415_), .Y(new_n5416_));
  AND2X1   g02980(.A(pi0159), .B(pi0158), .Y(new_n5417_));
  INVX1    g02981(.A(new_n5414_), .Y(new_n5418_));
  AOI21X1  g02982(.A0(new_n5412_), .A1(pi0970), .B0(new_n2953_), .Y(new_n5419_));
  OAI21X1  g02983(.A0(new_n5196_), .A1(new_n5192_), .B0(new_n5033_), .Y(new_n5420_));
  OAI21X1  g02984(.A0(new_n5420_), .A1(new_n5418_), .B0(new_n5419_), .Y(new_n5421_));
  NAND3X1  g02985(.A(pi0299), .B(pi0159), .C(pi0158), .Y(new_n5422_));
  MX2X1    g02986(.A(new_n5212_), .B(new_n5198_), .S0(new_n5130_), .Y(new_n5423_));
  NAND2X1  g02987(.A(new_n5423_), .B(new_n5033_), .Y(new_n5424_));
  OAI22X1  g02988(.A0(new_n5424_), .A1(new_n5418_), .B0(new_n5413_), .B1(new_n5410_), .Y(new_n5425_));
  AOI22X1  g02989(.A0(new_n5425_), .A1(new_n5417_), .B0(new_n5422_), .B1(new_n5421_), .Y(new_n5426_));
  AOI21X1  g02990(.A0(new_n5222_), .A1(new_n5033_), .B0(new_n5228_), .Y(new_n5427_));
  NAND3X1  g02991(.A(new_n5232_), .B(new_n5033_), .C(new_n3013_), .Y(new_n5428_));
  OAI21X1  g02992(.A0(new_n5220_), .A1(new_n5192_), .B0(new_n5230_), .Y(new_n5429_));
  AND2X1   g02993(.A(new_n5429_), .B(new_n5413_), .Y(new_n5430_));
  AOI21X1  g02994(.A0(new_n5430_), .A1(new_n5428_), .B0(new_n5427_), .Y(new_n5431_));
  AOI21X1  g02995(.A0(new_n5431_), .A1(pi0967), .B0(pi0299), .Y(new_n5432_));
  OR2X1    g02996(.A(new_n5432_), .B(new_n5237_), .Y(new_n5433_));
  AND2X1   g02997(.A(new_n5222_), .B(new_n5033_), .Y(new_n5434_));
  AOI21X1  g02998(.A0(new_n5434_), .A1(pi0967), .B0(pi0299), .Y(new_n5435_));
  NAND2X1  g02999(.A(new_n5421_), .B(new_n5237_), .Y(new_n5436_));
  OAI22X1  g03000(.A0(new_n5436_), .A1(new_n5435_), .B0(new_n5433_), .B1(new_n5426_), .Y(new_n5437_));
  AND2X1   g03001(.A(pi0970), .B(pi0299), .Y(new_n5438_));
  NOR3X1   g03002(.A(new_n5263_), .B(new_n5242_), .C(new_n5057_), .Y(new_n5439_));
  OR2X1    g03003(.A(new_n5439_), .B(pi0228), .Y(new_n5440_));
  AND2X1   g03004(.A(pi0967), .B(new_n2953_), .Y(new_n5441_));
  OAI21X1  g03005(.A0(new_n5269_), .A1(new_n5057_), .B0(new_n3013_), .Y(new_n5442_));
  AOI22X1  g03006(.A0(new_n5442_), .A1(new_n5441_), .B0(new_n5440_), .B1(new_n5438_), .Y(new_n5443_));
  AOI21X1  g03007(.A0(new_n5033_), .A1(pi0030), .B0(new_n3013_), .Y(new_n5444_));
  OR2X1    g03008(.A(new_n5444_), .B(new_n2959_), .Y(new_n5445_));
  OAI21X1  g03009(.A0(new_n5445_), .A1(new_n5443_), .B0(new_n2996_), .Y(new_n5446_));
  AOI21X1  g03010(.A0(new_n5437_), .A1(new_n2959_), .B0(new_n5446_), .Y(new_n5447_));
  INVX1    g03011(.A(new_n5046_), .Y(new_n5448_));
  AOI21X1  g03012(.A0(new_n5448_), .A1(new_n3013_), .B0(new_n5444_), .Y(new_n5449_));
  AOI21X1  g03013(.A0(new_n5449_), .A1(pi0967), .B0(pi0299), .Y(new_n5450_));
  OAI21X1  g03014(.A0(new_n5418_), .A1(new_n5448_), .B0(new_n5419_), .Y(new_n5451_));
  NAND2X1  g03015(.A(new_n5451_), .B(new_n2959_), .Y(new_n5452_));
  NOR2X1   g03016(.A(new_n5452_), .B(new_n5450_), .Y(new_n5453_));
  OAI21X1  g03017(.A0(new_n5441_), .A1(new_n5438_), .B0(new_n5412_), .Y(new_n5454_));
  OAI21X1  g03018(.A0(new_n5454_), .A1(new_n2959_), .B0(pi0038), .Y(new_n5455_));
  NOR2X1   g03019(.A(new_n5455_), .B(new_n5453_), .Y(new_n5456_));
  OAI21X1  g03020(.A0(new_n5456_), .A1(new_n5447_), .B0(new_n3026_), .Y(new_n5457_));
  NOR2X1   g03021(.A(new_n5289_), .B(new_n5081_), .Y(new_n5458_));
  NOR3X1   g03022(.A(new_n5284_), .B(new_n5082_), .C(new_n5057_), .Y(new_n5459_));
  NOR3X1   g03023(.A(new_n5459_), .B(new_n5458_), .C(pi0228), .Y(new_n5460_));
  NOR2X1   g03024(.A(new_n5460_), .B(new_n5444_), .Y(new_n5461_));
  AND2X1   g03025(.A(new_n5461_), .B(pi0967), .Y(new_n5462_));
  AND2X1   g03026(.A(new_n5289_), .B(new_n3056_), .Y(new_n5463_));
  AOI21X1  g03027(.A0(new_n5283_), .A1(new_n5033_), .B0(new_n3056_), .Y(new_n5464_));
  OR4X1    g03028(.A(new_n5464_), .B(new_n5463_), .C(new_n5410_), .D(pi0228), .Y(new_n5465_));
  AOI21X1  g03029(.A0(new_n5465_), .A1(new_n5419_), .B0(new_n3066_), .Y(new_n5466_));
  OAI21X1  g03030(.A0(new_n5462_), .A1(pi0299), .B0(new_n5466_), .Y(new_n5467_));
  INVX1    g03031(.A(new_n5454_), .Y(new_n5468_));
  AOI21X1  g03032(.A0(new_n5468_), .A1(new_n3066_), .B0(new_n3026_), .Y(new_n5469_));
  AOI21X1  g03033(.A0(new_n5469_), .A1(new_n5467_), .B0(pi0087), .Y(new_n5470_));
  OAI21X1  g03034(.A0(new_n5454_), .A1(new_n3156_), .B0(new_n3095_), .Y(new_n5471_));
  AOI21X1  g03035(.A0(new_n5470_), .A1(new_n5457_), .B0(new_n5471_), .Y(new_n5472_));
  AOI22X1  g03036(.A0(new_n5468_), .A1(new_n3092_), .B0(new_n5453_), .B1(new_n3108_), .Y(new_n5473_));
  INVX1    g03037(.A(new_n5473_), .Y(new_n5474_));
  OAI21X1  g03038(.A0(new_n5474_), .A1(new_n3095_), .B0(new_n3100_), .Y(new_n5475_));
  NAND2X1  g03039(.A(new_n5473_), .B(new_n3095_), .Y(new_n5476_));
  AOI21X1  g03040(.A0(new_n5454_), .A1(pi0075), .B0(new_n3100_), .Y(new_n5477_));
  AOI21X1  g03041(.A0(new_n5477_), .A1(new_n5476_), .B0(pi0054), .Y(new_n5478_));
  OAI21X1  g03042(.A0(new_n5475_), .A1(new_n5472_), .B0(new_n5478_), .Y(new_n5479_));
  MX2X1    g03043(.A(new_n5473_), .B(new_n5454_), .S0(new_n5315_), .Y(new_n5480_));
  AOI21X1  g03044(.A0(new_n5480_), .A1(pi0054), .B0(pi0074), .Y(new_n5481_));
  NOR3X1   g03045(.A(new_n5474_), .B(new_n5315_), .C(pi0054), .Y(new_n5482_));
  OAI21X1  g03046(.A0(new_n5468_), .A1(new_n5319_), .B0(pi0074), .Y(new_n5483_));
  OAI21X1  g03047(.A0(new_n5483_), .A1(new_n5482_), .B0(new_n3128_), .Y(new_n5484_));
  AOI21X1  g03048(.A0(new_n5481_), .A1(new_n5479_), .B0(new_n5484_), .Y(new_n5485_));
  NOR4X1   g03049(.A(new_n5418_), .B(new_n5057_), .C(new_n3131_), .D(new_n3015_), .Y(new_n5486_));
  AND2X1   g03050(.A(new_n5412_), .B(pi0970), .Y(new_n5487_));
  OR2X1    g03051(.A(new_n5487_), .B(new_n3128_), .Y(new_n5488_));
  OAI21X1  g03052(.A0(new_n5488_), .A1(new_n5486_), .B0(new_n3148_), .Y(new_n5489_));
  AOI21X1  g03053(.A0(new_n5487_), .A1(new_n5324_), .B0(pi0059), .Y(new_n5490_));
  OAI21X1  g03054(.A0(new_n5489_), .A1(new_n5485_), .B0(new_n5490_), .Y(new_n5491_));
  NAND4X1  g03055(.A(new_n5414_), .B(new_n5327_), .C(new_n5046_), .D(new_n3130_), .Y(new_n5492_));
  AOI21X1  g03056(.A0(new_n5412_), .A1(pi0970), .B0(new_n3153_), .Y(new_n5493_));
  AOI21X1  g03057(.A0(new_n5493_), .A1(new_n5492_), .B0(pi0057), .Y(new_n5494_));
  AOI22X1  g03058(.A0(new_n5494_), .A1(new_n5491_), .B0(new_n5416_), .B1(pi0057), .Y(po0173));
  INVX1    g03059(.A(pi0972), .Y(new_n5496_));
  AND2X1   g03060(.A(pi0972), .B(new_n3013_), .Y(new_n5497_));
  NAND4X1  g03061(.A(new_n5497_), .B(new_n5117_), .C(new_n5046_), .D(new_n3130_), .Y(new_n5498_));
  OAI21X1  g03062(.A0(new_n5413_), .A1(new_n5496_), .B0(new_n5498_), .Y(new_n5499_));
  INVX1    g03063(.A(new_n5497_), .Y(new_n5500_));
  AOI21X1  g03064(.A0(new_n5412_), .A1(pi0972), .B0(new_n2953_), .Y(new_n5501_));
  OAI21X1  g03065(.A0(new_n5500_), .A1(new_n5420_), .B0(new_n5501_), .Y(new_n5502_));
  OAI22X1  g03066(.A0(new_n5500_), .A1(new_n5424_), .B0(new_n5413_), .B1(new_n5496_), .Y(new_n5503_));
  AOI22X1  g03067(.A0(new_n5503_), .A1(new_n5417_), .B0(new_n5502_), .B1(new_n5422_), .Y(new_n5504_));
  AOI21X1  g03068(.A0(new_n5431_), .A1(pi0961), .B0(pi0299), .Y(new_n5505_));
  OR2X1    g03069(.A(new_n5505_), .B(new_n5237_), .Y(new_n5506_));
  AOI21X1  g03070(.A0(new_n5434_), .A1(pi0961), .B0(pi0299), .Y(new_n5507_));
  NAND2X1  g03071(.A(new_n5502_), .B(new_n5237_), .Y(new_n5508_));
  OAI22X1  g03072(.A0(new_n5508_), .A1(new_n5507_), .B0(new_n5506_), .B1(new_n5504_), .Y(new_n5509_));
  AND2X1   g03073(.A(pi0961), .B(new_n2953_), .Y(new_n5510_));
  AND2X1   g03074(.A(pi0972), .B(pi0299), .Y(new_n5511_));
  AOI22X1  g03075(.A0(new_n5511_), .A1(new_n5440_), .B0(new_n5510_), .B1(new_n5442_), .Y(new_n5512_));
  OAI21X1  g03076(.A0(new_n5512_), .A1(new_n5445_), .B0(new_n2996_), .Y(new_n5513_));
  AOI21X1  g03077(.A0(new_n5509_), .A1(new_n2959_), .B0(new_n5513_), .Y(new_n5514_));
  AOI21X1  g03078(.A0(new_n5449_), .A1(pi0961), .B0(pi0299), .Y(new_n5515_));
  OAI21X1  g03079(.A0(new_n5500_), .A1(new_n5448_), .B0(new_n5501_), .Y(new_n5516_));
  NAND2X1  g03080(.A(new_n5516_), .B(new_n2959_), .Y(new_n5517_));
  NOR2X1   g03081(.A(new_n5517_), .B(new_n5515_), .Y(new_n5518_));
  OAI21X1  g03082(.A0(new_n5511_), .A1(new_n5510_), .B0(new_n5412_), .Y(new_n5519_));
  OAI21X1  g03083(.A0(new_n5519_), .A1(new_n2959_), .B0(pi0038), .Y(new_n5520_));
  NOR2X1   g03084(.A(new_n5520_), .B(new_n5518_), .Y(new_n5521_));
  OAI21X1  g03085(.A0(new_n5521_), .A1(new_n5514_), .B0(new_n3026_), .Y(new_n5522_));
  AND2X1   g03086(.A(new_n5461_), .B(pi0961), .Y(new_n5523_));
  OR4X1    g03087(.A(new_n5464_), .B(new_n5463_), .C(new_n5496_), .D(pi0228), .Y(new_n5524_));
  AOI21X1  g03088(.A0(new_n5524_), .A1(new_n5501_), .B0(new_n3066_), .Y(new_n5525_));
  OAI21X1  g03089(.A0(new_n5523_), .A1(pi0299), .B0(new_n5525_), .Y(new_n5526_));
  INVX1    g03090(.A(new_n5519_), .Y(new_n5527_));
  AOI21X1  g03091(.A0(new_n5527_), .A1(new_n3066_), .B0(new_n3026_), .Y(new_n5528_));
  AOI21X1  g03092(.A0(new_n5528_), .A1(new_n5526_), .B0(pi0087), .Y(new_n5529_));
  OAI21X1  g03093(.A0(new_n5519_), .A1(new_n3156_), .B0(new_n3095_), .Y(new_n5530_));
  AOI21X1  g03094(.A0(new_n5529_), .A1(new_n5522_), .B0(new_n5530_), .Y(new_n5531_));
  AOI22X1  g03095(.A0(new_n5527_), .A1(new_n3092_), .B0(new_n5518_), .B1(new_n3108_), .Y(new_n5532_));
  INVX1    g03096(.A(new_n5532_), .Y(new_n5533_));
  OAI21X1  g03097(.A0(new_n5533_), .A1(new_n3095_), .B0(new_n3100_), .Y(new_n5534_));
  NAND2X1  g03098(.A(new_n5532_), .B(new_n3095_), .Y(new_n5535_));
  AOI21X1  g03099(.A0(new_n5519_), .A1(pi0075), .B0(new_n3100_), .Y(new_n5536_));
  AOI21X1  g03100(.A0(new_n5536_), .A1(new_n5535_), .B0(pi0054), .Y(new_n5537_));
  OAI21X1  g03101(.A0(new_n5534_), .A1(new_n5531_), .B0(new_n5537_), .Y(new_n5538_));
  MX2X1    g03102(.A(new_n5532_), .B(new_n5519_), .S0(new_n5315_), .Y(new_n5539_));
  AOI21X1  g03103(.A0(new_n5539_), .A1(pi0054), .B0(pi0074), .Y(new_n5540_));
  NOR3X1   g03104(.A(new_n5533_), .B(new_n5315_), .C(pi0054), .Y(new_n5541_));
  OAI21X1  g03105(.A0(new_n5527_), .A1(new_n5319_), .B0(pi0074), .Y(new_n5542_));
  OAI21X1  g03106(.A0(new_n5542_), .A1(new_n5541_), .B0(new_n3128_), .Y(new_n5543_));
  AOI21X1  g03107(.A0(new_n5540_), .A1(new_n5538_), .B0(new_n5543_), .Y(new_n5544_));
  NOR4X1   g03108(.A(new_n5500_), .B(new_n5057_), .C(new_n3131_), .D(new_n3015_), .Y(new_n5545_));
  AND2X1   g03109(.A(new_n5412_), .B(pi0972), .Y(new_n5546_));
  OR2X1    g03110(.A(new_n5546_), .B(new_n3128_), .Y(new_n5547_));
  OAI21X1  g03111(.A0(new_n5547_), .A1(new_n5545_), .B0(new_n3148_), .Y(new_n5548_));
  AOI21X1  g03112(.A0(new_n5546_), .A1(new_n5324_), .B0(pi0059), .Y(new_n5549_));
  OAI21X1  g03113(.A0(new_n5548_), .A1(new_n5544_), .B0(new_n5549_), .Y(new_n5550_));
  NAND4X1  g03114(.A(new_n5497_), .B(new_n5327_), .C(new_n5046_), .D(new_n3130_), .Y(new_n5551_));
  AOI21X1  g03115(.A0(new_n5412_), .A1(pi0972), .B0(new_n3153_), .Y(new_n5552_));
  AOI21X1  g03116(.A0(new_n5552_), .A1(new_n5551_), .B0(pi0057), .Y(new_n5553_));
  AOI22X1  g03117(.A0(new_n5553_), .A1(new_n5550_), .B0(new_n5499_), .B1(pi0057), .Y(po0174));
  AND2X1   g03118(.A(pi0960), .B(new_n3013_), .Y(new_n5555_));
  NAND4X1  g03119(.A(new_n5555_), .B(new_n5117_), .C(new_n5046_), .D(new_n3130_), .Y(new_n5556_));
  OAI21X1  g03120(.A0(new_n5413_), .A1(new_n5066_), .B0(new_n5556_), .Y(new_n5557_));
  INVX1    g03121(.A(new_n5555_), .Y(new_n5558_));
  AOI21X1  g03122(.A0(new_n5412_), .A1(pi0960), .B0(new_n2953_), .Y(new_n5559_));
  OAI21X1  g03123(.A0(new_n5558_), .A1(new_n5420_), .B0(new_n5559_), .Y(new_n5560_));
  OAI22X1  g03124(.A0(new_n5558_), .A1(new_n5424_), .B0(new_n5413_), .B1(new_n5066_), .Y(new_n5561_));
  AOI22X1  g03125(.A0(new_n5561_), .A1(new_n5417_), .B0(new_n5560_), .B1(new_n5422_), .Y(new_n5562_));
  AOI21X1  g03126(.A0(new_n5431_), .A1(pi0977), .B0(pi0299), .Y(new_n5563_));
  OR2X1    g03127(.A(new_n5563_), .B(new_n5237_), .Y(new_n5564_));
  AOI21X1  g03128(.A0(new_n5434_), .A1(pi0977), .B0(pi0299), .Y(new_n5565_));
  NAND2X1  g03129(.A(new_n5560_), .B(new_n5237_), .Y(new_n5566_));
  OAI22X1  g03130(.A0(new_n5566_), .A1(new_n5565_), .B0(new_n5564_), .B1(new_n5562_), .Y(new_n5567_));
  AND2X1   g03131(.A(pi0977), .B(new_n2953_), .Y(new_n5568_));
  AND2X1   g03132(.A(pi0960), .B(pi0299), .Y(new_n5569_));
  AOI22X1  g03133(.A0(new_n5569_), .A1(new_n5440_), .B0(new_n5568_), .B1(new_n5442_), .Y(new_n5570_));
  OAI21X1  g03134(.A0(new_n5570_), .A1(new_n5445_), .B0(new_n2996_), .Y(new_n5571_));
  AOI21X1  g03135(.A0(new_n5567_), .A1(new_n2959_), .B0(new_n5571_), .Y(new_n5572_));
  AOI21X1  g03136(.A0(new_n5449_), .A1(pi0977), .B0(pi0299), .Y(new_n5573_));
  OAI21X1  g03137(.A0(new_n5558_), .A1(new_n5448_), .B0(new_n5559_), .Y(new_n5574_));
  NAND2X1  g03138(.A(new_n5574_), .B(new_n2959_), .Y(new_n5575_));
  NOR2X1   g03139(.A(new_n5575_), .B(new_n5573_), .Y(new_n5576_));
  OAI21X1  g03140(.A0(new_n5569_), .A1(new_n5568_), .B0(new_n5412_), .Y(new_n5577_));
  OAI21X1  g03141(.A0(new_n5577_), .A1(new_n2959_), .B0(pi0038), .Y(new_n5578_));
  NOR2X1   g03142(.A(new_n5578_), .B(new_n5576_), .Y(new_n5579_));
  OAI21X1  g03143(.A0(new_n5579_), .A1(new_n5572_), .B0(new_n3026_), .Y(new_n5580_));
  AND2X1   g03144(.A(new_n5461_), .B(pi0977), .Y(new_n5581_));
  OR4X1    g03145(.A(new_n5464_), .B(new_n5463_), .C(new_n5066_), .D(pi0228), .Y(new_n5582_));
  AOI21X1  g03146(.A0(new_n5582_), .A1(new_n5559_), .B0(new_n3066_), .Y(new_n5583_));
  OAI21X1  g03147(.A0(new_n5581_), .A1(pi0299), .B0(new_n5583_), .Y(new_n5584_));
  INVX1    g03148(.A(new_n5577_), .Y(new_n5585_));
  AOI21X1  g03149(.A0(new_n5585_), .A1(new_n3066_), .B0(new_n3026_), .Y(new_n5586_));
  AOI21X1  g03150(.A0(new_n5586_), .A1(new_n5584_), .B0(pi0087), .Y(new_n5587_));
  OAI21X1  g03151(.A0(new_n5577_), .A1(new_n3156_), .B0(new_n3095_), .Y(new_n5588_));
  AOI21X1  g03152(.A0(new_n5587_), .A1(new_n5580_), .B0(new_n5588_), .Y(new_n5589_));
  AOI22X1  g03153(.A0(new_n5585_), .A1(new_n3092_), .B0(new_n5576_), .B1(new_n3108_), .Y(new_n5590_));
  INVX1    g03154(.A(new_n5590_), .Y(new_n5591_));
  OAI21X1  g03155(.A0(new_n5591_), .A1(new_n3095_), .B0(new_n3100_), .Y(new_n5592_));
  NAND2X1  g03156(.A(new_n5590_), .B(new_n3095_), .Y(new_n5593_));
  AOI21X1  g03157(.A0(new_n5577_), .A1(pi0075), .B0(new_n3100_), .Y(new_n5594_));
  AOI21X1  g03158(.A0(new_n5594_), .A1(new_n5593_), .B0(pi0054), .Y(new_n5595_));
  OAI21X1  g03159(.A0(new_n5592_), .A1(new_n5589_), .B0(new_n5595_), .Y(new_n5596_));
  MX2X1    g03160(.A(new_n5590_), .B(new_n5577_), .S0(new_n5315_), .Y(new_n5597_));
  AOI21X1  g03161(.A0(new_n5597_), .A1(pi0054), .B0(pi0074), .Y(new_n5598_));
  NOR3X1   g03162(.A(new_n5591_), .B(new_n5315_), .C(pi0054), .Y(new_n5599_));
  OAI21X1  g03163(.A0(new_n5585_), .A1(new_n5319_), .B0(pi0074), .Y(new_n5600_));
  OAI21X1  g03164(.A0(new_n5600_), .A1(new_n5599_), .B0(new_n3128_), .Y(new_n5601_));
  AOI21X1  g03165(.A0(new_n5598_), .A1(new_n5596_), .B0(new_n5601_), .Y(new_n5602_));
  NOR4X1   g03166(.A(new_n5558_), .B(new_n5057_), .C(new_n3131_), .D(new_n3015_), .Y(new_n5603_));
  AND2X1   g03167(.A(new_n5412_), .B(pi0960), .Y(new_n5604_));
  OR2X1    g03168(.A(new_n5604_), .B(new_n3128_), .Y(new_n5605_));
  OAI21X1  g03169(.A0(new_n5605_), .A1(new_n5603_), .B0(new_n3148_), .Y(new_n5606_));
  AOI21X1  g03170(.A0(new_n5604_), .A1(new_n5324_), .B0(pi0059), .Y(new_n5607_));
  OAI21X1  g03171(.A0(new_n5606_), .A1(new_n5602_), .B0(new_n5607_), .Y(new_n5608_));
  NAND4X1  g03172(.A(new_n5555_), .B(new_n5327_), .C(new_n5046_), .D(new_n3130_), .Y(new_n5609_));
  AOI21X1  g03173(.A0(new_n5412_), .A1(pi0960), .B0(new_n3153_), .Y(new_n5610_));
  AOI21X1  g03174(.A0(new_n5610_), .A1(new_n5609_), .B0(pi0057), .Y(new_n5611_));
  AOI22X1  g03175(.A0(new_n5611_), .A1(new_n5608_), .B0(new_n5557_), .B1(pi0057), .Y(po0175));
  AND2X1   g03176(.A(pi0963), .B(new_n3013_), .Y(new_n5613_));
  NAND4X1  g03177(.A(new_n5613_), .B(new_n5117_), .C(new_n5046_), .D(new_n3130_), .Y(new_n5614_));
  OAI21X1  g03178(.A0(new_n5413_), .A1(new_n5067_), .B0(new_n5614_), .Y(new_n5615_));
  INVX1    g03179(.A(new_n5613_), .Y(new_n5616_));
  AOI21X1  g03180(.A0(new_n5412_), .A1(pi0963), .B0(new_n2953_), .Y(new_n5617_));
  OAI21X1  g03181(.A0(new_n5616_), .A1(new_n5420_), .B0(new_n5617_), .Y(new_n5618_));
  OAI22X1  g03182(.A0(new_n5616_), .A1(new_n5424_), .B0(new_n5413_), .B1(new_n5067_), .Y(new_n5619_));
  AOI22X1  g03183(.A0(new_n5619_), .A1(new_n5417_), .B0(new_n5618_), .B1(new_n5422_), .Y(new_n5620_));
  AOI21X1  g03184(.A0(new_n5431_), .A1(pi0969), .B0(pi0299), .Y(new_n5621_));
  OR2X1    g03185(.A(new_n5621_), .B(new_n5237_), .Y(new_n5622_));
  AOI21X1  g03186(.A0(new_n5434_), .A1(pi0969), .B0(pi0299), .Y(new_n5623_));
  NAND2X1  g03187(.A(new_n5618_), .B(new_n5237_), .Y(new_n5624_));
  OAI22X1  g03188(.A0(new_n5624_), .A1(new_n5623_), .B0(new_n5622_), .B1(new_n5620_), .Y(new_n5625_));
  AND2X1   g03189(.A(pi0969), .B(new_n2953_), .Y(new_n5626_));
  AND2X1   g03190(.A(pi0963), .B(pi0299), .Y(new_n5627_));
  AOI22X1  g03191(.A0(new_n5627_), .A1(new_n5440_), .B0(new_n5626_), .B1(new_n5442_), .Y(new_n5628_));
  OAI21X1  g03192(.A0(new_n5628_), .A1(new_n5445_), .B0(new_n2996_), .Y(new_n5629_));
  AOI21X1  g03193(.A0(new_n5625_), .A1(new_n2959_), .B0(new_n5629_), .Y(new_n5630_));
  AOI21X1  g03194(.A0(new_n5449_), .A1(pi0969), .B0(pi0299), .Y(new_n5631_));
  OAI21X1  g03195(.A0(new_n5616_), .A1(new_n5448_), .B0(new_n5617_), .Y(new_n5632_));
  NAND2X1  g03196(.A(new_n5632_), .B(new_n2959_), .Y(new_n5633_));
  NOR2X1   g03197(.A(new_n5633_), .B(new_n5631_), .Y(new_n5634_));
  OAI21X1  g03198(.A0(new_n5627_), .A1(new_n5626_), .B0(new_n5412_), .Y(new_n5635_));
  OAI21X1  g03199(.A0(new_n5635_), .A1(new_n2959_), .B0(pi0038), .Y(new_n5636_));
  NOR2X1   g03200(.A(new_n5636_), .B(new_n5634_), .Y(new_n5637_));
  OAI21X1  g03201(.A0(new_n5637_), .A1(new_n5630_), .B0(new_n3026_), .Y(new_n5638_));
  AND2X1   g03202(.A(new_n5461_), .B(pi0969), .Y(new_n5639_));
  OR4X1    g03203(.A(new_n5464_), .B(new_n5463_), .C(new_n5067_), .D(pi0228), .Y(new_n5640_));
  AOI21X1  g03204(.A0(new_n5640_), .A1(new_n5617_), .B0(new_n3066_), .Y(new_n5641_));
  OAI21X1  g03205(.A0(new_n5639_), .A1(pi0299), .B0(new_n5641_), .Y(new_n5642_));
  INVX1    g03206(.A(new_n5635_), .Y(new_n5643_));
  AOI21X1  g03207(.A0(new_n5643_), .A1(new_n3066_), .B0(new_n3026_), .Y(new_n5644_));
  AOI21X1  g03208(.A0(new_n5644_), .A1(new_n5642_), .B0(pi0087), .Y(new_n5645_));
  OAI21X1  g03209(.A0(new_n5635_), .A1(new_n3156_), .B0(new_n3095_), .Y(new_n5646_));
  AOI21X1  g03210(.A0(new_n5645_), .A1(new_n5638_), .B0(new_n5646_), .Y(new_n5647_));
  AOI22X1  g03211(.A0(new_n5643_), .A1(new_n3092_), .B0(new_n5634_), .B1(new_n3108_), .Y(new_n5648_));
  INVX1    g03212(.A(new_n5648_), .Y(new_n5649_));
  OAI21X1  g03213(.A0(new_n5649_), .A1(new_n3095_), .B0(new_n3100_), .Y(new_n5650_));
  NAND2X1  g03214(.A(new_n5648_), .B(new_n3095_), .Y(new_n5651_));
  AOI21X1  g03215(.A0(new_n5635_), .A1(pi0075), .B0(new_n3100_), .Y(new_n5652_));
  AOI21X1  g03216(.A0(new_n5652_), .A1(new_n5651_), .B0(pi0054), .Y(new_n5653_));
  OAI21X1  g03217(.A0(new_n5650_), .A1(new_n5647_), .B0(new_n5653_), .Y(new_n5654_));
  MX2X1    g03218(.A(new_n5648_), .B(new_n5635_), .S0(new_n5315_), .Y(new_n5655_));
  AOI21X1  g03219(.A0(new_n5655_), .A1(pi0054), .B0(pi0074), .Y(new_n5656_));
  NOR3X1   g03220(.A(new_n5649_), .B(new_n5315_), .C(pi0054), .Y(new_n5657_));
  OAI21X1  g03221(.A0(new_n5643_), .A1(new_n5319_), .B0(pi0074), .Y(new_n5658_));
  OAI21X1  g03222(.A0(new_n5658_), .A1(new_n5657_), .B0(new_n3128_), .Y(new_n5659_));
  AOI21X1  g03223(.A0(new_n5656_), .A1(new_n5654_), .B0(new_n5659_), .Y(new_n5660_));
  NOR4X1   g03224(.A(new_n5616_), .B(new_n5057_), .C(new_n3131_), .D(new_n3015_), .Y(new_n5661_));
  AND2X1   g03225(.A(new_n5412_), .B(pi0963), .Y(new_n5662_));
  OR2X1    g03226(.A(new_n5662_), .B(new_n3128_), .Y(new_n5663_));
  OAI21X1  g03227(.A0(new_n5663_), .A1(new_n5661_), .B0(new_n3148_), .Y(new_n5664_));
  AOI21X1  g03228(.A0(new_n5662_), .A1(new_n5324_), .B0(pi0059), .Y(new_n5665_));
  OAI21X1  g03229(.A0(new_n5664_), .A1(new_n5660_), .B0(new_n5665_), .Y(new_n5666_));
  NAND4X1  g03230(.A(new_n5613_), .B(new_n5327_), .C(new_n5046_), .D(new_n3130_), .Y(new_n5667_));
  AOI21X1  g03231(.A0(new_n5412_), .A1(pi0963), .B0(new_n3153_), .Y(new_n5668_));
  AOI21X1  g03232(.A0(new_n5668_), .A1(new_n5667_), .B0(pi0057), .Y(new_n5669_));
  AOI22X1  g03233(.A0(new_n5669_), .A1(new_n5666_), .B0(new_n5615_), .B1(pi0057), .Y(po0176));
  INVX1    g03234(.A(pi0975), .Y(new_n5671_));
  AND2X1   g03235(.A(pi0975), .B(new_n3013_), .Y(new_n5672_));
  NAND4X1  g03236(.A(new_n5672_), .B(new_n5117_), .C(new_n5046_), .D(new_n3130_), .Y(new_n5673_));
  OAI21X1  g03237(.A0(new_n5413_), .A1(new_n5671_), .B0(new_n5673_), .Y(new_n5674_));
  INVX1    g03238(.A(new_n5672_), .Y(new_n5675_));
  AOI21X1  g03239(.A0(new_n5412_), .A1(pi0975), .B0(new_n2953_), .Y(new_n5676_));
  OAI21X1  g03240(.A0(new_n5675_), .A1(new_n5420_), .B0(new_n5676_), .Y(new_n5677_));
  OAI22X1  g03241(.A0(new_n5675_), .A1(new_n5424_), .B0(new_n5413_), .B1(new_n5671_), .Y(new_n5678_));
  AOI22X1  g03242(.A0(new_n5678_), .A1(new_n5417_), .B0(new_n5677_), .B1(new_n5422_), .Y(new_n5679_));
  AOI21X1  g03243(.A0(new_n5431_), .A1(pi0971), .B0(pi0299), .Y(new_n5680_));
  OR2X1    g03244(.A(new_n5680_), .B(new_n5237_), .Y(new_n5681_));
  AOI21X1  g03245(.A0(new_n5434_), .A1(pi0971), .B0(pi0299), .Y(new_n5682_));
  NAND2X1  g03246(.A(new_n5677_), .B(new_n5237_), .Y(new_n5683_));
  OAI22X1  g03247(.A0(new_n5683_), .A1(new_n5682_), .B0(new_n5681_), .B1(new_n5679_), .Y(new_n5684_));
  AND2X1   g03248(.A(pi0971), .B(new_n2953_), .Y(new_n5685_));
  AND2X1   g03249(.A(pi0975), .B(pi0299), .Y(new_n5686_));
  AOI22X1  g03250(.A0(new_n5686_), .A1(new_n5440_), .B0(new_n5685_), .B1(new_n5442_), .Y(new_n5687_));
  OAI21X1  g03251(.A0(new_n5687_), .A1(new_n5445_), .B0(new_n2996_), .Y(new_n5688_));
  AOI21X1  g03252(.A0(new_n5684_), .A1(new_n2959_), .B0(new_n5688_), .Y(new_n5689_));
  AOI21X1  g03253(.A0(new_n5449_), .A1(pi0971), .B0(pi0299), .Y(new_n5690_));
  OAI21X1  g03254(.A0(new_n5675_), .A1(new_n5448_), .B0(new_n5676_), .Y(new_n5691_));
  NAND2X1  g03255(.A(new_n5691_), .B(new_n2959_), .Y(new_n5692_));
  NOR2X1   g03256(.A(new_n5692_), .B(new_n5690_), .Y(new_n5693_));
  OAI21X1  g03257(.A0(new_n5686_), .A1(new_n5685_), .B0(new_n5412_), .Y(new_n5694_));
  OAI21X1  g03258(.A0(new_n5694_), .A1(new_n2959_), .B0(pi0038), .Y(new_n5695_));
  NOR2X1   g03259(.A(new_n5695_), .B(new_n5693_), .Y(new_n5696_));
  OAI21X1  g03260(.A0(new_n5696_), .A1(new_n5689_), .B0(new_n3026_), .Y(new_n5697_));
  AND2X1   g03261(.A(new_n5461_), .B(pi0971), .Y(new_n5698_));
  OR4X1    g03262(.A(new_n5464_), .B(new_n5463_), .C(new_n5671_), .D(pi0228), .Y(new_n5699_));
  AOI21X1  g03263(.A0(new_n5699_), .A1(new_n5676_), .B0(new_n3066_), .Y(new_n5700_));
  OAI21X1  g03264(.A0(new_n5698_), .A1(pi0299), .B0(new_n5700_), .Y(new_n5701_));
  INVX1    g03265(.A(new_n5694_), .Y(new_n5702_));
  AOI21X1  g03266(.A0(new_n5702_), .A1(new_n3066_), .B0(new_n3026_), .Y(new_n5703_));
  AOI21X1  g03267(.A0(new_n5703_), .A1(new_n5701_), .B0(pi0087), .Y(new_n5704_));
  OAI21X1  g03268(.A0(new_n5694_), .A1(new_n3156_), .B0(new_n3095_), .Y(new_n5705_));
  AOI21X1  g03269(.A0(new_n5704_), .A1(new_n5697_), .B0(new_n5705_), .Y(new_n5706_));
  AOI22X1  g03270(.A0(new_n5702_), .A1(new_n3092_), .B0(new_n5693_), .B1(new_n3108_), .Y(new_n5707_));
  INVX1    g03271(.A(new_n5707_), .Y(new_n5708_));
  OAI21X1  g03272(.A0(new_n5708_), .A1(new_n3095_), .B0(new_n3100_), .Y(new_n5709_));
  NAND2X1  g03273(.A(new_n5707_), .B(new_n3095_), .Y(new_n5710_));
  AOI21X1  g03274(.A0(new_n5694_), .A1(pi0075), .B0(new_n3100_), .Y(new_n5711_));
  AOI21X1  g03275(.A0(new_n5711_), .A1(new_n5710_), .B0(pi0054), .Y(new_n5712_));
  OAI21X1  g03276(.A0(new_n5709_), .A1(new_n5706_), .B0(new_n5712_), .Y(new_n5713_));
  MX2X1    g03277(.A(new_n5707_), .B(new_n5694_), .S0(new_n5315_), .Y(new_n5714_));
  AOI21X1  g03278(.A0(new_n5714_), .A1(pi0054), .B0(pi0074), .Y(new_n5715_));
  NOR3X1   g03279(.A(new_n5708_), .B(new_n5315_), .C(pi0054), .Y(new_n5716_));
  OAI21X1  g03280(.A0(new_n5702_), .A1(new_n5319_), .B0(pi0074), .Y(new_n5717_));
  OAI21X1  g03281(.A0(new_n5717_), .A1(new_n5716_), .B0(new_n3128_), .Y(new_n5718_));
  AOI21X1  g03282(.A0(new_n5715_), .A1(new_n5713_), .B0(new_n5718_), .Y(new_n5719_));
  NOR4X1   g03283(.A(new_n5675_), .B(new_n5057_), .C(new_n3131_), .D(new_n3015_), .Y(new_n5720_));
  AND2X1   g03284(.A(new_n5412_), .B(pi0975), .Y(new_n5721_));
  OR2X1    g03285(.A(new_n5721_), .B(new_n3128_), .Y(new_n5722_));
  OAI21X1  g03286(.A0(new_n5722_), .A1(new_n5720_), .B0(new_n3148_), .Y(new_n5723_));
  AOI21X1  g03287(.A0(new_n5721_), .A1(new_n5324_), .B0(pi0059), .Y(new_n5724_));
  OAI21X1  g03288(.A0(new_n5723_), .A1(new_n5719_), .B0(new_n5724_), .Y(new_n5725_));
  NAND4X1  g03289(.A(new_n5672_), .B(new_n5327_), .C(new_n5046_), .D(new_n3130_), .Y(new_n5726_));
  AOI21X1  g03290(.A0(new_n5412_), .A1(pi0975), .B0(new_n3153_), .Y(new_n5727_));
  AOI21X1  g03291(.A0(new_n5727_), .A1(new_n5726_), .B0(pi0057), .Y(new_n5728_));
  AOI22X1  g03292(.A0(new_n5728_), .A1(new_n5725_), .B0(new_n5674_), .B1(pi0057), .Y(po0177));
  AND2X1   g03293(.A(new_n5412_), .B(pi0978), .Y(new_n5730_));
  INVX1    g03294(.A(pi0978), .Y(new_n5731_));
  OR2X1    g03295(.A(new_n5731_), .B(pi0228), .Y(new_n5732_));
  NOR4X1   g03296(.A(new_n5732_), .B(new_n5057_), .C(new_n3131_), .D(new_n3015_), .Y(new_n5733_));
  AND2X1   g03297(.A(new_n5733_), .B(new_n5117_), .Y(new_n5734_));
  OR2X1    g03298(.A(new_n5734_), .B(new_n5730_), .Y(new_n5735_));
  AOI21X1  g03299(.A0(new_n5033_), .A1(new_n3000_), .B0(pi0228), .Y(new_n5736_));
  AND2X1   g03300(.A(pi0978), .B(pi0299), .Y(new_n5737_));
  AOI21X1  g03301(.A0(pi0974), .A1(new_n2953_), .B0(new_n5737_), .Y(new_n5738_));
  NOR3X1   g03302(.A(new_n5738_), .B(new_n5736_), .C(new_n5444_), .Y(new_n5739_));
  NOR4X1   g03303(.A(new_n5738_), .B(new_n5057_), .C(new_n3013_), .D(new_n5411_), .Y(new_n5740_));
  INVX1    g03304(.A(new_n5740_), .Y(new_n5741_));
  OAI21X1  g03305(.A0(new_n5741_), .A1(new_n2959_), .B0(pi0038), .Y(new_n5742_));
  AOI21X1  g03306(.A0(new_n5739_), .A1(new_n2959_), .B0(new_n5742_), .Y(new_n5743_));
  AOI21X1  g03307(.A0(new_n5412_), .A1(pi0978), .B0(new_n2953_), .Y(new_n5744_));
  OAI21X1  g03308(.A0(new_n5732_), .A1(new_n5420_), .B0(new_n5744_), .Y(new_n5745_));
  OAI22X1  g03309(.A0(new_n5732_), .A1(new_n5424_), .B0(new_n5413_), .B1(new_n5731_), .Y(new_n5746_));
  AOI22X1  g03310(.A0(new_n5746_), .A1(new_n5417_), .B0(new_n5745_), .B1(new_n5422_), .Y(new_n5747_));
  AOI21X1  g03311(.A0(new_n5431_), .A1(pi0974), .B0(pi0299), .Y(new_n5748_));
  OR2X1    g03312(.A(new_n5748_), .B(new_n5237_), .Y(new_n5749_));
  AOI21X1  g03313(.A0(new_n5434_), .A1(pi0974), .B0(pi0299), .Y(new_n5750_));
  NAND2X1  g03314(.A(new_n5745_), .B(new_n5237_), .Y(new_n5751_));
  OAI22X1  g03315(.A0(new_n5751_), .A1(new_n5750_), .B0(new_n5749_), .B1(new_n5747_), .Y(new_n5752_));
  AND2X1   g03316(.A(pi0974), .B(new_n2953_), .Y(new_n5753_));
  AOI22X1  g03317(.A0(new_n5737_), .A1(new_n5440_), .B0(new_n5753_), .B1(new_n5442_), .Y(new_n5754_));
  OAI21X1  g03318(.A0(new_n5754_), .A1(new_n5445_), .B0(new_n2996_), .Y(new_n5755_));
  AOI21X1  g03319(.A0(new_n5752_), .A1(new_n2959_), .B0(new_n5755_), .Y(new_n5756_));
  OAI21X1  g03320(.A0(new_n5756_), .A1(new_n5743_), .B0(new_n3026_), .Y(new_n5757_));
  AND2X1   g03321(.A(new_n5461_), .B(pi0974), .Y(new_n5758_));
  OR4X1    g03322(.A(new_n5464_), .B(new_n5463_), .C(new_n5731_), .D(pi0228), .Y(new_n5759_));
  AOI21X1  g03323(.A0(new_n5759_), .A1(new_n5744_), .B0(new_n3066_), .Y(new_n5760_));
  OAI21X1  g03324(.A0(new_n5758_), .A1(pi0299), .B0(new_n5760_), .Y(new_n5761_));
  AOI21X1  g03325(.A0(new_n5740_), .A1(new_n3066_), .B0(new_n3026_), .Y(new_n5762_));
  AOI21X1  g03326(.A0(new_n5762_), .A1(new_n5761_), .B0(pi0087), .Y(new_n5763_));
  OAI21X1  g03327(.A0(new_n5741_), .A1(new_n3156_), .B0(new_n3095_), .Y(new_n5764_));
  AOI21X1  g03328(.A0(new_n5763_), .A1(new_n5757_), .B0(new_n5764_), .Y(new_n5765_));
  OAI21X1  g03329(.A0(new_n3091_), .A1(pi0228), .B0(new_n5739_), .Y(new_n5766_));
  INVX1    g03330(.A(new_n5766_), .Y(new_n5767_));
  OAI21X1  g03331(.A0(new_n5767_), .A1(new_n3095_), .B0(new_n3100_), .Y(new_n5768_));
  OAI21X1  g03332(.A0(new_n5740_), .A1(new_n3095_), .B0(pi0092), .Y(new_n5769_));
  AOI21X1  g03333(.A0(new_n5766_), .A1(new_n3095_), .B0(new_n5769_), .Y(new_n5770_));
  NOR2X1   g03334(.A(new_n5770_), .B(pi0054), .Y(new_n5771_));
  OAI21X1  g03335(.A0(new_n5768_), .A1(new_n5765_), .B0(new_n5771_), .Y(new_n5772_));
  MX2X1    g03336(.A(new_n5766_), .B(new_n5741_), .S0(new_n5315_), .Y(new_n5773_));
  AOI21X1  g03337(.A0(new_n5773_), .A1(pi0054), .B0(pi0074), .Y(new_n5774_));
  NOR3X1   g03338(.A(new_n5767_), .B(new_n5315_), .C(pi0054), .Y(new_n5775_));
  OAI21X1  g03339(.A0(new_n5740_), .A1(new_n5319_), .B0(pi0074), .Y(new_n5776_));
  OAI21X1  g03340(.A0(new_n5776_), .A1(new_n5775_), .B0(new_n3128_), .Y(new_n5777_));
  AOI21X1  g03341(.A0(new_n5774_), .A1(new_n5772_), .B0(new_n5777_), .Y(new_n5778_));
  OR2X1    g03342(.A(new_n5730_), .B(new_n3128_), .Y(new_n5779_));
  OAI21X1  g03343(.A0(new_n5779_), .A1(new_n5733_), .B0(new_n3148_), .Y(new_n5780_));
  AOI21X1  g03344(.A0(new_n5730_), .A1(new_n5324_), .B0(pi0059), .Y(new_n5781_));
  OAI21X1  g03345(.A0(new_n5780_), .A1(new_n5778_), .B0(new_n5781_), .Y(new_n5782_));
  NAND2X1  g03346(.A(new_n5733_), .B(new_n5327_), .Y(new_n5783_));
  AOI21X1  g03347(.A0(new_n5412_), .A1(pi0978), .B0(new_n3153_), .Y(new_n5784_));
  AOI21X1  g03348(.A0(new_n5784_), .A1(new_n5783_), .B0(pi0057), .Y(new_n5785_));
  AOI22X1  g03349(.A0(new_n5785_), .A1(new_n5782_), .B0(new_n5735_), .B1(pi0057), .Y(po0178));
  INVX1    g03350(.A(pi0024), .Y(new_n5787_));
  INVX1    g03351(.A(new_n3108_), .Y(new_n5788_));
  NOR4X1   g03352(.A(new_n5788_), .B(new_n3003_), .C(new_n2555_), .D(pi0039), .Y(new_n5789_));
  NOR2X1   g03353(.A(new_n5789_), .B(new_n3095_), .Y(new_n5790_));
  INVX1    g03354(.A(new_n5790_), .Y(new_n5791_));
  INVX1    g03355(.A(new_n3277_), .Y(new_n5792_));
  NOR4X1   g03356(.A(new_n3101_), .B(new_n5792_), .C(new_n3074_), .D(pi0039), .Y(new_n5793_));
  OR2X1    g03357(.A(new_n5793_), .B(new_n3100_), .Y(new_n5794_));
  AND2X1   g03358(.A(new_n5794_), .B(new_n5791_), .Y(new_n5795_));
  NOR4X1   g03359(.A(new_n5263_), .B(new_n5242_), .C(new_n5074_), .D(new_n2953_), .Y(new_n5796_));
  OR2X1    g03360(.A(new_n5058_), .B(pi0299), .Y(new_n5797_));
  OAI21X1  g03361(.A0(new_n5797_), .A1(new_n5269_), .B0(pi0039), .Y(new_n5798_));
  NAND3X1  g03362(.A(new_n5232_), .B(new_n5228_), .C(new_n5033_), .Y(new_n5799_));
  AOI21X1  g03363(.A0(new_n5221_), .A1(new_n5057_), .B0(pi0299), .Y(new_n5800_));
  NAND3X1  g03364(.A(new_n5800_), .B(new_n5799_), .C(new_n5429_), .Y(new_n5801_));
  INVX1    g03365(.A(new_n5423_), .Y(new_n5802_));
  AOI21X1  g03366(.A0(new_n5198_), .A1(new_n5057_), .B0(new_n5422_), .Y(new_n5803_));
  NAND2X1  g03367(.A(new_n5197_), .B(pi0299), .Y(new_n5804_));
  OAI21X1  g03368(.A0(new_n5804_), .A1(new_n5417_), .B0(pi0232), .Y(new_n5805_));
  AOI21X1  g03369(.A0(new_n5803_), .A1(new_n5802_), .B0(new_n5805_), .Y(new_n5806_));
  AND2X1   g03370(.A(new_n5806_), .B(new_n5801_), .Y(new_n5807_));
  NOR3X1   g03371(.A(new_n5220_), .B(new_n5192_), .C(pi0299), .Y(new_n5808_));
  NAND2X1  g03372(.A(new_n5804_), .B(new_n5237_), .Y(new_n5809_));
  OAI21X1  g03373(.A0(new_n5809_), .A1(new_n5808_), .B0(new_n2959_), .Y(new_n5810_));
  OAI22X1  g03374(.A0(new_n5810_), .A1(new_n5807_), .B0(new_n5798_), .B1(new_n5796_), .Y(new_n5811_));
  MX2X1    g03375(.A(new_n5811_), .B(new_n4996_), .S0(pi0038), .Y(new_n5812_));
  NOR4X1   g03376(.A(new_n3003_), .B(new_n2555_), .C(pi0039), .D(pi0038), .Y(new_n5813_));
  OAI21X1  g03377(.A0(new_n5813_), .A1(new_n3026_), .B0(new_n5102_), .Y(new_n5814_));
  AOI21X1  g03378(.A0(new_n5812_), .A1(new_n3026_), .B0(new_n5814_), .Y(new_n5815_));
  OAI21X1  g03379(.A0(new_n5815_), .A1(new_n5315_), .B0(new_n5795_), .Y(new_n5816_));
  AND2X1   g03380(.A(new_n5793_), .B(new_n3100_), .Y(new_n5817_));
  INVX1    g03381(.A(new_n5817_), .Y(new_n5818_));
  MX2X1    g03382(.A(new_n5818_), .B(new_n5816_), .S0(new_n3112_), .Y(new_n5819_));
  AOI21X1  g03383(.A0(new_n5819_), .A1(new_n4991_), .B0(new_n4993_), .Y(new_n5820_));
  NOR2X1   g03384(.A(new_n3139_), .B(new_n3136_), .Y(new_n5821_));
  AOI21X1  g03385(.A0(new_n4988_), .A1(new_n5821_), .B0(new_n3128_), .Y(new_n5822_));
  NOR3X1   g03386(.A(new_n5822_), .B(pi0062), .C(pi0056), .Y(new_n5823_));
  OAI21X1  g03387(.A0(new_n5820_), .A1(pi0055), .B0(new_n5823_), .Y(new_n5824_));
  AOI21X1  g03388(.A0(new_n5824_), .A1(new_n3246_), .B0(new_n4985_), .Y(po0195));
  MX2X1    g03389(.A(po0195), .B(new_n5787_), .S0(pi0954), .Y(po0182));
  NOR4X1   g03390(.A(new_n3138_), .B(new_n3003_), .C(new_n2555_), .D(pi0228), .Y(new_n5827_));
  AND2X1   g03391(.A(new_n5827_), .B(new_n3247_), .Y(new_n5828_));
  OAI21X1  g03392(.A0(new_n5828_), .A1(new_n3028_), .B0(pi0062), .Y(new_n5829_));
  NOR3X1   g03393(.A(new_n3204_), .B(pi0228), .C(pi0100), .Y(new_n5830_));
  OAI21X1  g03394(.A0(new_n5287_), .A1(new_n3074_), .B0(new_n2953_), .Y(new_n5831_));
  OAI21X1  g03395(.A0(new_n3220_), .A1(new_n2953_), .B0(new_n5831_), .Y(new_n5832_));
  OR4X1    g03396(.A(new_n3003_), .B(new_n2555_), .C(pi0228), .D(new_n3026_), .Y(new_n5833_));
  OAI21X1  g03397(.A0(new_n5833_), .A1(new_n5832_), .B0(new_n2959_), .Y(new_n5834_));
  NOR2X1   g03398(.A(new_n5834_), .B(new_n5830_), .Y(new_n5835_));
  NOR4X1   g03399(.A(new_n3003_), .B(new_n2555_), .C(pi0228), .D(pi0100), .Y(new_n5836_));
  OAI21X1  g03400(.A0(new_n5836_), .A1(new_n2959_), .B0(new_n2996_), .Y(new_n5837_));
  OAI21X1  g03401(.A0(new_n5837_), .A1(new_n5835_), .B0(new_n3030_), .Y(new_n5838_));
  OAI21X1  g03402(.A0(new_n5827_), .A1(new_n3028_), .B0(pi0087), .Y(new_n5839_));
  NAND2X1  g03403(.A(new_n5839_), .B(new_n3095_), .Y(new_n5840_));
  AOI21X1  g03404(.A0(new_n5838_), .A1(new_n3156_), .B0(new_n5840_), .Y(new_n5841_));
  OAI21X1  g03405(.A0(new_n3028_), .A1(new_n3095_), .B0(new_n3100_), .Y(new_n5842_));
  INVX1    g03406(.A(new_n3230_), .Y(new_n5843_));
  NOR4X1   g03407(.A(new_n5843_), .B(new_n3003_), .C(new_n2555_), .D(pi0228), .Y(new_n5844_));
  OAI21X1  g03408(.A0(new_n5844_), .A1(new_n3028_), .B0(pi0092), .Y(new_n5845_));
  AND2X1   g03409(.A(new_n5845_), .B(new_n3135_), .Y(new_n5846_));
  OAI21X1  g03410(.A0(new_n5842_), .A1(new_n5841_), .B0(new_n5846_), .Y(new_n5847_));
  AOI21X1  g03411(.A0(new_n3136_), .A1(new_n3030_), .B0(pi0055), .Y(new_n5848_));
  AND2X1   g03412(.A(new_n4992_), .B(new_n3137_), .Y(new_n5849_));
  INVX1    g03413(.A(new_n5849_), .Y(new_n5850_));
  NOR4X1   g03414(.A(new_n5850_), .B(new_n3003_), .C(new_n2555_), .D(pi0228), .Y(new_n5851_));
  AOI21X1  g03415(.A0(new_n5851_), .A1(new_n4991_), .B0(new_n3028_), .Y(new_n5852_));
  OAI21X1  g03416(.A0(new_n5852_), .A1(new_n3128_), .B0(new_n3143_), .Y(new_n5853_));
  AOI21X1  g03417(.A0(new_n5848_), .A1(new_n5847_), .B0(new_n5853_), .Y(new_n5854_));
  NOR4X1   g03418(.A(new_n3242_), .B(new_n3003_), .C(new_n2555_), .D(pi0228), .Y(new_n5855_));
  OR2X1    g03419(.A(new_n3028_), .B(new_n3143_), .Y(new_n5856_));
  OAI21X1  g03420(.A0(new_n5856_), .A1(new_n5855_), .B0(new_n3245_), .Y(new_n5857_));
  OAI21X1  g03421(.A0(new_n5857_), .A1(new_n5854_), .B0(new_n5829_), .Y(new_n5858_));
  MX2X1    g03422(.A(new_n5858_), .B(new_n3028_), .S0(new_n3393_), .Y(po0183));
  INVX1    g03423(.A(pi0468), .Y(new_n5860_));
  NAND2X1  g03424(.A(pi1056), .B(pi0119), .Y(new_n5861_));
  INVX1    g03425(.A(pi0119), .Y(new_n5862_));
  OAI21X1  g03426(.A0(new_n3053_), .A1(pi0228), .B0(new_n5862_), .Y(new_n5863_));
  NAND3X1  g03427(.A(new_n5863_), .B(new_n5861_), .C(new_n5860_), .Y(po0184));
  NAND2X1  g03428(.A(pi1077), .B(pi0119), .Y(new_n5865_));
  NAND3X1  g03429(.A(new_n5865_), .B(new_n5863_), .C(new_n5860_), .Y(po0185));
  NAND2X1  g03430(.A(pi1073), .B(pi0119), .Y(new_n5867_));
  NAND3X1  g03431(.A(new_n5867_), .B(new_n5863_), .C(new_n5860_), .Y(po0186));
  NAND2X1  g03432(.A(pi1041), .B(pi0119), .Y(new_n5869_));
  NAND3X1  g03433(.A(new_n5869_), .B(new_n5863_), .C(new_n5860_), .Y(po0187));
  XOR2X1   g03434(.A(pi0462), .B(pi0360), .Y(new_n5871_));
  INVX1    g03435(.A(pi0352), .Y(new_n5872_));
  XOR2X1   g03436(.A(pi0353), .B(new_n5872_), .Y(new_n5873_));
  XOR2X1   g03437(.A(new_n5873_), .B(new_n5871_), .Y(new_n5874_));
  XOR2X1   g03438(.A(new_n5874_), .B(pi0354), .Y(new_n5875_));
  INVX1    g03439(.A(new_n5875_), .Y(new_n5876_));
  INVX1    g03440(.A(pi0356), .Y(new_n5877_));
  INVX1    g03441(.A(pi0357), .Y(new_n5878_));
  INVX1    g03442(.A(pi0461), .Y(new_n5879_));
  XOR2X1   g03443(.A(pi0346), .B(pi0345), .Y(new_n5880_));
  XOR2X1   g03444(.A(new_n5880_), .B(pi0323), .Y(new_n5881_));
  INVX1    g03445(.A(pi0358), .Y(new_n5882_));
  XOR2X1   g03446(.A(pi0450), .B(new_n5882_), .Y(new_n5883_));
  XOR2X1   g03447(.A(new_n5883_), .B(new_n5881_), .Y(new_n5884_));
  XOR2X1   g03448(.A(pi0362), .B(pi0327), .Y(new_n5885_));
  XOR2X1   g03449(.A(pi0344), .B(pi0343), .Y(new_n5886_));
  XOR2X1   g03450(.A(new_n5886_), .B(new_n5885_), .Y(new_n5887_));
  INVX1    g03451(.A(new_n5887_), .Y(new_n5888_));
  INVX1    g03452(.A(pi1197), .Y(new_n5889_));
  AOI21X1  g03453(.A0(new_n5888_), .A1(new_n5884_), .B0(new_n5889_), .Y(new_n5890_));
  OAI21X1  g03454(.A0(new_n5888_), .A1(new_n5884_), .B0(new_n5890_), .Y(new_n5891_));
  INVX1    g03455(.A(new_n5891_), .Y(new_n5892_));
  NOR3X1   g03456(.A(pi0092), .B(pi0074), .C(pi0054), .Y(new_n5893_));
  NOR3X1   g03457(.A(new_n5041_), .B(new_n2755_), .C(new_n5096_), .Y(new_n5894_));
  INVX1    g03458(.A(new_n5894_), .Y(new_n5895_));
  INVX1    g03459(.A(new_n2869_), .Y(new_n5896_));
  NOR3X1   g03460(.A(new_n5012_), .B(pi0070), .C(pi0035), .Y(new_n5897_));
  NOR4X1   g03461(.A(new_n2484_), .B(new_n2480_), .C(pi0841), .D(new_n2701_), .Y(new_n5898_));
  NOR2X1   g03462(.A(new_n5898_), .B(pi0093), .Y(new_n5899_));
  INVX1    g03463(.A(new_n5899_), .Y(new_n5900_));
  AOI21X1  g03464(.A0(new_n5900_), .A1(new_n5897_), .B0(pi0051), .Y(new_n5901_));
  INVX1    g03465(.A(new_n5901_), .Y(new_n5902_));
  INVX1    g03466(.A(pi0098), .Y(new_n5903_));
  OR4X1    g03467(.A(new_n2579_), .B(pi0094), .C(pi0077), .D(pi0050), .Y(new_n5904_));
  NOR4X1   g03468(.A(new_n5904_), .B(new_n2476_), .C(new_n5903_), .D(pi0088), .Y(new_n5905_));
  NOR2X1   g03469(.A(new_n5905_), .B(pi0097), .Y(new_n5906_));
  NOR3X1   g03470(.A(pi0093), .B(pi0090), .C(pi0035), .Y(new_n5907_));
  INVX1    g03471(.A(new_n5907_), .Y(new_n5908_));
  NOR4X1   g03472(.A(new_n5908_), .B(new_n5906_), .C(new_n2506_), .D(pi0070), .Y(new_n5909_));
  OAI21X1  g03473(.A0(new_n5909_), .A1(new_n5902_), .B0(new_n5896_), .Y(new_n5910_));
  NAND2X1  g03474(.A(new_n3002_), .B(new_n2526_), .Y(new_n5911_));
  NOR3X1   g03475(.A(new_n5911_), .B(new_n5910_), .C(new_n5895_), .Y(new_n5912_));
  OAI21X1  g03476(.A0(new_n5258_), .A1(pi0122), .B0(new_n5912_), .Y(new_n5913_));
  AND2X1   g03477(.A(new_n5910_), .B(new_n2526_), .Y(new_n5914_));
  OR2X1    g03478(.A(new_n5194_), .B(new_n5193_), .Y(new_n5915_));
  AND2X1   g03479(.A(new_n5915_), .B(pi0096), .Y(new_n5916_));
  NOR4X1   g03480(.A(new_n2755_), .B(new_n5096_), .C(new_n5258_), .D(pi0122), .Y(new_n5917_));
  INVX1    g03481(.A(new_n5917_), .Y(new_n5918_));
  OR4X1    g03482(.A(new_n5918_), .B(new_n5916_), .C(new_n5914_), .D(new_n3256_), .Y(new_n5919_));
  AOI21X1  g03483(.A0(new_n5919_), .A1(new_n5913_), .B0(pi1093), .Y(new_n5920_));
  INVX1    g03484(.A(new_n5920_), .Y(new_n5921_));
  INVX1    g03485(.A(po0740), .Y(new_n5922_));
  NOR3X1   g03486(.A(new_n5922_), .B(new_n3003_), .C(new_n2555_), .Y(new_n5923_));
  NOR4X1   g03487(.A(pi0100), .B(pi0075), .C(pi0039), .D(pi0038), .Y(new_n5924_));
  OAI21X1  g03488(.A0(new_n5923_), .A1(new_n3156_), .B0(new_n5924_), .Y(new_n5925_));
  AOI21X1  g03489(.A0(new_n5921_), .A1(new_n3156_), .B0(new_n5925_), .Y(new_n5926_));
  OAI21X1  g03490(.A0(new_n5926_), .A1(pi0567), .B0(new_n5893_), .Y(new_n5927_));
  INVX1    g03491(.A(pi0567), .Y(new_n5928_));
  MX2X1    g03492(.A(new_n2980_), .B(new_n2451_), .S0(pi0299), .Y(new_n5929_));
  AND2X1   g03493(.A(new_n5033_), .B(pi0232), .Y(new_n5930_));
  AOI21X1  g03494(.A0(new_n5930_), .A1(new_n5929_), .B0(new_n3092_), .Y(new_n5931_));
  NOR4X1   g03495(.A(new_n3003_), .B(new_n2555_), .C(new_n3053_), .D(pi0024), .Y(new_n5932_));
  NOR4X1   g03496(.A(new_n5918_), .B(new_n5094_), .C(new_n2829_), .D(new_n2722_), .Y(new_n5933_));
  NAND4X1  g03497(.A(new_n5933_), .B(new_n5932_), .C(new_n5931_), .D(pi1093), .Y(new_n5934_));
  AND2X1   g03498(.A(new_n5934_), .B(pi0075), .Y(new_n5935_));
  INVX1    g03499(.A(new_n5935_), .Y(new_n5936_));
  AOI21X1  g03500(.A0(pi0957), .A1(new_n2721_), .B0(new_n2756_), .Y(new_n5937_));
  AND2X1   g03501(.A(new_n2783_), .B(pi0824), .Y(new_n5938_));
  INVX1    g03502(.A(new_n5938_), .Y(new_n5939_));
  NOR4X1   g03503(.A(new_n5939_), .B(new_n5911_), .C(new_n5901_), .D(new_n2869_), .Y(new_n5940_));
  NAND2X1  g03504(.A(new_n5940_), .B(new_n5258_), .Y(new_n5941_));
  AND2X1   g03505(.A(new_n2563_), .B(pi0091), .Y(new_n5942_));
  AND2X1   g03506(.A(new_n5942_), .B(new_n5787_), .Y(new_n5943_));
  NAND4X1  g03507(.A(new_n5199_), .B(new_n2576_), .C(pi0097), .D(new_n2694_), .Y(new_n5944_));
  NOR4X1   g03508(.A(new_n5944_), .B(new_n2582_), .C(new_n2586_), .D(pi0091), .Y(new_n5945_));
  OR2X1    g03509(.A(new_n5945_), .B(new_n5943_), .Y(new_n5946_));
  NAND3X1  g03510(.A(new_n5946_), .B(new_n5897_), .C(new_n2519_), .Y(new_n5947_));
  AOI21X1  g03511(.A0(new_n5947_), .A1(new_n5901_), .B0(new_n2869_), .Y(new_n5948_));
  NOR3X1   g03512(.A(new_n5916_), .B(new_n3256_), .C(new_n2785_), .Y(new_n5949_));
  OAI21X1  g03513(.A0(new_n5948_), .A1(pi0096), .B0(new_n5949_), .Y(new_n5950_));
  AOI21X1  g03514(.A0(new_n5950_), .A1(new_n5941_), .B0(pi0122), .Y(new_n5951_));
  INVX1    g03515(.A(pi0122), .Y(new_n5952_));
  OR4X1    g03516(.A(new_n5901_), .B(new_n3256_), .C(new_n2869_), .D(pi0096), .Y(new_n5953_));
  NOR3X1   g03517(.A(new_n5953_), .B(new_n5895_), .C(new_n5952_), .Y(new_n5954_));
  OAI21X1  g03518(.A0(new_n5954_), .A1(new_n5951_), .B0(new_n5937_), .Y(new_n5955_));
  OAI21X1  g03519(.A0(new_n5955_), .A1(new_n2722_), .B0(new_n5921_), .Y(new_n5956_));
  NOR2X1   g03520(.A(new_n5956_), .B(pi0039), .Y(new_n5957_));
  NOR4X1   g03521(.A(new_n5245_), .B(new_n5243_), .C(new_n2738_), .D(new_n2829_), .Y(new_n5958_));
  INVX1    g03522(.A(new_n5958_), .Y(new_n5959_));
  NOR4X1   g03523(.A(new_n5959_), .B(new_n5074_), .C(new_n2740_), .D(new_n2722_), .Y(new_n5960_));
  NAND3X1  g03524(.A(new_n5960_), .B(new_n5352_), .C(new_n2438_), .Y(new_n5961_));
  NOR4X1   g03525(.A(new_n5959_), .B(new_n5058_), .C(new_n2740_), .D(new_n2722_), .Y(new_n5962_));
  NOR4X1   g03526(.A(pi0299), .B(pi0224), .C(pi0223), .D(new_n2960_), .Y(new_n5963_));
  AOI21X1  g03527(.A0(new_n5963_), .A1(new_n5962_), .B0(new_n2959_), .Y(new_n5964_));
  AND2X1   g03528(.A(new_n5964_), .B(new_n5961_), .Y(new_n5965_));
  OR2X1    g03529(.A(new_n5965_), .B(pi0038), .Y(new_n5966_));
  OAI21X1  g03530(.A0(new_n5966_), .A1(new_n5957_), .B0(new_n3026_), .Y(new_n5967_));
  OR4X1    g03531(.A(new_n5965_), .B(new_n5953_), .C(new_n5248_), .D(pi0038), .Y(new_n5968_));
  AOI21X1  g03532(.A0(new_n5955_), .A1(pi1091), .B0(new_n5968_), .Y(new_n5969_));
  AND2X1   g03533(.A(new_n5930_), .B(new_n5929_), .Y(new_n5970_));
  AND2X1   g03534(.A(new_n5917_), .B(pi1093), .Y(new_n5971_));
  INVX1    g03535(.A(new_n5971_), .Y(new_n5972_));
  NOR3X1   g03536(.A(new_n5972_), .B(new_n5094_), .C(new_n2829_), .Y(new_n5973_));
  INVX1    g03537(.A(new_n5973_), .Y(new_n5974_));
  NOR4X1   g03538(.A(new_n5974_), .B(new_n3003_), .C(new_n2555_), .D(new_n2722_), .Y(new_n5975_));
  INVX1    g03539(.A(new_n5975_), .Y(new_n5976_));
  NOR4X1   g03540(.A(new_n5976_), .B(new_n5970_), .C(new_n3066_), .D(new_n3013_), .Y(new_n5977_));
  NOR2X1   g03541(.A(new_n5977_), .B(new_n3026_), .Y(new_n5978_));
  INVX1    g03542(.A(new_n5978_), .Y(new_n5979_));
  OAI21X1  g03543(.A0(new_n5969_), .A1(new_n5967_), .B0(new_n5979_), .Y(new_n5980_));
  NOR3X1   g03544(.A(new_n5939_), .B(new_n3003_), .C(new_n2555_), .Y(new_n5981_));
  AND2X1   g03545(.A(pi1093), .B(new_n2722_), .Y(new_n5982_));
  INVX1    g03546(.A(new_n5982_), .Y(new_n5983_));
  OR2X1    g03547(.A(new_n5983_), .B(new_n5981_), .Y(new_n5984_));
  NOR3X1   g03548(.A(new_n2756_), .B(new_n2780_), .C(pi0833), .Y(new_n5985_));
  NOR4X1   g03549(.A(new_n5985_), .B(new_n5895_), .C(new_n3003_), .D(new_n2555_), .Y(new_n5986_));
  NOR2X1   g03550(.A(new_n5986_), .B(new_n5982_), .Y(new_n5987_));
  NOR2X1   g03551(.A(new_n5987_), .B(new_n3157_), .Y(new_n5988_));
  AOI21X1  g03552(.A0(new_n5988_), .A1(new_n5984_), .B0(new_n3156_), .Y(new_n5989_));
  AOI21X1  g03553(.A0(new_n5980_), .A1(new_n3156_), .B0(new_n5989_), .Y(new_n5990_));
  OR2X1    g03554(.A(new_n5990_), .B(pi0075), .Y(new_n5991_));
  AOI21X1  g03555(.A0(new_n5991_), .A1(new_n5936_), .B0(new_n5928_), .Y(new_n5992_));
  NOR2X1   g03556(.A(new_n5992_), .B(new_n5927_), .Y(new_n5993_));
  INVX1    g03557(.A(new_n5927_), .Y(new_n5994_));
  NOR2X1   g03558(.A(new_n5978_), .B(pi0087), .Y(new_n5995_));
  AND2X1   g03559(.A(new_n5995_), .B(new_n5967_), .Y(new_n5996_));
  NOR2X1   g03560(.A(new_n5986_), .B(new_n2722_), .Y(new_n5997_));
  NOR2X1   g03561(.A(new_n5923_), .B(pi1091), .Y(new_n5998_));
  NAND3X1  g03562(.A(new_n3065_), .B(new_n3026_), .C(pi0087), .Y(new_n5999_));
  NOR3X1   g03563(.A(new_n5999_), .B(new_n5998_), .C(new_n5997_), .Y(new_n6000_));
  NOR3X1   g03564(.A(new_n6000_), .B(new_n5996_), .C(pi0075), .Y(new_n6001_));
  NOR2X1   g03565(.A(new_n6001_), .B(new_n5935_), .Y(new_n6002_));
  OAI21X1  g03566(.A0(new_n6002_), .A1(new_n5928_), .B0(new_n5994_), .Y(new_n6003_));
  INVX1    g03567(.A(new_n6003_), .Y(new_n6004_));
  MX2X1    g03568(.A(new_n6004_), .B(new_n5993_), .S0(pi0592), .Y(new_n6005_));
  INVX1    g03569(.A(new_n5993_), .Y(new_n6006_));
  OR2X1    g03570(.A(pi0592), .B(pi0350), .Y(new_n6007_));
  INVX1    g03571(.A(pi0321), .Y(new_n6008_));
  XOR2X1   g03572(.A(pi0347), .B(new_n6008_), .Y(new_n6009_));
  XOR2X1   g03573(.A(pi0349), .B(pi0316), .Y(new_n6010_));
  XOR2X1   g03574(.A(new_n6010_), .B(pi0348), .Y(new_n6011_));
  INVX1    g03575(.A(pi0315), .Y(new_n6012_));
  XOR2X1   g03576(.A(pi0359), .B(new_n6012_), .Y(new_n6013_));
  XOR2X1   g03577(.A(new_n6013_), .B(pi0322), .Y(new_n6014_));
  XOR2X1   g03578(.A(new_n6014_), .B(new_n6011_), .Y(new_n6015_));
  XOR2X1   g03579(.A(new_n6015_), .B(new_n6009_), .Y(new_n6016_));
  OAI21X1  g03580(.A0(new_n6004_), .A1(new_n6007_), .B0(new_n6016_), .Y(new_n6017_));
  AOI21X1  g03581(.A0(new_n6007_), .A1(new_n6006_), .B0(new_n6017_), .Y(new_n6018_));
  INVX1    g03582(.A(pi0350), .Y(new_n6019_));
  OR2X1    g03583(.A(pi0592), .B(new_n6019_), .Y(new_n6020_));
  INVX1    g03584(.A(new_n6016_), .Y(new_n6021_));
  OAI21X1  g03585(.A0(new_n6020_), .A1(new_n6004_), .B0(new_n6021_), .Y(new_n6022_));
  AOI21X1  g03586(.A0(new_n6020_), .A1(new_n6006_), .B0(new_n6022_), .Y(new_n6023_));
  INVX1    g03587(.A(pi0452), .Y(new_n6024_));
  XOR2X1   g03588(.A(pi0455), .B(new_n6024_), .Y(new_n6025_));
  XOR2X1   g03589(.A(new_n6025_), .B(pi0355), .Y(new_n6026_));
  XOR2X1   g03590(.A(pi0460), .B(pi0320), .Y(new_n6027_));
  XOR2X1   g03591(.A(new_n6027_), .B(pi0342), .Y(new_n6028_));
  INVX1    g03592(.A(pi0361), .Y(new_n6029_));
  XOR2X1   g03593(.A(pi0441), .B(new_n6029_), .Y(new_n6030_));
  XOR2X1   g03594(.A(new_n6030_), .B(new_n6028_), .Y(new_n6031_));
  XOR2X1   g03595(.A(new_n6031_), .B(pi0458), .Y(new_n6032_));
  XOR2X1   g03596(.A(new_n6032_), .B(new_n6026_), .Y(new_n6033_));
  AND2X1   g03597(.A(new_n6033_), .B(pi1196), .Y(new_n6034_));
  NOR3X1   g03598(.A(new_n6034_), .B(new_n6023_), .C(new_n6018_), .Y(new_n6035_));
  INVX1    g03599(.A(new_n6034_), .Y(new_n6036_));
  OAI21X1  g03600(.A0(new_n6005_), .A1(new_n6036_), .B0(pi1198), .Y(new_n6037_));
  INVX1    g03601(.A(pi0458), .Y(new_n6038_));
  INVX1    g03602(.A(pi0355), .Y(new_n6039_));
  MX2X1    g03603(.A(new_n6005_), .B(new_n5993_), .S0(pi0455), .Y(new_n6040_));
  INVX1    g03604(.A(pi0455), .Y(new_n6041_));
  MX2X1    g03605(.A(new_n6005_), .B(new_n5993_), .S0(new_n6041_), .Y(new_n6042_));
  MX2X1    g03606(.A(new_n6042_), .B(new_n6040_), .S0(new_n6024_), .Y(new_n6043_));
  MX2X1    g03607(.A(new_n6042_), .B(new_n6040_), .S0(pi0452), .Y(new_n6044_));
  MX2X1    g03608(.A(new_n6044_), .B(new_n6043_), .S0(new_n6039_), .Y(new_n6045_));
  NOR2X1   g03609(.A(new_n6045_), .B(new_n6038_), .Y(new_n6046_));
  MX2X1    g03610(.A(new_n6044_), .B(new_n6043_), .S0(pi0355), .Y(new_n6047_));
  OAI21X1  g03611(.A0(new_n6047_), .A1(pi0458), .B0(new_n6031_), .Y(new_n6048_));
  NOR2X1   g03612(.A(new_n6048_), .B(new_n6046_), .Y(new_n6049_));
  NOR2X1   g03613(.A(new_n6047_), .B(new_n6038_), .Y(new_n6050_));
  INVX1    g03614(.A(new_n6031_), .Y(new_n6051_));
  OAI21X1  g03615(.A0(new_n6045_), .A1(pi0458), .B0(new_n6051_), .Y(new_n6052_));
  OAI21X1  g03616(.A0(new_n6052_), .A1(new_n6050_), .B0(pi1196), .Y(new_n6053_));
  NOR2X1   g03617(.A(new_n6053_), .B(new_n6049_), .Y(new_n6054_));
  INVX1    g03618(.A(pi1198), .Y(new_n6055_));
  OAI21X1  g03619(.A0(new_n5993_), .A1(pi1196), .B0(new_n6055_), .Y(new_n6056_));
  OAI22X1  g03620(.A0(new_n6056_), .A1(new_n6054_), .B0(new_n6037_), .B1(new_n6035_), .Y(new_n6057_));
  MX2X1    g03621(.A(new_n6057_), .B(new_n6005_), .S0(new_n5892_), .Y(new_n6058_));
  INVX1    g03622(.A(pi0351), .Y(new_n6059_));
  AND2X1   g03623(.A(pi1199), .B(new_n6059_), .Y(new_n6060_));
  INVX1    g03624(.A(pi1199), .Y(new_n6061_));
  OR2X1    g03625(.A(new_n6005_), .B(new_n6061_), .Y(new_n6062_));
  OAI22X1  g03626(.A0(new_n6062_), .A1(pi0351), .B0(new_n6060_), .B1(new_n6058_), .Y(new_n6063_));
  AND2X1   g03627(.A(pi1199), .B(pi0351), .Y(new_n6064_));
  OAI22X1  g03628(.A0(new_n6064_), .A1(new_n6058_), .B0(new_n6062_), .B1(new_n6059_), .Y(new_n6065_));
  MX2X1    g03629(.A(new_n6065_), .B(new_n6063_), .S0(new_n5879_), .Y(new_n6066_));
  MX2X1    g03630(.A(new_n6065_), .B(new_n6063_), .S0(pi0461), .Y(new_n6067_));
  MX2X1    g03631(.A(new_n6067_), .B(new_n6066_), .S0(new_n5878_), .Y(new_n6068_));
  MX2X1    g03632(.A(new_n6067_), .B(new_n6066_), .S0(pi0357), .Y(new_n6069_));
  MX2X1    g03633(.A(new_n6069_), .B(new_n6068_), .S0(new_n5877_), .Y(new_n6070_));
  NAND2X1  g03634(.A(new_n6070_), .B(new_n5876_), .Y(new_n6071_));
  MX2X1    g03635(.A(new_n6069_), .B(new_n6068_), .S0(pi0356), .Y(new_n6072_));
  AOI21X1  g03636(.A0(new_n6072_), .A1(new_n5875_), .B0(pi0591), .Y(new_n6073_));
  INVX1    g03637(.A(pi0591), .Y(new_n6074_));
  OAI21X1  g03638(.A0(new_n6006_), .A1(new_n6074_), .B0(pi0590), .Y(new_n6075_));
  AOI21X1  g03639(.A0(new_n6073_), .A1(new_n6071_), .B0(new_n6075_), .Y(new_n6076_));
  NOR4X1   g03640(.A(pi0289), .B(pi0288), .C(pi0286), .D(pi0285), .Y(new_n6077_));
  INVX1    g03641(.A(pi0375), .Y(new_n6078_));
  INVX1    g03642(.A(pi0373), .Y(new_n6079_));
  INVX1    g03643(.A(pi0371), .Y(new_n6080_));
  INVX1    g03644(.A(pi0370), .Y(new_n6081_));
  INVX1    g03645(.A(pi0369), .Y(new_n6082_));
  XOR2X1   g03646(.A(pi0372), .B(pi0363), .Y(new_n6083_));
  XOR2X1   g03647(.A(new_n6083_), .B(pi0386), .Y(new_n6084_));
  XOR2X1   g03648(.A(pi0388), .B(pi0338), .Y(new_n6085_));
  XOR2X1   g03649(.A(pi0339), .B(pi0337), .Y(new_n6086_));
  XOR2X1   g03650(.A(new_n6086_), .B(pi0387), .Y(new_n6087_));
  XOR2X1   g03651(.A(new_n6087_), .B(pi0380), .Y(new_n6088_));
  XOR2X1   g03652(.A(new_n6088_), .B(new_n6085_), .Y(new_n6089_));
  XOR2X1   g03653(.A(new_n6089_), .B(new_n6084_), .Y(new_n6090_));
  AND2X1   g03654(.A(new_n6090_), .B(pi1196), .Y(new_n6091_));
  INVX1    g03655(.A(new_n6091_), .Y(new_n6092_));
  XOR2X1   g03656(.A(pi0389), .B(pi0368), .Y(new_n6093_));
  INVX1    g03657(.A(new_n6093_), .Y(new_n6094_));
  INVX1    g03658(.A(pi0367), .Y(new_n6095_));
  XOR2X1   g03659(.A(pi0447), .B(pi0365), .Y(new_n6096_));
  INVX1    g03660(.A(new_n6096_), .Y(new_n6097_));
  XOR2X1   g03661(.A(pi0383), .B(pi0336), .Y(new_n6098_));
  XOR2X1   g03662(.A(pi0366), .B(pi0364), .Y(new_n6099_));
  XOR2X1   g03663(.A(new_n6099_), .B(new_n6098_), .Y(new_n6100_));
  XOR2X1   g03664(.A(new_n6100_), .B(new_n6097_), .Y(new_n6101_));
  XOR2X1   g03665(.A(new_n6101_), .B(new_n6095_), .Y(new_n6102_));
  INVX1    g03666(.A(new_n6102_), .Y(new_n6103_));
  AOI21X1  g03667(.A0(new_n6103_), .A1(new_n6094_), .B0(new_n5889_), .Y(new_n6104_));
  OAI21X1  g03668(.A0(new_n6103_), .A1(new_n6094_), .B0(new_n6104_), .Y(new_n6105_));
  AND2X1   g03669(.A(new_n6105_), .B(new_n6092_), .Y(new_n6106_));
  AND2X1   g03670(.A(pi0592), .B(pi0377), .Y(new_n6107_));
  INVX1    g03671(.A(new_n6107_), .Y(new_n6108_));
  OAI21X1  g03672(.A0(new_n5992_), .A1(new_n5927_), .B0(new_n6108_), .Y(new_n6109_));
  XOR2X1   g03673(.A(pi0382), .B(pi0379), .Y(new_n6110_));
  XOR2X1   g03674(.A(pi0439), .B(pi0376), .Y(new_n6111_));
  XOR2X1   g03675(.A(new_n6111_), .B(pi0381), .Y(new_n6112_));
  INVX1    g03676(.A(pi0378), .Y(new_n6113_));
  XOR2X1   g03677(.A(pi0385), .B(pi0317), .Y(new_n6114_));
  XOR2X1   g03678(.A(new_n6114_), .B(new_n6113_), .Y(new_n6115_));
  XOR2X1   g03679(.A(new_n6115_), .B(new_n6112_), .Y(new_n6116_));
  XOR2X1   g03680(.A(new_n6116_), .B(new_n6110_), .Y(new_n6117_));
  INVX1    g03681(.A(new_n6117_), .Y(new_n6118_));
  AOI21X1  g03682(.A0(new_n6107_), .A1(new_n6003_), .B0(new_n6118_), .Y(new_n6119_));
  INVX1    g03683(.A(pi0592), .Y(new_n6120_));
  OAI22X1  g03684(.A0(new_n5992_), .A1(new_n5927_), .B0(new_n6120_), .B1(pi0377), .Y(new_n6121_));
  INVX1    g03685(.A(pi0377), .Y(new_n6122_));
  AND2X1   g03686(.A(pi0592), .B(new_n6122_), .Y(new_n6123_));
  AOI21X1  g03687(.A0(new_n6123_), .A1(new_n6003_), .B0(new_n6117_), .Y(new_n6124_));
  AOI22X1  g03688(.A0(new_n6124_), .A1(new_n6121_), .B0(new_n6119_), .B1(new_n6109_), .Y(new_n6125_));
  MX2X1    g03689(.A(new_n6003_), .B(new_n6006_), .S0(new_n6120_), .Y(new_n6126_));
  MX2X1    g03690(.A(new_n6126_), .B(new_n6125_), .S0(new_n6106_), .Y(new_n6127_));
  NAND2X1  g03691(.A(new_n6127_), .B(pi1199), .Y(new_n6128_));
  INVX1    g03692(.A(new_n6105_), .Y(new_n6129_));
  MX2X1    g03693(.A(new_n6006_), .B(new_n6126_), .S0(new_n6129_), .Y(new_n6130_));
  OR2X1    g03694(.A(new_n6130_), .B(new_n6090_), .Y(new_n6131_));
  INVX1    g03695(.A(pi1196), .Y(new_n6132_));
  AOI21X1  g03696(.A0(new_n6105_), .A1(new_n6132_), .B0(new_n6126_), .Y(new_n6133_));
  NOR4X1   g03697(.A(new_n6129_), .B(new_n5992_), .C(new_n5927_), .D(pi1196), .Y(new_n6134_));
  OAI21X1  g03698(.A0(new_n6134_), .A1(new_n6133_), .B0(new_n6090_), .Y(new_n6135_));
  NAND3X1  g03699(.A(new_n6135_), .B(new_n6131_), .C(new_n6061_), .Y(new_n6136_));
  AOI21X1  g03700(.A0(new_n6136_), .A1(new_n6128_), .B0(pi0374), .Y(new_n6137_));
  AND2X1   g03701(.A(pi1199), .B(new_n6055_), .Y(new_n6138_));
  AOI22X1  g03702(.A0(new_n6138_), .A1(new_n6127_), .B0(new_n6126_), .B1(pi1198), .Y(new_n6139_));
  OAI21X1  g03703(.A0(new_n6136_), .A1(pi1198), .B0(new_n6139_), .Y(new_n6140_));
  AOI21X1  g03704(.A0(new_n6140_), .A1(pi0374), .B0(new_n6137_), .Y(new_n6141_));
  OR2X1    g03705(.A(new_n6141_), .B(new_n6082_), .Y(new_n6142_));
  INVX1    g03706(.A(pi0374), .Y(new_n6143_));
  AOI21X1  g03707(.A0(new_n6136_), .A1(new_n6128_), .B0(new_n6143_), .Y(new_n6144_));
  AOI21X1  g03708(.A0(new_n6140_), .A1(new_n6143_), .B0(new_n6144_), .Y(new_n6145_));
  OAI21X1  g03709(.A0(new_n6145_), .A1(pi0369), .B0(new_n6142_), .Y(new_n6146_));
  AND2X1   g03710(.A(new_n6146_), .B(new_n6081_), .Y(new_n6147_));
  OR2X1    g03711(.A(new_n6141_), .B(pi0369), .Y(new_n6148_));
  OAI21X1  g03712(.A0(new_n6145_), .A1(new_n6082_), .B0(new_n6148_), .Y(new_n6149_));
  AOI21X1  g03713(.A0(new_n6149_), .A1(pi0370), .B0(new_n6147_), .Y(new_n6150_));
  OR2X1    g03714(.A(new_n6150_), .B(pi0371), .Y(new_n6151_));
  AND2X1   g03715(.A(new_n6149_), .B(new_n6081_), .Y(new_n6152_));
  AOI21X1  g03716(.A0(new_n6146_), .A1(pi0370), .B0(new_n6152_), .Y(new_n6153_));
  OAI21X1  g03717(.A0(new_n6153_), .A1(new_n6080_), .B0(new_n6151_), .Y(new_n6154_));
  AND2X1   g03718(.A(new_n6154_), .B(new_n6079_), .Y(new_n6155_));
  OR2X1    g03719(.A(new_n6153_), .B(pi0371), .Y(new_n6156_));
  OAI21X1  g03720(.A0(new_n6150_), .A1(new_n6080_), .B0(new_n6156_), .Y(new_n6157_));
  AOI21X1  g03721(.A0(new_n6157_), .A1(pi0373), .B0(new_n6155_), .Y(new_n6158_));
  XOR2X1   g03722(.A(pi0442), .B(pi0384), .Y(new_n6159_));
  XOR2X1   g03723(.A(new_n6159_), .B(pi0440), .Y(new_n6160_));
  MX2X1    g03724(.A(new_n6157_), .B(new_n6154_), .S0(pi0373), .Y(new_n6161_));
  OAI21X1  g03725(.A0(new_n6161_), .A1(new_n6078_), .B0(new_n6160_), .Y(new_n6162_));
  AOI21X1  g03726(.A0(new_n6158_), .A1(new_n6078_), .B0(new_n6162_), .Y(new_n6163_));
  INVX1    g03727(.A(new_n6160_), .Y(new_n6164_));
  OAI21X1  g03728(.A0(new_n6161_), .A1(pi0375), .B0(new_n6164_), .Y(new_n6165_));
  AOI21X1  g03729(.A0(new_n6158_), .A1(pi0375), .B0(new_n6165_), .Y(new_n6166_));
  NOR3X1   g03730(.A(new_n6166_), .B(new_n6163_), .C(pi0591), .Y(new_n6167_));
  INVX1    g03731(.A(pi0590), .Y(new_n6168_));
  INVX1    g03732(.A(pi0334), .Y(new_n6169_));
  INVX1    g03733(.A(pi0393), .Y(new_n6170_));
  INVX1    g03734(.A(pi0392), .Y(new_n6171_));
  INVX1    g03735(.A(pi0333), .Y(new_n6172_));
  INVX1    g03736(.A(pi0328), .Y(new_n6173_));
  XOR2X1   g03737(.A(pi0408), .B(new_n6173_), .Y(new_n6174_));
  XOR2X1   g03738(.A(pi0396), .B(pi0394), .Y(new_n6175_));
  XOR2X1   g03739(.A(new_n6175_), .B(new_n6174_), .Y(new_n6176_));
  INVX1    g03740(.A(pi0400), .Y(new_n6177_));
  XOR2X1   g03741(.A(pi0399), .B(pi0398), .Y(new_n6178_));
  XOR2X1   g03742(.A(new_n6178_), .B(pi0395), .Y(new_n6179_));
  XOR2X1   g03743(.A(new_n6179_), .B(pi0329), .Y(new_n6180_));
  XOR2X1   g03744(.A(new_n6180_), .B(new_n6177_), .Y(new_n6181_));
  XOR2X1   g03745(.A(new_n6181_), .B(new_n6176_), .Y(new_n6182_));
  AND2X1   g03746(.A(new_n6182_), .B(pi1198), .Y(new_n6183_));
  XOR2X1   g03747(.A(pi0410), .B(pi0390), .Y(new_n6184_));
  INVX1    g03748(.A(new_n6184_), .Y(new_n6185_));
  XOR2X1   g03749(.A(pi0412), .B(pi0397), .Y(new_n6186_));
  XOR2X1   g03750(.A(new_n6186_), .B(pi0404), .Y(new_n6187_));
  XOR2X1   g03751(.A(pi0324), .B(pi0319), .Y(new_n6188_));
  XOR2X1   g03752(.A(new_n6188_), .B(pi0456), .Y(new_n6189_));
  XOR2X1   g03753(.A(new_n6189_), .B(new_n6187_), .Y(new_n6190_));
  XOR2X1   g03754(.A(new_n6190_), .B(new_n6185_), .Y(new_n6191_));
  XOR2X1   g03755(.A(new_n6191_), .B(pi0411), .Y(new_n6192_));
  AOI21X1  g03756(.A0(new_n6192_), .A1(new_n5969_), .B0(new_n5967_), .Y(new_n6193_));
  NOR3X1   g03757(.A(new_n6193_), .B(new_n5978_), .C(pi0087), .Y(new_n6194_));
  AOI21X1  g03758(.A0(new_n6192_), .A1(new_n5981_), .B0(new_n5983_), .Y(new_n6195_));
  NOR3X1   g03759(.A(new_n6195_), .B(new_n5999_), .C(new_n5987_), .Y(new_n6196_));
  OR4X1    g03760(.A(new_n6196_), .B(new_n6132_), .C(pi0592), .D(pi0075), .Y(new_n6197_));
  OAI22X1  g03761(.A0(new_n6197_), .A1(new_n6194_), .B0(new_n5991_), .B1(pi1196), .Y(new_n6198_));
  AND2X1   g03762(.A(new_n6198_), .B(new_n6061_), .Y(new_n6199_));
  INVX1    g03763(.A(new_n6199_), .Y(new_n6200_));
  AND2X1   g03764(.A(new_n5955_), .B(pi1091), .Y(new_n6201_));
  XOR2X1   g03765(.A(pi0409), .B(pi0318), .Y(new_n6202_));
  INVX1    g03766(.A(pi0406), .Y(new_n6203_));
  XOR2X1   g03767(.A(pi0402), .B(pi0401), .Y(new_n6204_));
  XOR2X1   g03768(.A(new_n6204_), .B(new_n6203_), .Y(new_n6205_));
  XOR2X1   g03769(.A(pi0405), .B(pi0403), .Y(new_n6206_));
  XOR2X1   g03770(.A(pi0326), .B(pi0325), .Y(new_n6207_));
  XOR2X1   g03771(.A(new_n6207_), .B(new_n6206_), .Y(new_n6208_));
  XOR2X1   g03772(.A(new_n6208_), .B(new_n6205_), .Y(new_n6209_));
  XOR2X1   g03773(.A(new_n6209_), .B(new_n6202_), .Y(new_n6210_));
  INVX1    g03774(.A(new_n6210_), .Y(new_n6211_));
  NOR3X1   g03775(.A(new_n6192_), .B(new_n6132_), .C(pi0075), .Y(new_n6212_));
  NOR4X1   g03776(.A(new_n6212_), .B(new_n6211_), .C(new_n5968_), .D(new_n6201_), .Y(new_n6213_));
  OAI21X1  g03777(.A0(new_n6213_), .A1(new_n5967_), .B0(new_n5995_), .Y(new_n6214_));
  NOR2X1   g03778(.A(pi0592), .B(pi0075), .Y(new_n6215_));
  INVX1    g03779(.A(new_n6215_), .Y(new_n6216_));
  AOI21X1  g03780(.A0(new_n6210_), .A1(new_n5981_), .B0(new_n5983_), .Y(new_n6217_));
  NOR4X1   g03781(.A(new_n6217_), .B(new_n5999_), .C(new_n5987_), .D(pi1196), .Y(new_n6218_));
  NOR4X1   g03782(.A(new_n6217_), .B(new_n6195_), .C(new_n5999_), .D(new_n5987_), .Y(new_n6219_));
  NOR4X1   g03783(.A(new_n6219_), .B(new_n6218_), .C(new_n6216_), .D(new_n6061_), .Y(new_n6220_));
  AOI21X1  g03784(.A0(new_n5991_), .A1(new_n5936_), .B0(new_n6215_), .Y(new_n6221_));
  AOI21X1  g03785(.A0(new_n6220_), .A1(new_n6214_), .B0(new_n6221_), .Y(new_n6222_));
  AOI21X1  g03786(.A0(new_n6222_), .A1(new_n6200_), .B0(new_n5928_), .Y(new_n6223_));
  NOR3X1   g03787(.A(new_n6223_), .B(new_n6183_), .C(new_n5927_), .Y(new_n6224_));
  AOI21X1  g03788(.A0(new_n6183_), .A1(new_n6005_), .B0(new_n6224_), .Y(new_n6225_));
  INVX1    g03789(.A(new_n6225_), .Y(new_n6226_));
  MX2X1    g03790(.A(new_n6226_), .B(new_n6005_), .S0(pi1197), .Y(new_n6227_));
  MX2X1    g03791(.A(new_n6227_), .B(new_n6226_), .S0(new_n6172_), .Y(new_n6228_));
  MX2X1    g03792(.A(new_n6227_), .B(new_n6226_), .S0(pi0333), .Y(new_n6229_));
  MX2X1    g03793(.A(new_n6229_), .B(new_n6228_), .S0(pi0391), .Y(new_n6230_));
  INVX1    g03794(.A(pi0391), .Y(new_n6231_));
  MX2X1    g03795(.A(new_n6229_), .B(new_n6228_), .S0(new_n6231_), .Y(new_n6232_));
  MX2X1    g03796(.A(new_n6232_), .B(new_n6230_), .S0(new_n6171_), .Y(new_n6233_));
  MX2X1    g03797(.A(new_n6232_), .B(new_n6230_), .S0(pi0392), .Y(new_n6234_));
  MX2X1    g03798(.A(new_n6234_), .B(new_n6233_), .S0(new_n6170_), .Y(new_n6235_));
  XOR2X1   g03799(.A(pi0463), .B(pi0407), .Y(new_n6236_));
  INVX1    g03800(.A(pi0335), .Y(new_n6237_));
  XOR2X1   g03801(.A(pi0413), .B(new_n6237_), .Y(new_n6238_));
  XOR2X1   g03802(.A(new_n6238_), .B(new_n6236_), .Y(new_n6239_));
  INVX1    g03803(.A(new_n6239_), .Y(new_n6240_));
  OR2X1    g03804(.A(new_n6234_), .B(pi0393), .Y(new_n6241_));
  OAI21X1  g03805(.A0(new_n6233_), .A1(new_n6170_), .B0(new_n6241_), .Y(new_n6242_));
  OAI21X1  g03806(.A0(new_n6242_), .A1(new_n6169_), .B0(new_n6240_), .Y(new_n6243_));
  AOI21X1  g03807(.A0(new_n6235_), .A1(new_n6169_), .B0(new_n6243_), .Y(new_n6244_));
  NOR2X1   g03808(.A(new_n6242_), .B(pi0334), .Y(new_n6245_));
  AND2X1   g03809(.A(new_n6235_), .B(pi0334), .Y(new_n6246_));
  OR2X1    g03810(.A(new_n6246_), .B(new_n6240_), .Y(new_n6247_));
  OAI21X1  g03811(.A0(new_n6247_), .A1(new_n6245_), .B0(pi0591), .Y(new_n6248_));
  OAI21X1  g03812(.A0(new_n6248_), .A1(new_n6244_), .B0(new_n6168_), .Y(new_n6249_));
  OAI21X1  g03813(.A0(new_n6249_), .A1(new_n6167_), .B0(new_n6077_), .Y(new_n6250_));
  INVX1    g03814(.A(new_n6060_), .Y(new_n6251_));
  INVX1    g03815(.A(new_n5931_), .Y(new_n6252_));
  AOI21X1  g03816(.A0(new_n5973_), .A1(new_n5932_), .B0(new_n2722_), .Y(new_n6253_));
  NOR2X1   g03817(.A(new_n6253_), .B(new_n6252_), .Y(new_n6254_));
  INVX1    g03818(.A(new_n6254_), .Y(new_n6255_));
  AND2X1   g03819(.A(pi1093), .B(new_n5952_), .Y(new_n6256_));
  NOR4X1   g03820(.A(new_n2755_), .B(new_n5096_), .C(new_n5251_), .D(pi0098), .Y(new_n6257_));
  AOI21X1  g03821(.A0(new_n6257_), .A1(new_n6256_), .B0(pi1091), .Y(new_n6258_));
  INVX1    g03822(.A(new_n6256_), .Y(new_n6259_));
  NOR4X1   g03823(.A(new_n6259_), .B(new_n5939_), .C(pi1091), .D(pi0098), .Y(new_n6260_));
  AOI21X1  g03824(.A0(new_n6260_), .A1(new_n6252_), .B0(new_n3095_), .Y(new_n6261_));
  OAI21X1  g03825(.A0(new_n6258_), .A1(new_n6255_), .B0(new_n6261_), .Y(new_n6262_));
  AOI21X1  g03826(.A0(new_n6201_), .A1(new_n5921_), .B0(pi0039), .Y(new_n6263_));
  NOR2X1   g03827(.A(new_n5920_), .B(pi1091), .Y(new_n6264_));
  AND2X1   g03828(.A(new_n6257_), .B(new_n5952_), .Y(new_n6265_));
  AOI21X1  g03829(.A0(new_n5940_), .A1(pi0122), .B0(new_n6265_), .Y(new_n6266_));
  OAI21X1  g03830(.A0(new_n6266_), .A1(new_n2756_), .B0(new_n6264_), .Y(new_n6267_));
  AND2X1   g03831(.A(new_n6267_), .B(new_n6263_), .Y(new_n6268_));
  NOR2X1   g03832(.A(new_n5033_), .B(new_n5031_), .Y(new_n6269_));
  INVX1    g03833(.A(new_n6269_), .Y(new_n6270_));
  INVX1    g03834(.A(new_n6260_), .Y(new_n6271_));
  AOI21X1  g03835(.A0(new_n5958_), .A1(new_n2739_), .B0(new_n2722_), .Y(new_n6272_));
  OR2X1    g03836(.A(new_n6272_), .B(new_n6258_), .Y(new_n6273_));
  MX2X1    g03837(.A(new_n6273_), .B(new_n6271_), .S0(new_n6270_), .Y(new_n6274_));
  NAND2X1  g03838(.A(new_n6274_), .B(new_n5050_), .Y(new_n6275_));
  MX2X1    g03839(.A(new_n6273_), .B(new_n6271_), .S0(new_n5052_), .Y(new_n6276_));
  NOR3X1   g03840(.A(pi0224), .B(pi0223), .C(new_n2960_), .Y(new_n6277_));
  INVX1    g03841(.A(new_n6277_), .Y(new_n6278_));
  AOI21X1  g03842(.A0(new_n6276_), .A1(new_n5051_), .B0(new_n6278_), .Y(new_n6279_));
  OAI21X1  g03843(.A0(new_n6277_), .A1(new_n6271_), .B0(new_n2953_), .Y(new_n6280_));
  AOI21X1  g03844(.A0(new_n6279_), .A1(new_n6275_), .B0(new_n6280_), .Y(new_n6281_));
  NAND2X1  g03845(.A(new_n6274_), .B(new_n5070_), .Y(new_n6282_));
  NOR3X1   g03846(.A(new_n2437_), .B(pi0216), .C(pi0215), .Y(new_n6283_));
  INVX1    g03847(.A(new_n6283_), .Y(new_n6284_));
  AOI21X1  g03848(.A0(new_n6276_), .A1(new_n5071_), .B0(new_n6284_), .Y(new_n6285_));
  OAI21X1  g03849(.A0(new_n6283_), .A1(new_n6271_), .B0(pi0299), .Y(new_n6286_));
  AOI21X1  g03850(.A0(new_n6285_), .A1(new_n6282_), .B0(new_n6286_), .Y(new_n6287_));
  NOR3X1   g03851(.A(new_n6287_), .B(new_n6281_), .C(new_n2959_), .Y(new_n6288_));
  OAI21X1  g03852(.A0(new_n6288_), .A1(new_n6268_), .B0(new_n2996_), .Y(new_n6289_));
  AOI21X1  g03853(.A0(new_n6260_), .A1(pi0038), .B0(pi0100), .Y(new_n6290_));
  AOI21X1  g03854(.A0(new_n5930_), .A1(new_n5929_), .B0(new_n3013_), .Y(new_n6291_));
  OR4X1    g03855(.A(new_n5974_), .B(new_n3003_), .C(new_n2709_), .D(pi0070), .Y(new_n6292_));
  AND2X1   g03856(.A(new_n6257_), .B(new_n6256_), .Y(new_n6293_));
  INVX1    g03857(.A(new_n6293_), .Y(new_n6294_));
  MX2X1    g03858(.A(new_n6294_), .B(new_n6292_), .S0(pi1091), .Y(new_n6295_));
  OAI21X1  g03859(.A0(new_n6291_), .A1(new_n6260_), .B0(new_n3065_), .Y(new_n6296_));
  AOI21X1  g03860(.A0(new_n6295_), .A1(new_n6291_), .B0(new_n6296_), .Y(new_n6297_));
  OAI21X1  g03861(.A0(new_n6271_), .A1(new_n3065_), .B0(pi0100), .Y(new_n6298_));
  OAI21X1  g03862(.A0(new_n6298_), .A1(new_n6297_), .B0(new_n3156_), .Y(new_n6299_));
  AOI21X1  g03863(.A0(new_n6290_), .A1(new_n6289_), .B0(new_n6299_), .Y(new_n6300_));
  NOR4X1   g03864(.A(new_n5939_), .B(new_n3003_), .C(new_n2555_), .D(new_n5952_), .Y(new_n6301_));
  OAI21X1  g03865(.A0(new_n6301_), .A1(new_n6265_), .B0(pi1093), .Y(new_n6302_));
  NAND2X1  g03866(.A(new_n6302_), .B(new_n5998_), .Y(new_n6303_));
  NOR2X1   g03867(.A(new_n5997_), .B(new_n3157_), .Y(new_n6304_));
  AOI21X1  g03868(.A0(new_n6304_), .A1(new_n6303_), .B0(new_n6260_), .Y(new_n6305_));
  OAI21X1  g03869(.A0(new_n6305_), .A1(new_n3156_), .B0(new_n3095_), .Y(new_n6306_));
  OAI21X1  g03870(.A0(new_n6306_), .A1(new_n6300_), .B0(new_n6262_), .Y(new_n6307_));
  AOI21X1  g03871(.A0(new_n6307_), .A1(pi0567), .B0(new_n5927_), .Y(new_n6308_));
  INVX1    g03872(.A(new_n5893_), .Y(new_n6309_));
  AND2X1   g03873(.A(new_n6260_), .B(pi0567), .Y(new_n6310_));
  AND2X1   g03874(.A(new_n6310_), .B(new_n6309_), .Y(new_n6311_));
  NOR3X1   g03875(.A(new_n6311_), .B(new_n6308_), .C(new_n6120_), .Y(new_n6312_));
  AOI21X1  g03876(.A0(new_n6003_), .A1(new_n6120_), .B0(new_n6312_), .Y(new_n6313_));
  NOR2X1   g03877(.A(new_n6311_), .B(new_n6308_), .Y(new_n6314_));
  INVX1    g03878(.A(new_n6313_), .Y(new_n6315_));
  MX2X1    g03879(.A(new_n6315_), .B(new_n6314_), .S0(new_n6041_), .Y(new_n6316_));
  NAND2X1  g03880(.A(new_n6316_), .B(new_n6024_), .Y(new_n6317_));
  XOR2X1   g03881(.A(new_n6032_), .B(pi0355), .Y(new_n6318_));
  MX2X1    g03882(.A(new_n6315_), .B(new_n6314_), .S0(pi0455), .Y(new_n6319_));
  NAND2X1  g03883(.A(new_n6319_), .B(pi0452), .Y(new_n6320_));
  NAND3X1  g03884(.A(new_n6320_), .B(new_n6318_), .C(new_n6317_), .Y(new_n6321_));
  NAND2X1  g03885(.A(new_n6319_), .B(new_n6024_), .Y(new_n6322_));
  AOI21X1  g03886(.A0(new_n6316_), .A1(pi0452), .B0(new_n6318_), .Y(new_n6323_));
  AOI21X1  g03887(.A0(new_n6323_), .A1(new_n6322_), .B0(new_n6132_), .Y(new_n6324_));
  NOR3X1   g03888(.A(new_n6311_), .B(new_n6308_), .C(pi1196), .Y(new_n6325_));
  OR2X1    g03889(.A(new_n6325_), .B(pi1198), .Y(new_n6326_));
  AOI21X1  g03890(.A0(new_n6324_), .A1(new_n6321_), .B0(new_n6326_), .Y(new_n6327_));
  AOI21X1  g03891(.A0(new_n6314_), .A1(new_n6020_), .B0(new_n6022_), .Y(new_n6328_));
  AOI21X1  g03892(.A0(new_n6314_), .A1(new_n6007_), .B0(new_n6017_), .Y(new_n6329_));
  NOR3X1   g03893(.A(new_n6329_), .B(new_n6328_), .C(new_n6034_), .Y(new_n6330_));
  OAI21X1  g03894(.A0(new_n6313_), .A1(new_n6036_), .B0(pi1198), .Y(new_n6331_));
  OAI21X1  g03895(.A0(new_n6331_), .A1(new_n6330_), .B0(new_n5891_), .Y(new_n6332_));
  OAI22X1  g03896(.A0(new_n6332_), .A1(new_n6327_), .B0(new_n6313_), .B1(new_n5891_), .Y(new_n6333_));
  NOR3X1   g03897(.A(new_n6313_), .B(new_n6061_), .C(pi0351), .Y(new_n6334_));
  AOI21X1  g03898(.A0(new_n6333_), .A1(new_n6251_), .B0(new_n6334_), .Y(new_n6335_));
  INVX1    g03899(.A(new_n6064_), .Y(new_n6336_));
  NOR3X1   g03900(.A(new_n6313_), .B(new_n6061_), .C(new_n6059_), .Y(new_n6337_));
  AOI21X1  g03901(.A0(new_n6333_), .A1(new_n6336_), .B0(new_n6337_), .Y(new_n6338_));
  MX2X1    g03902(.A(new_n6338_), .B(new_n6335_), .S0(new_n5879_), .Y(new_n6339_));
  MX2X1    g03903(.A(new_n6338_), .B(new_n6335_), .S0(pi0461), .Y(new_n6340_));
  MX2X1    g03904(.A(new_n6340_), .B(new_n6339_), .S0(new_n5878_), .Y(new_n6341_));
  MX2X1    g03905(.A(new_n6340_), .B(new_n6339_), .S0(pi0357), .Y(new_n6342_));
  MX2X1    g03906(.A(new_n6342_), .B(new_n6341_), .S0(new_n5877_), .Y(new_n6343_));
  NOR2X1   g03907(.A(new_n6343_), .B(new_n5875_), .Y(new_n6344_));
  MX2X1    g03908(.A(new_n6342_), .B(new_n6341_), .S0(pi0356), .Y(new_n6345_));
  OAI21X1  g03909(.A0(new_n6345_), .A1(new_n5876_), .B0(new_n6074_), .Y(new_n6346_));
  INVX1    g03910(.A(new_n6314_), .Y(new_n6347_));
  AOI21X1  g03911(.A0(new_n6347_), .A1(pi0591), .B0(new_n6168_), .Y(new_n6348_));
  OAI21X1  g03912(.A0(new_n6346_), .A1(new_n6344_), .B0(new_n6348_), .Y(new_n6349_));
  XOR2X1   g03913(.A(new_n6160_), .B(pi0375), .Y(new_n6350_));
  XOR2X1   g03914(.A(new_n6350_), .B(new_n6079_), .Y(new_n6351_));
  INVX1    g03915(.A(new_n6106_), .Y(new_n6352_));
  AND2X1   g03916(.A(new_n6003_), .B(pi0592), .Y(new_n6353_));
  AOI21X1  g03917(.A0(new_n6314_), .A1(new_n6120_), .B0(new_n6353_), .Y(new_n6354_));
  AND2X1   g03918(.A(new_n6354_), .B(new_n6352_), .Y(new_n6355_));
  INVX1    g03919(.A(new_n6355_), .Y(new_n6356_));
  AOI21X1  g03920(.A0(new_n6347_), .A1(new_n6106_), .B0(pi1199), .Y(new_n6357_));
  OAI21X1  g03921(.A0(new_n6347_), .A1(new_n6123_), .B0(new_n6124_), .Y(new_n6358_));
  OAI21X1  g03922(.A0(new_n6347_), .A1(new_n6107_), .B0(new_n6119_), .Y(new_n6359_));
  AOI21X1  g03923(.A0(new_n6359_), .A1(new_n6358_), .B0(new_n6352_), .Y(new_n6360_));
  NOR3X1   g03924(.A(new_n6360_), .B(new_n6355_), .C(new_n6061_), .Y(new_n6361_));
  AOI21X1  g03925(.A0(new_n6357_), .A1(new_n6356_), .B0(new_n6361_), .Y(new_n6362_));
  MX2X1    g03926(.A(new_n6362_), .B(new_n6354_), .S0(pi1198), .Y(new_n6363_));
  MX2X1    g03927(.A(new_n6363_), .B(new_n6362_), .S0(new_n6143_), .Y(new_n6364_));
  MX2X1    g03928(.A(new_n6363_), .B(new_n6362_), .S0(pi0374), .Y(new_n6365_));
  MX2X1    g03929(.A(new_n6365_), .B(new_n6364_), .S0(pi0369), .Y(new_n6366_));
  MX2X1    g03930(.A(new_n6365_), .B(new_n6364_), .S0(new_n6082_), .Y(new_n6367_));
  MX2X1    g03931(.A(new_n6367_), .B(new_n6366_), .S0(new_n6081_), .Y(new_n6368_));
  MX2X1    g03932(.A(new_n6367_), .B(new_n6366_), .S0(pi0370), .Y(new_n6369_));
  MX2X1    g03933(.A(new_n6369_), .B(new_n6368_), .S0(new_n6080_), .Y(new_n6370_));
  OR2X1    g03934(.A(new_n6369_), .B(pi0371), .Y(new_n6371_));
  OAI21X1  g03935(.A0(new_n6368_), .A1(new_n6080_), .B0(new_n6371_), .Y(new_n6372_));
  AOI21X1  g03936(.A0(new_n6372_), .A1(new_n6351_), .B0(pi0591), .Y(new_n6373_));
  OAI21X1  g03937(.A0(new_n6370_), .A1(new_n6351_), .B0(new_n6373_), .Y(new_n6374_));
  XOR2X1   g03938(.A(new_n6239_), .B(pi0334), .Y(new_n6375_));
  XOR2X1   g03939(.A(new_n6375_), .B(pi0393), .Y(new_n6376_));
  AND2X1   g03940(.A(pi1196), .B(new_n6120_), .Y(new_n6377_));
  INVX1    g03941(.A(new_n6377_), .Y(new_n6378_));
  INVX1    g03942(.A(new_n6192_), .Y(new_n6379_));
  NOR3X1   g03943(.A(new_n6294_), .B(new_n6379_), .C(pi1091), .Y(new_n6380_));
  INVX1    g03944(.A(new_n6380_), .Y(new_n6381_));
  NOR3X1   g03945(.A(new_n6381_), .B(new_n5893_), .C(new_n5928_), .Y(new_n6382_));
  AND2X1   g03946(.A(new_n6257_), .B(new_n6210_), .Y(new_n6383_));
  AOI21X1  g03947(.A0(new_n6383_), .A1(new_n6382_), .B0(new_n6378_), .Y(new_n6384_));
  INVX1    g03948(.A(new_n6384_), .Y(new_n6385_));
  AOI21X1  g03949(.A0(new_n6380_), .A1(new_n6284_), .B0(new_n2953_), .Y(new_n6386_));
  NOR3X1   g03950(.A(new_n6294_), .B(new_n6211_), .C(pi1091), .Y(new_n6387_));
  AOI21X1  g03951(.A0(new_n6387_), .A1(new_n6284_), .B0(new_n2953_), .Y(new_n6388_));
  OR2X1    g03952(.A(new_n6388_), .B(new_n6386_), .Y(new_n6389_));
  NOR4X1   g03953(.A(new_n6294_), .B(new_n6211_), .C(new_n6379_), .D(pi1091), .Y(new_n6390_));
  NOR4X1   g03954(.A(new_n5959_), .B(new_n6270_), .C(new_n2740_), .D(new_n2722_), .Y(new_n6391_));
  NOR3X1   g03955(.A(new_n6391_), .B(new_n6390_), .C(new_n5071_), .Y(new_n6392_));
  NOR4X1   g03956(.A(new_n5959_), .B(new_n5052_), .C(new_n2740_), .D(new_n2722_), .Y(new_n6393_));
  NOR3X1   g03957(.A(new_n6393_), .B(new_n6390_), .C(new_n5070_), .Y(new_n6394_));
  OR4X1    g03958(.A(new_n6394_), .B(new_n6392_), .C(new_n5242_), .D(pi0216), .Y(new_n6395_));
  AND2X1   g03959(.A(new_n6395_), .B(new_n6389_), .Y(new_n6396_));
  AOI21X1  g03960(.A0(new_n6380_), .A1(new_n6278_), .B0(pi0299), .Y(new_n6397_));
  AOI21X1  g03961(.A0(new_n6387_), .A1(new_n6278_), .B0(pi0299), .Y(new_n6398_));
  OR2X1    g03962(.A(new_n6398_), .B(new_n6397_), .Y(new_n6399_));
  AND2X1   g03963(.A(new_n2961_), .B(pi0222), .Y(new_n6400_));
  INVX1    g03964(.A(new_n6400_), .Y(new_n6401_));
  NOR3X1   g03965(.A(new_n6391_), .B(new_n6390_), .C(new_n5051_), .Y(new_n6402_));
  NOR3X1   g03966(.A(new_n6393_), .B(new_n6390_), .C(new_n5050_), .Y(new_n6403_));
  OR4X1    g03967(.A(new_n6403_), .B(new_n6402_), .C(new_n6401_), .D(pi0223), .Y(new_n6404_));
  AND2X1   g03968(.A(new_n6404_), .B(new_n6399_), .Y(new_n6405_));
  NOR3X1   g03969(.A(new_n6405_), .B(new_n6396_), .C(new_n2959_), .Y(new_n6406_));
  NAND2X1  g03970(.A(new_n6379_), .B(new_n6264_), .Y(new_n6407_));
  NAND3X1  g03971(.A(new_n6407_), .B(new_n6267_), .C(new_n6263_), .Y(new_n6408_));
  INVX1    g03972(.A(new_n6408_), .Y(new_n6409_));
  AOI21X1  g03973(.A0(new_n6210_), .A1(new_n5940_), .B0(new_n5952_), .Y(new_n6410_));
  OAI21X1  g03974(.A0(new_n6383_), .A1(pi0122), .B0(pi1093), .Y(new_n6411_));
  OAI21X1  g03975(.A0(new_n6411_), .A1(new_n6410_), .B0(new_n6264_), .Y(new_n6412_));
  AOI21X1  g03976(.A0(new_n6412_), .A1(new_n6409_), .B0(new_n6406_), .Y(new_n6413_));
  AOI21X1  g03977(.A0(new_n6380_), .A1(pi0038), .B0(pi0100), .Y(new_n6414_));
  AOI21X1  g03978(.A0(new_n6387_), .A1(pi0038), .B0(pi0100), .Y(new_n6415_));
  OAI22X1  g03979(.A0(new_n6415_), .A1(new_n6414_), .B0(new_n6413_), .B1(pi0038), .Y(new_n6416_));
  NOR2X1   g03980(.A(new_n2980_), .B(pi0299), .Y(new_n6417_));
  AND2X1   g03981(.A(new_n6292_), .B(pi1091), .Y(new_n6418_));
  NOR2X1   g03982(.A(new_n2451_), .B(new_n2953_), .Y(new_n6419_));
  INVX1    g03983(.A(new_n6419_), .Y(new_n6420_));
  AOI21X1  g03984(.A0(new_n6420_), .A1(new_n5033_), .B0(new_n6417_), .Y(new_n6421_));
  INVX1    g03985(.A(new_n6421_), .Y(new_n6422_));
  NOR2X1   g03986(.A(new_n6390_), .B(pi1091), .Y(new_n6423_));
  NOR3X1   g03987(.A(new_n6423_), .B(new_n6422_), .C(new_n6418_), .Y(new_n6424_));
  AOI21X1  g03988(.A0(new_n5975_), .A1(new_n6417_), .B0(new_n6424_), .Y(new_n6425_));
  NOR2X1   g03989(.A(new_n6425_), .B(new_n3013_), .Y(new_n6426_));
  INVX1    g03990(.A(new_n6390_), .Y(new_n6427_));
  AND2X1   g03991(.A(new_n6421_), .B(pi0228), .Y(new_n6428_));
  OAI21X1  g03992(.A0(new_n6428_), .A1(new_n6427_), .B0(pi0232), .Y(new_n6429_));
  NOR2X1   g03993(.A(new_n6390_), .B(pi0232), .Y(new_n6430_));
  OAI21X1  g03994(.A0(new_n5976_), .A1(new_n3013_), .B0(new_n6430_), .Y(new_n6431_));
  AND2X1   g03995(.A(new_n6431_), .B(new_n3065_), .Y(new_n6432_));
  OAI21X1  g03996(.A0(new_n6429_), .A1(new_n6426_), .B0(new_n6432_), .Y(new_n6433_));
  AOI21X1  g03997(.A0(new_n6390_), .A1(new_n3066_), .B0(new_n3026_), .Y(new_n6434_));
  AND2X1   g03998(.A(new_n6434_), .B(new_n6433_), .Y(new_n6435_));
  INVX1    g03999(.A(new_n6435_), .Y(new_n6436_));
  AND2X1   g04000(.A(new_n6436_), .B(new_n6416_), .Y(new_n6437_));
  AOI21X1  g04001(.A0(new_n6380_), .A1(new_n3157_), .B0(new_n3156_), .Y(new_n6438_));
  AOI21X1  g04002(.A0(new_n6387_), .A1(new_n3157_), .B0(new_n3156_), .Y(new_n6439_));
  NOR3X1   g04003(.A(new_n6192_), .B(new_n5923_), .C(pi1091), .Y(new_n6440_));
  INVX1    g04004(.A(new_n5998_), .Y(new_n6441_));
  AND2X1   g04005(.A(new_n6304_), .B(new_n6303_), .Y(new_n6442_));
  OAI21X1  g04006(.A0(new_n6210_), .A1(new_n6441_), .B0(new_n6442_), .Y(new_n6443_));
  OAI22X1  g04007(.A0(new_n6443_), .A1(new_n6440_), .B0(new_n6439_), .B1(new_n6438_), .Y(new_n6444_));
  OAI21X1  g04008(.A0(new_n6437_), .A1(pi0087), .B0(new_n6444_), .Y(new_n6445_));
  AOI21X1  g04009(.A0(new_n6380_), .A1(new_n6252_), .B0(new_n3095_), .Y(new_n6446_));
  AOI21X1  g04010(.A0(new_n6387_), .A1(new_n6252_), .B0(new_n3095_), .Y(new_n6447_));
  OAI22X1  g04011(.A0(new_n6447_), .A1(new_n6446_), .B0(new_n6423_), .B1(new_n6255_), .Y(new_n6448_));
  INVX1    g04012(.A(new_n6448_), .Y(new_n6449_));
  AOI21X1  g04013(.A0(new_n6445_), .A1(new_n3095_), .B0(new_n6449_), .Y(new_n6450_));
  NOR2X1   g04014(.A(new_n6450_), .B(new_n6385_), .Y(new_n6451_));
  NOR4X1   g04015(.A(new_n6294_), .B(new_n6211_), .C(pi1091), .D(new_n5928_), .Y(new_n6452_));
  NOR2X1   g04016(.A(pi1196), .B(pi0592), .Y(new_n6453_));
  INVX1    g04017(.A(new_n6453_), .Y(new_n6454_));
  AOI21X1  g04018(.A0(new_n6452_), .A1(new_n6309_), .B0(new_n6454_), .Y(new_n6455_));
  INVX1    g04019(.A(new_n6455_), .Y(new_n6456_));
  AND2X1   g04020(.A(new_n6443_), .B(new_n6439_), .Y(new_n6457_));
  NOR3X1   g04021(.A(new_n6387_), .B(new_n5977_), .C(new_n3026_), .Y(new_n6458_));
  INVX1    g04022(.A(new_n6458_), .Y(new_n6459_));
  INVX1    g04023(.A(new_n6388_), .Y(new_n6460_));
  NOR3X1   g04024(.A(new_n6393_), .B(new_n6387_), .C(new_n5070_), .Y(new_n6461_));
  INVX1    g04025(.A(new_n6461_), .Y(new_n6462_));
  OR4X1    g04026(.A(new_n6391_), .B(new_n6387_), .C(new_n5069_), .D(new_n5065_), .Y(new_n6463_));
  AND2X1   g04027(.A(new_n6463_), .B(new_n6283_), .Y(new_n6464_));
  AOI21X1  g04028(.A0(new_n6464_), .A1(new_n6462_), .B0(new_n6460_), .Y(new_n6465_));
  INVX1    g04029(.A(new_n6398_), .Y(new_n6466_));
  NOR3X1   g04030(.A(new_n6393_), .B(new_n6387_), .C(new_n5050_), .Y(new_n6467_));
  NOR3X1   g04031(.A(new_n6391_), .B(new_n6387_), .C(new_n5051_), .Y(new_n6468_));
  NOR3X1   g04032(.A(new_n6468_), .B(new_n6467_), .C(new_n6278_), .Y(new_n6469_));
  NOR2X1   g04033(.A(new_n6469_), .B(new_n6466_), .Y(new_n6470_));
  NOR3X1   g04034(.A(new_n6470_), .B(new_n6465_), .C(new_n2959_), .Y(new_n6471_));
  AOI21X1  g04035(.A0(new_n6412_), .A1(new_n6263_), .B0(new_n6471_), .Y(new_n6472_));
  OAI21X1  g04036(.A0(new_n6472_), .A1(pi0038), .B0(new_n6415_), .Y(new_n6473_));
  AOI21X1  g04037(.A0(new_n6473_), .A1(new_n6459_), .B0(pi0087), .Y(new_n6474_));
  OAI21X1  g04038(.A0(new_n6474_), .A1(new_n6457_), .B0(new_n3095_), .Y(new_n6475_));
  AOI21X1  g04039(.A0(new_n6293_), .A1(new_n6210_), .B0(pi1091), .Y(new_n6476_));
  OAI21X1  g04040(.A0(new_n6476_), .A1(new_n6255_), .B0(new_n6447_), .Y(new_n6477_));
  AOI21X1  g04041(.A0(new_n6477_), .A1(new_n6475_), .B0(new_n6456_), .Y(new_n6478_));
  OAI21X1  g04042(.A0(new_n6478_), .A1(new_n6451_), .B0(pi0567), .Y(new_n6479_));
  OR2X1    g04043(.A(new_n6455_), .B(new_n6384_), .Y(new_n6480_));
  AOI21X1  g04044(.A0(new_n6480_), .A1(new_n5927_), .B0(new_n6061_), .Y(new_n6481_));
  AND2X1   g04045(.A(new_n6481_), .B(new_n6479_), .Y(new_n6482_));
  INVX1    g04046(.A(new_n6414_), .Y(new_n6483_));
  NOR3X1   g04047(.A(new_n6393_), .B(new_n6380_), .C(new_n5070_), .Y(new_n6484_));
  OR2X1    g04048(.A(new_n6391_), .B(new_n6380_), .Y(new_n6485_));
  OAI21X1  g04049(.A0(new_n6485_), .A1(new_n5071_), .B0(new_n6283_), .Y(new_n6486_));
  OAI21X1  g04050(.A0(new_n6486_), .A1(new_n6484_), .B0(new_n6386_), .Y(new_n6487_));
  NOR3X1   g04051(.A(new_n6393_), .B(new_n6380_), .C(new_n5050_), .Y(new_n6488_));
  OAI21X1  g04052(.A0(new_n6485_), .A1(new_n5051_), .B0(new_n6277_), .Y(new_n6489_));
  OAI21X1  g04053(.A0(new_n6489_), .A1(new_n6488_), .B0(new_n6397_), .Y(new_n6490_));
  NAND3X1  g04054(.A(new_n6490_), .B(new_n6487_), .C(pi0039), .Y(new_n6491_));
  AOI21X1  g04055(.A0(new_n6491_), .A1(new_n6408_), .B0(pi0038), .Y(new_n6492_));
  OAI22X1  g04056(.A0(new_n6492_), .A1(new_n6483_), .B0(new_n6380_), .B1(new_n5979_), .Y(new_n6493_));
  OAI21X1  g04057(.A0(new_n6192_), .A1(new_n6441_), .B0(new_n6442_), .Y(new_n6494_));
  AOI22X1  g04058(.A0(new_n6494_), .A1(new_n6438_), .B0(new_n6493_), .B1(new_n3156_), .Y(new_n6495_));
  AOI21X1  g04059(.A0(new_n6293_), .A1(new_n6192_), .B0(pi1091), .Y(new_n6496_));
  OAI21X1  g04060(.A0(new_n6496_), .A1(new_n6255_), .B0(new_n6446_), .Y(new_n6497_));
  OAI21X1  g04061(.A0(new_n6495_), .A1(pi0075), .B0(new_n6497_), .Y(new_n6498_));
  AOI21X1  g04062(.A0(new_n6498_), .A1(pi0567), .B0(new_n5927_), .Y(new_n6499_));
  NOR3X1   g04063(.A(new_n6499_), .B(new_n6382_), .C(new_n6378_), .Y(new_n6500_));
  NOR3X1   g04064(.A(new_n6500_), .B(new_n6325_), .C(pi1199), .Y(new_n6501_));
  NOR3X1   g04065(.A(new_n6501_), .B(new_n6482_), .C(new_n6183_), .Y(new_n6502_));
  AND2X1   g04066(.A(new_n6003_), .B(new_n6120_), .Y(new_n6503_));
  AND2X1   g04067(.A(new_n6183_), .B(new_n6503_), .Y(new_n6504_));
  NOR3X1   g04068(.A(new_n6504_), .B(new_n6502_), .C(new_n6312_), .Y(new_n6505_));
  MX2X1    g04069(.A(new_n6505_), .B(new_n6313_), .S0(pi1197), .Y(new_n6506_));
  MX2X1    g04070(.A(new_n6506_), .B(new_n6505_), .S0(pi0333), .Y(new_n6507_));
  MX2X1    g04071(.A(new_n6506_), .B(new_n6505_), .S0(new_n6172_), .Y(new_n6508_));
  MX2X1    g04072(.A(new_n6508_), .B(new_n6507_), .S0(new_n6231_), .Y(new_n6509_));
  MX2X1    g04073(.A(new_n6508_), .B(new_n6507_), .S0(pi0391), .Y(new_n6510_));
  MX2X1    g04074(.A(new_n6510_), .B(new_n6509_), .S0(new_n6171_), .Y(new_n6511_));
  OR2X1    g04075(.A(new_n6511_), .B(new_n6376_), .Y(new_n6512_));
  OR2X1    g04076(.A(new_n6510_), .B(pi0392), .Y(new_n6513_));
  OAI21X1  g04077(.A0(new_n6509_), .A1(new_n6171_), .B0(new_n6513_), .Y(new_n6514_));
  AOI21X1  g04078(.A0(new_n6514_), .A1(new_n6376_), .B0(new_n6074_), .Y(new_n6515_));
  AOI21X1  g04079(.A0(new_n6515_), .A1(new_n6512_), .B0(pi0590), .Y(new_n6516_));
  AOI21X1  g04080(.A0(new_n6516_), .A1(new_n6374_), .B0(new_n6077_), .Y(new_n6517_));
  AOI21X1  g04081(.A0(new_n6517_), .A1(new_n6349_), .B0(pi0588), .Y(new_n6518_));
  OAI21X1  g04082(.A0(new_n6250_), .A1(new_n6076_), .B0(new_n6518_), .Y(new_n6519_));
  AND2X1   g04083(.A(new_n5117_), .B(new_n2436_), .Y(new_n6520_));
  INVX1    g04084(.A(new_n6520_), .Y(po1038));
  INVX1    g04085(.A(pi0448), .Y(new_n6522_));
  INVX1    g04086(.A(pi0449), .Y(new_n6523_));
  XOR2X1   g04087(.A(pi0451), .B(pi0433), .Y(new_n6524_));
  XOR2X1   g04088(.A(new_n6524_), .B(new_n6523_), .Y(new_n6525_));
  XOR2X1   g04089(.A(new_n6525_), .B(new_n6522_), .Y(new_n6526_));
  INVX1    g04090(.A(pi0427), .Y(new_n6527_));
  INVX1    g04091(.A(pi0428), .Y(new_n6528_));
  INVX1    g04092(.A(new_n6005_), .Y(new_n6529_));
  XOR2X1   g04093(.A(pi0418), .B(pi0417), .Y(new_n6530_));
  XOR2X1   g04094(.A(new_n6530_), .B(pi0437), .Y(new_n6531_));
  INVX1    g04095(.A(pi0453), .Y(new_n6532_));
  XOR2X1   g04096(.A(pi0464), .B(new_n6532_), .Y(new_n6533_));
  XOR2X1   g04097(.A(new_n6533_), .B(new_n6531_), .Y(new_n6534_));
  XOR2X1   g04098(.A(pi0431), .B(pi0415), .Y(new_n6535_));
  INVX1    g04099(.A(pi0416), .Y(new_n6536_));
  XOR2X1   g04100(.A(pi0438), .B(new_n6536_), .Y(new_n6537_));
  XOR2X1   g04101(.A(new_n6537_), .B(new_n6535_), .Y(new_n6538_));
  AND2X1   g04102(.A(new_n6538_), .B(new_n6534_), .Y(new_n6539_));
  OAI21X1  g04103(.A0(new_n6538_), .A1(new_n6534_), .B0(pi1197), .Y(new_n6540_));
  XOR2X1   g04104(.A(pi0454), .B(pi0421), .Y(new_n6541_));
  XOR2X1   g04105(.A(pi0459), .B(pi0432), .Y(new_n6542_));
  XOR2X1   g04106(.A(new_n6542_), .B(new_n6541_), .Y(new_n6543_));
  XOR2X1   g04107(.A(pi0420), .B(pi0419), .Y(new_n6544_));
  XOR2X1   g04108(.A(pi0424), .B(pi0423), .Y(new_n6545_));
  XOR2X1   g04109(.A(new_n6545_), .B(new_n6544_), .Y(new_n6546_));
  XOR2X1   g04110(.A(new_n6546_), .B(new_n6543_), .Y(new_n6547_));
  AND2X1   g04111(.A(new_n6547_), .B(pi0425), .Y(new_n6548_));
  OAI21X1  g04112(.A0(new_n6547_), .A1(pi0425), .B0(pi1198), .Y(new_n6549_));
  OAI22X1  g04113(.A0(new_n6549_), .A1(new_n6548_), .B0(new_n6540_), .B1(new_n6539_), .Y(new_n6550_));
  NAND2X1  g04114(.A(new_n6550_), .B(new_n6005_), .Y(new_n6551_));
  INVX1    g04115(.A(pi0444), .Y(new_n6552_));
  NOR2X1   g04116(.A(pi0592), .B(pi0443), .Y(new_n6553_));
  MX2X1    g04117(.A(new_n5993_), .B(new_n6004_), .S0(new_n6553_), .Y(new_n6554_));
  AND2X1   g04118(.A(new_n6120_), .B(pi0443), .Y(new_n6555_));
  MX2X1    g04119(.A(new_n5993_), .B(new_n6004_), .S0(new_n6555_), .Y(new_n6556_));
  MX2X1    g04120(.A(new_n6556_), .B(new_n6554_), .S0(new_n6552_), .Y(new_n6557_));
  NOR2X1   g04121(.A(new_n6557_), .B(pi0436), .Y(new_n6558_));
  INVX1    g04122(.A(pi0436), .Y(new_n6559_));
  XOR2X1   g04123(.A(pi0435), .B(pi0429), .Y(new_n6560_));
  XOR2X1   g04124(.A(pi0446), .B(pi0434), .Y(new_n6561_));
  INVX1    g04125(.A(pi0414), .Y(new_n6562_));
  XOR2X1   g04126(.A(pi0422), .B(new_n6562_), .Y(new_n6563_));
  XOR2X1   g04127(.A(new_n6563_), .B(new_n6561_), .Y(new_n6564_));
  INVX1    g04128(.A(new_n6564_), .Y(new_n6565_));
  XOR2X1   g04129(.A(new_n6565_), .B(new_n6560_), .Y(new_n6566_));
  MX2X1    g04130(.A(new_n6556_), .B(new_n6554_), .S0(pi0444), .Y(new_n6567_));
  OAI21X1  g04131(.A0(new_n6567_), .A1(new_n6559_), .B0(new_n6566_), .Y(new_n6568_));
  NOR2X1   g04132(.A(new_n6568_), .B(new_n6558_), .Y(new_n6569_));
  NOR2X1   g04133(.A(new_n6567_), .B(pi0436), .Y(new_n6570_));
  INVX1    g04134(.A(new_n6566_), .Y(new_n6571_));
  OAI21X1  g04135(.A0(new_n6557_), .A1(new_n6559_), .B0(new_n6571_), .Y(new_n6572_));
  OAI21X1  g04136(.A0(new_n6572_), .A1(new_n6570_), .B0(pi1196), .Y(new_n6573_));
  AOI21X1  g04137(.A0(new_n6006_), .A1(new_n6132_), .B0(new_n6550_), .Y(new_n6574_));
  OAI21X1  g04138(.A0(new_n6573_), .A1(new_n6569_), .B0(new_n6574_), .Y(new_n6575_));
  AND2X1   g04139(.A(new_n6575_), .B(new_n6551_), .Y(new_n6576_));
  MX2X1    g04140(.A(new_n6576_), .B(new_n6529_), .S0(new_n6528_), .Y(new_n6577_));
  MX2X1    g04141(.A(new_n6576_), .B(new_n6529_), .S0(pi0428), .Y(new_n6578_));
  MX2X1    g04142(.A(new_n6578_), .B(new_n6577_), .S0(new_n6527_), .Y(new_n6579_));
  MX2X1    g04143(.A(new_n6578_), .B(new_n6577_), .S0(pi0427), .Y(new_n6580_));
  MX2X1    g04144(.A(new_n6580_), .B(new_n6579_), .S0(pi0430), .Y(new_n6581_));
  INVX1    g04145(.A(pi0430), .Y(new_n6582_));
  MX2X1    g04146(.A(new_n6580_), .B(new_n6579_), .S0(new_n6582_), .Y(new_n6583_));
  MX2X1    g04147(.A(new_n6583_), .B(new_n6581_), .S0(pi0426), .Y(new_n6584_));
  INVX1    g04148(.A(pi0426), .Y(new_n6585_));
  MX2X1    g04149(.A(new_n6583_), .B(new_n6581_), .S0(new_n6585_), .Y(new_n6586_));
  MX2X1    g04150(.A(new_n6586_), .B(new_n6584_), .S0(pi0445), .Y(new_n6587_));
  OR2X1    g04151(.A(new_n6587_), .B(new_n6526_), .Y(new_n6588_));
  INVX1    g04152(.A(pi0445), .Y(new_n6589_));
  OR2X1    g04153(.A(new_n6586_), .B(new_n6589_), .Y(new_n6590_));
  OAI21X1  g04154(.A0(new_n6584_), .A1(pi0445), .B0(new_n6590_), .Y(new_n6591_));
  AOI21X1  g04155(.A0(new_n6591_), .A1(new_n6526_), .B0(new_n6061_), .Y(new_n6592_));
  NOR2X1   g04156(.A(pi0591), .B(pi0590), .Y(new_n6593_));
  NAND3X1  g04157(.A(new_n6575_), .B(new_n6551_), .C(new_n6061_), .Y(new_n6594_));
  NAND2X1  g04158(.A(new_n6594_), .B(new_n6593_), .Y(new_n6595_));
  AOI21X1  g04159(.A0(new_n6592_), .A1(new_n6588_), .B0(new_n6595_), .Y(new_n6596_));
  OAI21X1  g04160(.A0(new_n6593_), .A1(new_n6006_), .B0(new_n6077_), .Y(new_n6597_));
  XOR2X1   g04161(.A(pi0444), .B(new_n6559_), .Y(new_n6598_));
  XOR2X1   g04162(.A(new_n6598_), .B(new_n6571_), .Y(new_n6599_));
  INVX1    g04163(.A(new_n6599_), .Y(new_n6600_));
  AOI21X1  g04164(.A0(new_n6553_), .A1(new_n6003_), .B0(new_n6600_), .Y(new_n6601_));
  OAI21X1  g04165(.A0(new_n6553_), .A1(new_n6347_), .B0(new_n6601_), .Y(new_n6602_));
  NOR3X1   g04166(.A(new_n6555_), .B(new_n6311_), .C(new_n6308_), .Y(new_n6603_));
  INVX1    g04167(.A(new_n6603_), .Y(new_n6604_));
  AOI21X1  g04168(.A0(new_n6555_), .A1(new_n6003_), .B0(new_n6599_), .Y(new_n6605_));
  AOI21X1  g04169(.A0(new_n6605_), .A1(new_n6604_), .B0(new_n6132_), .Y(new_n6606_));
  AOI21X1  g04170(.A0(new_n6606_), .A1(new_n6602_), .B0(new_n6325_), .Y(new_n6607_));
  MX2X1    g04171(.A(new_n6607_), .B(new_n6313_), .S0(new_n6550_), .Y(new_n6608_));
  OAI21X1  g04172(.A0(new_n6315_), .A1(pi0428), .B0(pi0427), .Y(new_n6609_));
  AOI21X1  g04173(.A0(new_n6608_), .A1(pi0428), .B0(new_n6609_), .Y(new_n6610_));
  OAI21X1  g04174(.A0(new_n6315_), .A1(new_n6528_), .B0(new_n6527_), .Y(new_n6611_));
  AOI21X1  g04175(.A0(new_n6608_), .A1(new_n6528_), .B0(new_n6611_), .Y(new_n6612_));
  OR2X1    g04176(.A(new_n6612_), .B(new_n6610_), .Y(new_n6613_));
  INVX1    g04177(.A(new_n6608_), .Y(new_n6614_));
  XOR2X1   g04178(.A(pi0428), .B(new_n6527_), .Y(new_n6615_));
  MX2X1    g04179(.A(new_n6614_), .B(new_n6315_), .S0(new_n6615_), .Y(new_n6616_));
  MX2X1    g04180(.A(new_n6616_), .B(new_n6613_), .S0(new_n6582_), .Y(new_n6617_));
  MX2X1    g04181(.A(new_n6616_), .B(new_n6613_), .S0(pi0430), .Y(new_n6618_));
  MX2X1    g04182(.A(new_n6618_), .B(new_n6617_), .S0(new_n6585_), .Y(new_n6619_));
  AND2X1   g04183(.A(new_n6619_), .B(new_n6589_), .Y(new_n6620_));
  MX2X1    g04184(.A(new_n6618_), .B(new_n6617_), .S0(pi0426), .Y(new_n6621_));
  AOI21X1  g04185(.A0(new_n6621_), .A1(pi0445), .B0(new_n6620_), .Y(new_n6622_));
  INVX1    g04186(.A(new_n6525_), .Y(new_n6623_));
  MX2X1    g04187(.A(new_n6621_), .B(new_n6619_), .S0(pi0445), .Y(new_n6624_));
  OAI21X1  g04188(.A0(new_n6624_), .A1(pi0448), .B0(new_n6623_), .Y(new_n6625_));
  AOI21X1  g04189(.A0(new_n6622_), .A1(pi0448), .B0(new_n6625_), .Y(new_n6626_));
  OAI21X1  g04190(.A0(new_n6624_), .A1(new_n6522_), .B0(new_n6525_), .Y(new_n6627_));
  AOI21X1  g04191(.A0(new_n6622_), .A1(new_n6522_), .B0(new_n6627_), .Y(new_n6628_));
  OAI21X1  g04192(.A0(new_n6628_), .A1(new_n6626_), .B0(pi1199), .Y(new_n6629_));
  INVX1    g04193(.A(new_n6593_), .Y(new_n6630_));
  AOI21X1  g04194(.A0(new_n6614_), .A1(new_n6061_), .B0(new_n6630_), .Y(new_n6631_));
  AND2X1   g04195(.A(new_n6631_), .B(new_n6629_), .Y(new_n6632_));
  INVX1    g04196(.A(new_n6077_), .Y(new_n6633_));
  OAI21X1  g04197(.A0(new_n6593_), .A1(new_n6314_), .B0(new_n6633_), .Y(new_n6634_));
  OAI22X1  g04198(.A0(new_n6634_), .A1(new_n6632_), .B0(new_n6597_), .B1(new_n6596_), .Y(new_n6635_));
  AOI21X1  g04199(.A0(new_n6635_), .A1(pi0588), .B0(po1038), .Y(new_n6636_));
  INVX1    g04200(.A(pi0217), .Y(new_n6637_));
  INVX1    g04201(.A(new_n6310_), .Y(new_n6638_));
  AND2X1   g04202(.A(new_n6033_), .B(new_n6120_), .Y(new_n6639_));
  NOR3X1   g04203(.A(new_n6639_), .B(new_n6638_), .C(new_n6028_), .Y(new_n6640_));
  INVX1    g04204(.A(new_n6640_), .Y(new_n6641_));
  INVX1    g04205(.A(pi0441), .Y(new_n6642_));
  XOR2X1   g04206(.A(pi0458), .B(new_n6029_), .Y(new_n6643_));
  XOR2X1   g04207(.A(new_n6643_), .B(new_n6026_), .Y(new_n6644_));
  NAND2X1  g04208(.A(new_n6644_), .B(new_n6642_), .Y(new_n6645_));
  OR2X1    g04209(.A(new_n6644_), .B(new_n6642_), .Y(new_n6646_));
  NAND3X1  g04210(.A(new_n6646_), .B(new_n6645_), .C(new_n6120_), .Y(new_n6647_));
  AND2X1   g04211(.A(new_n6310_), .B(new_n6028_), .Y(new_n6648_));
  AOI21X1  g04212(.A0(new_n6648_), .A1(new_n6647_), .B0(new_n6132_), .Y(new_n6649_));
  AOI21X1  g04213(.A0(new_n6649_), .A1(new_n6641_), .B0(pi1198), .Y(new_n6650_));
  INVX1    g04214(.A(new_n6650_), .Y(new_n6651_));
  XOR2X1   g04215(.A(new_n6016_), .B(new_n6019_), .Y(new_n6652_));
  AND2X1   g04216(.A(new_n6652_), .B(new_n6036_), .Y(new_n6653_));
  NAND4X1  g04217(.A(new_n6653_), .B(new_n6310_), .C(pi1198), .D(new_n6120_), .Y(new_n6654_));
  AOI21X1  g04218(.A0(new_n6654_), .A1(new_n6651_), .B0(new_n5892_), .Y(new_n6655_));
  INVX1    g04219(.A(new_n6655_), .Y(new_n6656_));
  AOI21X1  g04220(.A0(new_n6656_), .A1(new_n6120_), .B0(new_n6638_), .Y(new_n6657_));
  INVX1    g04221(.A(new_n6657_), .Y(new_n6658_));
  AOI21X1  g04222(.A0(new_n6310_), .A1(pi0592), .B0(new_n6061_), .Y(new_n6659_));
  AOI22X1  g04223(.A0(new_n6659_), .A1(pi0351), .B0(new_n6658_), .B1(new_n6336_), .Y(new_n6660_));
  AOI22X1  g04224(.A0(new_n6659_), .A1(new_n6059_), .B0(new_n6658_), .B1(new_n6251_), .Y(new_n6661_));
  MX2X1    g04225(.A(new_n6661_), .B(new_n6660_), .S0(new_n5879_), .Y(new_n6662_));
  MX2X1    g04226(.A(new_n6661_), .B(new_n6660_), .S0(pi0461), .Y(new_n6663_));
  MX2X1    g04227(.A(new_n6663_), .B(new_n6662_), .S0(new_n5878_), .Y(new_n6664_));
  OR2X1    g04228(.A(new_n6664_), .B(pi0356), .Y(new_n6665_));
  MX2X1    g04229(.A(new_n6663_), .B(new_n6662_), .S0(pi0357), .Y(new_n6666_));
  OR2X1    g04230(.A(new_n6666_), .B(new_n5877_), .Y(new_n6667_));
  NAND3X1  g04231(.A(new_n6667_), .B(new_n6665_), .C(new_n5875_), .Y(new_n6668_));
  OR2X1    g04232(.A(new_n6666_), .B(pi0356), .Y(new_n6669_));
  OR2X1    g04233(.A(new_n6664_), .B(new_n5877_), .Y(new_n6670_));
  NAND3X1  g04234(.A(new_n6670_), .B(new_n6669_), .C(new_n5876_), .Y(new_n6671_));
  AND2X1   g04235(.A(new_n6671_), .B(new_n6668_), .Y(new_n6672_));
  NAND3X1  g04236(.A(new_n6260_), .B(new_n6120_), .C(pi0567), .Y(new_n6673_));
  AND2X1   g04237(.A(new_n6310_), .B(pi0592), .Y(new_n6674_));
  XOR2X1   g04238(.A(new_n6117_), .B(pi0377), .Y(new_n6675_));
  AND2X1   g04239(.A(new_n6675_), .B(new_n6106_), .Y(new_n6676_));
  OAI21X1  g04240(.A0(new_n6676_), .A1(new_n6120_), .B0(new_n6310_), .Y(new_n6677_));
  AOI22X1  g04241(.A0(new_n6677_), .A1(pi1199), .B0(new_n6352_), .B1(pi0592), .Y(new_n6678_));
  NAND3X1  g04242(.A(new_n6678_), .B(new_n6674_), .C(new_n6055_), .Y(new_n6679_));
  XOR2X1   g04243(.A(pi0374), .B(pi0369), .Y(new_n6680_));
  XOR2X1   g04244(.A(new_n6680_), .B(pi0370), .Y(new_n6681_));
  XOR2X1   g04245(.A(new_n6681_), .B(pi0371), .Y(new_n6682_));
  XOR2X1   g04246(.A(new_n6682_), .B(pi0373), .Y(new_n6683_));
  XOR2X1   g04247(.A(new_n6683_), .B(new_n6078_), .Y(new_n6684_));
  XOR2X1   g04248(.A(new_n6684_), .B(new_n6160_), .Y(new_n6685_));
  NAND3X1  g04249(.A(new_n6685_), .B(new_n6678_), .C(new_n6674_), .Y(new_n6686_));
  NAND3X1  g04250(.A(new_n6686_), .B(new_n6679_), .C(new_n6673_), .Y(new_n6687_));
  AOI21X1  g04251(.A0(new_n6687_), .A1(new_n6168_), .B0(pi0591), .Y(new_n6688_));
  OAI21X1  g04252(.A0(new_n6672_), .A1(new_n6168_), .B0(new_n6688_), .Y(new_n6689_));
  OR2X1    g04253(.A(new_n6674_), .B(new_n5889_), .Y(new_n6690_));
  INVX1    g04254(.A(new_n6452_), .Y(new_n6691_));
  OAI21X1  g04255(.A0(new_n6192_), .A1(new_n6132_), .B0(new_n6120_), .Y(new_n6692_));
  OAI21X1  g04256(.A0(new_n6692_), .A1(new_n6691_), .B0(new_n6659_), .Y(new_n6693_));
  NAND4X1  g04257(.A(new_n6293_), .B(new_n6192_), .C(new_n2722_), .D(pi0567), .Y(new_n6694_));
  AOI21X1  g04258(.A0(new_n6378_), .A1(new_n6310_), .B0(pi1199), .Y(new_n6695_));
  OAI21X1  g04259(.A0(new_n6694_), .A1(new_n6378_), .B0(new_n6695_), .Y(new_n6696_));
  AND2X1   g04260(.A(new_n6696_), .B(new_n6693_), .Y(new_n6697_));
  OAI21X1  g04261(.A0(new_n6697_), .A1(pi1197), .B0(new_n6690_), .Y(new_n6698_));
  AND2X1   g04262(.A(new_n6698_), .B(pi0333), .Y(new_n6699_));
  INVX1    g04263(.A(new_n6182_), .Y(new_n6700_));
  AOI21X1  g04264(.A0(new_n6310_), .A1(pi0592), .B0(new_n6055_), .Y(new_n6701_));
  INVX1    g04265(.A(new_n6701_), .Y(new_n6702_));
  AND2X1   g04266(.A(new_n6702_), .B(new_n6697_), .Y(new_n6703_));
  OAI22X1  g04267(.A0(new_n6703_), .A1(new_n6700_), .B0(new_n6697_), .B1(pi0333), .Y(new_n6704_));
  OR2X1    g04268(.A(new_n6704_), .B(new_n6699_), .Y(new_n6705_));
  AND2X1   g04269(.A(new_n6698_), .B(new_n6172_), .Y(new_n6706_));
  OAI21X1  g04270(.A0(new_n6702_), .A1(new_n6700_), .B0(new_n6697_), .Y(new_n6707_));
  OR2X1    g04271(.A(new_n6707_), .B(new_n6706_), .Y(new_n6708_));
  MX2X1    g04272(.A(new_n6708_), .B(new_n6705_), .S0(new_n6231_), .Y(new_n6709_));
  MX2X1    g04273(.A(new_n6708_), .B(new_n6705_), .S0(pi0391), .Y(new_n6710_));
  MX2X1    g04274(.A(new_n6710_), .B(new_n6709_), .S0(new_n6171_), .Y(new_n6711_));
  NAND2X1  g04275(.A(new_n6711_), .B(new_n6170_), .Y(new_n6712_));
  INVX1    g04276(.A(new_n6375_), .Y(new_n6713_));
  MX2X1    g04277(.A(new_n6710_), .B(new_n6709_), .S0(pi0392), .Y(new_n6714_));
  AOI21X1  g04278(.A0(new_n6714_), .A1(pi0393), .B0(new_n6713_), .Y(new_n6715_));
  NAND2X1  g04279(.A(new_n6714_), .B(new_n6170_), .Y(new_n6716_));
  AOI21X1  g04280(.A0(new_n6711_), .A1(pi0393), .B0(new_n6375_), .Y(new_n6717_));
  AOI22X1  g04281(.A0(new_n6717_), .A1(new_n6716_), .B0(new_n6715_), .B1(new_n6712_), .Y(new_n6718_));
  AOI21X1  g04282(.A0(new_n6310_), .A1(pi0590), .B0(new_n6074_), .Y(new_n6719_));
  OAI21X1  g04283(.A0(new_n6718_), .A1(pi0590), .B0(new_n6719_), .Y(new_n6720_));
  AOI21X1  g04284(.A0(new_n6720_), .A1(new_n6689_), .B0(pi0588), .Y(new_n6721_));
  AOI21X1  g04285(.A0(new_n5117_), .A1(new_n2436_), .B0(new_n6077_), .Y(new_n6722_));
  XOR2X1   g04286(.A(pi0443), .B(pi0436), .Y(new_n6723_));
  XOR2X1   g04287(.A(new_n6723_), .B(new_n6552_), .Y(new_n6724_));
  OAI21X1  g04288(.A0(new_n6724_), .A1(new_n6571_), .B0(new_n6377_), .Y(new_n6725_));
  AOI21X1  g04289(.A0(new_n6724_), .A1(new_n6571_), .B0(new_n6725_), .Y(new_n6726_));
  NOR3X1   g04290(.A(new_n6726_), .B(new_n6673_), .C(new_n6550_), .Y(new_n6727_));
  XOR2X1   g04291(.A(new_n6615_), .B(new_n6582_), .Y(new_n6728_));
  XOR2X1   g04292(.A(new_n6728_), .B(pi0426), .Y(new_n6729_));
  XOR2X1   g04293(.A(new_n6729_), .B(pi0445), .Y(new_n6730_));
  XOR2X1   g04294(.A(new_n6730_), .B(new_n6522_), .Y(new_n6731_));
  AOI21X1  g04295(.A0(new_n6731_), .A1(new_n6727_), .B0(new_n6674_), .Y(new_n6732_));
  OR2X1    g04296(.A(new_n6732_), .B(new_n6623_), .Y(new_n6733_));
  NOR4X1   g04297(.A(new_n6731_), .B(new_n6726_), .C(new_n6673_), .D(new_n6550_), .Y(new_n6734_));
  OAI21X1  g04298(.A0(new_n6734_), .A1(new_n6674_), .B0(new_n6623_), .Y(new_n6735_));
  AND2X1   g04299(.A(new_n6735_), .B(pi1199), .Y(new_n6736_));
  OR2X1    g04300(.A(new_n6674_), .B(pi1199), .Y(new_n6737_));
  OAI21X1  g04301(.A0(new_n6737_), .A1(new_n6727_), .B0(new_n6593_), .Y(new_n6738_));
  AOI21X1  g04302(.A0(new_n6736_), .A1(new_n6733_), .B0(new_n6738_), .Y(new_n6739_));
  OAI21X1  g04303(.A0(new_n6593_), .A1(new_n6638_), .B0(pi0588), .Y(new_n6740_));
  OAI21X1  g04304(.A0(new_n6740_), .A1(new_n6739_), .B0(new_n6722_), .Y(new_n6741_));
  OAI21X1  g04305(.A0(new_n6741_), .A1(new_n6721_), .B0(new_n6637_), .Y(new_n6742_));
  AOI21X1  g04306(.A0(new_n6636_), .A1(new_n6519_), .B0(new_n6742_), .Y(new_n6743_));
  OAI21X1  g04307(.A0(new_n6347_), .A1(new_n6077_), .B0(new_n6520_), .Y(new_n6744_));
  AOI21X1  g04308(.A0(new_n6077_), .A1(new_n6006_), .B0(new_n6744_), .Y(new_n6745_));
  INVX1    g04309(.A(new_n6722_), .Y(new_n6746_));
  OAI21X1  g04310(.A0(new_n6746_), .A1(new_n6638_), .B0(pi0217), .Y(new_n6747_));
  NOR3X1   g04311(.A(pi1163), .B(pi1162), .C(pi1161), .Y(new_n6748_));
  OAI21X1  g04312(.A0(new_n6747_), .A1(new_n6745_), .B0(new_n6748_), .Y(new_n6749_));
  INVX1    g04313(.A(pi0031), .Y(new_n6750_));
  INVX1    g04314(.A(pi1161), .Y(new_n6751_));
  NOR4X1   g04315(.A(pi1163), .B(new_n6751_), .C(new_n2756_), .D(new_n2755_), .Y(new_n6752_));
  NAND3X1  g04316(.A(new_n6752_), .B(pi1162), .C(new_n6750_), .Y(new_n6753_));
  OAI21X1  g04317(.A0(new_n6749_), .A1(new_n6743_), .B0(new_n6753_), .Y(po0189));
  OR2X1    g04318(.A(pi0074), .B(pi0055), .Y(new_n6755_));
  NOR4X1   g04319(.A(new_n6755_), .B(new_n5107_), .C(new_n3393_), .D(new_n5324_), .Y(new_n6756_));
  AND2X1   g04320(.A(new_n3065_), .B(pi0100), .Y(new_n6757_));
  INVX1    g04321(.A(new_n5094_), .Y(po1057));
  NOR4X1   g04322(.A(new_n5098_), .B(po1057), .C(new_n5083_), .D(new_n3074_), .Y(new_n6759_));
  NAND2X1  g04323(.A(new_n6759_), .B(new_n2453_), .Y(new_n6760_));
  NOR3X1   g04324(.A(new_n3003_), .B(new_n2555_), .C(new_n5095_), .Y(new_n6761_));
  INVX1    g04325(.A(new_n6761_), .Y(new_n6762_));
  NOR2X1   g04326(.A(new_n5970_), .B(new_n5094_), .Y(new_n6763_));
  OR4X1    g04327(.A(new_n6763_), .B(new_n5084_), .C(new_n3053_), .D(pi0137), .Y(new_n6764_));
  OAI21X1  g04328(.A0(new_n6764_), .A1(new_n6762_), .B0(new_n6760_), .Y(new_n6765_));
  INVX1    g04329(.A(new_n2476_), .Y(new_n6766_));
  NOR4X1   g04330(.A(new_n2579_), .B(new_n2577_), .C(pi0077), .D(new_n2580_), .Y(new_n6767_));
  NOR4X1   g04331(.A(new_n2511_), .B(new_n2477_), .C(pi0094), .D(pi0046), .Y(new_n6768_));
  AND2X1   g04332(.A(new_n6768_), .B(new_n2483_), .Y(new_n6769_));
  NAND4X1  g04333(.A(new_n6769_), .B(new_n6767_), .C(new_n6766_), .D(new_n2531_), .Y(new_n6770_));
  OR4X1    g04334(.A(new_n6770_), .B(new_n5020_), .C(pi0090), .D(pi0024), .Y(new_n6771_));
  NOR4X1   g04335(.A(pi1093), .B(new_n2755_), .C(new_n5096_), .D(new_n5258_), .Y(new_n6772_));
  AOI21X1  g04336(.A0(new_n2757_), .A1(new_n2723_), .B0(new_n6772_), .Y(new_n6773_));
  AOI21X1  g04337(.A0(new_n6773_), .A1(new_n6633_), .B0(pi0137), .Y(new_n6774_));
  INVX1    g04338(.A(pi0084), .Y(new_n6775_));
  NOR4X1   g04339(.A(pi0073), .B(pi0068), .C(pi0066), .D(pi0049), .Y(new_n6776_));
  NAND4X1  g04340(.A(new_n6776_), .B(new_n5142_), .C(new_n6775_), .D(pi0076), .Y(new_n6777_));
  OR4X1    g04341(.A(pi0102), .B(pi0089), .C(pi0077), .D(pi0050), .Y(new_n6778_));
  OR4X1    g04342(.A(new_n6778_), .B(new_n2472_), .C(pi0081), .D(pi0064), .Y(new_n6779_));
  OR4X1    g04343(.A(pi0098), .B(pi0088), .C(pi0067), .D(pi0036), .Y(new_n6780_));
  OR4X1    g04344(.A(new_n6780_), .B(pi0106), .C(pi0103), .D(pi0085), .Y(new_n6781_));
  OR4X1    g04345(.A(pi0083), .B(pi0071), .C(pi0069), .D(pi0065), .Y(new_n6782_));
  OR2X1    g04346(.A(pi0048), .B(pi0045), .Y(new_n6783_));
  OR4X1    g04347(.A(new_n6783_), .B(new_n6782_), .C(pi0104), .D(pi0061), .Y(new_n6784_));
  NOR4X1   g04348(.A(new_n6784_), .B(new_n6781_), .C(new_n6779_), .D(new_n6777_), .Y(new_n6785_));
  NOR2X1   g04349(.A(new_n2484_), .B(new_n2478_), .Y(new_n6786_));
  OAI21X1  g04350(.A0(new_n6785_), .A1(new_n6767_), .B0(new_n6786_), .Y(new_n6787_));
  AND2X1   g04351(.A(new_n6787_), .B(new_n5787_), .Y(new_n6788_));
  INVX1    g04352(.A(new_n6769_), .Y(new_n6789_));
  OR4X1    g04353(.A(new_n6784_), .B(new_n6781_), .C(new_n6779_), .D(new_n6777_), .Y(new_n6790_));
  NOR3X1   g04354(.A(new_n6790_), .B(new_n6789_), .C(new_n2476_), .Y(new_n6791_));
  NAND3X1  g04355(.A(new_n2767_), .B(new_n5134_), .C(new_n2516_), .Y(new_n6792_));
  OR4X1    g04356(.A(new_n6792_), .B(new_n2492_), .C(pi0137), .D(pi0035), .Y(new_n6793_));
  AOI21X1  g04357(.A0(new_n6773_), .A1(new_n6633_), .B0(new_n6793_), .Y(new_n6794_));
  OAI21X1  g04358(.A0(new_n6791_), .A1(new_n5787_), .B0(new_n6794_), .Y(new_n6795_));
  OAI22X1  g04359(.A0(new_n6795_), .A1(new_n6788_), .B0(new_n6774_), .B1(new_n6771_), .Y(new_n6796_));
  AOI21X1  g04360(.A0(new_n2726_), .A1(new_n5787_), .B0(new_n2456_), .Y(new_n6797_));
  AOI22X1  g04361(.A0(new_n6797_), .A1(new_n2488_), .B0(new_n6796_), .B1(new_n2456_), .Y(new_n6798_));
  AND2X1   g04362(.A(new_n6771_), .B(new_n2456_), .Y(new_n6799_));
  OAI21X1  g04363(.A0(new_n5021_), .A1(new_n2456_), .B0(new_n5019_), .Y(new_n6800_));
  OAI22X1  g04364(.A0(new_n6800_), .A1(new_n6799_), .B0(new_n6798_), .B1(new_n5019_), .Y(new_n6801_));
  NOR4X1   g04365(.A(pi0100), .B(pi0095), .C(pi0039), .D(pi0038), .Y(new_n6802_));
  AOI22X1  g04366(.A0(new_n6802_), .A1(new_n6801_), .B0(new_n6765_), .B1(new_n6757_), .Y(new_n6803_));
  INVX1    g04367(.A(new_n6773_), .Y(po0840));
  OR4X1    g04368(.A(new_n2542_), .B(new_n2513_), .C(new_n2520_), .D(pi0024), .Y(new_n6805_));
  NOR2X1   g04369(.A(new_n3256_), .B(new_n2725_), .Y(new_n6806_));
  INVX1    g04370(.A(new_n6806_), .Y(new_n6807_));
  OR4X1    g04371(.A(new_n6807_), .B(new_n6805_), .C(po0840), .D(pi0051), .Y(new_n6808_));
  NOR2X1   g04372(.A(new_n5094_), .B(new_n5083_), .Y(new_n6809_));
  NOR2X1   g04373(.A(new_n6763_), .B(new_n3053_), .Y(new_n6810_));
  NOR4X1   g04374(.A(new_n3066_), .B(pi0100), .C(pi0087), .D(new_n3095_), .Y(new_n6811_));
  INVX1    g04375(.A(new_n6811_), .Y(new_n6812_));
  OR4X1    g04376(.A(new_n6812_), .B(new_n6810_), .C(new_n6809_), .D(pi0137), .Y(new_n6813_));
  OAI22X1  g04377(.A0(new_n6813_), .A1(new_n6808_), .B0(new_n6803_), .B1(new_n3101_), .Y(new_n6814_));
  AND2X1   g04378(.A(new_n6814_), .B(new_n6756_), .Y(po0190));
  INVX1    g04379(.A(pi0079), .Y(new_n6816_));
  INVX1    g04380(.A(pi0118), .Y(new_n6817_));
  NOR4X1   g04381(.A(pi0196), .B(pi0195), .C(pi0139), .D(pi0138), .Y(new_n6818_));
  NAND3X1  g04382(.A(new_n6818_), .B(new_n6817_), .C(new_n6816_), .Y(new_n6819_));
  NOR2X1   g04383(.A(new_n6819_), .B(pi0034), .Y(new_n6820_));
  NOR2X1   g04384(.A(new_n6820_), .B(pi0033), .Y(new_n6821_));
  NOR2X1   g04385(.A(pi0157), .B(pi0149), .Y(new_n6822_));
  NOR3X1   g04386(.A(new_n6822_), .B(pi0468), .C(pi0332), .Y(new_n6823_));
  INVX1    g04387(.A(new_n6823_), .Y(new_n6824_));
  AOI21X1  g04388(.A0(pi0157), .A1(pi0149), .B0(new_n6824_), .Y(new_n6825_));
  INVX1    g04389(.A(new_n6825_), .Y(new_n6826_));
  OAI22X1  g04390(.A0(new_n6826_), .A1(new_n5237_), .B0(pi0100), .B1(pi0075), .Y(new_n6827_));
  NOR2X1   g04391(.A(pi0100), .B(pi0075), .Y(new_n6828_));
  NAND4X1  g04392(.A(new_n6828_), .B(new_n5033_), .C(pi0232), .D(pi0164), .Y(new_n6829_));
  AOI21X1  g04393(.A0(new_n6829_), .A1(new_n6827_), .B0(pi0074), .Y(new_n6830_));
  INVX1    g04394(.A(new_n6827_), .Y(new_n6831_));
  INVX1    g04395(.A(new_n6828_), .Y(new_n6832_));
  NOR4X1   g04396(.A(new_n6832_), .B(new_n5057_), .C(new_n5237_), .D(new_n4210_), .Y(new_n6833_));
  OAI21X1  g04397(.A0(new_n6833_), .A1(new_n6831_), .B0(pi0074), .Y(new_n6834_));
  NAND2X1  g04398(.A(new_n6834_), .B(new_n3393_), .Y(new_n6835_));
  NOR2X1   g04399(.A(new_n6835_), .B(new_n6830_), .Y(new_n6836_));
  OR2X1    g04400(.A(pi0183), .B(pi0178), .Y(new_n6837_));
  NAND2X1  g04401(.A(new_n6837_), .B(new_n5033_), .Y(new_n6838_));
  AOI21X1  g04402(.A0(pi0183), .A1(pi0178), .B0(new_n6838_), .Y(new_n6839_));
  OAI21X1  g04403(.A0(new_n6839_), .A1(pi0299), .B0(pi0232), .Y(new_n6840_));
  AOI21X1  g04404(.A0(new_n6826_), .A1(pi0299), .B0(new_n6840_), .Y(new_n6841_));
  NOR2X1   g04405(.A(new_n6841_), .B(new_n3026_), .Y(new_n6842_));
  NOR2X1   g04406(.A(new_n6841_), .B(new_n3095_), .Y(new_n6843_));
  INVX1    g04407(.A(pi0191), .Y(new_n6844_));
  MX2X1    g04408(.A(new_n6844_), .B(new_n4210_), .S0(pi0299), .Y(new_n6845_));
  NOR4X1   g04409(.A(new_n6845_), .B(new_n6832_), .C(new_n5057_), .D(new_n5237_), .Y(new_n6846_));
  NOR3X1   g04410(.A(new_n6846_), .B(new_n6843_), .C(new_n6842_), .Y(new_n6847_));
  OAI21X1  g04411(.A0(new_n6847_), .A1(new_n4991_), .B0(new_n3128_), .Y(new_n6848_));
  MX2X1    g04412(.A(pi0186), .B(pi0164), .S0(pi0299), .Y(new_n6849_));
  NAND3X1  g04413(.A(new_n6849_), .B(new_n5033_), .C(pi0232), .Y(new_n6850_));
  NOR2X1   g04414(.A(new_n6850_), .B(new_n6832_), .Y(new_n6851_));
  NOR3X1   g04415(.A(new_n6851_), .B(new_n6843_), .C(new_n6842_), .Y(new_n6852_));
  NOR2X1   g04416(.A(new_n6852_), .B(new_n3112_), .Y(new_n6853_));
  INVX1    g04417(.A(new_n6853_), .Y(new_n6854_));
  INVX1    g04418(.A(new_n5930_), .Y(new_n6855_));
  NOR3X1   g04419(.A(new_n6855_), .B(new_n4995_), .C(new_n2953_), .Y(new_n6856_));
  NOR3X1   g04420(.A(new_n3003_), .B(new_n2555_), .C(pi0039), .Y(new_n6857_));
  OAI21X1  g04421(.A0(new_n6855_), .A1(new_n6857_), .B0(pi0186), .Y(new_n6858_));
  AND2X1   g04422(.A(new_n6858_), .B(pi0164), .Y(new_n6859_));
  OAI21X1  g04423(.A0(new_n6856_), .A1(pi0186), .B0(new_n6859_), .Y(new_n6860_));
  INVX1    g04424(.A(pi0186), .Y(new_n6861_));
  NAND3X1  g04425(.A(new_n5033_), .B(new_n2953_), .C(pi0232), .Y(new_n6862_));
  NOR4X1   g04426(.A(new_n6862_), .B(new_n4995_), .C(new_n6861_), .D(pi0164), .Y(new_n6863_));
  INVX1    g04427(.A(new_n6863_), .Y(new_n6864_));
  AOI21X1  g04428(.A0(new_n6864_), .A1(new_n6860_), .B0(new_n2996_), .Y(new_n6865_));
  INVX1    g04429(.A(pi0176), .Y(new_n6866_));
  AND2X1   g04430(.A(pi0232), .B(new_n6866_), .Y(new_n6867_));
  INVX1    g04431(.A(new_n6867_), .Y(new_n6868_));
  NOR3X1   g04432(.A(pi0107), .B(pi0063), .C(pi0040), .Y(new_n6869_));
  INVX1    g04433(.A(new_n6869_), .Y(new_n6870_));
  NOR2X1   g04434(.A(pi0081), .B(pi0064), .Y(new_n6871_));
  NAND2X1  g04435(.A(new_n6871_), .B(new_n2578_), .Y(new_n6872_));
  OR4X1    g04436(.A(new_n6872_), .B(new_n2459_), .C(pi0071), .D(pi0065), .Y(new_n6873_));
  OR2X1    g04437(.A(new_n6873_), .B(new_n2471_), .Y(new_n6874_));
  NAND2X1  g04438(.A(new_n2505_), .B(new_n2497_), .Y(new_n6875_));
  OR4X1    g04439(.A(new_n6875_), .B(new_n6874_), .C(pi0060), .D(pi0053), .Y(new_n6876_));
  NOR3X1   g04440(.A(new_n6876_), .B(new_n5908_), .C(pi0058), .Y(new_n6877_));
  NAND3X1  g04441(.A(new_n6877_), .B(new_n2543_), .C(new_n2456_), .Y(new_n6878_));
  NOR2X1   g04442(.A(new_n6878_), .B(pi0095), .Y(new_n6879_));
  INVX1    g04443(.A(new_n6879_), .Y(new_n6880_));
  INVX1    g04444(.A(new_n5246_), .Y(new_n6881_));
  NOR4X1   g04445(.A(new_n5260_), .B(new_n6881_), .C(new_n5040_), .D(new_n2755_), .Y(new_n6882_));
  INVX1    g04446(.A(new_n6882_), .Y(new_n6883_));
  AOI21X1  g04447(.A0(new_n6883_), .A1(new_n5060_), .B0(new_n6880_), .Y(new_n6884_));
  AOI21X1  g04448(.A0(new_n6884_), .A1(new_n6269_), .B0(new_n6870_), .Y(new_n6885_));
  NOR3X1   g04449(.A(new_n2961_), .B(pi0223), .C(new_n2960_), .Y(new_n6886_));
  NOR2X1   g04450(.A(new_n6886_), .B(new_n6870_), .Y(new_n6887_));
  INVX1    g04451(.A(new_n6887_), .Y(new_n6888_));
  OR4X1    g04452(.A(new_n6883_), .B(new_n6878_), .C(new_n5057_), .D(pi0095), .Y(new_n6889_));
  AOI21X1  g04453(.A0(new_n6889_), .A1(new_n6869_), .B0(new_n5050_), .Y(new_n6890_));
  NAND3X1  g04454(.A(new_n6890_), .B(new_n6888_), .C(pi0174), .Y(new_n6891_));
  OAI21X1  g04455(.A0(new_n6887_), .A1(new_n6885_), .B0(new_n6891_), .Y(new_n6892_));
  NOR3X1   g04456(.A(new_n2437_), .B(new_n2438_), .C(pi0215), .Y(new_n6893_));
  OR2X1    g04457(.A(new_n6893_), .B(new_n6870_), .Y(new_n6894_));
  AND2X1   g04458(.A(new_n6894_), .B(pi0299), .Y(new_n6895_));
  INVX1    g04459(.A(new_n6885_), .Y(new_n6896_));
  INVX1    g04460(.A(new_n6884_), .Y(new_n6897_));
  OAI21X1  g04461(.A0(new_n6897_), .A1(new_n5057_), .B0(new_n6869_), .Y(new_n6898_));
  AOI21X1  g04462(.A0(new_n6898_), .A1(new_n5071_), .B0(new_n6896_), .Y(new_n6899_));
  INVX1    g04463(.A(pi0152), .Y(new_n6900_));
  NOR3X1   g04464(.A(new_n6878_), .B(new_n5060_), .C(pi0095), .Y(new_n6901_));
  AOI21X1  g04465(.A0(new_n6901_), .A1(new_n5053_), .B0(new_n6870_), .Y(new_n6902_));
  NAND3X1  g04466(.A(new_n6902_), .B(new_n5033_), .C(new_n6900_), .Y(new_n6903_));
  NAND2X1  g04467(.A(new_n6903_), .B(new_n3158_), .Y(new_n6904_));
  INVX1    g04468(.A(new_n6893_), .Y(new_n6905_));
  NOR2X1   g04469(.A(new_n5070_), .B(new_n5057_), .Y(new_n6906_));
  NOR3X1   g04470(.A(new_n6883_), .B(new_n6878_), .C(pi0095), .Y(new_n6907_));
  OAI21X1  g04471(.A0(new_n6907_), .A1(new_n6870_), .B0(new_n6906_), .Y(new_n6908_));
  OAI21X1  g04472(.A0(new_n6908_), .A1(new_n6900_), .B0(new_n6885_), .Y(new_n6909_));
  AOI21X1  g04473(.A0(new_n6909_), .A1(pi0154), .B0(new_n6905_), .Y(new_n6910_));
  OAI21X1  g04474(.A0(new_n6904_), .A1(new_n6899_), .B0(new_n6910_), .Y(new_n6911_));
  AOI22X1  g04475(.A0(new_n6911_), .A1(new_n6895_), .B0(new_n6892_), .B1(new_n2953_), .Y(new_n6912_));
  INVX1    g04476(.A(new_n6886_), .Y(new_n6913_));
  OR2X1    g04477(.A(new_n5050_), .B(new_n5057_), .Y(new_n6914_));
  OR4X1    g04478(.A(new_n6878_), .B(new_n5060_), .C(new_n6914_), .D(pi0095), .Y(new_n6915_));
  OAI21X1  g04479(.A0(new_n6915_), .A1(new_n6913_), .B0(new_n6869_), .Y(new_n6916_));
  NAND2X1  g04480(.A(new_n6916_), .B(new_n2953_), .Y(new_n6917_));
  AOI21X1  g04481(.A0(new_n6917_), .A1(new_n6912_), .B0(new_n6868_), .Y(new_n6918_));
  AND2X1   g04482(.A(pi0232), .B(pi0176), .Y(new_n6919_));
  INVX1    g04483(.A(new_n6919_), .Y(new_n6920_));
  NOR2X1   g04484(.A(new_n6920_), .B(new_n6912_), .Y(new_n6921_));
  INVX1    g04485(.A(new_n6895_), .Y(new_n6922_));
  AND2X1   g04486(.A(new_n6898_), .B(new_n5051_), .Y(new_n6923_));
  OAI21X1  g04487(.A0(new_n6923_), .A1(new_n6896_), .B0(new_n6888_), .Y(new_n6924_));
  OAI22X1  g04488(.A0(new_n6924_), .A1(pi0299), .B0(new_n6899_), .B1(new_n6922_), .Y(new_n6925_));
  AND2X1   g04489(.A(new_n6925_), .B(new_n5237_), .Y(new_n6926_));
  OR4X1    g04490(.A(new_n6926_), .B(new_n6921_), .C(new_n6918_), .D(new_n2959_), .Y(new_n6927_));
  INVX1    g04491(.A(pi0183), .Y(new_n6928_));
  NOR2X1   g04492(.A(new_n6869_), .B(new_n2540_), .Y(new_n6929_));
  NOR2X1   g04493(.A(pi0479), .B(pi0040), .Y(new_n6930_));
  INVX1    g04494(.A(new_n6930_), .Y(new_n6931_));
  AND2X1   g04495(.A(new_n6878_), .B(new_n2607_), .Y(new_n6932_));
  INVX1    g04496(.A(new_n6932_), .Y(new_n6933_));
  OAI22X1  g04497(.A0(new_n6933_), .A1(new_n6931_), .B0(new_n6929_), .B1(new_n2455_), .Y(new_n6934_));
  INVX1    g04498(.A(new_n6934_), .Y(new_n6935_));
  OR2X1    g04499(.A(new_n6869_), .B(new_n2456_), .Y(new_n6936_));
  NOR2X1   g04500(.A(pi0096), .B(pi0072), .Y(new_n6937_));
  INVX1    g04501(.A(new_n6937_), .Y(new_n6938_));
  OAI21X1  g04502(.A0(new_n6877_), .A1(new_n2472_), .B0(pi0070), .Y(new_n6939_));
  INVX1    g04503(.A(new_n6939_), .Y(new_n6940_));
  AOI21X1  g04504(.A0(new_n6876_), .A1(new_n2607_), .B0(new_n2502_), .Y(new_n6941_));
  NOR3X1   g04505(.A(new_n6873_), .B(new_n2471_), .C(pi0060), .Y(new_n6942_));
  AOI21X1  g04506(.A0(new_n6767_), .A1(new_n2494_), .B0(new_n2745_), .Y(new_n6943_));
  INVX1    g04507(.A(new_n6943_), .Y(new_n6944_));
  OAI21X1  g04508(.A0(new_n6942_), .A1(new_n2493_), .B0(new_n6944_), .Y(new_n6945_));
  OR4X1    g04509(.A(pi0111), .B(pi0103), .C(pi0083), .D(pi0036), .Y(new_n6946_));
  OR4X1    g04510(.A(new_n6946_), .B(pi0069), .C(pi0068), .D(pi0067), .Y(new_n6947_));
  INVX1    g04511(.A(pi0073), .Y(new_n6948_));
  OR4X1    g04512(.A(pi0084), .B(pi0082), .C(new_n6948_), .D(pi0066), .Y(new_n6949_));
  NOR4X1   g04513(.A(new_n6949_), .B(new_n6947_), .C(new_n6873_), .D(new_n2642_), .Y(new_n6950_));
  AOI21X1  g04514(.A0(new_n6950_), .A1(new_n2475_), .B0(new_n2472_), .Y(new_n6951_));
  AOI21X1  g04515(.A0(new_n6951_), .A1(new_n6945_), .B0(new_n2498_), .Y(new_n6952_));
  INVX1    g04516(.A(new_n6952_), .Y(new_n6953_));
  INVX1    g04517(.A(new_n2505_), .Y(new_n6954_));
  AOI21X1  g04518(.A0(new_n2498_), .A1(new_n2472_), .B0(new_n6954_), .Y(new_n6955_));
  OAI21X1  g04519(.A0(new_n2505_), .A1(new_n2472_), .B0(new_n2502_), .Y(new_n6956_));
  AOI21X1  g04520(.A0(new_n6955_), .A1(new_n6953_), .B0(new_n6956_), .Y(new_n6957_));
  OAI21X1  g04521(.A0(new_n6957_), .A1(new_n6941_), .B0(new_n2701_), .Y(new_n6958_));
  NOR3X1   g04522(.A(new_n6876_), .B(pi0841), .C(pi0058), .Y(new_n6959_));
  OAI21X1  g04523(.A0(new_n6959_), .A1(new_n2472_), .B0(pi0090), .Y(new_n6960_));
  AND2X1   g04524(.A(new_n6960_), .B(new_n2541_), .Y(new_n6961_));
  AOI21X1  g04525(.A0(new_n2542_), .A1(new_n2607_), .B0(pi0070), .Y(new_n6962_));
  INVX1    g04526(.A(new_n6962_), .Y(new_n6963_));
  AOI21X1  g04527(.A0(new_n6961_), .A1(new_n6958_), .B0(new_n6963_), .Y(new_n6964_));
  OAI21X1  g04528(.A0(new_n6964_), .A1(new_n6940_), .B0(new_n2516_), .Y(new_n6965_));
  AOI21X1  g04529(.A0(new_n2472_), .A1(pi0051), .B0(new_n6938_), .Y(new_n6966_));
  AOI22X1  g04530(.A0(new_n6966_), .A1(new_n6965_), .B0(new_n6938_), .B1(new_n2607_), .Y(new_n6967_));
  OAI21X1  g04531(.A0(new_n6967_), .A1(pi0040), .B0(new_n2456_), .Y(new_n6968_));
  AOI21X1  g04532(.A0(new_n6968_), .A1(new_n6936_), .B0(pi0095), .Y(new_n6969_));
  NOR2X1   g04533(.A(new_n6969_), .B(new_n6935_), .Y(new_n6970_));
  OR2X1    g04534(.A(pi0093), .B(pi0072), .Y(new_n6971_));
  NOR3X1   g04535(.A(new_n6971_), .B(new_n2485_), .C(pi0090), .Y(new_n6972_));
  AOI21X1  g04536(.A0(new_n6972_), .A1(new_n6959_), .B0(new_n6870_), .Y(new_n6973_));
  NOR2X1   g04537(.A(new_n6973_), .B(new_n2456_), .Y(new_n6974_));
  INVX1    g04538(.A(new_n6974_), .Y(new_n6975_));
  AOI21X1  g04539(.A0(new_n6975_), .A1(new_n6968_), .B0(pi0095), .Y(new_n6976_));
  NAND2X1  g04540(.A(new_n6976_), .B(new_n2973_), .Y(new_n6977_));
  AND2X1   g04541(.A(new_n6977_), .B(new_n6970_), .Y(new_n6978_));
  AND2X1   g04542(.A(new_n6978_), .B(new_n5057_), .Y(new_n6979_));
  OAI21X1  g04543(.A0(new_n6945_), .A1(new_n6875_), .B0(new_n2607_), .Y(new_n6980_));
  AOI21X1  g04544(.A0(new_n6980_), .A1(new_n2502_), .B0(new_n6941_), .Y(new_n6981_));
  OAI21X1  g04545(.A0(new_n6981_), .A1(pi0090), .B0(new_n6961_), .Y(new_n6982_));
  AOI21X1  g04546(.A0(new_n6982_), .A1(new_n6962_), .B0(new_n6940_), .Y(new_n6983_));
  OAI21X1  g04547(.A0(new_n6983_), .A1(pi0051), .B0(new_n6966_), .Y(new_n6984_));
  OAI21X1  g04548(.A0(new_n6937_), .A1(new_n2472_), .B0(new_n6984_), .Y(new_n6985_));
  AND2X1   g04549(.A(new_n6985_), .B(new_n2549_), .Y(new_n6986_));
  OR2X1    g04550(.A(new_n6986_), .B(pi0032), .Y(new_n6987_));
  AOI21X1  g04551(.A0(new_n6987_), .A1(new_n6975_), .B0(pi0095), .Y(new_n6988_));
  AND2X1   g04552(.A(new_n6988_), .B(new_n2973_), .Y(new_n6989_));
  AOI21X1  g04553(.A0(new_n6987_), .A1(new_n6936_), .B0(pi0095), .Y(new_n6990_));
  NOR4X1   g04554(.A(new_n6990_), .B(new_n6989_), .C(new_n6929_), .D(new_n5057_), .Y(new_n6991_));
  OR2X1    g04555(.A(new_n6991_), .B(new_n6979_), .Y(new_n6992_));
  INVX1    g04556(.A(new_n6978_), .Y(new_n6993_));
  NOR2X1   g04557(.A(new_n6929_), .B(new_n5057_), .Y(new_n6994_));
  AOI21X1  g04558(.A0(new_n2472_), .A1(pi0032), .B0(pi0040), .Y(new_n6995_));
  INVX1    g04559(.A(new_n6995_), .Y(new_n6996_));
  AND2X1   g04560(.A(new_n2543_), .B(new_n2518_), .Y(new_n6997_));
  INVX1    g04561(.A(new_n6997_), .Y(new_n6998_));
  AOI21X1  g04562(.A0(new_n6998_), .A1(new_n2607_), .B0(pi0032), .Y(new_n6999_));
  AOI21X1  g04563(.A0(new_n2472_), .A1(pi0093), .B0(new_n6998_), .Y(new_n7000_));
  OAI21X1  g04564(.A0(new_n6941_), .A1(new_n2472_), .B0(new_n2701_), .Y(new_n7001_));
  AND2X1   g04565(.A(new_n7001_), .B(new_n6960_), .Y(new_n7002_));
  OAI21X1  g04566(.A0(new_n7002_), .A1(pi0093), .B0(new_n7000_), .Y(new_n7003_));
  AOI21X1  g04567(.A0(new_n7003_), .A1(new_n6999_), .B0(new_n6996_), .Y(new_n7004_));
  OAI21X1  g04568(.A0(new_n7004_), .A1(pi0095), .B0(new_n6994_), .Y(new_n7005_));
  OAI21X1  g04569(.A0(new_n6993_), .A1(new_n5033_), .B0(new_n7005_), .Y(new_n7006_));
  MX2X1    g04570(.A(new_n7006_), .B(new_n6992_), .S0(new_n6928_), .Y(new_n7007_));
  INVX1    g04571(.A(pi0174), .Y(new_n7008_));
  AND2X1   g04572(.A(new_n6934_), .B(new_n7008_), .Y(new_n7009_));
  OAI21X1  g04573(.A0(new_n7007_), .A1(pi0095), .B0(new_n7009_), .Y(new_n7010_));
  AND2X1   g04574(.A(new_n5033_), .B(pi0183), .Y(new_n7011_));
  NAND3X1  g04575(.A(new_n6950_), .B(new_n6786_), .C(new_n2701_), .Y(new_n7012_));
  AND2X1   g04576(.A(new_n7012_), .B(new_n7002_), .Y(new_n7013_));
  OAI21X1  g04577(.A0(new_n7013_), .A1(pi0093), .B0(new_n7000_), .Y(new_n7014_));
  AOI21X1  g04578(.A0(new_n7014_), .A1(new_n6999_), .B0(new_n6996_), .Y(new_n7015_));
  NOR2X1   g04579(.A(new_n7015_), .B(pi0095), .Y(new_n7016_));
  OAI21X1  g04580(.A0(new_n7016_), .A1(new_n6935_), .B0(new_n5033_), .Y(new_n7017_));
  INVX1    g04581(.A(new_n7017_), .Y(new_n7018_));
  AOI21X1  g04582(.A0(new_n7018_), .A1(pi0183), .B0(new_n7008_), .Y(new_n7019_));
  OAI21X1  g04583(.A0(new_n7011_), .A1(new_n6978_), .B0(new_n7019_), .Y(new_n7020_));
  AND2X1   g04584(.A(new_n7020_), .B(new_n5225_), .Y(new_n7021_));
  NAND2X1  g04585(.A(new_n7007_), .B(new_n7008_), .Y(new_n7022_));
  NOR3X1   g04586(.A(new_n7016_), .B(new_n6929_), .C(new_n5057_), .Y(new_n7023_));
  OR2X1    g04587(.A(new_n7023_), .B(new_n6979_), .Y(new_n7024_));
  NOR3X1   g04588(.A(pi0468), .B(pi0332), .C(pi0040), .Y(new_n7025_));
  NOR2X1   g04589(.A(new_n6969_), .B(new_n6929_), .Y(new_n7026_));
  NAND3X1  g04590(.A(new_n7026_), .B(new_n7025_), .C(new_n6977_), .Y(new_n7027_));
  OAI21X1  g04591(.A0(new_n6993_), .A1(new_n5033_), .B0(new_n7027_), .Y(new_n7028_));
  MX2X1    g04592(.A(new_n7028_), .B(new_n7024_), .S0(pi0183), .Y(new_n7029_));
  AOI21X1  g04593(.A0(new_n7029_), .A1(pi0174), .B0(new_n5225_), .Y(new_n7030_));
  AOI22X1  g04594(.A0(new_n7030_), .A1(new_n7022_), .B0(new_n7021_), .B1(new_n7010_), .Y(new_n7031_));
  AOI21X1  g04595(.A0(new_n2472_), .A1(new_n2549_), .B0(new_n2456_), .Y(new_n7032_));
  INVX1    g04596(.A(new_n7032_), .Y(new_n7033_));
  INVX1    g04597(.A(new_n6966_), .Y(new_n7034_));
  OR4X1    g04598(.A(pi0093), .B(pi0090), .C(pi0058), .D(pi0035), .Y(new_n7035_));
  AND2X1   g04599(.A(new_n7035_), .B(new_n2472_), .Y(new_n7036_));
  AOI21X1  g04600(.A0(new_n6957_), .A1(new_n5907_), .B0(new_n7036_), .Y(new_n7037_));
  OAI21X1  g04601(.A0(new_n7037_), .A1(pi0070), .B0(new_n6939_), .Y(new_n7038_));
  AOI21X1  g04602(.A0(new_n7038_), .A1(new_n2516_), .B0(new_n7034_), .Y(new_n7039_));
  OAI21X1  g04603(.A0(new_n6937_), .A1(new_n2472_), .B0(new_n2549_), .Y(new_n7040_));
  OAI21X1  g04604(.A0(new_n7040_), .A1(new_n7039_), .B0(new_n2456_), .Y(new_n7041_));
  AOI22X1  g04605(.A0(new_n7041_), .A1(new_n7033_), .B0(new_n6870_), .B1(new_n2768_), .Y(new_n7042_));
  NOR2X1   g04606(.A(new_n7042_), .B(pi0095), .Y(new_n7043_));
  NOR2X1   g04607(.A(new_n7043_), .B(new_n6935_), .Y(new_n7044_));
  INVX1    g04608(.A(new_n7044_), .Y(new_n7045_));
  NOR3X1   g04609(.A(new_n6869_), .B(pi0468), .C(pi0332), .Y(new_n7046_));
  INVX1    g04610(.A(new_n7046_), .Y(new_n7047_));
  MX2X1    g04611(.A(new_n7042_), .B(new_n6869_), .S0(pi0095), .Y(new_n7048_));
  AOI21X1  g04612(.A0(new_n2472_), .A1(new_n2549_), .B0(new_n2540_), .Y(new_n7049_));
  OAI21X1  g04613(.A0(new_n6973_), .A1(pi0040), .B0(pi0032), .Y(new_n7050_));
  AOI21X1  g04614(.A0(new_n7050_), .A1(new_n7041_), .B0(pi0095), .Y(new_n7051_));
  OR2X1    g04615(.A(new_n7051_), .B(new_n7049_), .Y(new_n7052_));
  AND2X1   g04616(.A(new_n7052_), .B(new_n7048_), .Y(new_n7053_));
  OAI21X1  g04617(.A0(new_n7053_), .A1(pi0198), .B0(new_n5033_), .Y(new_n7054_));
  AOI21X1  g04618(.A0(new_n7054_), .A1(new_n7047_), .B0(new_n7045_), .Y(new_n7055_));
  OAI21X1  g04619(.A0(new_n7055_), .A1(new_n6979_), .B0(new_n6928_), .Y(new_n7056_));
  OR4X1    g04620(.A(new_n6998_), .B(new_n2492_), .C(new_n2484_), .D(new_n2478_), .Y(new_n7057_));
  NOR2X1   g04621(.A(new_n7057_), .B(pi0032), .Y(new_n7058_));
  AOI21X1  g04622(.A0(new_n7058_), .A1(new_n6950_), .B0(new_n6870_), .Y(new_n7059_));
  NOR2X1   g04623(.A(new_n7059_), .B(pi0095), .Y(new_n7060_));
  NOR3X1   g04624(.A(new_n7060_), .B(new_n6935_), .C(new_n5057_), .Y(new_n7061_));
  OAI21X1  g04625(.A0(new_n7061_), .A1(new_n6979_), .B0(pi0183), .Y(new_n7062_));
  AND2X1   g04626(.A(new_n7062_), .B(pi0174), .Y(new_n7063_));
  AOI21X1  g04627(.A0(new_n6977_), .A1(new_n6970_), .B0(new_n5033_), .Y(new_n7064_));
  INVX1    g04628(.A(new_n7036_), .Y(new_n7065_));
  NAND3X1  g04629(.A(new_n6980_), .B(new_n5907_), .C(new_n2502_), .Y(new_n7066_));
  AOI21X1  g04630(.A0(new_n7066_), .A1(new_n7065_), .B0(pi0070), .Y(new_n7067_));
  OAI21X1  g04631(.A0(new_n7067_), .A1(new_n6940_), .B0(new_n2516_), .Y(new_n7068_));
  AOI22X1  g04632(.A0(new_n7068_), .A1(new_n6966_), .B0(new_n6938_), .B1(new_n2607_), .Y(new_n7069_));
  OAI21X1  g04633(.A0(new_n7069_), .A1(pi0040), .B0(new_n2456_), .Y(new_n7070_));
  AOI21X1  g04634(.A0(new_n7070_), .A1(new_n6936_), .B0(pi0095), .Y(new_n7071_));
  NOR2X1   g04635(.A(new_n7071_), .B(new_n6935_), .Y(new_n7072_));
  AOI21X1  g04636(.A0(new_n7070_), .A1(new_n6975_), .B0(pi0095), .Y(new_n7073_));
  NAND2X1  g04637(.A(new_n7073_), .B(new_n2973_), .Y(new_n7074_));
  NAND2X1  g04638(.A(new_n7074_), .B(new_n7072_), .Y(new_n7075_));
  AOI21X1  g04639(.A0(new_n7075_), .A1(new_n5033_), .B0(new_n7064_), .Y(new_n7076_));
  AND2X1   g04640(.A(new_n7076_), .B(new_n6928_), .Y(new_n7077_));
  AOI21X1  g04641(.A0(new_n6870_), .A1(new_n2540_), .B0(new_n6935_), .Y(new_n7078_));
  AOI21X1  g04642(.A0(new_n7078_), .A1(new_n5033_), .B0(new_n6979_), .Y(new_n7079_));
  OAI21X1  g04643(.A0(new_n7079_), .A1(new_n6928_), .B0(new_n7008_), .Y(new_n7080_));
  OAI21X1  g04644(.A0(new_n7080_), .A1(new_n7077_), .B0(new_n5225_), .Y(new_n7081_));
  AOI21X1  g04645(.A0(new_n7063_), .A1(new_n7056_), .B0(new_n7081_), .Y(new_n7082_));
  INVX1    g04646(.A(pi0193), .Y(new_n7083_));
  INVX1    g04647(.A(new_n7048_), .Y(new_n7084_));
  OAI22X1  g04648(.A0(new_n7054_), .A1(new_n7084_), .B0(new_n6993_), .B1(new_n5033_), .Y(new_n7085_));
  AND2X1   g04649(.A(new_n7085_), .B(new_n6928_), .Y(new_n7086_));
  INVX1    g04650(.A(new_n6979_), .Y(new_n7087_));
  OAI21X1  g04651(.A0(new_n7059_), .A1(pi0095), .B0(new_n6994_), .Y(new_n7088_));
  AOI21X1  g04652(.A0(new_n7088_), .A1(new_n7087_), .B0(new_n6928_), .Y(new_n7089_));
  NOR3X1   g04653(.A(new_n7089_), .B(new_n7086_), .C(new_n7008_), .Y(new_n7090_));
  NOR3X1   g04654(.A(new_n7064_), .B(new_n7046_), .C(new_n6928_), .Y(new_n7091_));
  INVX1    g04655(.A(new_n7025_), .Y(new_n7092_));
  INVX1    g04656(.A(new_n7049_), .Y(new_n7093_));
  AOI21X1  g04657(.A0(new_n7069_), .A1(new_n2549_), .B0(pi0032), .Y(new_n7094_));
  OAI21X1  g04658(.A0(new_n7094_), .A1(new_n7032_), .B0(new_n2540_), .Y(new_n7095_));
  AOI21X1  g04659(.A0(new_n7095_), .A1(new_n7093_), .B0(new_n2973_), .Y(new_n7096_));
  INVX1    g04660(.A(new_n7050_), .Y(new_n7097_));
  OAI21X1  g04661(.A0(new_n7094_), .A1(new_n7097_), .B0(new_n2540_), .Y(new_n7098_));
  AOI21X1  g04662(.A0(new_n7098_), .A1(new_n7093_), .B0(pi0198), .Y(new_n7099_));
  NOR2X1   g04663(.A(new_n7099_), .B(new_n7096_), .Y(new_n7100_));
  OAI22X1  g04664(.A0(new_n7100_), .A1(new_n7092_), .B0(new_n6993_), .B1(new_n5033_), .Y(new_n7101_));
  AND2X1   g04665(.A(new_n7101_), .B(new_n6928_), .Y(new_n7102_));
  NOR3X1   g04666(.A(new_n7102_), .B(new_n7091_), .C(pi0174), .Y(new_n7103_));
  NOR3X1   g04667(.A(new_n7103_), .B(new_n7090_), .C(new_n5225_), .Y(new_n7104_));
  OR2X1    g04668(.A(new_n7104_), .B(new_n7083_), .Y(new_n7105_));
  OAI22X1  g04669(.A0(new_n7105_), .A1(new_n7082_), .B0(new_n7031_), .B1(pi0193), .Y(new_n7106_));
  AND2X1   g04670(.A(pi0299), .B(pi0158), .Y(new_n7107_));
  AND2X1   g04671(.A(new_n6976_), .B(new_n2766_), .Y(new_n7108_));
  NOR4X1   g04672(.A(new_n7108_), .B(new_n6969_), .C(new_n6935_), .D(new_n5033_), .Y(new_n7109_));
  AND2X1   g04673(.A(new_n6988_), .B(new_n2766_), .Y(new_n7110_));
  NOR4X1   g04674(.A(new_n7110_), .B(new_n6990_), .C(new_n6929_), .D(new_n5057_), .Y(new_n7111_));
  NOR2X1   g04675(.A(new_n7111_), .B(new_n7109_), .Y(new_n7112_));
  NOR2X1   g04676(.A(new_n7112_), .B(pi0152), .Y(new_n7113_));
  NOR3X1   g04677(.A(new_n7108_), .B(new_n6969_), .C(new_n6935_), .Y(new_n7114_));
  INVX1    g04678(.A(new_n7026_), .Y(new_n7115_));
  OAI21X1  g04679(.A0(new_n7108_), .A1(new_n7115_), .B0(new_n5033_), .Y(new_n7116_));
  OAI21X1  g04680(.A0(new_n7114_), .A1(new_n5033_), .B0(new_n7116_), .Y(new_n7117_));
  OAI21X1  g04681(.A0(new_n7117_), .A1(new_n6900_), .B0(new_n3601_), .Y(new_n7118_));
  INVX1    g04682(.A(new_n7109_), .Y(new_n7119_));
  OAI21X1  g04683(.A0(new_n7053_), .A1(pi0210), .B0(new_n5033_), .Y(new_n7120_));
  OAI21X1  g04684(.A0(new_n7120_), .A1(new_n7084_), .B0(new_n7119_), .Y(new_n7121_));
  AND2X1   g04685(.A(new_n7121_), .B(pi0152), .Y(new_n7122_));
  OAI21X1  g04686(.A0(new_n7073_), .A1(new_n6929_), .B0(new_n2766_), .Y(new_n7123_));
  NAND2X1  g04687(.A(new_n7123_), .B(new_n5033_), .Y(new_n7124_));
  NOR3X1   g04688(.A(new_n7124_), .B(new_n7071_), .C(new_n6929_), .Y(new_n7125_));
  OAI21X1  g04689(.A0(new_n7125_), .A1(new_n7109_), .B0(new_n6900_), .Y(new_n7126_));
  NAND2X1  g04690(.A(new_n7126_), .B(pi0172), .Y(new_n7127_));
  OAI22X1  g04691(.A0(new_n7127_), .A1(new_n7122_), .B0(new_n7118_), .B1(new_n7113_), .Y(new_n7128_));
  INVX1    g04692(.A(pi0149), .Y(new_n7129_));
  AOI21X1  g04693(.A0(new_n7120_), .A1(new_n7047_), .B0(new_n7045_), .Y(new_n7130_));
  INVX1    g04694(.A(new_n7130_), .Y(new_n7131_));
  INVX1    g04695(.A(new_n7072_), .Y(new_n7132_));
  AOI21X1  g04696(.A0(new_n7124_), .A1(new_n7047_), .B0(new_n7132_), .Y(new_n7133_));
  OAI21X1  g04697(.A0(new_n7133_), .A1(pi0152), .B0(pi0172), .Y(new_n7134_));
  AOI21X1  g04698(.A0(new_n7131_), .A1(pi0152), .B0(new_n7134_), .Y(new_n7135_));
  NOR4X1   g04699(.A(new_n7110_), .B(new_n6990_), .C(new_n6935_), .D(new_n5057_), .Y(new_n7136_));
  NOR2X1   g04700(.A(new_n7136_), .B(pi0152), .Y(new_n7137_));
  OAI21X1  g04701(.A0(new_n7114_), .A1(new_n6900_), .B0(new_n3601_), .Y(new_n7138_));
  AND2X1   g04702(.A(pi0299), .B(new_n5128_), .Y(new_n7139_));
  INVX1    g04703(.A(new_n7139_), .Y(new_n7140_));
  NOR2X1   g04704(.A(new_n7140_), .B(new_n7109_), .Y(new_n7141_));
  OAI21X1  g04705(.A0(new_n7138_), .A1(new_n7137_), .B0(new_n7141_), .Y(new_n7142_));
  OAI21X1  g04706(.A0(new_n7142_), .A1(new_n7135_), .B0(new_n7129_), .Y(new_n7143_));
  AOI21X1  g04707(.A0(new_n7128_), .A1(new_n7107_), .B0(new_n7143_), .Y(new_n7144_));
  OR2X1    g04708(.A(new_n7109_), .B(new_n7023_), .Y(new_n7145_));
  NOR2X1   g04709(.A(new_n7004_), .B(pi0095), .Y(new_n7146_));
  INVX1    g04710(.A(new_n7146_), .Y(new_n7147_));
  AOI21X1  g04711(.A0(new_n7147_), .A1(new_n6994_), .B0(new_n7109_), .Y(new_n7148_));
  OAI21X1  g04712(.A0(new_n7148_), .A1(pi0152), .B0(new_n3601_), .Y(new_n7149_));
  AOI21X1  g04713(.A0(new_n7145_), .A1(pi0152), .B0(new_n7149_), .Y(new_n7150_));
  NAND2X1  g04714(.A(new_n7119_), .B(new_n7088_), .Y(new_n7151_));
  OAI21X1  g04715(.A0(new_n7114_), .A1(new_n5033_), .B0(new_n7047_), .Y(new_n7152_));
  OAI21X1  g04716(.A0(new_n7152_), .A1(pi0152), .B0(pi0172), .Y(new_n7153_));
  AOI21X1  g04717(.A0(new_n7151_), .A1(pi0152), .B0(new_n7153_), .Y(new_n7154_));
  OAI21X1  g04718(.A0(new_n7154_), .A1(new_n7150_), .B0(new_n7107_), .Y(new_n7155_));
  OR2X1    g04719(.A(new_n7109_), .B(new_n7061_), .Y(new_n7156_));
  AND2X1   g04720(.A(new_n7156_), .B(pi0152), .Y(new_n7157_));
  AOI21X1  g04721(.A0(new_n7078_), .A1(new_n5033_), .B0(new_n7109_), .Y(new_n7158_));
  OAI21X1  g04722(.A0(new_n7158_), .A1(pi0152), .B0(pi0172), .Y(new_n7159_));
  NOR2X1   g04723(.A(new_n7114_), .B(new_n5033_), .Y(new_n7160_));
  AOI21X1  g04724(.A0(new_n7147_), .A1(new_n6934_), .B0(new_n5057_), .Y(new_n7161_));
  NOR3X1   g04725(.A(new_n7161_), .B(new_n7160_), .C(pi0152), .Y(new_n7162_));
  OAI21X1  g04726(.A0(new_n7114_), .A1(new_n5033_), .B0(new_n7017_), .Y(new_n7163_));
  OAI21X1  g04727(.A0(new_n7163_), .A1(new_n6900_), .B0(new_n3601_), .Y(new_n7164_));
  OAI22X1  g04728(.A0(new_n7164_), .A1(new_n7162_), .B0(new_n7159_), .B1(new_n7157_), .Y(new_n7165_));
  AOI21X1  g04729(.A0(new_n7165_), .A1(new_n7139_), .B0(new_n7129_), .Y(new_n7166_));
  AOI21X1  g04730(.A0(new_n7166_), .A1(new_n7155_), .B0(new_n7144_), .Y(new_n7167_));
  AOI21X1  g04731(.A0(new_n7106_), .A1(new_n2953_), .B0(new_n7167_), .Y(new_n7168_));
  INVX1    g04732(.A(new_n5019_), .Y(new_n7169_));
  AND2X1   g04733(.A(new_n6976_), .B(new_n7169_), .Y(new_n7170_));
  NOR3X1   g04734(.A(new_n7170_), .B(new_n6969_), .C(new_n6935_), .Y(new_n7171_));
  NOR2X1   g04735(.A(new_n7171_), .B(pi0232), .Y(new_n7172_));
  NOR2X1   g04736(.A(new_n7172_), .B(pi0039), .Y(new_n7173_));
  OAI21X1  g04737(.A0(new_n7168_), .A1(new_n5237_), .B0(new_n7173_), .Y(new_n7174_));
  AOI21X1  g04738(.A0(new_n7174_), .A1(new_n6927_), .B0(pi0038), .Y(new_n7175_));
  OAI21X1  g04739(.A0(new_n7175_), .A1(new_n6865_), .B0(new_n3026_), .Y(new_n7176_));
  NOR2X1   g04740(.A(new_n6842_), .B(pi0087), .Y(new_n7177_));
  NOR2X1   g04741(.A(new_n6850_), .B(new_n2996_), .Y(new_n7178_));
  AOI21X1  g04742(.A0(new_n7178_), .A1(new_n3026_), .B0(new_n6842_), .Y(new_n7179_));
  AND2X1   g04743(.A(new_n6869_), .B(new_n3277_), .Y(new_n7180_));
  INVX1    g04744(.A(new_n7180_), .Y(new_n7181_));
  NAND3X1  g04745(.A(new_n7181_), .B(new_n7179_), .C(pi0087), .Y(new_n7182_));
  NAND2X1  g04746(.A(new_n7182_), .B(new_n3105_), .Y(new_n7183_));
  AOI21X1  g04747(.A0(new_n7177_), .A1(new_n7176_), .B0(new_n7183_), .Y(new_n7184_));
  AND2X1   g04748(.A(pi0092), .B(new_n3095_), .Y(new_n7185_));
  INVX1    g04749(.A(new_n7185_), .Y(new_n7186_));
  INVX1    g04750(.A(new_n7179_), .Y(new_n7187_));
  OR2X1    g04751(.A(pi0087), .B(pi0039), .Y(new_n7188_));
  AOI21X1  g04752(.A0(pi0299), .A1(new_n3158_), .B0(new_n5237_), .Y(new_n7189_));
  NOR2X1   g04753(.A(pi0299), .B(pi0176), .Y(new_n7190_));
  NOR3X1   g04754(.A(new_n7190_), .B(pi0468), .C(pi0332), .Y(new_n7191_));
  AND2X1   g04755(.A(new_n7191_), .B(new_n7189_), .Y(new_n7192_));
  OR4X1    g04756(.A(new_n7192_), .B(new_n6878_), .C(new_n7188_), .D(pi0095), .Y(new_n7193_));
  AOI21X1  g04757(.A0(new_n7193_), .A1(new_n7180_), .B0(new_n7187_), .Y(new_n7194_));
  OAI22X1  g04758(.A0(new_n7194_), .A1(new_n7186_), .B0(new_n6841_), .B1(new_n3095_), .Y(new_n7195_));
  OAI21X1  g04759(.A0(new_n7195_), .A1(new_n7184_), .B0(new_n3112_), .Y(new_n7196_));
  AOI21X1  g04760(.A0(new_n7196_), .A1(new_n6854_), .B0(pi0074), .Y(new_n7197_));
  AND2X1   g04761(.A(new_n6834_), .B(pi0055), .Y(new_n7198_));
  AOI21X1  g04762(.A0(new_n6829_), .A1(new_n6827_), .B0(new_n3112_), .Y(new_n7199_));
  AND2X1   g04763(.A(new_n6825_), .B(pi0232), .Y(new_n7200_));
  OAI21X1  g04764(.A0(new_n7200_), .A1(new_n3095_), .B0(new_n3100_), .Y(new_n7201_));
  INVX1    g04765(.A(new_n7201_), .Y(new_n7202_));
  AOI21X1  g04766(.A0(new_n5930_), .A1(pi0164), .B0(new_n2996_), .Y(new_n7203_));
  NOR2X1   g04767(.A(new_n7203_), .B(new_n3124_), .Y(new_n7204_));
  INVX1    g04768(.A(new_n7204_), .Y(new_n7205_));
  OAI21X1  g04769(.A0(new_n6855_), .A1(new_n7129_), .B0(new_n2959_), .Y(new_n7206_));
  OAI21X1  g04770(.A0(new_n7206_), .A1(new_n6880_), .B0(new_n6869_), .Y(new_n7207_));
  AOI21X1  g04771(.A0(new_n7207_), .A1(new_n2996_), .B0(new_n7205_), .Y(new_n7208_));
  AOI21X1  g04772(.A0(new_n6825_), .A1(pi0232), .B0(new_n3026_), .Y(new_n7209_));
  NOR2X1   g04773(.A(new_n6869_), .B(pi0038), .Y(new_n7210_));
  NOR4X1   g04774(.A(new_n7210_), .B(new_n7203_), .C(pi0100), .D(new_n3156_), .Y(new_n7211_));
  OR2X1    g04775(.A(new_n7211_), .B(new_n7209_), .Y(new_n7212_));
  OAI21X1  g04776(.A0(new_n7212_), .A1(new_n7208_), .B0(new_n3095_), .Y(new_n7213_));
  NOR4X1   g04777(.A(new_n7210_), .B(new_n7203_), .C(pi0100), .D(pi0075), .Y(new_n7214_));
  NAND2X1  g04778(.A(new_n6827_), .B(pi0092), .Y(new_n7215_));
  OAI21X1  g04779(.A0(new_n7215_), .A1(new_n7214_), .B0(new_n3112_), .Y(new_n7216_));
  AOI21X1  g04780(.A0(new_n7213_), .A1(new_n7202_), .B0(new_n7216_), .Y(new_n7217_));
  OAI21X1  g04781(.A0(new_n7217_), .A1(new_n7199_), .B0(new_n4991_), .Y(new_n7218_));
  AOI21X1  g04782(.A0(new_n7218_), .A1(new_n7198_), .B0(new_n5324_), .Y(new_n7219_));
  OAI21X1  g04783(.A0(new_n7197_), .A1(new_n6848_), .B0(new_n7219_), .Y(new_n7220_));
  INVX1    g04784(.A(new_n6834_), .Y(new_n7221_));
  INVX1    g04785(.A(new_n7199_), .Y(new_n7222_));
  INVX1    g04786(.A(pi0164), .Y(new_n7223_));
  NOR4X1   g04787(.A(new_n5057_), .B(new_n5237_), .C(new_n7223_), .D(new_n2996_), .Y(new_n7224_));
  AOI21X1  g04788(.A0(new_n7224_), .A1(new_n6828_), .B0(new_n6831_), .Y(new_n7225_));
  AOI21X1  g04789(.A0(new_n7225_), .A1(new_n7222_), .B0(pi0074), .Y(new_n7226_));
  OAI21X1  g04790(.A0(new_n7226_), .A1(new_n7221_), .B0(new_n5324_), .Y(new_n7227_));
  NAND2X1  g04791(.A(new_n7227_), .B(new_n3246_), .Y(new_n7228_));
  NOR4X1   g04792(.A(pi0107), .B(pi0063), .C(pi0040), .D(pi0038), .Y(new_n7229_));
  INVX1    g04793(.A(new_n7229_), .Y(new_n7230_));
  NOR4X1   g04794(.A(new_n7230_), .B(new_n6832_), .C(new_n3148_), .D(new_n3136_), .Y(new_n7231_));
  NOR2X1   g04795(.A(new_n7231_), .B(new_n7228_), .Y(new_n7232_));
  AOI21X1  g04796(.A0(new_n7232_), .A1(new_n7220_), .B0(new_n6836_), .Y(new_n7233_));
  INVX1    g04797(.A(new_n6848_), .Y(new_n7234_));
  NOR3X1   g04798(.A(new_n5257_), .B(new_n5070_), .C(new_n5057_), .Y(new_n7235_));
  NOR2X1   g04799(.A(new_n7235_), .B(new_n3158_), .Y(new_n7236_));
  AND2X1   g04800(.A(new_n5261_), .B(new_n6906_), .Y(new_n7237_));
  OAI21X1  g04801(.A0(new_n7237_), .A1(pi0154), .B0(new_n6900_), .Y(new_n7238_));
  AND2X1   g04802(.A(new_n5958_), .B(new_n2739_), .Y(new_n7239_));
  INVX1    g04803(.A(new_n7239_), .Y(new_n7240_));
  NOR4X1   g04804(.A(new_n7240_), .B(new_n5070_), .C(new_n5057_), .D(new_n2722_), .Y(new_n7241_));
  NAND3X1  g04805(.A(new_n7241_), .B(pi0154), .C(pi0152), .Y(new_n7242_));
  OAI21X1  g04806(.A0(new_n7238_), .A1(new_n7236_), .B0(new_n7242_), .Y(new_n7243_));
  AOI21X1  g04807(.A0(new_n7243_), .A1(new_n6893_), .B0(new_n2953_), .Y(new_n7244_));
  NAND4X1  g04808(.A(new_n6886_), .B(new_n5261_), .C(new_n5051_), .D(new_n5033_), .Y(new_n7245_));
  OAI21X1  g04809(.A0(new_n7245_), .A1(pi0174), .B0(new_n2953_), .Y(new_n7246_));
  OR4X1    g04810(.A(new_n6913_), .B(new_n5257_), .C(new_n6914_), .D(pi0174), .Y(new_n7247_));
  NOR4X1   g04811(.A(new_n6913_), .B(new_n7240_), .C(new_n6914_), .D(new_n2722_), .Y(new_n7248_));
  AOI21X1  g04812(.A0(new_n7248_), .A1(pi0174), .B0(pi0299), .Y(new_n7249_));
  AOI21X1  g04813(.A0(new_n7249_), .A1(new_n7247_), .B0(new_n6920_), .Y(new_n7250_));
  AOI21X1  g04814(.A0(new_n7246_), .A1(new_n6867_), .B0(new_n7250_), .Y(new_n7251_));
  NOR3X1   g04815(.A(new_n7251_), .B(new_n7244_), .C(new_n2959_), .Y(new_n7252_));
  AOI21X1  g04816(.A0(new_n2550_), .A1(new_n2726_), .B0(new_n2701_), .Y(new_n7253_));
  NOR3X1   g04817(.A(new_n7253_), .B(new_n5000_), .C(new_n2542_), .Y(new_n7254_));
  INVX1    g04818(.A(new_n7254_), .Y(new_n7255_));
  NOR4X1   g04819(.A(new_n2542_), .B(new_n2506_), .C(new_n2501_), .D(pi0090), .Y(new_n7256_));
  AND2X1   g04820(.A(new_n7256_), .B(new_n2607_), .Y(new_n7257_));
  AOI21X1  g04821(.A0(new_n7257_), .A1(new_n6952_), .B0(pi0070), .Y(new_n7258_));
  NOR3X1   g04822(.A(new_n3256_), .B(new_n2894_), .C(new_n2870_), .Y(new_n7259_));
  INVX1    g04823(.A(new_n7259_), .Y(new_n7260_));
  AOI21X1  g04824(.A0(new_n7258_), .A1(new_n7255_), .B0(new_n7260_), .Y(new_n7261_));
  INVX1    g04825(.A(new_n7261_), .Y(new_n7262_));
  NOR2X1   g04826(.A(new_n5195_), .B(pi0095), .Y(new_n7263_));
  NOR2X1   g04827(.A(new_n7260_), .B(new_n7258_), .Y(new_n7264_));
  NOR2X1   g04828(.A(new_n7264_), .B(new_n7263_), .Y(new_n7265_));
  OAI21X1  g04829(.A0(new_n7265_), .A1(pi0198), .B0(new_n7262_), .Y(new_n7266_));
  NOR3X1   g04830(.A(new_n7253_), .B(new_n6971_), .C(new_n2485_), .Y(new_n7267_));
  NAND3X1  g04831(.A(new_n6950_), .B(new_n6786_), .C(new_n2607_), .Y(new_n7268_));
  NAND2X1  g04832(.A(new_n7268_), .B(new_n5000_), .Y(new_n7269_));
  AND2X1   g04833(.A(new_n7269_), .B(new_n7267_), .Y(new_n7270_));
  NOR2X1   g04834(.A(pi0095), .B(pi0032), .Y(new_n7271_));
  INVX1    g04835(.A(new_n7271_), .Y(new_n7272_));
  NOR3X1   g04836(.A(new_n5057_), .B(new_n7272_), .C(pi0040), .Y(new_n7273_));
  AND2X1   g04837(.A(new_n7273_), .B(new_n7270_), .Y(new_n7274_));
  INVX1    g04838(.A(new_n7274_), .Y(new_n7275_));
  OAI21X1  g04839(.A0(new_n7275_), .A1(pi0183), .B0(new_n7008_), .Y(new_n7276_));
  AOI21X1  g04840(.A0(new_n7266_), .A1(new_n7011_), .B0(new_n7276_), .Y(new_n7277_));
  AOI21X1  g04841(.A0(new_n7256_), .A1(new_n6944_), .B0(pi0070), .Y(new_n7278_));
  AOI21X1  g04842(.A0(new_n7278_), .A1(new_n7255_), .B0(new_n7260_), .Y(new_n7279_));
  OAI21X1  g04843(.A0(new_n7279_), .A1(new_n5220_), .B0(new_n5033_), .Y(new_n7280_));
  OR2X1    g04844(.A(new_n7280_), .B(new_n6928_), .Y(new_n7281_));
  NOR4X1   g04845(.A(new_n7253_), .B(new_n6971_), .C(new_n5000_), .D(new_n2485_), .Y(new_n7282_));
  AND2X1   g04846(.A(new_n7282_), .B(new_n7273_), .Y(new_n7283_));
  AOI21X1  g04847(.A0(new_n7283_), .A1(new_n6928_), .B0(new_n7008_), .Y(new_n7284_));
  AND2X1   g04848(.A(new_n7284_), .B(new_n7281_), .Y(new_n7285_));
  OAI21X1  g04849(.A0(new_n7285_), .A1(new_n7277_), .B0(pi0193), .Y(new_n7286_));
  NOR3X1   g04850(.A(new_n7264_), .B(new_n5220_), .C(pi0174), .Y(new_n7287_));
  NOR2X1   g04851(.A(new_n7278_), .B(new_n7260_), .Y(new_n7288_));
  NOR3X1   g04852(.A(new_n7288_), .B(new_n5220_), .C(new_n7008_), .Y(new_n7289_));
  OR4X1    g04853(.A(new_n7289_), .B(new_n7287_), .C(new_n5057_), .D(new_n6928_), .Y(new_n7290_));
  NAND4X1  g04854(.A(new_n6972_), .B(new_n6950_), .C(new_n6786_), .D(new_n2607_), .Y(new_n7291_));
  NOR3X1   g04855(.A(new_n7291_), .B(new_n7092_), .C(new_n7272_), .Y(new_n7292_));
  NAND3X1  g04856(.A(new_n7292_), .B(new_n6928_), .C(new_n7008_), .Y(new_n7293_));
  NAND3X1  g04857(.A(new_n7293_), .B(new_n7290_), .C(new_n7083_), .Y(new_n7294_));
  AND2X1   g04858(.A(new_n5033_), .B(new_n2901_), .Y(new_n7295_));
  INVX1    g04859(.A(new_n7295_), .Y(new_n7296_));
  OAI21X1  g04860(.A0(new_n7296_), .A1(new_n5225_), .B0(new_n2953_), .Y(new_n7297_));
  AOI21X1  g04861(.A0(new_n7294_), .A1(new_n7286_), .B0(new_n7297_), .Y(new_n7298_));
  AND2X1   g04862(.A(pi0232), .B(new_n2959_), .Y(new_n7299_));
  INVX1    g04863(.A(new_n7299_), .Y(new_n7300_));
  NOR3X1   g04864(.A(new_n7264_), .B(new_n5196_), .C(pi0152), .Y(new_n7301_));
  OAI21X1  g04865(.A0(new_n7262_), .A1(new_n3601_), .B0(new_n7301_), .Y(new_n7302_));
  NOR2X1   g04866(.A(new_n7288_), .B(new_n5196_), .Y(new_n7303_));
  AOI21X1  g04867(.A0(new_n7279_), .A1(pi0172), .B0(new_n6900_), .Y(new_n7304_));
  NAND2X1  g04868(.A(new_n5033_), .B(pi0149), .Y(new_n7305_));
  AOI21X1  g04869(.A0(new_n7304_), .A1(new_n7303_), .B0(new_n7305_), .Y(new_n7306_));
  INVX1    g04870(.A(new_n7283_), .Y(new_n7307_));
  OAI21X1  g04871(.A0(new_n7275_), .A1(pi0152), .B0(new_n7307_), .Y(new_n7308_));
  NOR2X1   g04872(.A(pi0172), .B(pi0152), .Y(new_n7309_));
  AOI22X1  g04873(.A0(new_n7309_), .A1(new_n7292_), .B0(new_n7308_), .B1(pi0172), .Y(new_n7310_));
  AOI21X1  g04874(.A0(new_n7295_), .A1(pi0158), .B0(new_n2953_), .Y(new_n7311_));
  OAI21X1  g04875(.A0(new_n7310_), .A1(pi0149), .B0(new_n7311_), .Y(new_n7312_));
  AOI21X1  g04876(.A0(new_n7306_), .A1(new_n7302_), .B0(new_n7312_), .Y(new_n7313_));
  NOR3X1   g04877(.A(new_n7313_), .B(new_n7300_), .C(new_n7298_), .Y(new_n7314_));
  OAI21X1  g04878(.A0(new_n7314_), .A1(new_n7252_), .B0(new_n2996_), .Y(new_n7315_));
  NOR2X1   g04879(.A(new_n6865_), .B(pi0087), .Y(new_n7316_));
  OAI21X1  g04880(.A0(new_n7178_), .A1(new_n3156_), .B0(new_n3026_), .Y(new_n7317_));
  AOI21X1  g04881(.A0(new_n7316_), .A1(new_n7315_), .B0(new_n7317_), .Y(new_n7318_));
  OAI21X1  g04882(.A0(new_n7318_), .A1(new_n6842_), .B0(new_n3105_), .Y(new_n7319_));
  NOR2X1   g04883(.A(pi0087), .B(pi0038), .Y(new_n7320_));
  NAND4X1  g04884(.A(new_n7320_), .B(new_n7192_), .C(new_n4995_), .D(new_n3026_), .Y(new_n7321_));
  AOI21X1  g04885(.A0(new_n7321_), .A1(new_n7179_), .B0(new_n7186_), .Y(new_n7322_));
  NOR2X1   g04886(.A(new_n7322_), .B(new_n6843_), .Y(new_n7323_));
  AOI21X1  g04887(.A0(new_n7323_), .A1(new_n7319_), .B0(pi0054), .Y(new_n7324_));
  OAI21X1  g04888(.A0(new_n7324_), .A1(new_n6853_), .B0(new_n4991_), .Y(new_n7325_));
  INVX1    g04889(.A(new_n7198_), .Y(new_n7326_));
  NOR4X1   g04890(.A(new_n6855_), .B(new_n3015_), .C(new_n7129_), .D(pi0039), .Y(new_n7327_));
  OAI21X1  g04891(.A0(new_n7327_), .A1(pi0038), .B0(new_n7204_), .Y(new_n7328_));
  AND2X1   g04892(.A(new_n3026_), .B(pi0087), .Y(new_n7329_));
  AOI21X1  g04893(.A0(new_n7224_), .A1(new_n7329_), .B0(new_n7209_), .Y(new_n7330_));
  AOI21X1  g04894(.A0(new_n7330_), .A1(new_n7328_), .B0(pi0075), .Y(new_n7331_));
  AOI21X1  g04895(.A0(new_n7225_), .A1(pi0092), .B0(pi0054), .Y(new_n7332_));
  OAI21X1  g04896(.A0(new_n7331_), .A1(new_n7201_), .B0(new_n7332_), .Y(new_n7333_));
  AOI21X1  g04897(.A0(new_n7333_), .A1(new_n7222_), .B0(pi0074), .Y(new_n7334_));
  OAI21X1  g04898(.A0(new_n7334_), .A1(new_n7326_), .B0(new_n3148_), .Y(new_n7335_));
  AOI21X1  g04899(.A0(new_n7325_), .A1(new_n7234_), .B0(new_n7335_), .Y(new_n7336_));
  OAI22X1  g04900(.A0(new_n7336_), .A1(new_n7228_), .B0(new_n6835_), .B1(new_n6830_), .Y(new_n7337_));
  AOI21X1  g04901(.A0(new_n7337_), .A1(new_n6821_), .B0(pi0954), .Y(new_n7338_));
  OAI21X1  g04902(.A0(new_n7233_), .A1(new_n6821_), .B0(new_n7338_), .Y(new_n7339_));
  INVX1    g04903(.A(pi0954), .Y(po1110));
  AOI21X1  g04904(.A0(new_n7337_), .A1(pi0033), .B0(po1110), .Y(new_n7341_));
  OAI21X1  g04905(.A0(new_n7233_), .A1(pi0033), .B0(new_n7341_), .Y(new_n7342_));
  AND2X1   g04906(.A(new_n7342_), .B(new_n7339_), .Y(po0191));
  XOR2X1   g04907(.A(new_n6822_), .B(pi0197), .Y(new_n7344_));
  NAND2X1  g04908(.A(new_n5033_), .B(pi0162), .Y(new_n7345_));
  NAND2X1  g04909(.A(new_n7345_), .B(new_n7344_), .Y(new_n7346_));
  INVX1    g04910(.A(pi0197), .Y(new_n7347_));
  NOR4X1   g04911(.A(new_n7345_), .B(new_n7347_), .C(pi0157), .D(pi0149), .Y(new_n7348_));
  INVX1    g04912(.A(pi0162), .Y(new_n7349_));
  AOI21X1  g04913(.A0(new_n7347_), .A1(new_n7349_), .B0(new_n6824_), .Y(new_n7350_));
  NOR3X1   g04914(.A(new_n7350_), .B(new_n7348_), .C(new_n5057_), .Y(new_n7351_));
  OAI21X1  g04915(.A0(new_n7351_), .A1(new_n7344_), .B0(new_n7346_), .Y(new_n7352_));
  NOR3X1   g04916(.A(new_n7352_), .B(new_n6828_), .C(new_n5237_), .Y(new_n7353_));
  INVX1    g04917(.A(pi0167), .Y(new_n7354_));
  NOR4X1   g04918(.A(pi0468), .B(pi0332), .C(new_n5237_), .D(new_n7354_), .Y(new_n7355_));
  AOI21X1  g04919(.A0(new_n7355_), .A1(new_n6828_), .B0(new_n7353_), .Y(new_n7356_));
  NOR4X1   g04920(.A(new_n6832_), .B(new_n5057_), .C(new_n5237_), .D(new_n4036_), .Y(new_n7357_));
  NOR3X1   g04921(.A(new_n7357_), .B(new_n7353_), .C(new_n4991_), .Y(new_n7358_));
  AOI21X1  g04922(.A0(new_n7356_), .A1(new_n4991_), .B0(new_n7358_), .Y(new_n7359_));
  NAND2X1  g04923(.A(new_n7359_), .B(new_n3393_), .Y(new_n7360_));
  NAND4X1  g04924(.A(new_n6828_), .B(new_n5033_), .C(pi0232), .D(pi0167), .Y(new_n7361_));
  NOR2X1   g04925(.A(new_n7353_), .B(pi0054), .Y(new_n7362_));
  OAI21X1  g04926(.A0(new_n7361_), .A1(new_n2996_), .B0(new_n7362_), .Y(new_n7363_));
  OAI21X1  g04927(.A0(new_n7363_), .A1(pi0074), .B0(new_n7359_), .Y(new_n7364_));
  AOI21X1  g04928(.A0(new_n7364_), .A1(new_n5324_), .B0(new_n3393_), .Y(new_n7365_));
  AND2X1   g04929(.A(new_n7229_), .B(new_n6828_), .Y(new_n7366_));
  AND2X1   g04930(.A(new_n7366_), .B(new_n3135_), .Y(new_n7367_));
  INVX1    g04931(.A(new_n7367_), .Y(new_n7368_));
  AOI21X1  g04932(.A0(new_n7368_), .A1(new_n5324_), .B0(new_n3393_), .Y(new_n7369_));
  NOR2X1   g04933(.A(new_n7369_), .B(new_n7365_), .Y(new_n7370_));
  AND2X1   g04934(.A(pi0145), .B(pi0140), .Y(new_n7371_));
  NOR2X1   g04935(.A(pi0145), .B(pi0140), .Y(new_n7372_));
  NOR4X1   g04936(.A(new_n7372_), .B(new_n7371_), .C(new_n6837_), .D(new_n5057_), .Y(new_n7373_));
  XOR2X1   g04937(.A(pi0145), .B(pi0140), .Y(new_n7374_));
  OAI21X1  g04938(.A0(new_n7374_), .A1(new_n6838_), .B0(new_n2953_), .Y(new_n7375_));
  OAI21X1  g04939(.A0(new_n7375_), .A1(new_n7373_), .B0(pi0232), .Y(new_n7376_));
  AOI21X1  g04940(.A0(new_n7352_), .A1(pi0299), .B0(new_n7376_), .Y(new_n7377_));
  NOR2X1   g04941(.A(new_n7377_), .B(new_n3026_), .Y(new_n7378_));
  NOR2X1   g04942(.A(new_n7377_), .B(new_n3095_), .Y(new_n7379_));
  NOR2X1   g04943(.A(new_n7379_), .B(new_n7378_), .Y(new_n7380_));
  INVX1    g04944(.A(new_n7380_), .Y(new_n7381_));
  INVX1    g04945(.A(pi0141), .Y(new_n7382_));
  MX2X1    g04946(.A(new_n4036_), .B(new_n7382_), .S0(new_n2953_), .Y(new_n7383_));
  NOR3X1   g04947(.A(new_n7383_), .B(new_n5057_), .C(new_n5237_), .Y(new_n7384_));
  INVX1    g04948(.A(new_n7384_), .Y(new_n7385_));
  AOI21X1  g04949(.A0(new_n7385_), .A1(new_n6828_), .B0(new_n7381_), .Y(new_n7386_));
  OAI21X1  g04950(.A0(new_n7386_), .A1(new_n4991_), .B0(new_n3128_), .Y(new_n7387_));
  INVX1    g04951(.A(new_n7387_), .Y(new_n7388_));
  INVX1    g04952(.A(pi0188), .Y(new_n7389_));
  MX2X1    g04953(.A(new_n7389_), .B(new_n7354_), .S0(pi0299), .Y(new_n7390_));
  NOR3X1   g04954(.A(new_n7390_), .B(new_n5057_), .C(new_n5237_), .Y(new_n7391_));
  NOR3X1   g04955(.A(new_n7391_), .B(pi0100), .C(pi0075), .Y(new_n7392_));
  OAI21X1  g04956(.A0(new_n7392_), .A1(new_n7381_), .B0(pi0054), .Y(new_n7393_));
  INVX1    g04957(.A(new_n7393_), .Y(new_n7394_));
  OAI21X1  g04958(.A0(new_n7055_), .A1(new_n6979_), .B0(new_n2972_), .Y(new_n7395_));
  AOI21X1  g04959(.A0(new_n6978_), .A1(pi0142), .B0(pi0140), .Y(new_n7396_));
  AND2X1   g04960(.A(new_n7396_), .B(new_n7395_), .Y(new_n7397_));
  INVX1    g04961(.A(pi0140), .Y(new_n7398_));
  INVX1    g04962(.A(new_n7061_), .Y(new_n7399_));
  AOI21X1  g04963(.A0(new_n7399_), .A1(new_n7087_), .B0(pi0142), .Y(new_n7400_));
  NOR3X1   g04964(.A(new_n7064_), .B(new_n7018_), .C(new_n2972_), .Y(new_n7401_));
  NOR3X1   g04965(.A(new_n7401_), .B(new_n7400_), .C(new_n7398_), .Y(new_n7402_));
  OAI21X1  g04966(.A0(new_n7402_), .A1(new_n7397_), .B0(new_n5226_), .Y(new_n7403_));
  NAND2X1  g04967(.A(new_n7085_), .B(new_n2972_), .Y(new_n7404_));
  AOI21X1  g04968(.A0(new_n7028_), .A1(pi0142), .B0(pi0140), .Y(new_n7405_));
  AND2X1   g04969(.A(new_n7405_), .B(new_n7404_), .Y(new_n7406_));
  AND2X1   g04970(.A(new_n7024_), .B(pi0142), .Y(new_n7407_));
  AOI21X1  g04971(.A0(new_n7088_), .A1(new_n7087_), .B0(pi0142), .Y(new_n7408_));
  NOR3X1   g04972(.A(new_n7408_), .B(new_n7407_), .C(new_n7398_), .Y(new_n7409_));
  OAI21X1  g04973(.A0(new_n7409_), .A1(new_n7406_), .B0(pi0181), .Y(new_n7410_));
  NAND3X1  g04974(.A(new_n7410_), .B(new_n7403_), .C(pi0144), .Y(new_n7411_));
  OAI21X1  g04975(.A0(new_n6991_), .A1(new_n6979_), .B0(pi0142), .Y(new_n7412_));
  AOI21X1  g04976(.A0(new_n7101_), .A1(new_n2972_), .B0(pi0140), .Y(new_n7413_));
  NOR2X1   g04977(.A(new_n7064_), .B(new_n7046_), .Y(new_n7414_));
  NAND2X1  g04978(.A(new_n7414_), .B(new_n2972_), .Y(new_n7415_));
  AOI21X1  g04979(.A0(new_n7006_), .A1(pi0142), .B0(new_n7398_), .Y(new_n7416_));
  AOI22X1  g04980(.A0(new_n7416_), .A1(new_n7415_), .B0(new_n7413_), .B1(new_n7412_), .Y(new_n7417_));
  AND2X1   g04981(.A(new_n7076_), .B(new_n2972_), .Y(new_n7418_));
  NOR3X1   g04982(.A(new_n6990_), .B(new_n6989_), .C(new_n6935_), .Y(new_n7419_));
  OAI21X1  g04983(.A0(new_n7419_), .A1(new_n5057_), .B0(pi0142), .Y(new_n7420_));
  OAI21X1  g04984(.A0(new_n7420_), .A1(new_n7064_), .B0(new_n7398_), .Y(new_n7421_));
  NOR2X1   g04985(.A(new_n7079_), .B(pi0142), .Y(new_n7422_));
  OR2X1    g04986(.A(new_n7161_), .B(new_n2972_), .Y(new_n7423_));
  OAI21X1  g04987(.A0(new_n7423_), .A1(new_n7064_), .B0(pi0140), .Y(new_n7424_));
  OAI22X1  g04988(.A0(new_n7424_), .A1(new_n7422_), .B0(new_n7421_), .B1(new_n7418_), .Y(new_n7425_));
  AOI21X1  g04989(.A0(new_n7425_), .A1(new_n5226_), .B0(pi0144), .Y(new_n7426_));
  OAI21X1  g04990(.A0(new_n7417_), .A1(new_n5226_), .B0(new_n7426_), .Y(new_n7427_));
  NAND3X1  g04991(.A(new_n7427_), .B(new_n7411_), .C(new_n2953_), .Y(new_n7428_));
  AND2X1   g04992(.A(pi0299), .B(new_n5129_), .Y(new_n7429_));
  OR2X1    g04993(.A(new_n7161_), .B(new_n7160_), .Y(new_n7430_));
  OR2X1    g04994(.A(new_n7430_), .B(new_n2800_), .Y(new_n7431_));
  OR2X1    g04995(.A(new_n7158_), .B(pi0146), .Y(new_n7432_));
  AND2X1   g04996(.A(new_n7432_), .B(new_n4613_), .Y(new_n7433_));
  OR2X1    g04997(.A(new_n7163_), .B(new_n2800_), .Y(new_n7434_));
  AOI21X1  g04998(.A0(new_n7156_), .A1(new_n2800_), .B0(new_n4613_), .Y(new_n7435_));
  AOI22X1  g04999(.A0(new_n7435_), .A1(new_n7434_), .B0(new_n7433_), .B1(new_n7431_), .Y(new_n7436_));
  OAI21X1  g05000(.A0(new_n7133_), .A1(pi0161), .B0(new_n2800_), .Y(new_n7437_));
  AOI21X1  g05001(.A0(new_n7131_), .A1(pi0161), .B0(new_n7437_), .Y(new_n7438_));
  NOR2X1   g05002(.A(new_n7136_), .B(pi0161), .Y(new_n7439_));
  OAI21X1  g05003(.A0(new_n7114_), .A1(new_n4613_), .B0(pi0146), .Y(new_n7440_));
  NOR2X1   g05004(.A(new_n7109_), .B(pi0162), .Y(new_n7441_));
  OAI21X1  g05005(.A0(new_n7440_), .A1(new_n7439_), .B0(new_n7441_), .Y(new_n7442_));
  OAI22X1  g05006(.A0(new_n7442_), .A1(new_n7438_), .B0(new_n7436_), .B1(new_n7349_), .Y(new_n7443_));
  AND2X1   g05007(.A(new_n7121_), .B(new_n2800_), .Y(new_n7444_));
  OAI21X1  g05008(.A0(new_n7117_), .A1(new_n2800_), .B0(pi0161), .Y(new_n7445_));
  OAI21X1  g05009(.A0(new_n7111_), .A1(new_n7109_), .B0(pi0146), .Y(new_n7446_));
  OAI21X1  g05010(.A0(new_n7125_), .A1(new_n7109_), .B0(new_n2800_), .Y(new_n7447_));
  NAND3X1  g05011(.A(new_n7447_), .B(new_n7446_), .C(new_n4613_), .Y(new_n7448_));
  AND2X1   g05012(.A(new_n7448_), .B(new_n7349_), .Y(new_n7449_));
  OAI21X1  g05013(.A0(new_n7445_), .A1(new_n7444_), .B0(new_n7449_), .Y(new_n7450_));
  NOR2X1   g05014(.A(new_n7152_), .B(pi0146), .Y(new_n7451_));
  OAI21X1  g05015(.A0(new_n7148_), .A1(new_n2800_), .B0(new_n4613_), .Y(new_n7452_));
  OR2X1    g05016(.A(new_n7452_), .B(new_n7451_), .Y(new_n7453_));
  OAI21X1  g05017(.A0(new_n7109_), .A1(new_n7023_), .B0(pi0146), .Y(new_n7454_));
  AOI21X1  g05018(.A0(new_n7151_), .A1(new_n2800_), .B0(new_n4613_), .Y(new_n7455_));
  AOI21X1  g05019(.A0(new_n7455_), .A1(new_n7454_), .B0(new_n7349_), .Y(new_n7456_));
  AND2X1   g05020(.A(pi0299), .B(pi0159), .Y(new_n7457_));
  INVX1    g05021(.A(new_n7457_), .Y(new_n7458_));
  AOI21X1  g05022(.A0(new_n7456_), .A1(new_n7453_), .B0(new_n7458_), .Y(new_n7459_));
  AOI22X1  g05023(.A0(new_n7459_), .A1(new_n7450_), .B0(new_n7443_), .B1(new_n7429_), .Y(new_n7460_));
  AOI21X1  g05024(.A0(new_n7460_), .A1(new_n7428_), .B0(new_n5237_), .Y(new_n7461_));
  OAI21X1  g05025(.A0(new_n7461_), .A1(new_n7172_), .B0(new_n3065_), .Y(new_n7462_));
  AND2X1   g05026(.A(new_n6924_), .B(pi0144), .Y(new_n7463_));
  NOR2X1   g05027(.A(pi0299), .B(pi0177), .Y(new_n7464_));
  INVX1    g05028(.A(new_n6916_), .Y(new_n7465_));
  AOI21X1  g05029(.A0(new_n6888_), .A1(new_n6896_), .B0(pi0144), .Y(new_n7466_));
  NAND2X1  g05030(.A(new_n7466_), .B(new_n7465_), .Y(new_n7467_));
  NAND2X1  g05031(.A(new_n7467_), .B(new_n7464_), .Y(new_n7468_));
  INVX1    g05032(.A(pi0177), .Y(new_n7469_));
  OAI21X1  g05033(.A0(new_n6890_), .A1(new_n6896_), .B0(new_n6888_), .Y(new_n7470_));
  OR4X1    g05034(.A(new_n7470_), .B(new_n7466_), .C(pi0299), .D(new_n7469_), .Y(new_n7471_));
  OAI21X1  g05035(.A0(new_n7468_), .A1(new_n7463_), .B0(new_n7471_), .Y(new_n7472_));
  AOI21X1  g05036(.A0(new_n7472_), .A1(pi0232), .B0(new_n6926_), .Y(new_n7473_));
  INVX1    g05037(.A(new_n6902_), .Y(new_n7474_));
  NOR3X1   g05038(.A(new_n7474_), .B(new_n5057_), .C(pi0161), .Y(new_n7475_));
  OAI21X1  g05039(.A0(new_n7475_), .A1(new_n6899_), .B0(new_n6893_), .Y(new_n7476_));
  NOR2X1   g05040(.A(pi0155), .B(pi0038), .Y(new_n7477_));
  AND2X1   g05041(.A(new_n7477_), .B(new_n6895_), .Y(new_n7478_));
  NOR2X1   g05042(.A(new_n6908_), .B(new_n4613_), .Y(new_n7479_));
  NOR3X1   g05043(.A(new_n7479_), .B(new_n6905_), .C(new_n6896_), .Y(new_n7480_));
  AND2X1   g05044(.A(pi0155), .B(new_n2996_), .Y(new_n7481_));
  INVX1    g05045(.A(new_n7481_), .Y(new_n7482_));
  NOR3X1   g05046(.A(new_n7482_), .B(new_n7480_), .C(new_n6922_), .Y(new_n7483_));
  AOI21X1  g05047(.A0(new_n7478_), .A1(new_n7476_), .B0(new_n7483_), .Y(new_n7484_));
  OAI22X1  g05048(.A0(new_n7484_), .A1(new_n5237_), .B0(new_n7473_), .B1(pi0038), .Y(new_n7485_));
  AOI21X1  g05049(.A0(new_n3000_), .A1(new_n2959_), .B0(new_n6862_), .Y(new_n7486_));
  INVX1    g05050(.A(new_n7486_), .Y(new_n7487_));
  OAI21X1  g05051(.A0(new_n7487_), .A1(new_n7389_), .B0(new_n7354_), .Y(new_n7488_));
  INVX1    g05052(.A(new_n6856_), .Y(new_n7489_));
  NOR2X1   g05053(.A(new_n6855_), .B(new_n6857_), .Y(new_n7490_));
  NOR3X1   g05054(.A(new_n7490_), .B(new_n7389_), .C(new_n7354_), .Y(new_n7491_));
  AOI21X1  g05055(.A0(new_n7489_), .A1(new_n7389_), .B0(new_n7491_), .Y(new_n7492_));
  AOI21X1  g05056(.A0(new_n7492_), .A1(new_n7488_), .B0(new_n2996_), .Y(new_n7493_));
  OR2X1    g05057(.A(new_n7493_), .B(pi0087), .Y(new_n7494_));
  AOI21X1  g05058(.A0(new_n7485_), .A1(pi0039), .B0(new_n7494_), .Y(new_n7495_));
  INVX1    g05059(.A(new_n7391_), .Y(new_n7496_));
  MX2X1    g05060(.A(new_n7496_), .B(new_n6870_), .S0(new_n2996_), .Y(new_n7497_));
  OAI21X1  g05061(.A0(new_n7497_), .A1(new_n3156_), .B0(new_n3026_), .Y(new_n7498_));
  AOI21X1  g05062(.A0(new_n7495_), .A1(new_n7462_), .B0(new_n7498_), .Y(new_n7499_));
  OAI21X1  g05063(.A0(new_n7499_), .A1(new_n7378_), .B0(new_n3105_), .Y(new_n7500_));
  INVX1    g05064(.A(new_n7378_), .Y(new_n7501_));
  NOR3X1   g05065(.A(new_n6878_), .B(new_n7188_), .C(pi0095), .Y(new_n7502_));
  MX2X1    g05066(.A(pi0177), .B(pi0155), .S0(pi0299), .Y(new_n7503_));
  OAI21X1  g05067(.A0(new_n7503_), .A1(pi0038), .B0(new_n5930_), .Y(new_n7504_));
  AOI21X1  g05068(.A0(new_n7504_), .A1(new_n7502_), .B0(new_n7497_), .Y(new_n7505_));
  OAI21X1  g05069(.A0(new_n7505_), .A1(pi0100), .B0(new_n7501_), .Y(new_n7506_));
  AOI21X1  g05070(.A0(new_n7506_), .A1(new_n7185_), .B0(new_n7379_), .Y(new_n7507_));
  AOI21X1  g05071(.A0(new_n7507_), .A1(new_n7500_), .B0(pi0054), .Y(new_n7508_));
  OAI21X1  g05072(.A0(new_n7508_), .A1(new_n7394_), .B0(new_n4991_), .Y(new_n7509_));
  NOR2X1   g05073(.A(new_n7358_), .B(new_n3128_), .Y(new_n7510_));
  INVX1    g05074(.A(new_n7510_), .Y(new_n7511_));
  AND2X1   g05075(.A(new_n7356_), .B(pi0054), .Y(new_n7512_));
  INVX1    g05076(.A(new_n7512_), .Y(new_n7513_));
  OAI21X1  g05077(.A0(new_n7363_), .A1(new_n7366_), .B0(new_n5107_), .Y(new_n7514_));
  OAI21X1  g05078(.A0(new_n7352_), .A1(new_n5237_), .B0(pi0100), .Y(new_n7515_));
  INVX1    g05079(.A(new_n7355_), .Y(new_n7516_));
  AOI21X1  g05080(.A0(new_n7345_), .A1(new_n7502_), .B0(new_n7230_), .Y(new_n7517_));
  OR4X1    g05081(.A(new_n6878_), .B(new_n7188_), .C(pi0232), .D(pi0095), .Y(new_n7518_));
  OAI21X1  g05082(.A0(new_n7517_), .A1(pi0100), .B0(new_n7518_), .Y(new_n7519_));
  OAI21X1  g05083(.A0(new_n7516_), .A1(new_n2996_), .B0(new_n7519_), .Y(new_n7520_));
  AOI21X1  g05084(.A0(new_n7520_), .A1(new_n7515_), .B0(pi0075), .Y(new_n7521_));
  OAI21X1  g05085(.A0(new_n7352_), .A1(new_n5237_), .B0(pi0075), .Y(new_n7522_));
  NAND2X1  g05086(.A(new_n7522_), .B(new_n3100_), .Y(new_n7523_));
  OAI21X1  g05087(.A0(new_n7523_), .A1(new_n7521_), .B0(new_n7514_), .Y(new_n7524_));
  AOI21X1  g05088(.A0(new_n7524_), .A1(new_n7513_), .B0(pi0074), .Y(new_n7525_));
  OAI21X1  g05089(.A0(new_n7525_), .A1(new_n7511_), .B0(new_n3148_), .Y(new_n7526_));
  AOI21X1  g05090(.A0(new_n7509_), .A1(new_n7388_), .B0(new_n7526_), .Y(new_n7527_));
  OAI21X1  g05091(.A0(new_n7527_), .A1(new_n7370_), .B0(new_n7360_), .Y(new_n7528_));
  AOI21X1  g05092(.A0(new_n7273_), .A1(new_n7270_), .B0(pi0146), .Y(new_n7529_));
  OAI21X1  g05093(.A0(new_n7292_), .A1(new_n2800_), .B0(new_n4613_), .Y(new_n7530_));
  NAND4X1  g05094(.A(new_n7282_), .B(new_n7273_), .C(pi0161), .D(new_n2800_), .Y(new_n7531_));
  OAI21X1  g05095(.A0(new_n7530_), .A1(new_n7529_), .B0(new_n7531_), .Y(new_n7532_));
  AOI21X1  g05096(.A0(new_n7295_), .A1(new_n7349_), .B0(new_n7458_), .Y(new_n7533_));
  OAI21X1  g05097(.A0(new_n7533_), .A1(new_n7429_), .B0(new_n7345_), .Y(new_n7534_));
  NOR2X1   g05098(.A(new_n7264_), .B(new_n5196_), .Y(new_n7535_));
  NAND2X1  g05099(.A(new_n7261_), .B(new_n2800_), .Y(new_n7536_));
  AOI21X1  g05100(.A0(new_n7536_), .A1(new_n7535_), .B0(pi0161), .Y(new_n7537_));
  NAND2X1  g05101(.A(new_n7279_), .B(new_n2800_), .Y(new_n7538_));
  AOI21X1  g05102(.A0(new_n7538_), .A1(new_n7303_), .B0(new_n4613_), .Y(new_n7539_));
  AND2X1   g05103(.A(new_n2901_), .B(pi0159), .Y(new_n7540_));
  OR4X1    g05104(.A(new_n7540_), .B(new_n7539_), .C(new_n7537_), .D(new_n2953_), .Y(new_n7541_));
  AOI22X1  g05105(.A0(new_n7541_), .A1(new_n7534_), .B0(new_n7532_), .B1(new_n7349_), .Y(new_n7542_));
  AOI21X1  g05106(.A0(new_n7292_), .A1(pi0142), .B0(pi0140), .Y(new_n7543_));
  OAI21X1  g05107(.A0(new_n7275_), .A1(pi0142), .B0(new_n7543_), .Y(new_n7544_));
  NOR3X1   g05108(.A(new_n7264_), .B(new_n5220_), .C(new_n7398_), .Y(new_n7545_));
  OAI21X1  g05109(.A0(new_n7262_), .A1(pi0142), .B0(new_n7545_), .Y(new_n7546_));
  AOI21X1  g05110(.A0(new_n7546_), .A1(new_n7544_), .B0(pi0144), .Y(new_n7547_));
  INVX1    g05111(.A(pi0144), .Y(new_n7548_));
  NOR2X1   g05112(.A(new_n7288_), .B(new_n5220_), .Y(new_n7549_));
  AOI21X1  g05113(.A0(new_n7283_), .A1(new_n2972_), .B0(pi0140), .Y(new_n7550_));
  AOI21X1  g05114(.A0(new_n7279_), .A1(new_n2972_), .B0(new_n7398_), .Y(new_n7551_));
  AOI21X1  g05115(.A0(new_n7551_), .A1(new_n7549_), .B0(new_n7550_), .Y(new_n7552_));
  OAI22X1  g05116(.A0(new_n7552_), .A1(new_n7548_), .B0(new_n5033_), .B1(new_n7398_), .Y(new_n7553_));
  NOR2X1   g05117(.A(new_n7553_), .B(new_n7547_), .Y(new_n7554_));
  OAI21X1  g05118(.A0(new_n7296_), .A1(new_n5226_), .B0(new_n2953_), .Y(new_n7555_));
  OAI21X1  g05119(.A0(new_n7555_), .A1(new_n7554_), .B0(pi0232), .Y(new_n7556_));
  OAI21X1  g05120(.A0(new_n7556_), .A1(new_n7542_), .B0(new_n3065_), .Y(new_n7557_));
  NOR2X1   g05121(.A(new_n7241_), .B(new_n4613_), .Y(new_n7558_));
  OAI21X1  g05122(.A0(new_n7235_), .A1(pi0161), .B0(new_n6893_), .Y(new_n7559_));
  OR2X1    g05123(.A(new_n7559_), .B(new_n7558_), .Y(new_n7560_));
  NAND4X1  g05124(.A(new_n6893_), .B(new_n5261_), .C(new_n6906_), .D(new_n4613_), .Y(new_n7561_));
  AOI22X1  g05125(.A0(new_n7561_), .A1(new_n7477_), .B0(new_n7560_), .B1(new_n7481_), .Y(new_n7562_));
  OR4X1    g05126(.A(new_n6913_), .B(new_n5257_), .C(new_n6914_), .D(pi0144), .Y(new_n7563_));
  AND2X1   g05127(.A(new_n2953_), .B(pi0177), .Y(new_n7564_));
  INVX1    g05128(.A(new_n7564_), .Y(new_n7565_));
  AOI21X1  g05129(.A0(new_n7248_), .A1(pi0144), .B0(new_n7565_), .Y(new_n7566_));
  OAI21X1  g05130(.A0(new_n7245_), .A1(pi0144), .B0(new_n7464_), .Y(new_n7567_));
  NAND2X1  g05131(.A(new_n7567_), .B(pi0232), .Y(new_n7568_));
  AOI21X1  g05132(.A0(new_n7566_), .A1(new_n7563_), .B0(new_n7568_), .Y(new_n7569_));
  OAI22X1  g05133(.A0(new_n7569_), .A1(pi0038), .B0(new_n7562_), .B1(new_n2953_), .Y(new_n7570_));
  AOI21X1  g05134(.A0(new_n7570_), .A1(pi0039), .B0(new_n7493_), .Y(new_n7571_));
  AOI21X1  g05135(.A0(new_n7571_), .A1(new_n7557_), .B0(pi0100), .Y(new_n7572_));
  OAI21X1  g05136(.A0(new_n7572_), .A1(new_n7378_), .B0(new_n3156_), .Y(new_n7573_));
  OAI21X1  g05137(.A0(new_n7496_), .A1(new_n2996_), .B0(new_n3026_), .Y(new_n7574_));
  OAI21X1  g05138(.A0(new_n7377_), .A1(new_n3026_), .B0(new_n7574_), .Y(new_n7575_));
  AND2X1   g05139(.A(new_n7575_), .B(pi0087), .Y(new_n7576_));
  INVX1    g05140(.A(new_n7576_), .Y(new_n7577_));
  AOI21X1  g05141(.A0(new_n7577_), .A1(new_n7573_), .B0(new_n5315_), .Y(new_n7578_));
  OR2X1    g05142(.A(new_n7390_), .B(new_n2996_), .Y(new_n7579_));
  NAND3X1  g05143(.A(new_n7503_), .B(new_n3065_), .C(new_n3000_), .Y(new_n7580_));
  AOI21X1  g05144(.A0(new_n7580_), .A1(new_n7579_), .B0(new_n6855_), .Y(new_n7581_));
  OAI21X1  g05145(.A0(new_n7581_), .A1(pi0100), .B0(new_n7501_), .Y(new_n7582_));
  AOI21X1  g05146(.A0(new_n7582_), .A1(new_n3156_), .B0(new_n7576_), .Y(new_n7583_));
  OAI22X1  g05147(.A0(new_n7583_), .A1(new_n7186_), .B0(new_n7377_), .B1(new_n3095_), .Y(new_n7584_));
  OAI21X1  g05148(.A0(new_n7584_), .A1(new_n7578_), .B0(new_n3112_), .Y(new_n7585_));
  AOI21X1  g05149(.A0(new_n7585_), .A1(new_n7393_), .B0(pi0074), .Y(new_n7586_));
  INVX1    g05150(.A(new_n7362_), .Y(new_n7587_));
  NAND4X1  g05151(.A(new_n7320_), .B(new_n7299_), .C(pi0162), .D(new_n3100_), .Y(new_n7588_));
  OAI22X1  g05152(.A0(new_n7588_), .A1(new_n5448_), .B0(new_n7516_), .B1(new_n2996_), .Y(new_n7589_));
  AOI21X1  g05153(.A0(new_n7589_), .A1(new_n6828_), .B0(new_n7587_), .Y(new_n7590_));
  OAI21X1  g05154(.A0(new_n7590_), .A1(new_n7512_), .B0(new_n4991_), .Y(new_n7591_));
  AOI21X1  g05155(.A0(new_n7591_), .A1(new_n7510_), .B0(new_n5324_), .Y(new_n7592_));
  OAI21X1  g05156(.A0(new_n7586_), .A1(new_n7387_), .B0(new_n7592_), .Y(new_n7593_));
  AOI22X1  g05157(.A0(new_n7593_), .A1(new_n7365_), .B0(new_n7359_), .B1(new_n3393_), .Y(new_n7594_));
  NOR2X1   g05158(.A(pi0954), .B(pi0033), .Y(new_n7595_));
  AOI21X1  g05159(.A0(new_n7594_), .A1(pi0034), .B0(new_n7595_), .Y(new_n7596_));
  OAI21X1  g05160(.A0(new_n7528_), .A1(pi0034), .B0(new_n7596_), .Y(new_n7597_));
  INVX1    g05161(.A(pi0034), .Y(new_n7598_));
  AND2X1   g05162(.A(new_n6819_), .B(new_n7598_), .Y(new_n7599_));
  OR2X1    g05163(.A(pi0954), .B(pi0033), .Y(new_n7600_));
  AOI21X1  g05164(.A0(new_n7599_), .A1(new_n7594_), .B0(new_n7600_), .Y(new_n7601_));
  OAI21X1  g05165(.A0(new_n7599_), .A1(new_n7528_), .B0(new_n7601_), .Y(new_n7602_));
  AND2X1   g05166(.A(new_n7602_), .B(new_n7597_), .Y(po0192));
  NOR3X1   g05167(.A(new_n6807_), .B(new_n6805_), .C(pi0051), .Y(new_n7604_));
  INVX1    g05168(.A(new_n7604_), .Y(new_n7605_));
  AND2X1   g05169(.A(pi0252), .B(new_n2453_), .Y(new_n7606_));
  NOR4X1   g05170(.A(new_n2756_), .B(new_n2722_), .C(new_n2780_), .D(pi0833), .Y(new_n7607_));
  NOR3X1   g05171(.A(new_n7607_), .B(new_n5252_), .C(new_n5251_), .Y(new_n7608_));
  INVX1    g05172(.A(new_n7608_), .Y(new_n7609_));
  NOR2X1   g05173(.A(new_n5094_), .B(new_n3053_), .Y(new_n7610_));
  OAI21X1  g05174(.A0(new_n7609_), .A1(new_n5088_), .B0(new_n7610_), .Y(new_n7611_));
  NAND2X1  g05175(.A(new_n6417_), .B(pi0142), .Y(new_n7612_));
  OAI21X1  g05176(.A0(new_n6420_), .A1(new_n2800_), .B0(new_n7612_), .Y(new_n7613_));
  OR2X1    g05177(.A(new_n7613_), .B(new_n5929_), .Y(new_n7614_));
  AOI21X1  g05178(.A0(new_n7614_), .A1(new_n7611_), .B0(new_n5970_), .Y(new_n7615_));
  NAND3X1  g05179(.A(new_n7611_), .B(new_n6763_), .C(new_n5083_), .Y(new_n7616_));
  OAI21X1  g05180(.A0(new_n7615_), .A1(new_n7606_), .B0(new_n7616_), .Y(new_n7617_));
  AOI22X1  g05181(.A0(new_n7617_), .A1(new_n6761_), .B0(new_n6759_), .B1(pi0137), .Y(new_n7618_));
  NOR3X1   g05182(.A(new_n7618_), .B(new_n3066_), .C(new_n3026_), .Y(new_n7619_));
  AOI21X1  g05183(.A0(new_n4999_), .A1(new_n2701_), .B0(pi0093), .Y(new_n7620_));
  OAI21X1  g05184(.A0(new_n7620_), .A1(new_n5012_), .B0(new_n2518_), .Y(new_n7621_));
  AOI21X1  g05185(.A0(new_n2727_), .A1(pi0035), .B0(new_n6792_), .Y(new_n7622_));
  NAND2X1  g05186(.A(new_n7622_), .B(new_n7621_), .Y(new_n7623_));
  OR2X1    g05187(.A(pi0093), .B(new_n2456_), .Y(new_n7624_));
  NOR4X1   g05188(.A(new_n7624_), .B(new_n5020_), .C(pi0090), .D(pi0024), .Y(new_n7625_));
  NAND3X1  g05189(.A(new_n7625_), .B(new_n2550_), .C(new_n2726_), .Y(new_n7626_));
  OAI21X1  g05190(.A0(new_n7623_), .A1(pi0032), .B0(new_n7626_), .Y(new_n7627_));
  NAND3X1  g05191(.A(new_n7627_), .B(new_n7169_), .C(new_n2540_), .Y(new_n7628_));
  NAND2X1  g05192(.A(new_n7621_), .B(new_n5019_), .Y(new_n7629_));
  AND2X1   g05193(.A(new_n5971_), .B(new_n2723_), .Y(new_n7630_));
  AOI21X1  g05194(.A0(new_n7169_), .A1(new_n2453_), .B0(new_n6077_), .Y(new_n7631_));
  NOR2X1   g05195(.A(po0740), .B(pi0122), .Y(new_n7632_));
  AOI21X1  g05196(.A0(new_n7169_), .A1(new_n2453_), .B0(new_n6633_), .Y(new_n7633_));
  AOI22X1  g05197(.A0(new_n7633_), .A1(new_n7632_), .B0(new_n7631_), .B1(new_n7630_), .Y(new_n7634_));
  NAND2X1  g05198(.A(new_n7634_), .B(new_n7629_), .Y(new_n7635_));
  NOR4X1   g05199(.A(new_n6790_), .B(new_n6789_), .C(new_n2492_), .D(new_n2476_), .Y(new_n7636_));
  OR2X1    g05200(.A(new_n7636_), .B(new_n7621_), .Y(new_n7637_));
  NAND4X1  g05201(.A(new_n7637_), .B(new_n7635_), .C(new_n7622_), .D(new_n7271_), .Y(new_n7638_));
  NAND2X1  g05202(.A(new_n2545_), .B(pi0040), .Y(new_n7639_));
  NAND2X1  g05203(.A(new_n7623_), .B(new_n7639_), .Y(new_n7640_));
  AND2X1   g05204(.A(new_n7271_), .B(pi1082), .Y(new_n7641_));
  AOI21X1  g05205(.A0(new_n7641_), .A1(new_n7640_), .B0(pi0038), .Y(new_n7642_));
  NAND3X1  g05206(.A(new_n7642_), .B(new_n7638_), .C(new_n7628_), .Y(new_n7643_));
  OR2X1    g05207(.A(pi0100), .B(pi0039), .Y(new_n7644_));
  AOI21X1  g05208(.A0(new_n7605_), .A1(pi0038), .B0(new_n7644_), .Y(new_n7645_));
  AOI21X1  g05209(.A0(new_n7645_), .A1(new_n7643_), .B0(new_n7619_), .Y(new_n7646_));
  NOR3X1   g05210(.A(po0840), .B(new_n6809_), .C(new_n2453_), .Y(new_n7647_));
  OAI21X1  g05211(.A0(new_n7647_), .A1(new_n6810_), .B0(new_n6811_), .Y(new_n7648_));
  OAI22X1  g05212(.A0(new_n7648_), .A1(new_n7605_), .B0(new_n7646_), .B1(new_n3101_), .Y(new_n7649_));
  AOI21X1  g05213(.A0(new_n7649_), .A1(new_n3100_), .B0(pi0054), .Y(new_n7650_));
  AOI21X1  g05214(.A0(new_n5817_), .A1(new_n5787_), .B0(new_n3112_), .Y(new_n7651_));
  OR4X1    g05215(.A(new_n7651_), .B(new_n7650_), .C(new_n6755_), .D(new_n5324_), .Y(new_n7652_));
  NOR4X1   g05216(.A(new_n7605_), .B(new_n5324_), .C(new_n3131_), .D(pi0055), .Y(new_n7653_));
  OAI21X1  g05217(.A0(new_n7653_), .A1(new_n3153_), .B0(new_n2436_), .Y(new_n7654_));
  AOI21X1  g05218(.A0(new_n7652_), .A1(new_n3153_), .B0(new_n7654_), .Y(po0193));
  NOR2X1   g05219(.A(new_n2582_), .B(new_n2506_), .Y(new_n7656_));
  INVX1    g05220(.A(new_n7656_), .Y(new_n7657_));
  INVX1    g05221(.A(pi0069), .Y(new_n7658_));
  AND2X1   g05222(.A(new_n2660_), .B(new_n2614_), .Y(new_n7659_));
  NOR4X1   g05223(.A(new_n6872_), .B(new_n2472_), .C(new_n2577_), .D(pi0065), .Y(new_n7660_));
  NOR4X1   g05224(.A(pi0103), .B(pi0071), .C(pi0067), .D(new_n2658_), .Y(new_n7661_));
  NAND4X1  g05225(.A(new_n7661_), .B(new_n7660_), .C(new_n7659_), .D(new_n7658_), .Y(new_n7662_));
  NOR2X1   g05226(.A(new_n7662_), .B(new_n7657_), .Y(new_n7663_));
  NOR4X1   g05227(.A(new_n3255_), .B(new_n2530_), .C(pi0058), .D(pi0024), .Y(new_n7664_));
  NOR2X1   g05228(.A(new_n7664_), .B(new_n7663_), .Y(new_n7665_));
  INVX1    g05229(.A(new_n5189_), .Y(new_n7666_));
  NOR4X1   g05230(.A(new_n7666_), .B(new_n2544_), .C(new_n2492_), .D(pi0035), .Y(new_n7667_));
  NOR4X1   g05231(.A(po1038), .B(new_n5843_), .C(new_n3136_), .D(pi0092), .Y(new_n7668_));
  AND2X1   g05232(.A(new_n7668_), .B(new_n7667_), .Y(new_n7669_));
  INVX1    g05233(.A(new_n7669_), .Y(new_n7670_));
  NOR3X1   g05234(.A(new_n7670_), .B(new_n7665_), .C(new_n5922_), .Y(po0194));
  INVX1    g05235(.A(new_n2551_), .Y(new_n7672_));
  NAND2X1  g05236(.A(new_n3002_), .B(new_n2959_), .Y(new_n7673_));
  NOR3X1   g05237(.A(new_n7673_), .B(new_n7672_), .C(new_n5787_), .Y(new_n7674_));
  INVX1    g05238(.A(new_n7674_), .Y(new_n7675_));
  OR4X1    g05239(.A(new_n2472_), .B(new_n2466_), .C(pi0104), .D(pi0071), .Y(new_n7676_));
  OR4X1    g05240(.A(pi0073), .B(pi0066), .C(pi0049), .D(pi0045), .Y(new_n7677_));
  OR2X1    g05241(.A(pi0065), .B(pi0048), .Y(new_n7678_));
  OR4X1    g05242(.A(new_n7678_), .B(new_n2635_), .C(pi0084), .D(pi0082), .Y(new_n7679_));
  NOR4X1   g05243(.A(new_n7679_), .B(new_n7677_), .C(new_n7676_), .D(new_n6947_), .Y(new_n7680_));
  AOI21X1  g05244(.A0(new_n7680_), .A1(pi0332), .B0(pi0064), .Y(new_n7681_));
  NAND4X1  g05245(.A(new_n5189_), .B(new_n2541_), .C(new_n2512_), .D(new_n2519_), .Y(new_n7682_));
  NOR2X1   g05246(.A(new_n7682_), .B(new_n2544_), .Y(new_n7683_));
  NAND4X1  g05247(.A(new_n7683_), .B(new_n2460_), .C(new_n2726_), .D(new_n2959_), .Y(new_n7684_));
  NOR4X1   g05248(.A(new_n7684_), .B(new_n7681_), .C(new_n2608_), .D(pi0081), .Y(new_n7685_));
  AND2X1   g05249(.A(new_n6520_), .B(new_n3129_), .Y(new_n7686_));
  OAI21X1  g05250(.A0(new_n7685_), .A1(pi0038), .B0(new_n7686_), .Y(new_n7687_));
  AOI21X1  g05251(.A0(new_n7675_), .A1(pi0038), .B0(new_n7687_), .Y(po0196));
  AND2X1   g05252(.A(new_n7686_), .B(new_n2996_), .Y(new_n7689_));
  INVX1    g05253(.A(new_n7689_), .Y(new_n7690_));
  NOR2X1   g05254(.A(new_n5037_), .B(new_n5034_), .Y(new_n7691_));
  INVX1    g05255(.A(new_n7691_), .Y(new_n7692_));
  OR2X1    g05256(.A(new_n2783_), .B(pi0984), .Y(new_n7693_));
  AOI21X1  g05257(.A0(new_n7693_), .A1(pi0835), .B0(new_n5037_), .Y(new_n7694_));
  NOR4X1   g05258(.A(new_n7694_), .B(new_n5043_), .C(new_n5041_), .D(new_n2756_), .Y(new_n7695_));
  NOR4X1   g05259(.A(new_n7695_), .B(new_n5243_), .C(new_n7692_), .D(pi0223), .Y(new_n7696_));
  NOR2X1   g05260(.A(new_n5043_), .B(new_n5041_), .Y(new_n7697_));
  INVX1    g05261(.A(new_n7697_), .Y(new_n7698_));
  NOR3X1   g05262(.A(new_n7694_), .B(new_n6270_), .C(new_n7698_), .Y(new_n7699_));
  NOR4X1   g05263(.A(new_n7699_), .B(new_n5243_), .C(new_n5051_), .D(new_n7692_), .Y(new_n7700_));
  NOR4X1   g05264(.A(new_n7694_), .B(new_n5052_), .C(new_n5043_), .D(new_n5041_), .Y(new_n7701_));
  NOR4X1   g05265(.A(new_n7701_), .B(new_n5243_), .C(new_n5050_), .D(new_n7692_), .Y(new_n7702_));
  NOR4X1   g05266(.A(new_n7702_), .B(new_n7700_), .C(new_n7696_), .D(pi0299), .Y(new_n7703_));
  INVX1    g05267(.A(pi0786), .Y(new_n7704_));
  NOR4X1   g05268(.A(new_n7695_), .B(new_n5243_), .C(new_n7692_), .D(pi0215), .Y(new_n7705_));
  OR4X1    g05269(.A(new_n7699_), .B(new_n5243_), .C(new_n5071_), .D(new_n7692_), .Y(new_n7706_));
  NOR4X1   g05270(.A(new_n7701_), .B(new_n5243_), .C(new_n5070_), .D(new_n7692_), .Y(new_n7707_));
  NOR2X1   g05271(.A(new_n7707_), .B(new_n2953_), .Y(new_n7708_));
  AND2X1   g05272(.A(new_n7708_), .B(new_n7706_), .Y(new_n7709_));
  INVX1    g05273(.A(new_n7709_), .Y(new_n7710_));
  OAI22X1  g05274(.A0(new_n7710_), .A1(new_n7705_), .B0(pi1082), .B1(new_n7704_), .Y(new_n7711_));
  INVX1    g05275(.A(pi1082), .Y(new_n7712_));
  INVX1    g05276(.A(new_n4898_), .Y(new_n7713_));
  OAI22X1  g05277(.A0(new_n5074_), .A1(new_n7713_), .B0(new_n5058_), .B1(new_n4781_), .Y(new_n7714_));
  NAND4X1  g05278(.A(new_n7714_), .B(po0740), .C(new_n7712_), .D(pi0786), .Y(new_n7715_));
  OR4X1    g05279(.A(new_n7715_), .B(new_n5245_), .C(new_n3074_), .D(pi0287), .Y(new_n7716_));
  OAI21X1  g05280(.A0(new_n7711_), .A1(new_n7703_), .B0(new_n7716_), .Y(new_n7717_));
  NOR2X1   g05281(.A(pi0095), .B(pi0039), .Y(new_n7718_));
  AOI21X1  g05282(.A0(new_n2583_), .A1(pi0108), .B0(new_n2504_), .Y(new_n7719_));
  OR4X1    g05283(.A(new_n6780_), .B(new_n6778_), .C(new_n2463_), .D(pi0111), .Y(new_n7720_));
  OR4X1    g05284(.A(pi0084), .B(pi0081), .C(pi0066), .D(pi0064), .Y(new_n7721_));
  OR2X1    g05285(.A(pi0069), .B(pi0065), .Y(new_n7722_));
  NOR2X1   g05286(.A(new_n7722_), .B(new_n7721_), .Y(new_n7723_));
  INVX1    g05287(.A(new_n7723_), .Y(new_n7724_));
  INVX1    g05288(.A(pi0045), .Y(new_n7725_));
  NOR4X1   g05289(.A(pi0082), .B(pi0068), .C(pi0049), .D(new_n2629_), .Y(new_n7726_));
  NAND3X1  g05290(.A(new_n7726_), .B(new_n6948_), .C(new_n7725_), .Y(new_n7727_));
  OR4X1    g05291(.A(new_n7727_), .B(new_n7724_), .C(new_n7720_), .D(new_n7676_), .Y(new_n7728_));
  NAND4X1  g05292(.A(new_n2497_), .B(new_n2475_), .C(new_n2726_), .D(new_n2880_), .Y(new_n7729_));
  NOR2X1   g05293(.A(new_n7729_), .B(new_n7728_), .Y(new_n7730_));
  NAND2X1  g05294(.A(new_n2503_), .B(pi0108), .Y(new_n7731_));
  OAI21X1  g05295(.A0(new_n7731_), .A1(new_n2583_), .B0(new_n2567_), .Y(new_n7732_));
  AOI21X1  g05296(.A0(new_n7730_), .A1(new_n7719_), .B0(new_n7732_), .Y(new_n7733_));
  INVX1    g05297(.A(pi0314), .Y(new_n7734_));
  OR2X1    g05298(.A(po0740), .B(pi0986), .Y(new_n7735_));
  AND2X1   g05299(.A(new_n7735_), .B(pi0252), .Y(new_n7736_));
  OR4X1    g05300(.A(new_n7736_), .B(new_n2570_), .C(new_n5007_), .D(new_n7734_), .Y(new_n7737_));
  NOR3X1   g05301(.A(new_n7728_), .B(pi0841), .C(pi0047), .Y(new_n7738_));
  AOI21X1  g05302(.A0(new_n2568_), .A1(pi0047), .B0(new_n7738_), .Y(new_n7739_));
  NOR3X1   g05303(.A(new_n5007_), .B(new_n2511_), .C(new_n2478_), .Y(new_n7740_));
  OAI21X1  g05304(.A0(new_n7736_), .A1(new_n7734_), .B0(new_n7740_), .Y(new_n7741_));
  OAI22X1  g05305(.A0(new_n7741_), .A1(new_n7739_), .B0(new_n7737_), .B1(new_n7733_), .Y(new_n7742_));
  AOI21X1  g05306(.A0(new_n7742_), .A1(new_n2491_), .B0(pi0035), .Y(new_n7743_));
  AOI21X1  g05307(.A0(new_n5194_), .A1(pi0035), .B0(new_n2544_), .Y(new_n7744_));
  NAND2X1  g05308(.A(new_n7744_), .B(new_n2715_), .Y(new_n7745_));
  OAI22X1  g05309(.A0(new_n7745_), .A1(new_n7743_), .B0(new_n5195_), .B1(new_n7169_), .Y(new_n7746_));
  AOI22X1  g05310(.A0(new_n7746_), .A1(new_n7718_), .B0(new_n7717_), .B1(pi0039), .Y(new_n7747_));
  NOR2X1   g05311(.A(new_n7747_), .B(new_n7690_), .Y(po0197));
  INVX1    g05312(.A(new_n7668_), .Y(new_n7749_));
  OAI21X1  g05313(.A0(new_n2545_), .A1(new_n2549_), .B0(new_n7271_), .Y(new_n7750_));
  INVX1    g05314(.A(new_n7750_), .Y(new_n7751_));
  INVX1    g05315(.A(new_n2512_), .Y(new_n7752_));
  OR4X1    g05316(.A(new_n2520_), .B(new_n2459_), .C(new_n2578_), .D(pi0093), .Y(new_n7753_));
  NOR4X1   g05317(.A(new_n7753_), .B(new_n6998_), .C(new_n7752_), .D(new_n2527_), .Y(new_n7754_));
  OR2X1    g05318(.A(new_n7754_), .B(pi0040), .Y(new_n7755_));
  AOI21X1  g05319(.A0(new_n7755_), .A1(new_n7751_), .B0(pi1082), .Y(new_n7756_));
  AOI21X1  g05320(.A0(new_n7754_), .A1(new_n5189_), .B0(new_n7712_), .Y(new_n7757_));
  NOR3X1   g05321(.A(new_n7757_), .B(new_n7756_), .C(new_n7749_), .Y(po0198));
  NOR2X1   g05322(.A(pi0072), .B(pi0041), .Y(new_n7759_));
  NOR2X1   g05323(.A(new_n7759_), .B(new_n6291_), .Y(new_n7760_));
  INVX1    g05324(.A(new_n6291_), .Y(new_n7761_));
  AOI21X1  g05325(.A0(new_n7759_), .A1(new_n2724_), .B0(new_n7761_), .Y(new_n7762_));
  INVX1    g05326(.A(new_n7762_), .Y(new_n7763_));
  INVX1    g05327(.A(new_n5932_), .Y(new_n7764_));
  OR4X1    g05328(.A(new_n3003_), .B(new_n2555_), .C(pi0101), .D(pi0044), .Y(new_n7765_));
  NOR2X1   g05329(.A(new_n7765_), .B(new_n5972_), .Y(new_n7766_));
  INVX1    g05330(.A(new_n7766_), .Y(new_n7767_));
  OAI21X1  g05331(.A0(new_n7767_), .A1(new_n7764_), .B0(pi0041), .Y(new_n7768_));
  OAI21X1  g05332(.A0(new_n2548_), .A1(pi0041), .B0(new_n2723_), .Y(new_n7769_));
  INVX1    g05333(.A(pi0099), .Y(new_n7770_));
  NAND2X1  g05334(.A(new_n5092_), .B(new_n7770_), .Y(new_n7771_));
  AOI21X1  g05335(.A0(pi0101), .A1(new_n2548_), .B0(pi0041), .Y(new_n7772_));
  INVX1    g05336(.A(new_n7772_), .Y(new_n7773_));
  NOR4X1   g05337(.A(new_n2487_), .B(new_n2484_), .C(new_n2480_), .D(pi0024), .Y(new_n7774_));
  NAND4X1  g05338(.A(new_n7774_), .B(new_n5971_), .C(new_n5189_), .D(pi0252), .Y(new_n7775_));
  NOR3X1   g05339(.A(new_n7775_), .B(new_n7773_), .C(pi0044), .Y(new_n7776_));
  AOI21X1  g05340(.A0(new_n7776_), .A1(new_n7771_), .B0(new_n7769_), .Y(new_n7777_));
  AOI21X1  g05341(.A0(new_n7777_), .A1(new_n7768_), .B0(new_n7763_), .Y(new_n7778_));
  OAI21X1  g05342(.A0(new_n7778_), .A1(new_n7760_), .B0(new_n2959_), .Y(new_n7779_));
  NOR3X1   g05343(.A(pi0468), .B(pi0332), .C(pi0189), .Y(new_n7780_));
  AND2X1   g05344(.A(new_n7780_), .B(pi0144), .Y(new_n7781_));
  AOI21X1  g05345(.A0(new_n7781_), .A1(new_n7008_), .B0(pi0299), .Y(new_n7782_));
  NOR3X1   g05346(.A(pi0468), .B(pi0332), .C(pi0166), .Y(new_n7783_));
  INVX1    g05347(.A(new_n7783_), .Y(new_n7784_));
  NOR3X1   g05348(.A(new_n7784_), .B(new_n4613_), .C(pi0152), .Y(new_n7785_));
  OAI21X1  g05349(.A0(new_n7785_), .A1(new_n6417_), .B0(pi0232), .Y(new_n7786_));
  NOR2X1   g05350(.A(new_n7786_), .B(new_n7782_), .Y(new_n7787_));
  INVX1    g05351(.A(new_n7787_), .Y(new_n7788_));
  AOI21X1  g05352(.A0(new_n7788_), .A1(new_n2548_), .B0(new_n2959_), .Y(new_n7789_));
  NOR2X1   g05353(.A(new_n7789_), .B(new_n5788_), .Y(new_n7790_));
  NOR2X1   g05354(.A(new_n7759_), .B(pi0039), .Y(new_n7791_));
  NOR2X1   g05355(.A(new_n7791_), .B(new_n7789_), .Y(new_n7792_));
  INVX1    g05356(.A(new_n7792_), .Y(new_n7793_));
  OAI21X1  g05357(.A0(new_n7793_), .A1(new_n3108_), .B0(pi0075), .Y(new_n7794_));
  AOI21X1  g05358(.A0(new_n7790_), .A1(new_n7779_), .B0(new_n7794_), .Y(new_n7795_));
  NOR2X1   g05359(.A(new_n5911_), .B(new_n5910_), .Y(new_n7796_));
  NAND2X1  g05360(.A(new_n5919_), .B(new_n2756_), .Y(new_n7797_));
  AOI21X1  g05361(.A0(new_n5918_), .A1(new_n7796_), .B0(new_n7797_), .Y(new_n7798_));
  NOR2X1   g05362(.A(new_n7798_), .B(pi0044), .Y(new_n7799_));
  OR4X1    g05363(.A(new_n5917_), .B(new_n5910_), .C(new_n3256_), .D(pi0096), .Y(new_n7800_));
  NOR2X1   g05364(.A(new_n5906_), .B(new_n2748_), .Y(new_n7801_));
  AOI21X1  g05365(.A0(new_n7801_), .A1(new_n2743_), .B0(new_n5943_), .Y(new_n7802_));
  OAI21X1  g05366(.A0(new_n7802_), .A1(new_n2520_), .B0(new_n5899_), .Y(new_n7803_));
  AOI21X1  g05367(.A0(new_n7803_), .A1(new_n5897_), .B0(pi0051), .Y(new_n7804_));
  OAI21X1  g05368(.A0(new_n7804_), .A1(new_n2869_), .B0(new_n2526_), .Y(new_n7805_));
  AOI21X1  g05369(.A0(new_n5915_), .A1(pi0096), .B0(new_n7666_), .Y(new_n7806_));
  NAND4X1  g05370(.A(new_n7806_), .B(new_n7805_), .C(new_n5917_), .D(new_n2548_), .Y(new_n7807_));
  NAND2X1  g05371(.A(new_n7807_), .B(new_n7800_), .Y(new_n7808_));
  OAI21X1  g05372(.A0(new_n7808_), .A1(new_n2756_), .B0(new_n7799_), .Y(new_n7809_));
  OAI21X1  g05373(.A0(new_n7809_), .A1(pi0101), .B0(pi0041), .Y(new_n7810_));
  INVX1    g05374(.A(pi0101), .Y(new_n7811_));
  NOR3X1   g05375(.A(new_n5917_), .B(new_n7796_), .C(pi0072), .Y(new_n7812_));
  NOR3X1   g05376(.A(new_n5916_), .B(new_n5914_), .C(new_n7666_), .Y(new_n7813_));
  NOR3X1   g05377(.A(new_n7813_), .B(new_n5918_), .C(pi0072), .Y(new_n7814_));
  NOR3X1   g05378(.A(new_n7814_), .B(new_n7812_), .C(pi1093), .Y(new_n7815_));
  NAND3X1  g05379(.A(new_n7807_), .B(new_n7800_), .C(new_n2548_), .Y(new_n7816_));
  AOI21X1  g05380(.A0(new_n7816_), .A1(pi1093), .B0(new_n7815_), .Y(new_n7817_));
  MX2X1    g05381(.A(new_n7817_), .B(new_n2548_), .S0(pi0044), .Y(new_n7818_));
  AOI21X1  g05382(.A0(new_n7818_), .A1(new_n7811_), .B0(new_n7773_), .Y(new_n7819_));
  NOR2X1   g05383(.A(new_n7819_), .B(new_n2724_), .Y(new_n7820_));
  NOR3X1   g05384(.A(new_n7815_), .B(new_n7796_), .C(pi0072), .Y(new_n7821_));
  MX2X1    g05385(.A(new_n7821_), .B(new_n2548_), .S0(pi0044), .Y(new_n7822_));
  AOI21X1  g05386(.A0(new_n7822_), .A1(new_n7811_), .B0(new_n7773_), .Y(new_n7823_));
  INVX1    g05387(.A(pi0041), .Y(new_n7824_));
  NOR2X1   g05388(.A(new_n7796_), .B(new_n2756_), .Y(new_n7825_));
  NOR4X1   g05389(.A(new_n7825_), .B(new_n7798_), .C(pi0101), .D(pi0044), .Y(new_n7826_));
  OAI21X1  g05390(.A0(new_n7826_), .A1(new_n7824_), .B0(new_n2724_), .Y(new_n7827_));
  OAI21X1  g05391(.A0(new_n7827_), .A1(new_n7823_), .B0(pi0228), .Y(new_n7828_));
  AOI21X1  g05392(.A0(new_n7820_), .A1(new_n7810_), .B0(new_n7828_), .Y(new_n7829_));
  INVX1    g05393(.A(pi0480), .Y(new_n7830_));
  AND2X1   g05394(.A(pi0949), .B(new_n7830_), .Y(new_n7831_));
  NAND3X1  g05395(.A(new_n2594_), .B(new_n2505_), .C(new_n2502_), .Y(new_n7832_));
  OR4X1    g05396(.A(new_n7832_), .B(new_n7831_), .C(new_n2485_), .D(new_n2492_), .Y(new_n7833_));
  NOR4X1   g05397(.A(pi0109), .B(pi0108), .C(pi0097), .D(pi0046), .Y(new_n7834_));
  NAND4X1  g05398(.A(new_n7834_), .B(new_n2597_), .C(pi0094), .D(new_n2474_), .Y(new_n7835_));
  NAND2X1  g05399(.A(new_n7835_), .B(new_n2482_), .Y(new_n7836_));
  NAND2X1  g05400(.A(new_n7831_), .B(new_n2486_), .Y(new_n7837_));
  NOR4X1   g05401(.A(new_n7837_), .B(new_n2566_), .C(new_n5007_), .D(pi0047), .Y(new_n7838_));
  INVX1    g05402(.A(pi0959), .Y(new_n7839_));
  NAND2X1  g05403(.A(new_n7839_), .B(pi0901), .Y(new_n7840_));
  AOI21X1  g05404(.A0(new_n7838_), .A1(new_n7836_), .B0(new_n7840_), .Y(new_n7841_));
  INVX1    g05405(.A(new_n2483_), .Y(new_n7842_));
  NOR4X1   g05406(.A(new_n7842_), .B(new_n2480_), .C(new_n2482_), .D(pi0109), .Y(new_n7843_));
  INVX1    g05407(.A(new_n7843_), .Y(new_n7844_));
  OAI21X1  g05408(.A0(new_n7844_), .A1(new_n7837_), .B0(new_n7840_), .Y(new_n7845_));
  INVX1    g05409(.A(pi0250), .Y(new_n7846_));
  AND2X1   g05410(.A(pi0252), .B(new_n7846_), .Y(new_n7847_));
  NAND3X1  g05411(.A(new_n7847_), .B(new_n7845_), .C(new_n5189_), .Y(new_n7848_));
  AOI21X1  g05412(.A0(new_n7841_), .A1(new_n7833_), .B0(new_n7848_), .Y(new_n7849_));
  AND2X1   g05413(.A(new_n7843_), .B(new_n7667_), .Y(new_n7850_));
  INVX1    g05414(.A(new_n7847_), .Y(new_n7851_));
  AND2X1   g05415(.A(new_n7851_), .B(new_n7831_), .Y(new_n7852_));
  AOI22X1  g05416(.A0(new_n7852_), .A1(new_n7850_), .B0(new_n7849_), .B1(new_n2548_), .Y(new_n7853_));
  OR2X1    g05417(.A(new_n7853_), .B(pi0044), .Y(new_n7854_));
  OR2X1    g05418(.A(new_n7854_), .B(pi0101), .Y(new_n7855_));
  NOR4X1   g05419(.A(new_n7847_), .B(new_n7844_), .C(new_n7837_), .D(new_n7666_), .Y(new_n7856_));
  NOR3X1   g05420(.A(new_n7856_), .B(new_n7849_), .C(pi0072), .Y(new_n7857_));
  MX2X1    g05421(.A(new_n7857_), .B(new_n2548_), .S0(pi0044), .Y(new_n7858_));
  AOI21X1  g05422(.A0(new_n7858_), .A1(new_n7811_), .B0(new_n7773_), .Y(new_n7859_));
  AOI21X1  g05423(.A0(new_n7855_), .A1(pi0041), .B0(new_n7859_), .Y(new_n7860_));
  OAI21X1  g05424(.A0(new_n7860_), .A1(pi0228), .B0(new_n2959_), .Y(new_n7861_));
  INVX1    g05425(.A(pi0287), .Y(new_n7862_));
  NOR3X1   g05426(.A(new_n3003_), .B(new_n2555_), .C(new_n7862_), .Y(new_n7863_));
  MX2X1    g05427(.A(new_n7863_), .B(new_n2548_), .S0(new_n7788_), .Y(new_n7864_));
  AOI21X1  g05428(.A0(new_n7864_), .A1(pi0039), .B0(new_n5792_), .Y(new_n7865_));
  OAI21X1  g05429(.A0(new_n7861_), .A1(new_n7829_), .B0(new_n7865_), .Y(new_n7866_));
  INVX1    g05430(.A(new_n7789_), .Y(new_n7867_));
  INVX1    g05431(.A(pi0044), .Y(new_n7868_));
  NAND4X1  g05432(.A(new_n5189_), .B(new_n2486_), .C(new_n2550_), .D(new_n7868_), .Y(new_n7869_));
  NOR2X1   g05433(.A(new_n7869_), .B(new_n7773_), .Y(new_n7870_));
  AOI21X1  g05434(.A0(pi0072), .A1(new_n7824_), .B0(new_n7870_), .Y(new_n7871_));
  AOI21X1  g05435(.A0(new_n5972_), .A1(new_n2548_), .B0(new_n7871_), .Y(new_n7872_));
  AND2X1   g05436(.A(new_n7771_), .B(new_n2723_), .Y(new_n7873_));
  INVX1    g05437(.A(new_n7873_), .Y(new_n7874_));
  AOI22X1  g05438(.A0(new_n7874_), .A1(new_n7769_), .B0(new_n7872_), .B1(new_n7771_), .Y(new_n7875_));
  OAI21X1  g05439(.A0(new_n7766_), .A1(new_n7824_), .B0(new_n7875_), .Y(new_n7876_));
  AOI21X1  g05440(.A0(new_n7876_), .A1(new_n7762_), .B0(new_n7760_), .Y(new_n7877_));
  OAI21X1  g05441(.A0(new_n7877_), .A1(pi0039), .B0(new_n7867_), .Y(new_n7878_));
  OAI21X1  g05442(.A0(new_n7792_), .A1(new_n2996_), .B0(new_n3156_), .Y(new_n7879_));
  AOI21X1  g05443(.A0(new_n7878_), .A1(new_n5085_), .B0(new_n7879_), .Y(new_n7880_));
  NAND2X1  g05444(.A(new_n7765_), .B(pi0041), .Y(new_n7881_));
  NAND3X1  g05445(.A(new_n7881_), .B(new_n7871_), .C(pi0228), .Y(new_n7882_));
  AOI21X1  g05446(.A0(new_n7759_), .A1(new_n3013_), .B0(new_n3157_), .Y(new_n7883_));
  AOI21X1  g05447(.A0(new_n7791_), .A1(new_n5792_), .B0(new_n3156_), .Y(new_n7884_));
  NAND2X1  g05448(.A(new_n7884_), .B(new_n7867_), .Y(new_n7885_));
  AOI21X1  g05449(.A0(new_n7883_), .A1(new_n7882_), .B0(new_n7885_), .Y(new_n7886_));
  OR2X1    g05450(.A(new_n7886_), .B(pi0075), .Y(new_n7887_));
  AOI21X1  g05451(.A0(new_n7880_), .A1(new_n7866_), .B0(new_n7887_), .Y(new_n7888_));
  OAI21X1  g05452(.A0(new_n7888_), .A1(new_n7795_), .B0(new_n5893_), .Y(new_n7889_));
  AOI21X1  g05453(.A0(new_n7793_), .A1(new_n6309_), .B0(po1038), .Y(new_n7890_));
  AND2X1   g05454(.A(pi0232), .B(pi0039), .Y(new_n7891_));
  INVX1    g05455(.A(new_n7891_), .Y(new_n7892_));
  NOR4X1   g05456(.A(new_n7892_), .B(new_n7784_), .C(new_n4613_), .D(pi0152), .Y(new_n7893_));
  NOR4X1   g05457(.A(new_n7893_), .B(new_n7791_), .C(new_n6520_), .D(pi0072), .Y(new_n7894_));
  AOI21X1  g05458(.A0(new_n7890_), .A1(new_n7889_), .B0(new_n7894_), .Y(po0199));
  AND2X1   g05459(.A(pi0208), .B(pi0207), .Y(new_n7896_));
  INVX1    g05460(.A(new_n7896_), .Y(new_n7897_));
  INVX1    g05461(.A(pi0115), .Y(new_n7898_));
  AND2X1   g05462(.A(new_n2723_), .B(new_n7898_), .Y(new_n7899_));
  INVX1    g05463(.A(pi0042), .Y(new_n7900_));
  OR2X1    g05464(.A(pi0114), .B(new_n7900_), .Y(new_n7901_));
  NOR2X1   g05465(.A(pi0099), .B(pi0041), .Y(new_n7902_));
  INVX1    g05466(.A(new_n7902_), .Y(new_n7903_));
  AOI22X1  g05467(.A0(new_n7819_), .A1(new_n7770_), .B0(new_n7903_), .B1(pi0072), .Y(new_n7904_));
  MX2X1    g05468(.A(new_n7904_), .B(new_n2548_), .S0(pi0113), .Y(new_n7905_));
  MX2X1    g05469(.A(new_n7905_), .B(new_n2548_), .S0(pi0116), .Y(new_n7906_));
  INVX1    g05470(.A(pi0114), .Y(new_n7907_));
  AOI21X1  g05471(.A0(new_n2548_), .A1(pi0042), .B0(new_n7907_), .Y(new_n7908_));
  OR2X1    g05472(.A(pi0116), .B(pi0113), .Y(new_n7909_));
  NOR4X1   g05473(.A(new_n7809_), .B(new_n7909_), .C(new_n7903_), .D(pi0101), .Y(new_n7910_));
  INVX1    g05474(.A(new_n7910_), .Y(new_n7911_));
  AOI21X1  g05475(.A0(new_n7911_), .A1(new_n7900_), .B0(new_n7908_), .Y(new_n7912_));
  OAI21X1  g05476(.A0(new_n7906_), .A1(new_n7901_), .B0(new_n7912_), .Y(new_n7913_));
  AND2X1   g05477(.A(new_n7913_), .B(new_n7899_), .Y(new_n7914_));
  INVX1    g05478(.A(new_n7908_), .Y(new_n7915_));
  NOR2X1   g05479(.A(new_n2723_), .B(pi0115), .Y(new_n7916_));
  INVX1    g05480(.A(new_n7916_), .Y(new_n7917_));
  AOI22X1  g05481(.A0(new_n7823_), .A1(new_n7770_), .B0(new_n7903_), .B1(pi0072), .Y(new_n7918_));
  MX2X1    g05482(.A(new_n7918_), .B(new_n2548_), .S0(pi0113), .Y(new_n7919_));
  MX2X1    g05483(.A(new_n7919_), .B(new_n2548_), .S0(pi0116), .Y(new_n7920_));
  INVX1    g05484(.A(new_n7920_), .Y(new_n7921_));
  INVX1    g05485(.A(new_n7826_), .Y(new_n7922_));
  NOR3X1   g05486(.A(new_n7922_), .B(new_n7909_), .C(new_n7903_), .Y(new_n7923_));
  AOI21X1  g05487(.A0(new_n7923_), .A1(new_n7900_), .B0(pi0114), .Y(new_n7924_));
  OAI21X1  g05488(.A0(new_n7921_), .A1(new_n7900_), .B0(new_n7924_), .Y(new_n7925_));
  AOI21X1  g05489(.A0(new_n7925_), .A1(new_n7915_), .B0(new_n7917_), .Y(new_n7926_));
  AOI21X1  g05490(.A0(new_n2548_), .A1(pi0042), .B0(new_n7898_), .Y(new_n7927_));
  NOR4X1   g05491(.A(new_n7927_), .B(new_n7926_), .C(new_n7914_), .D(new_n3013_), .Y(new_n7928_));
  AOI22X1  g05492(.A0(new_n7859_), .A1(new_n7770_), .B0(new_n7903_), .B1(pi0072), .Y(new_n7929_));
  MX2X1    g05493(.A(new_n7929_), .B(new_n2548_), .S0(pi0113), .Y(new_n7930_));
  MX2X1    g05494(.A(new_n7930_), .B(new_n2548_), .S0(pi0116), .Y(new_n7931_));
  NOR4X1   g05495(.A(new_n7855_), .B(new_n7903_), .C(pi0116), .D(pi0113), .Y(new_n7932_));
  OR2X1    g05496(.A(new_n7932_), .B(pi0042), .Y(new_n7933_));
  AND2X1   g05497(.A(new_n7933_), .B(new_n7915_), .Y(new_n7934_));
  OAI21X1  g05498(.A0(new_n7931_), .A1(new_n7901_), .B0(new_n7934_), .Y(new_n7935_));
  AND2X1   g05499(.A(new_n7935_), .B(new_n7898_), .Y(new_n7936_));
  NOR3X1   g05500(.A(new_n7936_), .B(new_n7927_), .C(pi0228), .Y(new_n7937_));
  NOR2X1   g05501(.A(new_n7937_), .B(pi0039), .Y(new_n7938_));
  INVX1    g05502(.A(new_n7938_), .Y(new_n7939_));
  NOR2X1   g05503(.A(new_n7939_), .B(new_n7928_), .Y(new_n7940_));
  INVX1    g05504(.A(pi0199), .Y(new_n7941_));
  INVX1    g05505(.A(pi0189), .Y(new_n7942_));
  NOR2X1   g05506(.A(new_n7780_), .B(pi0072), .Y(new_n7943_));
  NOR4X1   g05507(.A(new_n5057_), .B(new_n3003_), .C(new_n2555_), .D(new_n7862_), .Y(new_n7944_));
  AOI21X1  g05508(.A0(new_n7944_), .A1(new_n7942_), .B0(new_n7943_), .Y(new_n7945_));
  AND2X1   g05509(.A(new_n2953_), .B(pi0232), .Y(new_n7946_));
  OAI21X1  g05510(.A0(new_n7945_), .A1(new_n7941_), .B0(new_n7946_), .Y(new_n7947_));
  NOR4X1   g05511(.A(new_n7784_), .B(new_n3003_), .C(new_n2555_), .D(new_n7862_), .Y(new_n7948_));
  AOI21X1  g05512(.A0(new_n5930_), .A1(new_n4464_), .B0(pi0072), .Y(new_n7949_));
  NOR4X1   g05513(.A(new_n7949_), .B(new_n7948_), .C(new_n2953_), .D(new_n5237_), .Y(new_n7950_));
  AOI21X1  g05514(.A0(pi0199), .A1(new_n2548_), .B0(pi0232), .Y(new_n7951_));
  OAI21X1  g05515(.A0(pi0232), .A1(new_n2548_), .B0(pi0299), .Y(new_n7952_));
  AND2X1   g05516(.A(new_n7952_), .B(new_n7951_), .Y(new_n7953_));
  NOR2X1   g05517(.A(new_n7953_), .B(new_n7950_), .Y(new_n7954_));
  AOI21X1  g05518(.A0(new_n7954_), .A1(new_n7947_), .B0(new_n2959_), .Y(new_n7955_));
  OAI21X1  g05519(.A0(new_n7955_), .A1(new_n7940_), .B0(new_n3277_), .Y(new_n7956_));
  AND2X1   g05520(.A(new_n2548_), .B(pi0042), .Y(new_n7957_));
  NOR2X1   g05521(.A(new_n7957_), .B(new_n6291_), .Y(new_n7958_));
  INVX1    g05522(.A(new_n7957_), .Y(new_n7959_));
  OAI21X1  g05523(.A0(new_n7959_), .A1(new_n7899_), .B0(new_n6291_), .Y(new_n7960_));
  NOR4X1   g05524(.A(new_n7908_), .B(new_n2829_), .C(new_n2722_), .D(pi0115), .Y(new_n7961_));
  NOR3X1   g05525(.A(pi0052), .B(pi0043), .C(pi0042), .Y(new_n7962_));
  NOR4X1   g05526(.A(new_n7765_), .B(new_n5972_), .C(new_n7909_), .D(new_n7903_), .Y(new_n7963_));
  INVX1    g05527(.A(new_n7963_), .Y(new_n7964_));
  OR4X1    g05528(.A(new_n7964_), .B(new_n7962_), .C(pi0114), .D(pi0042), .Y(new_n7965_));
  NOR3X1   g05529(.A(new_n7869_), .B(new_n7909_), .C(new_n5090_), .Y(new_n7966_));
  INVX1    g05530(.A(new_n7966_), .Y(new_n7967_));
  OAI21X1  g05531(.A0(new_n7967_), .A1(new_n5972_), .B0(new_n2548_), .Y(new_n7968_));
  OR2X1    g05532(.A(new_n7968_), .B(new_n7900_), .Y(new_n7969_));
  NAND3X1  g05533(.A(new_n7969_), .B(new_n7965_), .C(new_n7907_), .Y(new_n7970_));
  AOI21X1  g05534(.A0(new_n7970_), .A1(new_n7961_), .B0(new_n7960_), .Y(new_n7971_));
  OAI21X1  g05535(.A0(new_n7971_), .A1(new_n7958_), .B0(new_n2959_), .Y(new_n7972_));
  NOR2X1   g05536(.A(new_n7951_), .B(pi0299), .Y(new_n7973_));
  NOR3X1   g05537(.A(new_n7780_), .B(new_n7941_), .C(pi0072), .Y(new_n7974_));
  OAI21X1  g05538(.A0(new_n7974_), .A1(new_n5237_), .B0(new_n7973_), .Y(new_n7975_));
  AOI21X1  g05539(.A0(new_n7949_), .A1(pi0299), .B0(new_n2959_), .Y(new_n7976_));
  AND2X1   g05540(.A(new_n7976_), .B(new_n7975_), .Y(new_n7977_));
  INVX1    g05541(.A(new_n7977_), .Y(new_n7978_));
  AOI21X1  g05542(.A0(new_n7978_), .A1(new_n7972_), .B0(new_n5086_), .Y(new_n7979_));
  AOI22X1  g05543(.A0(new_n7976_), .A1(new_n7975_), .B0(new_n7959_), .B1(new_n2959_), .Y(new_n7980_));
  OAI21X1  g05544(.A0(new_n7980_), .A1(new_n2996_), .B0(new_n3156_), .Y(new_n7981_));
  NOR2X1   g05545(.A(new_n7981_), .B(new_n7979_), .Y(new_n7982_));
  NOR4X1   g05546(.A(new_n7765_), .B(new_n7909_), .C(new_n7903_), .D(new_n3013_), .Y(new_n7983_));
  AND2X1   g05547(.A(new_n7983_), .B(new_n7898_), .Y(new_n7984_));
  AND2X1   g05548(.A(new_n7984_), .B(new_n7907_), .Y(new_n7985_));
  NOR4X1   g05549(.A(new_n7869_), .B(new_n5091_), .C(new_n5090_), .D(new_n3013_), .Y(new_n7986_));
  OAI21X1  g05550(.A0(new_n7986_), .A1(new_n7959_), .B0(new_n3085_), .Y(new_n7987_));
  AOI21X1  g05551(.A0(new_n7985_), .A1(new_n7900_), .B0(new_n7987_), .Y(new_n7988_));
  OAI21X1  g05552(.A0(pi0072), .A1(new_n7900_), .B0(new_n2959_), .Y(new_n7989_));
  OAI21X1  g05553(.A0(new_n7989_), .A1(new_n3277_), .B0(pi0087), .Y(new_n7990_));
  NOR3X1   g05554(.A(new_n7990_), .B(new_n7988_), .C(new_n7977_), .Y(new_n7991_));
  OR2X1    g05555(.A(new_n7991_), .B(pi0075), .Y(new_n7992_));
  AOI21X1  g05556(.A0(new_n7982_), .A1(new_n7956_), .B0(new_n7992_), .Y(new_n7993_));
  INVX1    g05557(.A(new_n7899_), .Y(new_n7994_));
  NOR4X1   g05558(.A(new_n7964_), .B(new_n7764_), .C(new_n7962_), .D(pi0114), .Y(new_n7995_));
  OR4X1    g05559(.A(new_n7775_), .B(new_n5090_), .C(pi0113), .D(pi0044), .Y(new_n7996_));
  OAI21X1  g05560(.A0(new_n7996_), .A1(pi0116), .B0(new_n7957_), .Y(new_n7997_));
  NAND2X1  g05561(.A(new_n7997_), .B(new_n7907_), .Y(new_n7998_));
  AOI21X1  g05562(.A0(new_n7995_), .A1(new_n7900_), .B0(new_n7998_), .Y(new_n7999_));
  NOR3X1   g05563(.A(new_n7999_), .B(new_n7908_), .C(new_n7994_), .Y(new_n8000_));
  NOR2X1   g05564(.A(new_n7958_), .B(new_n5788_), .Y(new_n8001_));
  OAI21X1  g05565(.A0(new_n8000_), .A1(new_n7960_), .B0(new_n8001_), .Y(new_n8002_));
  AOI21X1  g05566(.A0(new_n7957_), .A1(new_n5788_), .B0(pi0039), .Y(new_n8003_));
  AOI21X1  g05567(.A0(new_n8003_), .A1(new_n8002_), .B0(new_n7977_), .Y(new_n8004_));
  OAI21X1  g05568(.A0(new_n8004_), .A1(new_n3095_), .B0(new_n5893_), .Y(new_n8005_));
  OAI21X1  g05569(.A0(new_n8005_), .A1(new_n7993_), .B0(new_n7897_), .Y(new_n8006_));
  AOI21X1  g05570(.A0(pi0200), .A1(new_n2548_), .B0(pi0232), .Y(new_n8007_));
  NOR2X1   g05571(.A(new_n8007_), .B(pi0299), .Y(new_n8008_));
  INVX1    g05572(.A(pi0200), .Y(new_n8009_));
  NOR3X1   g05573(.A(new_n7780_), .B(new_n8009_), .C(pi0072), .Y(new_n8010_));
  OAI21X1  g05574(.A0(new_n8010_), .A1(new_n5237_), .B0(new_n8008_), .Y(new_n8011_));
  AND2X1   g05575(.A(new_n8011_), .B(pi0039), .Y(new_n8012_));
  AOI22X1  g05576(.A0(new_n8012_), .A1(new_n7975_), .B0(new_n7959_), .B1(new_n2959_), .Y(new_n8013_));
  AOI21X1  g05577(.A0(new_n8013_), .A1(new_n6309_), .B0(new_n7897_), .Y(new_n8014_));
  OR2X1    g05578(.A(new_n7945_), .B(new_n7941_), .Y(new_n8015_));
  OR2X1    g05579(.A(new_n7945_), .B(new_n8009_), .Y(new_n8016_));
  NAND4X1  g05580(.A(new_n8016_), .B(new_n8015_), .C(new_n2953_), .D(pi0232), .Y(new_n8017_));
  OR2X1    g05581(.A(new_n8009_), .B(pi0072), .Y(new_n8018_));
  AOI21X1  g05582(.A0(new_n8018_), .A1(new_n7953_), .B0(new_n7950_), .Y(new_n8019_));
  AOI21X1  g05583(.A0(new_n8019_), .A1(new_n8017_), .B0(new_n2959_), .Y(new_n8020_));
  OAI21X1  g05584(.A0(new_n8020_), .A1(new_n7940_), .B0(new_n3277_), .Y(new_n8021_));
  INVX1    g05585(.A(new_n8012_), .Y(new_n8022_));
  OAI21X1  g05586(.A0(new_n8022_), .A1(new_n7978_), .B0(new_n7972_), .Y(new_n8023_));
  OAI21X1  g05587(.A0(new_n8013_), .A1(new_n2996_), .B0(new_n3156_), .Y(new_n8024_));
  AOI22X1  g05588(.A0(new_n8024_), .A1(new_n7981_), .B0(new_n8023_), .B1(new_n5085_), .Y(new_n8025_));
  AND2X1   g05589(.A(new_n8012_), .B(new_n7977_), .Y(new_n8026_));
  OR2X1    g05590(.A(new_n8026_), .B(new_n7990_), .Y(new_n8027_));
  OAI21X1  g05591(.A0(new_n8027_), .A1(new_n7988_), .B0(new_n3095_), .Y(new_n8028_));
  AOI21X1  g05592(.A0(new_n8025_), .A1(new_n8021_), .B0(new_n8028_), .Y(new_n8029_));
  AOI21X1  g05593(.A0(new_n8003_), .A1(new_n8002_), .B0(new_n8026_), .Y(new_n8030_));
  OAI21X1  g05594(.A0(new_n8030_), .A1(new_n3095_), .B0(new_n5893_), .Y(new_n8031_));
  OAI21X1  g05595(.A0(new_n8031_), .A1(new_n8029_), .B0(new_n8014_), .Y(new_n8032_));
  AND2X1   g05596(.A(pi0214), .B(pi0211), .Y(new_n8033_));
  AOI21X1  g05597(.A0(new_n8033_), .A1(pi0212), .B0(pi0219), .Y(new_n8034_));
  AND2X1   g05598(.A(new_n7980_), .B(new_n6309_), .Y(new_n8035_));
  OR2X1    g05599(.A(new_n8035_), .B(new_n8034_), .Y(new_n8036_));
  AOI21X1  g05600(.A0(new_n8032_), .A1(new_n8006_), .B0(new_n8036_), .Y(new_n8037_));
  INVX1    g05601(.A(new_n8034_), .Y(new_n8038_));
  INVX1    g05602(.A(new_n7940_), .Y(new_n8039_));
  INVX1    g05603(.A(new_n7973_), .Y(new_n8040_));
  AND2X1   g05604(.A(new_n8015_), .B(pi0232), .Y(new_n8041_));
  OAI21X1  g05605(.A0(new_n8041_), .A1(new_n8040_), .B0(pi0039), .Y(new_n8042_));
  AOI21X1  g05606(.A0(new_n8042_), .A1(new_n8039_), .B0(new_n5792_), .Y(new_n8043_));
  AND2X1   g05607(.A(new_n7975_), .B(pi0039), .Y(new_n8044_));
  INVX1    g05608(.A(new_n8044_), .Y(new_n8045_));
  AOI21X1  g05609(.A0(new_n8045_), .A1(new_n7972_), .B0(new_n5086_), .Y(new_n8046_));
  AOI21X1  g05610(.A0(new_n7959_), .A1(new_n2959_), .B0(new_n8044_), .Y(new_n8047_));
  OAI21X1  g05611(.A0(new_n8047_), .A1(new_n2996_), .B0(new_n3156_), .Y(new_n8048_));
  OR2X1    g05612(.A(new_n8048_), .B(new_n8046_), .Y(new_n8049_));
  NOR2X1   g05613(.A(new_n7990_), .B(new_n7988_), .Y(new_n8050_));
  AOI21X1  g05614(.A0(new_n8045_), .A1(new_n8050_), .B0(pi0075), .Y(new_n8051_));
  OAI21X1  g05615(.A0(new_n8049_), .A1(new_n8043_), .B0(new_n8051_), .Y(new_n8052_));
  AND2X1   g05616(.A(new_n8003_), .B(new_n8002_), .Y(new_n8053_));
  OAI21X1  g05617(.A0(new_n8044_), .A1(new_n8053_), .B0(pi0075), .Y(new_n8054_));
  NAND3X1  g05618(.A(new_n8054_), .B(new_n8052_), .C(new_n5893_), .Y(new_n8055_));
  AOI21X1  g05619(.A0(new_n8047_), .A1(new_n6309_), .B0(new_n7896_), .Y(new_n8056_));
  NOR2X1   g05620(.A(new_n8008_), .B(new_n7973_), .Y(new_n8057_));
  AOI21X1  g05621(.A0(new_n8016_), .A1(new_n8041_), .B0(new_n8057_), .Y(new_n8058_));
  OR2X1    g05622(.A(new_n8058_), .B(new_n2959_), .Y(new_n8059_));
  AOI21X1  g05623(.A0(new_n8059_), .A1(new_n8039_), .B0(new_n5792_), .Y(new_n8060_));
  AND2X1   g05624(.A(new_n8012_), .B(new_n7975_), .Y(new_n8061_));
  INVX1    g05625(.A(new_n8061_), .Y(new_n8062_));
  AOI21X1  g05626(.A0(new_n8062_), .A1(new_n7972_), .B0(new_n5086_), .Y(new_n8063_));
  OR2X1    g05627(.A(new_n8063_), .B(new_n8024_), .Y(new_n8064_));
  AOI21X1  g05628(.A0(new_n8062_), .A1(new_n8050_), .B0(pi0075), .Y(new_n8065_));
  OAI21X1  g05629(.A0(new_n8064_), .A1(new_n8060_), .B0(new_n8065_), .Y(new_n8066_));
  OAI21X1  g05630(.A0(new_n8061_), .A1(new_n8053_), .B0(pi0075), .Y(new_n8067_));
  NAND3X1  g05631(.A(new_n8067_), .B(new_n8066_), .C(new_n5893_), .Y(new_n8068_));
  AOI22X1  g05632(.A0(new_n8068_), .A1(new_n8014_), .B0(new_n8056_), .B1(new_n8055_), .Y(new_n8069_));
  OAI21X1  g05633(.A0(new_n8069_), .A1(new_n8038_), .B0(new_n6520_), .Y(new_n8070_));
  AOI21X1  g05634(.A0(new_n8038_), .A1(new_n7949_), .B0(new_n2959_), .Y(new_n8071_));
  OAI21X1  g05635(.A0(new_n5118_), .A1(pi0057), .B0(new_n7989_), .Y(new_n8072_));
  OAI22X1  g05636(.A0(new_n8072_), .A1(new_n8071_), .B0(new_n8070_), .B1(new_n8037_), .Y(po0200));
  AND2X1   g05637(.A(pi0214), .B(pi0212), .Y(new_n8074_));
  NOR2X1   g05638(.A(pi0219), .B(pi0211), .Y(new_n8075_));
  MX2X1    g05639(.A(pi0211), .B(new_n8075_), .S0(new_n8074_), .Y(new_n8076_));
  MX2X1    g05640(.A(new_n7920_), .B(new_n7906_), .S0(new_n2723_), .Y(new_n8077_));
  OR2X1    g05641(.A(new_n7931_), .B(pi0228), .Y(new_n8078_));
  OAI21X1  g05642(.A0(new_n8077_), .A1(new_n3013_), .B0(new_n8078_), .Y(new_n8079_));
  NOR3X1   g05643(.A(pi0115), .B(pi0114), .C(pi0042), .Y(new_n8080_));
  NAND3X1  g05644(.A(new_n8080_), .B(new_n8079_), .C(pi0043), .Y(new_n8081_));
  INVX1    g05645(.A(pi0043), .Y(new_n8082_));
  NOR3X1   g05646(.A(new_n7809_), .B(new_n7903_), .C(pi0101), .Y(new_n8083_));
  OAI21X1  g05647(.A0(new_n7922_), .A1(new_n7903_), .B0(new_n2724_), .Y(new_n8084_));
  OAI21X1  g05648(.A0(new_n8083_), .A1(new_n2724_), .B0(new_n8084_), .Y(new_n8085_));
  NOR2X1   g05649(.A(new_n8085_), .B(new_n7909_), .Y(new_n8086_));
  MX2X1    g05650(.A(new_n8086_), .B(new_n7932_), .S0(new_n3013_), .Y(new_n8087_));
  INVX1    g05651(.A(new_n8087_), .Y(new_n8088_));
  AOI21X1  g05652(.A0(new_n2548_), .A1(pi0043), .B0(new_n8080_), .Y(new_n8089_));
  AOI21X1  g05653(.A0(new_n8088_), .A1(new_n8082_), .B0(new_n8089_), .Y(new_n8090_));
  AOI21X1  g05654(.A0(new_n8090_), .A1(new_n8081_), .B0(pi0039), .Y(new_n8091_));
  OAI21X1  g05655(.A0(new_n7945_), .A1(new_n8009_), .B0(pi0232), .Y(new_n8092_));
  AOI21X1  g05656(.A0(new_n8092_), .A1(new_n8008_), .B0(new_n2959_), .Y(new_n8093_));
  OAI21X1  g05657(.A0(new_n8093_), .A1(new_n8091_), .B0(new_n3277_), .Y(new_n8094_));
  AOI21X1  g05658(.A0(new_n2548_), .A1(pi0043), .B0(new_n6291_), .Y(new_n8095_));
  AND2X1   g05659(.A(new_n8080_), .B(new_n2723_), .Y(new_n8096_));
  OR2X1    g05660(.A(pi0072), .B(new_n8082_), .Y(new_n8097_));
  OAI21X1  g05661(.A0(new_n8096_), .A1(new_n8097_), .B0(new_n6291_), .Y(new_n8098_));
  NAND3X1  g05662(.A(new_n7963_), .B(pi0052), .C(new_n8082_), .Y(new_n8099_));
  OAI21X1  g05663(.A0(new_n7968_), .A1(new_n8082_), .B0(new_n8099_), .Y(new_n8100_));
  AOI21X1  g05664(.A0(new_n8100_), .A1(new_n8096_), .B0(new_n8098_), .Y(new_n8101_));
  OAI21X1  g05665(.A0(new_n8101_), .A1(new_n8095_), .B0(new_n2959_), .Y(new_n8102_));
  AOI21X1  g05666(.A0(new_n8102_), .A1(new_n8022_), .B0(new_n5086_), .Y(new_n8103_));
  AOI21X1  g05667(.A0(new_n2548_), .A1(pi0043), .B0(pi0039), .Y(new_n8104_));
  AOI21X1  g05668(.A0(new_n8011_), .A1(pi0039), .B0(new_n8104_), .Y(new_n8105_));
  OAI21X1  g05669(.A0(new_n8105_), .A1(new_n2996_), .B0(new_n3156_), .Y(new_n8106_));
  NOR2X1   g05670(.A(new_n8106_), .B(new_n8103_), .Y(new_n8107_));
  NOR3X1   g05671(.A(new_n7765_), .B(new_n7909_), .C(new_n7903_), .Y(new_n8108_));
  NOR2X1   g05672(.A(new_n8108_), .B(pi0043), .Y(new_n8109_));
  NOR2X1   g05673(.A(new_n7966_), .B(pi0072), .Y(new_n8110_));
  AND2X1   g05674(.A(new_n8080_), .B(pi0228), .Y(new_n8111_));
  OAI21X1  g05675(.A0(new_n8110_), .A1(new_n8082_), .B0(new_n8111_), .Y(new_n8112_));
  NOR2X1   g05676(.A(new_n8112_), .B(new_n8109_), .Y(new_n8113_));
  OAI21X1  g05677(.A0(new_n8111_), .A1(new_n8097_), .B0(new_n3085_), .Y(new_n8114_));
  AOI21X1  g05678(.A0(new_n8104_), .A1(new_n5792_), .B0(new_n3156_), .Y(new_n8115_));
  OAI21X1  g05679(.A0(new_n8114_), .A1(new_n8113_), .B0(new_n8115_), .Y(new_n8116_));
  OAI21X1  g05680(.A0(new_n8116_), .A1(new_n8012_), .B0(new_n3095_), .Y(new_n8117_));
  AOI21X1  g05681(.A0(new_n8107_), .A1(new_n8094_), .B0(new_n8117_), .Y(new_n8118_));
  INVX1    g05682(.A(new_n8104_), .Y(new_n8119_));
  OAI21X1  g05683(.A0(new_n7996_), .A1(pi0116), .B0(new_n2548_), .Y(new_n8120_));
  NAND4X1  g05684(.A(new_n7963_), .B(new_n5932_), .C(pi0052), .D(new_n8082_), .Y(new_n8121_));
  OAI21X1  g05685(.A0(new_n8120_), .A1(new_n8082_), .B0(new_n8121_), .Y(new_n8122_));
  AOI21X1  g05686(.A0(new_n8122_), .A1(new_n8096_), .B0(new_n8098_), .Y(new_n8123_));
  OAI21X1  g05687(.A0(new_n8123_), .A1(new_n8095_), .B0(new_n2959_), .Y(new_n8124_));
  MX2X1    g05688(.A(new_n8124_), .B(new_n8119_), .S0(new_n5788_), .Y(new_n8125_));
  AOI21X1  g05689(.A0(new_n8125_), .A1(new_n8022_), .B0(new_n3095_), .Y(new_n8126_));
  OR2X1    g05690(.A(new_n8126_), .B(new_n6309_), .Y(new_n8127_));
  AOI21X1  g05691(.A0(new_n8105_), .A1(new_n6309_), .B0(new_n7896_), .Y(new_n8128_));
  OAI21X1  g05692(.A0(new_n8127_), .A1(new_n8118_), .B0(new_n8128_), .Y(new_n8129_));
  NOR2X1   g05693(.A(pi0200), .B(pi0199), .Y(new_n8130_));
  NOR2X1   g05694(.A(new_n8130_), .B(pi0299), .Y(new_n8131_));
  INVX1    g05695(.A(new_n8131_), .Y(new_n8132_));
  AOI21X1  g05696(.A0(new_n8132_), .A1(new_n2548_), .B0(pi0232), .Y(new_n8133_));
  NOR2X1   g05697(.A(new_n8133_), .B(pi0299), .Y(new_n8134_));
  INVX1    g05698(.A(new_n8130_), .Y(new_n8135_));
  OAI21X1  g05699(.A0(new_n8135_), .A1(new_n7945_), .B0(pi0232), .Y(new_n8136_));
  AOI21X1  g05700(.A0(new_n8136_), .A1(new_n8134_), .B0(new_n2959_), .Y(new_n8137_));
  OAI21X1  g05701(.A0(new_n8137_), .A1(new_n8091_), .B0(new_n3277_), .Y(new_n8138_));
  AOI21X1  g05702(.A0(new_n8130_), .A1(new_n7943_), .B0(new_n5237_), .Y(new_n8139_));
  NOR3X1   g05703(.A(new_n8139_), .B(new_n8133_), .C(pi0299), .Y(new_n8140_));
  NOR2X1   g05704(.A(new_n8140_), .B(new_n2959_), .Y(new_n8141_));
  INVX1    g05705(.A(new_n8141_), .Y(new_n8142_));
  AOI21X1  g05706(.A0(new_n8142_), .A1(new_n8102_), .B0(new_n5086_), .Y(new_n8143_));
  NOR2X1   g05707(.A(new_n8141_), .B(new_n8104_), .Y(new_n8144_));
  OAI21X1  g05708(.A0(new_n8144_), .A1(new_n2996_), .B0(new_n3156_), .Y(new_n8145_));
  NOR2X1   g05709(.A(new_n8145_), .B(new_n8143_), .Y(new_n8146_));
  NOR2X1   g05710(.A(new_n8144_), .B(new_n3137_), .Y(new_n8147_));
  OAI21X1  g05711(.A0(new_n8147_), .A1(new_n8116_), .B0(new_n3095_), .Y(new_n8148_));
  AOI21X1  g05712(.A0(new_n8146_), .A1(new_n8138_), .B0(new_n8148_), .Y(new_n8149_));
  AOI21X1  g05713(.A0(new_n8142_), .A1(new_n8125_), .B0(new_n3095_), .Y(new_n8150_));
  OR2X1    g05714(.A(new_n8150_), .B(new_n6309_), .Y(new_n8151_));
  AOI21X1  g05715(.A0(new_n8144_), .A1(new_n6309_), .B0(new_n7897_), .Y(new_n8152_));
  OAI21X1  g05716(.A0(new_n8151_), .A1(new_n8149_), .B0(new_n8152_), .Y(new_n8153_));
  AOI21X1  g05717(.A0(new_n8153_), .A1(new_n8129_), .B0(new_n8076_), .Y(new_n8154_));
  INVX1    g05718(.A(new_n8076_), .Y(new_n8155_));
  OAI21X1  g05719(.A0(new_n7945_), .A1(new_n8009_), .B0(new_n7946_), .Y(new_n8156_));
  AOI21X1  g05720(.A0(new_n8007_), .A1(new_n7952_), .B0(new_n7950_), .Y(new_n8157_));
  AOI21X1  g05721(.A0(new_n8157_), .A1(new_n8156_), .B0(new_n2959_), .Y(new_n8158_));
  OAI21X1  g05722(.A0(new_n8158_), .A1(new_n8091_), .B0(new_n3277_), .Y(new_n8159_));
  AND2X1   g05723(.A(new_n8011_), .B(new_n7976_), .Y(new_n8160_));
  INVX1    g05724(.A(new_n8160_), .Y(new_n8161_));
  AOI21X1  g05725(.A0(new_n8161_), .A1(new_n8102_), .B0(new_n5086_), .Y(new_n8162_));
  AOI21X1  g05726(.A0(new_n8011_), .A1(new_n7976_), .B0(new_n8104_), .Y(new_n8163_));
  OAI21X1  g05727(.A0(new_n8163_), .A1(new_n2996_), .B0(new_n3156_), .Y(new_n8164_));
  NOR2X1   g05728(.A(new_n8164_), .B(new_n8162_), .Y(new_n8165_));
  OAI21X1  g05729(.A0(new_n8160_), .A1(new_n8116_), .B0(new_n3095_), .Y(new_n8166_));
  AOI21X1  g05730(.A0(new_n8165_), .A1(new_n8159_), .B0(new_n8166_), .Y(new_n8167_));
  AOI21X1  g05731(.A0(new_n8161_), .A1(new_n8125_), .B0(new_n3095_), .Y(new_n8168_));
  OR4X1    g05732(.A(new_n8168_), .B(new_n8167_), .C(new_n5107_), .D(pi0074), .Y(new_n8169_));
  AOI21X1  g05733(.A0(new_n8163_), .A1(new_n6309_), .B0(new_n7896_), .Y(new_n8170_));
  OAI21X1  g05734(.A0(new_n8135_), .A1(new_n7945_), .B0(new_n7946_), .Y(new_n8171_));
  NOR2X1   g05735(.A(new_n8133_), .B(new_n7950_), .Y(new_n8172_));
  AOI21X1  g05736(.A0(new_n8172_), .A1(new_n8171_), .B0(new_n2959_), .Y(new_n8173_));
  OAI21X1  g05737(.A0(new_n8173_), .A1(new_n8091_), .B0(new_n3277_), .Y(new_n8174_));
  NAND2X1  g05738(.A(new_n7949_), .B(pi0299), .Y(new_n8175_));
  AND2X1   g05739(.A(new_n8141_), .B(new_n8175_), .Y(new_n8176_));
  INVX1    g05740(.A(new_n8176_), .Y(new_n8177_));
  AOI21X1  g05741(.A0(new_n8177_), .A1(new_n8102_), .B0(new_n5086_), .Y(new_n8178_));
  AOI21X1  g05742(.A0(new_n8141_), .A1(new_n8175_), .B0(new_n8104_), .Y(new_n8179_));
  OAI21X1  g05743(.A0(new_n8179_), .A1(new_n2996_), .B0(new_n3156_), .Y(new_n8180_));
  NOR2X1   g05744(.A(new_n8180_), .B(new_n8178_), .Y(new_n8181_));
  OAI21X1  g05745(.A0(new_n8176_), .A1(new_n8116_), .B0(new_n3095_), .Y(new_n8182_));
  AOI21X1  g05746(.A0(new_n8181_), .A1(new_n8174_), .B0(new_n8182_), .Y(new_n8183_));
  AOI21X1  g05747(.A0(new_n8177_), .A1(new_n8125_), .B0(new_n3095_), .Y(new_n8184_));
  OR4X1    g05748(.A(new_n8184_), .B(new_n8183_), .C(new_n5107_), .D(pi0074), .Y(new_n8185_));
  AOI21X1  g05749(.A0(new_n8179_), .A1(new_n6309_), .B0(new_n7897_), .Y(new_n8186_));
  AOI22X1  g05750(.A0(new_n8186_), .A1(new_n8185_), .B0(new_n8170_), .B1(new_n8169_), .Y(new_n8187_));
  OAI21X1  g05751(.A0(new_n8187_), .A1(new_n8155_), .B0(new_n6520_), .Y(new_n8188_));
  AOI21X1  g05752(.A0(new_n8076_), .A1(new_n7949_), .B0(new_n2959_), .Y(new_n8189_));
  OR2X1    g05753(.A(new_n8104_), .B(new_n6520_), .Y(new_n8190_));
  OAI22X1  g05754(.A0(new_n8190_), .A1(new_n8189_), .B0(new_n8188_), .B1(new_n8154_), .Y(po0201));
  AND2X1   g05755(.A(new_n2548_), .B(pi0044), .Y(new_n8192_));
  INVX1    g05756(.A(new_n8192_), .Y(new_n8193_));
  AOI21X1  g05757(.A0(new_n8193_), .A1(new_n7761_), .B0(pi0039), .Y(new_n8194_));
  AOI21X1  g05758(.A0(new_n8192_), .A1(new_n2724_), .B0(new_n7761_), .Y(new_n8195_));
  AND2X1   g05759(.A(pi0072), .B(pi0044), .Y(new_n8196_));
  NOR4X1   g05760(.A(new_n8196_), .B(new_n5094_), .C(new_n2829_), .D(new_n2722_), .Y(new_n8197_));
  INVX1    g05761(.A(new_n8197_), .Y(new_n8198_));
  NOR4X1   g05762(.A(new_n5972_), .B(new_n3003_), .C(new_n2555_), .D(pi0044), .Y(new_n8199_));
  AND2X1   g05763(.A(new_n8199_), .B(new_n5932_), .Y(new_n8200_));
  AOI21X1  g05764(.A0(new_n7775_), .A1(pi0044), .B0(new_n8200_), .Y(new_n8201_));
  OAI21X1  g05765(.A0(new_n8201_), .A1(new_n8198_), .B0(new_n8195_), .Y(new_n8202_));
  NAND3X1  g05766(.A(new_n5930_), .B(new_n5929_), .C(pi0039), .Y(new_n8203_));
  NOR2X1   g05767(.A(new_n8203_), .B(pi0072), .Y(new_n8204_));
  AOI21X1  g05768(.A0(new_n8202_), .A1(new_n8194_), .B0(new_n8204_), .Y(new_n8205_));
  AOI21X1  g05769(.A0(new_n5970_), .A1(new_n2548_), .B0(new_n2959_), .Y(new_n8206_));
  AOI21X1  g05770(.A0(new_n8193_), .A1(new_n2959_), .B0(new_n8206_), .Y(new_n8207_));
  AOI21X1  g05771(.A0(new_n8207_), .A1(new_n5788_), .B0(new_n3095_), .Y(new_n8208_));
  OAI21X1  g05772(.A0(new_n8205_), .A1(new_n5788_), .B0(new_n8208_), .Y(new_n8209_));
  NAND2X1  g05773(.A(new_n7809_), .B(new_n2723_), .Y(new_n8210_));
  AOI21X1  g05774(.A0(new_n7817_), .A1(pi0044), .B0(new_n8210_), .Y(new_n8211_));
  NOR3X1   g05775(.A(new_n7825_), .B(new_n7798_), .C(pi0044), .Y(new_n8212_));
  NOR4X1   g05776(.A(new_n7815_), .B(new_n7796_), .C(pi0072), .D(new_n7868_), .Y(new_n8213_));
  NOR3X1   g05777(.A(new_n8213_), .B(new_n8212_), .C(new_n2723_), .Y(new_n8214_));
  OAI21X1  g05778(.A0(new_n8214_), .A1(new_n8211_), .B0(pi0228), .Y(new_n8215_));
  AOI21X1  g05779(.A0(new_n7857_), .A1(pi0044), .B0(pi0228), .Y(new_n8216_));
  AOI21X1  g05780(.A0(new_n8216_), .A1(new_n7854_), .B0(pi0039), .Y(new_n8217_));
  NOR4X1   g05781(.A(new_n7666_), .B(new_n2487_), .C(new_n2484_), .D(new_n2480_), .Y(new_n8218_));
  AOI21X1  g05782(.A0(new_n8218_), .A1(pi0287), .B0(pi0072), .Y(new_n8219_));
  INVX1    g05783(.A(new_n8219_), .Y(new_n8220_));
  OAI21X1  g05784(.A0(new_n8220_), .A1(new_n8203_), .B0(new_n3277_), .Y(new_n8221_));
  AOI21X1  g05785(.A0(new_n8217_), .A1(new_n8215_), .B0(new_n8221_), .Y(new_n8222_));
  NAND4X1  g05786(.A(new_n5971_), .B(new_n5189_), .C(new_n2486_), .D(new_n2550_), .Y(new_n8223_));
  AOI21X1  g05787(.A0(new_n8223_), .A1(pi0044), .B0(new_n8199_), .Y(new_n8224_));
  OAI21X1  g05788(.A0(new_n8224_), .A1(new_n8198_), .B0(new_n8195_), .Y(new_n8225_));
  OAI21X1  g05789(.A0(new_n8203_), .A1(pi0072), .B0(new_n5085_), .Y(new_n8226_));
  AOI21X1  g05790(.A0(new_n8225_), .A1(new_n8194_), .B0(new_n8226_), .Y(new_n8227_));
  OAI21X1  g05791(.A0(new_n8207_), .A1(new_n2996_), .B0(new_n3156_), .Y(new_n8228_));
  OR2X1    g05792(.A(new_n8228_), .B(new_n8227_), .Y(new_n8229_));
  NAND2X1  g05793(.A(new_n3277_), .B(pi0228), .Y(new_n8230_));
  OR4X1    g05794(.A(new_n8230_), .B(new_n3003_), .C(new_n2555_), .D(pi0044), .Y(new_n8231_));
  NAND3X1  g05795(.A(new_n8218_), .B(new_n3277_), .C(pi0228), .Y(new_n8232_));
  AOI21X1  g05796(.A0(new_n8232_), .A1(new_n8192_), .B0(pi0039), .Y(new_n8233_));
  NAND2X1  g05797(.A(new_n8233_), .B(new_n8231_), .Y(new_n8234_));
  NOR2X1   g05798(.A(new_n8206_), .B(new_n3156_), .Y(new_n8235_));
  AOI21X1  g05799(.A0(new_n8235_), .A1(new_n8234_), .B0(pi0075), .Y(new_n8236_));
  OAI21X1  g05800(.A0(new_n8229_), .A1(new_n8222_), .B0(new_n8236_), .Y(new_n8237_));
  AOI21X1  g05801(.A0(new_n8237_), .A1(new_n8209_), .B0(new_n6309_), .Y(new_n8238_));
  OAI21X1  g05802(.A0(new_n8207_), .A1(new_n5893_), .B0(new_n6520_), .Y(new_n8239_));
  AND2X1   g05803(.A(new_n5930_), .B(new_n2451_), .Y(new_n8240_));
  AOI21X1  g05804(.A0(new_n8240_), .A1(new_n2548_), .B0(new_n2959_), .Y(new_n8241_));
  OAI22X1  g05805(.A0(new_n8192_), .A1(pi0039), .B0(new_n5118_), .B1(pi0057), .Y(new_n8242_));
  OAI22X1  g05806(.A0(new_n8242_), .A1(new_n8241_), .B0(new_n8239_), .B1(new_n8238_), .Y(po0202));
  AND2X1   g05807(.A(pi0039), .B(new_n2996_), .Y(new_n8244_));
  NAND3X1  g05808(.A(new_n8244_), .B(new_n6520_), .C(new_n3129_), .Y(new_n8245_));
  NOR3X1   g05809(.A(new_n8245_), .B(new_n5243_), .C(new_n5035_), .Y(po0203));
  NOR3X1   g05810(.A(pi0111), .B(pi0104), .C(pi0102), .Y(new_n8247_));
  OR4X1    g05811(.A(pi0076), .B(pi0073), .C(pi0068), .D(pi0049), .Y(new_n8248_));
  NOR3X1   g05812(.A(new_n8248_), .B(new_n2472_), .C(pi0071), .Y(new_n8249_));
  AND2X1   g05813(.A(new_n8249_), .B(new_n8247_), .Y(new_n8250_));
  NOR2X1   g05814(.A(pi0077), .B(pi0050), .Y(new_n8251_));
  INVX1    g05815(.A(new_n8251_), .Y(new_n8252_));
  NAND4X1  g05816(.A(new_n2635_), .B(new_n2614_), .C(new_n2648_), .D(pi0061), .Y(new_n8253_));
  NOR4X1   g05817(.A(new_n8253_), .B(new_n6783_), .C(new_n6781_), .D(new_n8252_), .Y(new_n8254_));
  NAND4X1  g05818(.A(new_n8254_), .B(new_n8250_), .C(new_n7723_), .D(new_n6786_), .Y(new_n8255_));
  OR4X1    g05819(.A(new_n2587_), .B(new_n2484_), .C(new_n2477_), .D(new_n2694_), .Y(new_n8256_));
  OAI22X1  g05820(.A0(new_n8256_), .A1(new_n5787_), .B0(new_n8255_), .B1(pi0841), .Y(new_n8257_));
  AND2X1   g05821(.A(new_n8257_), .B(new_n7669_), .Y(po0204));
  INVX1    g05822(.A(new_n5985_), .Y(new_n8259_));
  AOI21X1  g05823(.A0(new_n2682_), .A1(pi0088), .B0(new_n8252_), .Y(new_n8260_));
  INVX1    g05824(.A(new_n8260_), .Y(new_n8261_));
  NOR2X1   g05825(.A(new_n2660_), .B(new_n2658_), .Y(new_n8262_));
  NAND3X1  g05826(.A(new_n2620_), .B(pi0104), .C(new_n6775_), .Y(new_n8263_));
  NOR4X1   g05827(.A(new_n8263_), .B(new_n7677_), .C(new_n2628_), .D(pi0082), .Y(new_n8264_));
  OR4X1    g05828(.A(pi0107), .B(pi0103), .C(pi0067), .D(pi0063), .Y(new_n8265_));
  NOR4X1   g05829(.A(new_n8265_), .B(new_n6872_), .C(new_n6782_), .D(pi0098), .Y(new_n8266_));
  OAI21X1  g05830(.A0(new_n8264_), .A1(pi0036), .B0(new_n8266_), .Y(new_n8267_));
  OAI21X1  g05831(.A0(new_n8267_), .A1(new_n8262_), .B0(new_n2681_), .Y(new_n8268_));
  NAND2X1  g05832(.A(new_n8268_), .B(new_n2528_), .Y(new_n8269_));
  NOR3X1   g05833(.A(new_n8269_), .B(new_n8261_), .C(new_n5007_), .Y(new_n8270_));
  OAI21X1  g05834(.A0(new_n8270_), .A1(new_n7664_), .B0(new_n7667_), .Y(new_n8271_));
  INVX1    g05835(.A(new_n8271_), .Y(new_n8272_));
  INVX1    g05836(.A(new_n2829_), .Y(new_n8273_));
  OR2X1    g05837(.A(new_n8271_), .B(new_n2783_), .Y(new_n8274_));
  NAND3X1  g05838(.A(new_n8266_), .B(new_n8264_), .C(new_n2658_), .Y(new_n8275_));
  AOI21X1  g05839(.A0(new_n8275_), .A1(new_n2681_), .B0(new_n8261_), .Y(new_n8276_));
  AND2X1   g05840(.A(new_n8276_), .B(new_n7683_), .Y(new_n8277_));
  AND2X1   g05841(.A(new_n2783_), .B(new_n5251_), .Y(new_n8278_));
  AOI21X1  g05842(.A0(new_n8278_), .A1(new_n8277_), .B0(new_n5258_), .Y(new_n8279_));
  NAND3X1  g05843(.A(new_n8279_), .B(new_n8274_), .C(new_n8273_), .Y(new_n8280_));
  OAI21X1  g05844(.A0(new_n8272_), .A1(new_n8259_), .B0(new_n8280_), .Y(new_n8281_));
  OR2X1    g05845(.A(new_n8271_), .B(new_n5938_), .Y(new_n8282_));
  AOI22X1  g05846(.A0(new_n8282_), .A1(new_n5258_), .B0(new_n8279_), .B1(new_n8274_), .Y(new_n8283_));
  INVX1    g05847(.A(new_n7667_), .Y(new_n8284_));
  NOR3X1   g05848(.A(new_n8284_), .B(new_n7665_), .C(new_n5939_), .Y(new_n8285_));
  AOI21X1  g05849(.A0(new_n5983_), .A1(new_n5259_), .B0(new_n8285_), .Y(new_n8286_));
  AOI21X1  g05850(.A0(new_n8286_), .A1(new_n8282_), .B0(new_n7749_), .Y(new_n8287_));
  OAI21X1  g05851(.A0(new_n8283_), .A1(pi1093), .B0(new_n8287_), .Y(new_n8288_));
  AOI21X1  g05852(.A0(new_n8281_), .A1(pi1091), .B0(new_n8288_), .Y(po0205));
  OR4X1    g05853(.A(new_n2725_), .B(new_n2726_), .C(pi0072), .D(pi0051), .Y(new_n8290_));
  NOR4X1   g05854(.A(new_n8290_), .B(new_n7728_), .C(new_n7682_), .D(new_n7749_), .Y(po0206));
  NOR4X1   g05855(.A(new_n2466_), .B(pi0089), .C(pi0082), .D(pi0048), .Y(new_n8292_));
  INVX1    g05856(.A(new_n8292_), .Y(new_n8293_));
  OR2X1    g05857(.A(new_n2472_), .B(new_n2459_), .Y(new_n8294_));
  OR4X1    g05858(.A(new_n7721_), .B(pi0103), .C(pi0067), .D(pi0036), .Y(new_n8295_));
  OR4X1    g05859(.A(new_n8295_), .B(new_n6782_), .C(pi0073), .D(pi0068), .Y(new_n8296_));
  NAND3X1  g05860(.A(new_n8247_), .B(pi0049), .C(new_n7725_), .Y(new_n8297_));
  NOR4X1   g05861(.A(new_n8297_), .B(new_n8296_), .C(new_n8294_), .D(new_n8293_), .Y(new_n8298_));
  NOR4X1   g05862(.A(new_n2484_), .B(new_n2478_), .C(pi0051), .D(pi0035), .Y(new_n8299_));
  AND2X1   g05863(.A(new_n8299_), .B(new_n8298_), .Y(new_n8300_));
  OR4X1    g05864(.A(new_n2726_), .B(pi0096), .C(pi0072), .D(pi0070), .Y(new_n8301_));
  NOR3X1   g05865(.A(new_n8301_), .B(new_n7666_), .C(new_n2492_), .Y(new_n8302_));
  AOI21X1  g05866(.A0(new_n8302_), .A1(new_n8300_), .B0(pi0074), .Y(new_n8303_));
  OR4X1    g05867(.A(new_n8303_), .B(new_n5850_), .C(new_n5118_), .D(pi0057), .Y(new_n8304_));
  AOI21X1  g05868(.A0(new_n7605_), .A1(pi0074), .B0(new_n8304_), .Y(po0207));
  INVX1    g05869(.A(new_n6756_), .Y(new_n8306_));
  NAND3X1  g05870(.A(new_n6768_), .B(new_n2483_), .C(pi0024), .Y(new_n8307_));
  NAND2X1  g05871(.A(new_n8307_), .B(new_n7832_), .Y(new_n8308_));
  NAND2X1  g05872(.A(new_n6767_), .B(new_n6766_), .Y(new_n8309_));
  NAND3X1  g05873(.A(new_n8309_), .B(new_n2590_), .C(pi0024), .Y(new_n8310_));
  MX2X1    g05874(.A(po0840), .B(new_n6763_), .S0(new_n3053_), .Y(new_n8311_));
  NAND4X1  g05875(.A(new_n8311_), .B(new_n8310_), .C(new_n8308_), .D(new_n7667_), .Y(new_n8312_));
  NOR2X1   g05876(.A(new_n5911_), .B(new_n5193_), .Y(new_n8313_));
  INVX1    g05877(.A(new_n8313_), .Y(new_n8314_));
  OR4X1    g05878(.A(new_n8314_), .B(new_n8311_), .C(pi0090), .D(new_n5787_), .Y(new_n8315_));
  OR2X1    g05879(.A(new_n8315_), .B(new_n6770_), .Y(new_n8316_));
  AOI21X1  g05880(.A0(new_n8316_), .A1(new_n8312_), .B0(pi0100), .Y(new_n8317_));
  NOR3X1   g05881(.A(new_n5284_), .B(new_n5083_), .C(new_n3026_), .Y(new_n8318_));
  NOR4X1   g05882(.A(pi0087), .B(pi0075), .C(pi0039), .D(pi0038), .Y(new_n8319_));
  OAI21X1  g05883(.A0(new_n8318_), .A1(new_n8317_), .B0(new_n8319_), .Y(new_n8320_));
  NAND4X1  g05884(.A(new_n6811_), .B(new_n7604_), .C(new_n6773_), .D(new_n6809_), .Y(new_n8321_));
  AOI21X1  g05885(.A0(new_n8321_), .A1(new_n8320_), .B0(new_n8306_), .Y(po0208));
  NOR4X1   g05886(.A(new_n7749_), .B(new_n8284_), .C(new_n2529_), .D(new_n5007_), .Y(new_n8323_));
  INVX1    g05887(.A(new_n8323_), .Y(new_n8324_));
  OR4X1    g05888(.A(new_n8294_), .B(new_n6872_), .C(pi0071), .D(pi0065), .Y(new_n8325_));
  OR4X1    g05889(.A(new_n8325_), .B(new_n5141_), .C(new_n2463_), .D(pi0069), .Y(new_n8326_));
  NOR3X1   g05890(.A(new_n8326_), .B(new_n8324_), .C(new_n2655_), .Y(po0209));
  OR2X1    g05891(.A(new_n8074_), .B(pi0211), .Y(new_n8328_));
  OR2X1    g05892(.A(new_n8328_), .B(pi0219), .Y(new_n8329_));
  INVX1    g05893(.A(pi0052), .Y(new_n8330_));
  NOR3X1   g05894(.A(pi0072), .B(new_n8330_), .C(pi0039), .Y(new_n8331_));
  AND2X1   g05895(.A(new_n2548_), .B(pi0052), .Y(new_n8332_));
  NOR4X1   g05896(.A(pi0115), .B(pi0114), .C(pi0043), .D(pi0042), .Y(new_n8333_));
  NAND2X1  g05897(.A(new_n8333_), .B(pi0228), .Y(new_n8334_));
  MX2X1    g05898(.A(new_n8110_), .B(new_n8108_), .S0(new_n8330_), .Y(new_n8335_));
  MX2X1    g05899(.A(new_n8335_), .B(new_n8332_), .S0(new_n8334_), .Y(new_n8336_));
  MX2X1    g05900(.A(new_n8336_), .B(new_n8331_), .S0(pi0038), .Y(new_n8337_));
  NOR2X1   g05901(.A(new_n8331_), .B(new_n3026_), .Y(new_n8338_));
  NOR3X1   g05902(.A(pi0100), .B(new_n2959_), .C(pi0038), .Y(new_n8339_));
  OR2X1    g05903(.A(new_n8339_), .B(new_n3156_), .Y(new_n8340_));
  NOR2X1   g05904(.A(new_n8340_), .B(new_n8338_), .Y(new_n8341_));
  OAI21X1  g05905(.A0(new_n8337_), .A1(pi0100), .B0(new_n8341_), .Y(new_n8342_));
  NOR3X1   g05906(.A(pi0114), .B(pi0043), .C(pi0042), .Y(new_n8343_));
  INVX1    g05907(.A(new_n8343_), .Y(new_n8344_));
  NAND2X1  g05908(.A(new_n7906_), .B(pi0052), .Y(new_n8345_));
  AOI21X1  g05909(.A0(new_n7910_), .A1(new_n8330_), .B0(new_n7994_), .Y(new_n8346_));
  INVX1    g05910(.A(new_n7923_), .Y(new_n8347_));
  OAI21X1  g05911(.A0(new_n8347_), .A1(pi0052), .B0(new_n7916_), .Y(new_n8348_));
  AOI21X1  g05912(.A0(new_n7920_), .A1(pi0052), .B0(new_n8348_), .Y(new_n8349_));
  AOI21X1  g05913(.A0(new_n8346_), .A1(new_n8345_), .B0(new_n8349_), .Y(new_n8350_));
  INVX1    g05914(.A(new_n8332_), .Y(new_n8351_));
  INVX1    g05915(.A(new_n8333_), .Y(new_n8352_));
  AOI21X1  g05916(.A0(new_n8352_), .A1(new_n8351_), .B0(new_n3013_), .Y(new_n8353_));
  OAI21X1  g05917(.A0(new_n8350_), .A1(new_n8344_), .B0(new_n8353_), .Y(new_n8354_));
  INVX1    g05918(.A(new_n7931_), .Y(new_n8355_));
  AOI21X1  g05919(.A0(new_n7932_), .A1(new_n8330_), .B0(new_n8352_), .Y(new_n8356_));
  OAI21X1  g05920(.A0(new_n8355_), .A1(new_n8330_), .B0(new_n8356_), .Y(new_n8357_));
  AOI21X1  g05921(.A0(new_n8352_), .A1(new_n8351_), .B0(pi0228), .Y(new_n8358_));
  AOI21X1  g05922(.A0(new_n8358_), .A1(new_n8357_), .B0(pi0039), .Y(new_n8359_));
  NAND3X1  g05923(.A(new_n8359_), .B(new_n8354_), .C(new_n3026_), .Y(new_n8360_));
  NAND4X1  g05924(.A(new_n8343_), .B(new_n7899_), .C(new_n6291_), .D(new_n5971_), .Y(new_n8361_));
  OAI21X1  g05925(.A0(new_n8361_), .A1(new_n7967_), .B0(new_n8332_), .Y(new_n8362_));
  AOI21X1  g05926(.A0(new_n8362_), .A1(pi0100), .B0(pi0039), .Y(new_n8363_));
  AOI21X1  g05927(.A0(new_n8363_), .A1(new_n8360_), .B0(pi0038), .Y(new_n8364_));
  OAI21X1  g05928(.A0(new_n8331_), .A1(new_n2996_), .B0(new_n3156_), .Y(new_n8365_));
  OAI21X1  g05929(.A0(new_n8365_), .A1(new_n8364_), .B0(new_n8342_), .Y(new_n8366_));
  AND2X1   g05930(.A(new_n7899_), .B(new_n6291_), .Y(new_n8367_));
  INVX1    g05931(.A(new_n8367_), .Y(new_n8368_));
  OR4X1    g05932(.A(new_n8368_), .B(new_n8344_), .C(new_n7996_), .D(pi0116), .Y(new_n8369_));
  OAI21X1  g05933(.A0(new_n8369_), .A1(new_n5788_), .B0(new_n8331_), .Y(new_n8370_));
  OAI21X1  g05934(.A0(new_n8370_), .A1(new_n3095_), .B0(new_n5893_), .Y(new_n8371_));
  AOI21X1  g05935(.A0(new_n8366_), .A1(new_n3095_), .B0(new_n8371_), .Y(new_n8372_));
  OAI21X1  g05936(.A0(new_n8331_), .A1(new_n5893_), .B0(new_n7896_), .Y(new_n8373_));
  AND2X1   g05937(.A(new_n8359_), .B(new_n8354_), .Y(new_n8374_));
  OAI21X1  g05938(.A0(new_n8374_), .A1(new_n8137_), .B0(new_n3277_), .Y(new_n8375_));
  AND2X1   g05939(.A(new_n8362_), .B(new_n2959_), .Y(new_n8376_));
  OAI21X1  g05940(.A0(new_n8376_), .A1(new_n8141_), .B0(new_n5085_), .Y(new_n8377_));
  MX2X1    g05941(.A(new_n8332_), .B(new_n8140_), .S0(pi0039), .Y(new_n8378_));
  OR2X1    g05942(.A(new_n8378_), .B(new_n2996_), .Y(new_n8379_));
  AND2X1   g05943(.A(new_n8379_), .B(new_n3156_), .Y(new_n8380_));
  AND2X1   g05944(.A(new_n8380_), .B(new_n8377_), .Y(new_n8381_));
  OR2X1    g05945(.A(new_n8336_), .B(pi0039), .Y(new_n8382_));
  NOR2X1   g05946(.A(new_n8141_), .B(new_n5792_), .Y(new_n8383_));
  AOI22X1  g05947(.A0(new_n8383_), .A1(new_n8382_), .B0(new_n8378_), .B1(new_n5792_), .Y(new_n8384_));
  OAI21X1  g05948(.A0(new_n8384_), .A1(new_n3156_), .B0(new_n3095_), .Y(new_n8385_));
  AOI21X1  g05949(.A0(new_n8381_), .A1(new_n8375_), .B0(new_n8385_), .Y(new_n8386_));
  AOI21X1  g05950(.A0(new_n8369_), .A1(new_n8332_), .B0(pi0039), .Y(new_n8387_));
  OAI21X1  g05951(.A0(new_n8140_), .A1(new_n2959_), .B0(new_n3108_), .Y(new_n8388_));
  AOI21X1  g05952(.A0(new_n8378_), .A1(new_n5788_), .B0(new_n3095_), .Y(new_n8389_));
  OAI21X1  g05953(.A0(new_n8388_), .A1(new_n8387_), .B0(new_n8389_), .Y(new_n8390_));
  NAND3X1  g05954(.A(new_n8390_), .B(new_n7897_), .C(new_n5893_), .Y(new_n8391_));
  OAI22X1  g05955(.A0(new_n8391_), .A1(new_n8386_), .B0(new_n8373_), .B1(new_n8372_), .Y(new_n8392_));
  NAND2X1  g05956(.A(new_n8392_), .B(new_n8329_), .Y(new_n8393_));
  INVX1    g05957(.A(new_n8374_), .Y(new_n8394_));
  OAI21X1  g05958(.A0(new_n7952_), .A1(new_n7950_), .B0(pi0039), .Y(new_n8395_));
  AOI21X1  g05959(.A0(new_n8395_), .A1(new_n8394_), .B0(new_n5792_), .Y(new_n8396_));
  AOI21X1  g05960(.A0(new_n8351_), .A1(new_n2959_), .B0(new_n7976_), .Y(new_n8397_));
  AOI21X1  g05961(.A0(new_n8362_), .A1(new_n2959_), .B0(new_n7976_), .Y(new_n8398_));
  OAI22X1  g05962(.A0(new_n8398_), .A1(new_n5086_), .B0(new_n8397_), .B1(new_n2996_), .Y(new_n8399_));
  OAI21X1  g05963(.A0(new_n8399_), .A1(new_n8396_), .B0(new_n3156_), .Y(new_n8400_));
  AOI21X1  g05964(.A0(new_n8397_), .A1(new_n5792_), .B0(new_n3156_), .Y(new_n8401_));
  NOR2X1   g05965(.A(new_n7976_), .B(new_n5792_), .Y(new_n8402_));
  OAI21X1  g05966(.A0(new_n8336_), .A1(pi0039), .B0(new_n8402_), .Y(new_n8403_));
  AOI21X1  g05967(.A0(new_n8403_), .A1(new_n8401_), .B0(new_n7897_), .Y(new_n8404_));
  AOI21X1  g05968(.A0(new_n8359_), .A1(new_n8354_), .B0(new_n8173_), .Y(new_n8405_));
  NOR2X1   g05969(.A(new_n8405_), .B(new_n5792_), .Y(new_n8406_));
  AOI21X1  g05970(.A0(new_n8362_), .A1(new_n2959_), .B0(new_n8176_), .Y(new_n8407_));
  OAI22X1  g05971(.A0(new_n8407_), .A1(new_n5086_), .B0(new_n8397_), .B1(new_n8379_), .Y(new_n8408_));
  OAI21X1  g05972(.A0(new_n8408_), .A1(new_n8406_), .B0(new_n3156_), .Y(new_n8409_));
  NAND3X1  g05973(.A(new_n8382_), .B(new_n8177_), .C(new_n3277_), .Y(new_n8410_));
  NAND2X1  g05974(.A(new_n8378_), .B(new_n5792_), .Y(new_n8411_));
  AND2X1   g05975(.A(new_n8401_), .B(new_n8411_), .Y(new_n8412_));
  AOI21X1  g05976(.A0(new_n8412_), .A1(new_n8410_), .B0(new_n7896_), .Y(new_n8413_));
  AOI22X1  g05977(.A0(new_n8413_), .A1(new_n8409_), .B0(new_n8404_), .B1(new_n8400_), .Y(new_n8414_));
  AOI21X1  g05978(.A0(new_n7976_), .A1(new_n7896_), .B0(new_n3095_), .Y(new_n8415_));
  OAI21X1  g05979(.A0(new_n8177_), .A1(new_n7896_), .B0(new_n8415_), .Y(new_n8416_));
  AOI21X1  g05980(.A0(new_n8370_), .A1(new_n2959_), .B0(new_n8416_), .Y(new_n8417_));
  NOR2X1   g05981(.A(new_n8417_), .B(new_n6309_), .Y(new_n8418_));
  OAI21X1  g05982(.A0(new_n8414_), .A1(pi0075), .B0(new_n8418_), .Y(new_n8419_));
  NOR2X1   g05983(.A(new_n8397_), .B(new_n5893_), .Y(new_n8420_));
  NOR2X1   g05984(.A(new_n8420_), .B(new_n8329_), .Y(new_n8421_));
  NAND3X1  g05985(.A(new_n8378_), .B(new_n7897_), .C(new_n6309_), .Y(new_n8422_));
  NAND2X1  g05986(.A(new_n8422_), .B(new_n6520_), .Y(new_n8423_));
  AOI21X1  g05987(.A0(new_n8421_), .A1(new_n8419_), .B0(new_n8423_), .Y(new_n8424_));
  NOR4X1   g05988(.A(new_n8074_), .B(pi0219), .C(pi0211), .D(new_n2959_), .Y(new_n8425_));
  OR2X1    g05989(.A(new_n8331_), .B(new_n6520_), .Y(new_n8426_));
  AOI21X1  g05990(.A0(new_n8425_), .A1(new_n7949_), .B0(new_n8426_), .Y(new_n8427_));
  AOI21X1  g05991(.A0(new_n8424_), .A1(new_n8393_), .B0(new_n8427_), .Y(po0210));
  AND2X1   g05992(.A(new_n7667_), .B(pi0024), .Y(new_n8429_));
  NOR4X1   g05993(.A(new_n2506_), .B(new_n2499_), .C(new_n2498_), .D(new_n2493_), .Y(new_n8430_));
  AOI21X1  g05994(.A0(new_n8430_), .A1(new_n8429_), .B0(pi0039), .Y(new_n8431_));
  NOR2X1   g05995(.A(pi0979), .B(pi0287), .Y(new_n8432_));
  AOI21X1  g05996(.A0(new_n8432_), .A1(new_n5034_), .B0(new_n2959_), .Y(new_n8433_));
  NOR4X1   g05997(.A(new_n8433_), .B(new_n8431_), .C(new_n7690_), .D(new_n3193_), .Y(po0211));
  NOR3X1   g05998(.A(new_n6755_), .B(new_n3393_), .C(new_n5324_), .Y(new_n8435_));
  INVX1    g05999(.A(new_n8435_), .Y(new_n8436_));
  AOI21X1  g06000(.A0(new_n7674_), .A1(new_n3109_), .B0(new_n3112_), .Y(new_n8437_));
  NAND4X1  g06001(.A(new_n6769_), .B(new_n2505_), .C(new_n2497_), .D(new_n2493_), .Y(new_n8438_));
  INVX1    g06002(.A(pi0106), .Y(new_n8439_));
  OR2X1    g06003(.A(pi0085), .B(pi0060), .Y(new_n8440_));
  OR4X1    g06004(.A(pi0111), .B(pi0102), .C(pi0089), .D(pi0082), .Y(new_n8441_));
  OR4X1    g06005(.A(new_n8441_), .B(new_n8440_), .C(new_n8248_), .D(new_n8439_), .Y(new_n8442_));
  OR4X1    g06006(.A(new_n8442_), .B(new_n8295_), .C(new_n8294_), .D(new_n6784_), .Y(new_n8443_));
  NOR2X1   g06007(.A(new_n8443_), .B(new_n8438_), .Y(new_n8444_));
  OR4X1    g06008(.A(new_n3256_), .B(new_n2725_), .C(new_n2492_), .D(pi0841), .Y(new_n8445_));
  NOR4X1   g06009(.A(new_n8445_), .B(new_n3107_), .C(pi0051), .D(pi0035), .Y(new_n8446_));
  AOI21X1  g06010(.A0(new_n8446_), .A1(new_n8444_), .B0(pi0054), .Y(new_n8447_));
  NOR3X1   g06011(.A(new_n8447_), .B(new_n8437_), .C(new_n8436_), .Y(po0212));
  NAND3X1  g06012(.A(new_n7674_), .B(new_n3109_), .C(new_n3112_), .Y(new_n8449_));
  NOR2X1   g06013(.A(new_n8449_), .B(pi0074), .Y(new_n8450_));
  NOR2X1   g06014(.A(new_n8450_), .B(new_n3128_), .Y(new_n8451_));
  OR4X1    g06015(.A(new_n2472_), .B(pi0111), .C(pi0082), .D(new_n7725_), .Y(new_n8452_));
  OR4X1    g06016(.A(new_n8452_), .B(new_n8296_), .C(new_n2467_), .D(pi0104), .Y(new_n8453_));
  OR2X1    g06017(.A(new_n7057_), .B(new_n7666_), .Y(new_n8454_));
  NOR4X1   g06018(.A(new_n8454_), .B(new_n8453_), .C(new_n3131_), .D(new_n2461_), .Y(new_n8455_));
  NOR2X1   g06019(.A(new_n8455_), .B(pi0055), .Y(new_n8456_));
  NOR4X1   g06020(.A(new_n8456_), .B(new_n8451_), .C(new_n3393_), .D(new_n5324_), .Y(po0213));
  OR2X1    g06021(.A(pi0062), .B(new_n3143_), .Y(new_n8458_));
  NAND4X1  g06022(.A(new_n7604_), .B(new_n3148_), .C(new_n3130_), .D(pi0055), .Y(new_n8459_));
  NOR4X1   g06023(.A(new_n5020_), .B(new_n3242_), .C(new_n7272_), .D(new_n2727_), .Y(new_n8460_));
  OAI21X1  g06024(.A0(new_n8460_), .A1(new_n3143_), .B0(new_n3246_), .Y(new_n8461_));
  AOI21X1  g06025(.A0(new_n8459_), .A1(new_n8458_), .B0(new_n8461_), .Y(po0214));
  AOI21X1  g06026(.A0(new_n8450_), .A1(new_n5327_), .B0(new_n2436_), .Y(new_n8463_));
  NOR4X1   g06027(.A(new_n5915_), .B(new_n3242_), .C(new_n7272_), .D(new_n2768_), .Y(new_n8464_));
  INVX1    g06028(.A(pi0924), .Y(new_n8465_));
  NAND3X1  g06029(.A(new_n8465_), .B(pi0062), .C(new_n3143_), .Y(new_n8466_));
  NAND2X1  g06030(.A(new_n8466_), .B(new_n8458_), .Y(new_n8467_));
  AOI21X1  g06031(.A0(new_n8467_), .A1(new_n8464_), .B0(pi0057), .Y(new_n8468_));
  NOR3X1   g06032(.A(new_n8468_), .B(new_n8463_), .C(pi0059), .Y(po0215));
  NOR3X1   g06033(.A(new_n8314_), .B(new_n7749_), .C(pi0093), .Y(new_n8470_));
  AND2X1   g06034(.A(new_n8470_), .B(new_n5898_), .Y(po0216));
  AOI21X1  g06035(.A0(new_n8450_), .A1(new_n5327_), .B0(new_n3153_), .Y(new_n8472_));
  NOR3X1   g06036(.A(new_n8465_), .B(new_n3245_), .C(pi0056), .Y(new_n8473_));
  AOI21X1  g06037(.A0(new_n8473_), .A1(new_n8464_), .B0(pi0059), .Y(new_n8474_));
  NOR3X1   g06038(.A(new_n8474_), .B(new_n8472_), .C(pi0057), .Y(po0217));
  OR4X1    g06039(.A(new_n5036_), .B(new_n5034_), .C(pi0979), .D(new_n2959_), .Y(new_n8476_));
  OR4X1    g06040(.A(new_n8476_), .B(new_n3003_), .C(new_n2555_), .D(pi0287), .Y(new_n8477_));
  OR4X1    g06041(.A(new_n8438_), .B(new_n8284_), .C(pi0039), .D(new_n5787_), .Y(new_n8478_));
  OR2X1    g06042(.A(new_n8478_), .B(new_n2495_), .Y(new_n8479_));
  AOI21X1  g06043(.A0(new_n8479_), .A1(new_n8477_), .B0(new_n7690_), .Y(po0218));
  OR2X1    g06044(.A(new_n8438_), .B(pi0024), .Y(new_n8481_));
  OAI22X1  g06045(.A0(new_n8481_), .A1(new_n2495_), .B0(new_n8255_), .B1(new_n2726_), .Y(new_n8482_));
  AND2X1   g06046(.A(new_n8482_), .B(new_n7669_), .Y(po0219));
  NOR2X1   g06047(.A(new_n7653_), .B(new_n2436_), .Y(new_n8484_));
  AND2X1   g06048(.A(pi0062), .B(new_n3143_), .Y(new_n8485_));
  AOI21X1  g06049(.A0(new_n8485_), .A1(new_n8460_), .B0(pi0057), .Y(new_n8486_));
  NOR3X1   g06050(.A(new_n8486_), .B(new_n8484_), .C(pi0059), .Y(po0220));
  INVX1    g06051(.A(pi0999), .Y(new_n8488_));
  INVX1    g06052(.A(new_n6786_), .Y(new_n8489_));
  OR4X1    g06053(.A(new_n6874_), .B(new_n8489_), .C(pi0107), .D(new_n2674_), .Y(new_n8490_));
  OAI22X1  g06054(.A0(new_n8490_), .A1(new_n8488_), .B0(new_n8256_), .B1(pi0024), .Y(new_n8491_));
  AND2X1   g06055(.A(new_n8491_), .B(new_n7669_), .Y(po0221));
  OR4X1    g06056(.A(new_n2471_), .B(new_n2462_), .C(new_n2609_), .D(pi0063), .Y(new_n8493_));
  AND2X1   g06057(.A(new_n8493_), .B(new_n2605_), .Y(new_n8494_));
  OR4X1    g06058(.A(new_n8494_), .B(new_n2608_), .C(new_n2461_), .D(pi0081), .Y(new_n8495_));
  NOR4X1   g06059(.A(new_n6873_), .B(new_n2471_), .C(new_n2609_), .D(pi0063), .Y(new_n8496_));
  OAI21X1  g06060(.A0(new_n8496_), .A1(pi0841), .B0(new_n8323_), .Y(new_n8497_));
  AOI21X1  g06061(.A0(new_n8495_), .A1(pi0841), .B0(new_n8497_), .Y(po0222));
  NOR3X1   g06062(.A(new_n7702_), .B(new_n7700_), .C(pi0299), .Y(new_n8499_));
  NAND3X1  g06063(.A(new_n7712_), .B(pi0786), .C(pi0039), .Y(new_n8500_));
  NOR4X1   g06064(.A(new_n8500_), .B(new_n7709_), .C(new_n8499_), .D(new_n7690_), .Y(po0223));
  NOR2X1   g06065(.A(pi0299), .B(pi0199), .Y(new_n8502_));
  INVX1    g06066(.A(new_n8502_), .Y(new_n8503_));
  OR4X1    g06067(.A(new_n7057_), .B(new_n7666_), .C(new_n2459_), .D(new_n7734_), .Y(new_n8504_));
  NOR4X1   g06068(.A(new_n8504_), .B(new_n2473_), .C(pi0102), .D(new_n2509_), .Y(new_n8505_));
  NAND3X1  g06069(.A(new_n8505_), .B(new_n8503_), .C(new_n3130_), .Y(new_n8506_));
  AND2X1   g06070(.A(new_n8506_), .B(pi0219), .Y(new_n8507_));
  NAND3X1  g06071(.A(new_n3135_), .B(new_n3105_), .C(new_n3277_), .Y(new_n8508_));
  NOR4X1   g06072(.A(new_n8508_), .B(new_n7188_), .C(pi0299), .D(new_n7941_), .Y(new_n8509_));
  AOI21X1  g06073(.A0(new_n8509_), .A1(new_n8505_), .B0(pi0219), .Y(new_n8510_));
  NOR3X1   g06074(.A(new_n8510_), .B(new_n8507_), .C(po1038), .Y(po0224));
  INVX1    g06075(.A(new_n2616_), .Y(new_n8512_));
  OR4X1    g06076(.A(new_n8325_), .B(new_n7749_), .C(pi0103), .D(new_n2614_), .Y(new_n8513_));
  NOR3X1   g06077(.A(new_n8513_), .B(new_n8504_), .C(new_n8512_), .Y(po0225));
  INVX1    g06078(.A(new_n5074_), .Y(new_n8515_));
  NOR4X1   g06079(.A(new_n2953_), .B(pi0221), .C(new_n2438_), .D(pi0215), .Y(new_n8516_));
  NAND3X1  g06080(.A(new_n8516_), .B(new_n5261_), .C(new_n8515_), .Y(new_n8517_));
  INVX1    g06081(.A(new_n5058_), .Y(new_n8518_));
  NOR4X1   g06082(.A(pi0299), .B(new_n2961_), .C(pi0223), .D(pi0222), .Y(new_n8519_));
  NAND3X1  g06083(.A(new_n8519_), .B(new_n5261_), .C(new_n8518_), .Y(new_n8520_));
  AOI21X1  g06084(.A0(new_n8520_), .A1(new_n8517_), .B0(new_n8245_), .Y(po0226));
  NOR4X1   g06085(.A(pi0103), .B(new_n7658_), .C(pi0067), .D(pi0036), .Y(new_n8522_));
  AOI21X1  g06086(.A0(new_n8522_), .A1(new_n7659_), .B0(pi0071), .Y(new_n8523_));
  OR4X1    g06087(.A(new_n2459_), .B(pi0314), .C(pi0102), .D(pi0081), .Y(new_n8524_));
  OR4X1    g06088(.A(new_n8524_), .B(new_n8523_), .C(po1049), .D(new_n2611_), .Y(new_n8525_));
  NAND4X1  g06089(.A(new_n7660_), .B(new_n8251_), .C(pi0314), .D(pi0071), .Y(new_n8526_));
  OR2X1    g06090(.A(new_n8526_), .B(new_n2471_), .Y(new_n8527_));
  AOI21X1  g06091(.A0(new_n8527_), .A1(new_n8525_), .B0(new_n8324_), .Y(po0227));
  OR4X1    g06092(.A(new_n2709_), .B(pi0096), .C(new_n5134_), .D(pi0051), .Y(new_n8529_));
  OR4X1    g06093(.A(new_n8529_), .B(new_n3256_), .C(pi0039), .D(new_n5787_), .Y(new_n8530_));
  AND2X1   g06094(.A(pi0589), .B(pi0198), .Y(new_n8531_));
  NOR2X1   g06095(.A(new_n5058_), .B(new_n3285_), .Y(new_n8532_));
  AND2X1   g06096(.A(pi0589), .B(pi0210), .Y(new_n8533_));
  NAND3X1  g06097(.A(pi0299), .B(new_n2437_), .C(new_n2954_), .Y(new_n8534_));
  NOR3X1   g06098(.A(new_n8534_), .B(new_n5074_), .C(pi0216), .Y(new_n8535_));
  AOI22X1  g06099(.A0(new_n8535_), .A1(new_n8533_), .B0(new_n8532_), .B1(new_n8531_), .Y(new_n8536_));
  NOR4X1   g06100(.A(new_n8536_), .B(new_n5255_), .C(new_n5245_), .D(pi0593), .Y(new_n8537_));
  OAI21X1  g06101(.A0(new_n8537_), .A1(pi0287), .B0(pi0039), .Y(new_n8538_));
  OR2X1    g06102(.A(new_n8538_), .B(new_n3074_), .Y(new_n8539_));
  AOI21X1  g06103(.A0(new_n8539_), .A1(new_n8530_), .B0(new_n7690_), .Y(po0228));
  OR4X1    g06104(.A(new_n7842_), .B(new_n2511_), .C(new_n2478_), .D(pi0050), .Y(new_n8541_));
  NOR4X1   g06105(.A(new_n8541_), .B(new_n5162_), .C(new_n2577_), .D(pi0077), .Y(new_n8542_));
  INVX1    g06106(.A(new_n8542_), .Y(new_n8543_));
  INVX1    g06107(.A(new_n5146_), .Y(new_n8544_));
  OR4X1    g06108(.A(new_n8265_), .B(new_n8544_), .C(new_n2469_), .D(new_n2465_), .Y(new_n8545_));
  NOR3X1   g06109(.A(new_n8545_), .B(new_n6782_), .C(pi0064), .Y(new_n8546_));
  NOR3X1   g06110(.A(pi0299), .B(new_n8009_), .C(pi0199), .Y(new_n8547_));
  INVX1    g06111(.A(pi0211), .Y(new_n8548_));
  NOR3X1   g06112(.A(new_n2953_), .B(pi0219), .C(new_n8548_), .Y(new_n8549_));
  NOR2X1   g06113(.A(new_n8549_), .B(new_n8547_), .Y(new_n8550_));
  NOR3X1   g06114(.A(new_n8550_), .B(new_n8284_), .C(new_n7734_), .Y(new_n8551_));
  OAI21X1  g06115(.A0(new_n8546_), .A1(pi0081), .B0(new_n8551_), .Y(new_n8552_));
  INVX1    g06116(.A(new_n8550_), .Y(new_n8553_));
  OR4X1    g06117(.A(new_n8553_), .B(new_n8504_), .C(new_n6872_), .D(new_n6782_), .Y(new_n8554_));
  OAI22X1  g06118(.A0(new_n8554_), .A1(new_n8545_), .B0(new_n8552_), .B1(new_n8543_), .Y(new_n8555_));
  AND2X1   g06119(.A(new_n8555_), .B(new_n7668_), .Y(po0229));
  NAND3X1  g06120(.A(new_n2486_), .B(new_n2550_), .C(pi0024), .Y(new_n8557_));
  NOR2X1   g06121(.A(new_n8557_), .B(new_n2548_), .Y(new_n8558_));
  INVX1    g06122(.A(new_n6972_), .Y(new_n8559_));
  OR4X1    g06123(.A(pi0077), .B(pi0060), .C(pi0053), .D(pi0050), .Y(new_n8560_));
  OR4X1    g06124(.A(new_n8560_), .B(new_n2506_), .C(new_n2498_), .D(new_n2681_), .Y(new_n8561_));
  NOR4X1   g06125(.A(new_n8561_), .B(new_n8559_), .C(new_n5254_), .D(new_n2682_), .Y(new_n8562_));
  OAI21X1  g06126(.A0(new_n8562_), .A1(new_n8558_), .B0(new_n5189_), .Y(new_n8563_));
  NAND2X1  g06127(.A(new_n8563_), .B(new_n2959_), .Y(new_n8564_));
  NOR4X1   g06128(.A(new_n5353_), .B(new_n5262_), .C(new_n5074_), .D(pi0216), .Y(new_n8565_));
  INVX1    g06129(.A(new_n8565_), .Y(new_n8566_));
  AND2X1   g06130(.A(new_n5261_), .B(new_n8518_), .Y(new_n8567_));
  AOI21X1  g06131(.A0(new_n8567_), .A1(new_n5963_), .B0(new_n2959_), .Y(new_n8568_));
  AOI21X1  g06132(.A0(new_n8568_), .A1(new_n8566_), .B0(new_n7690_), .Y(new_n8569_));
  AND2X1   g06133(.A(new_n8569_), .B(new_n8564_), .Y(po0230));
  AND2X1   g06134(.A(new_n8567_), .B(new_n6886_), .Y(new_n8571_));
  NAND3X1  g06135(.A(new_n6893_), .B(new_n5261_), .C(new_n8515_), .Y(new_n8572_));
  AND2X1   g06136(.A(new_n8572_), .B(pi0299), .Y(new_n8573_));
  INVX1    g06137(.A(new_n8573_), .Y(new_n8574_));
  OAI21X1  g06138(.A0(new_n8571_), .A1(pi0299), .B0(new_n8574_), .Y(new_n8575_));
  INVX1    g06139(.A(pi1050), .Y(new_n8576_));
  NAND4X1  g06140(.A(new_n7667_), .B(new_n6950_), .C(new_n6786_), .D(new_n2607_), .Y(new_n8577_));
  NOR3X1   g06141(.A(new_n8577_), .B(new_n8576_), .C(pi0314), .Y(new_n8578_));
  OAI21X1  g06142(.A0(new_n8578_), .A1(pi0039), .B0(new_n7689_), .Y(new_n8579_));
  AOI21X1  g06143(.A0(new_n8575_), .A1(pi0039), .B0(new_n8579_), .Y(po0231));
  NAND4X1  g06144(.A(new_n7674_), .B(new_n3109_), .C(pi0074), .D(new_n3112_), .Y(new_n8581_));
  OR4X1    g06145(.A(new_n5944_), .B(new_n2582_), .C(new_n2586_), .D(new_n2533_), .Y(new_n8582_));
  AND2X1   g06146(.A(new_n8582_), .B(new_n2526_), .Y(new_n8583_));
  NAND4X1  g06147(.A(new_n2783_), .B(new_n2756_), .C(pi0824), .D(new_n2526_), .Y(new_n8584_));
  AND2X1   g06148(.A(new_n5893_), .B(new_n3230_), .Y(new_n8585_));
  OAI21X1  g06149(.A0(new_n5019_), .A1(pi0096), .B0(pi0479), .Y(new_n8586_));
  NAND4X1  g06150(.A(new_n8586_), .B(new_n8585_), .C(new_n8584_), .D(new_n6773_), .Y(new_n8587_));
  OR4X1    g06151(.A(new_n8587_), .B(new_n8583_), .C(new_n5916_), .D(new_n3256_), .Y(new_n8588_));
  AOI21X1  g06152(.A0(new_n8588_), .A1(new_n8581_), .B0(po1038), .Y(po0232));
  OAI22X1  g06153(.A0(new_n8583_), .A1(new_n2782_), .B0(pi1093), .B1(new_n2526_), .Y(new_n8590_));
  NAND3X1  g06154(.A(new_n8590_), .B(new_n5949_), .C(new_n3091_), .Y(new_n8591_));
  NOR4X1   g06155(.A(new_n7673_), .B(new_n5788_), .C(new_n7672_), .D(new_n5787_), .Y(new_n8592_));
  OAI21X1  g06156(.A0(new_n8592_), .A1(new_n3095_), .B0(new_n6756_), .Y(new_n8593_));
  AOI21X1  g06157(.A0(new_n8591_), .A1(new_n3095_), .B0(new_n8593_), .Y(po0233));
  NOR4X1   g06158(.A(new_n2755_), .B(new_n5096_), .C(new_n5258_), .D(new_n3053_), .Y(new_n8595_));
  NOR4X1   g06159(.A(new_n8595_), .B(new_n7832_), .C(new_n3256_), .D(new_n2487_), .Y(new_n8596_));
  AND2X1   g06160(.A(new_n8596_), .B(new_n2453_), .Y(new_n8597_));
  AND2X1   g06161(.A(new_n2723_), .B(new_n2453_), .Y(new_n8598_));
  OAI21X1  g06162(.A0(new_n6790_), .A1(new_n2476_), .B0(new_n2590_), .Y(new_n8599_));
  NAND2X1  g06163(.A(new_n8599_), .B(new_n7667_), .Y(new_n8600_));
  AOI21X1  g06164(.A0(new_n7832_), .A1(new_n6789_), .B0(new_n8600_), .Y(new_n8601_));
  NOR2X1   g06165(.A(new_n8601_), .B(new_n2784_), .Y(new_n8602_));
  NOR4X1   g06166(.A(new_n7682_), .B(new_n6790_), .C(new_n2544_), .D(new_n3053_), .Y(new_n8603_));
  OR2X1    g06167(.A(new_n8603_), .B(new_n2785_), .Y(new_n8604_));
  AOI21X1  g06168(.A0(new_n8601_), .A1(new_n3053_), .B0(new_n8604_), .Y(new_n8605_));
  NOR2X1   g06169(.A(new_n8605_), .B(new_n8602_), .Y(new_n8606_));
  NOR2X1   g06170(.A(new_n8606_), .B(new_n5952_), .Y(new_n8607_));
  INVX1    g06171(.A(new_n8607_), .Y(new_n8608_));
  NOR3X1   g06172(.A(new_n8601_), .B(new_n5939_), .C(new_n2784_), .Y(new_n8609_));
  NOR3X1   g06173(.A(new_n7832_), .B(new_n3256_), .C(new_n2487_), .Y(new_n8610_));
  NOR2X1   g06174(.A(new_n8610_), .B(new_n5894_), .Y(new_n8611_));
  NOR3X1   g06175(.A(new_n8611_), .B(new_n8609_), .C(new_n8605_), .Y(new_n8612_));
  OAI21X1  g06176(.A0(new_n8612_), .A1(pi0122), .B0(new_n8608_), .Y(new_n8613_));
  OAI21X1  g06177(.A0(new_n8596_), .A1(pi0122), .B0(new_n8608_), .Y(new_n8614_));
  MX2X1    g06178(.A(new_n8614_), .B(new_n8613_), .S0(new_n2756_), .Y(new_n8615_));
  AOI21X1  g06179(.A0(new_n8615_), .A1(new_n2723_), .B0(new_n8598_), .Y(new_n8616_));
  NOR2X1   g06180(.A(new_n8601_), .B(new_n2756_), .Y(new_n8617_));
  NOR2X1   g06181(.A(new_n8617_), .B(new_n6256_), .Y(new_n8618_));
  AOI21X1  g06182(.A0(new_n8610_), .A1(new_n5952_), .B0(new_n8618_), .Y(new_n8619_));
  AOI21X1  g06183(.A0(new_n8613_), .A1(new_n2756_), .B0(new_n8619_), .Y(new_n8620_));
  NOR2X1   g06184(.A(new_n8620_), .B(new_n2723_), .Y(new_n8621_));
  AOI21X1  g06185(.A0(new_n2724_), .A1(new_n2453_), .B0(new_n8621_), .Y(new_n8622_));
  NAND2X1  g06186(.A(pi1092), .B(pi0252), .Y(new_n8623_));
  NOR2X1   g06187(.A(new_n8623_), .B(pi1093), .Y(new_n8624_));
  INVX1    g06188(.A(new_n8624_), .Y(new_n8625_));
  OAI21X1  g06189(.A0(new_n8625_), .A1(new_n2738_), .B0(new_n2453_), .Y(new_n8626_));
  NOR4X1   g06190(.A(new_n8626_), .B(new_n7832_), .C(new_n3256_), .D(new_n2487_), .Y(new_n8627_));
  OAI22X1  g06191(.A0(new_n8627_), .A1(new_n8622_), .B0(new_n8616_), .B1(new_n8597_), .Y(new_n8628_));
  OR4X1    g06192(.A(new_n7682_), .B(new_n7632_), .C(new_n6790_), .D(new_n2544_), .Y(new_n8629_));
  NOR2X1   g06193(.A(new_n5094_), .B(pi0137), .Y(new_n8630_));
  AOI21X1  g06194(.A0(new_n8629_), .A1(po1057), .B0(new_n8630_), .Y(new_n8631_));
  INVX1    g06195(.A(new_n8631_), .Y(new_n8632_));
  AOI21X1  g06196(.A0(new_n8628_), .A1(new_n5094_), .B0(new_n8632_), .Y(new_n8633_));
  AND2X1   g06197(.A(new_n8615_), .B(new_n2723_), .Y(new_n8634_));
  OR2X1    g06198(.A(new_n8621_), .B(new_n8634_), .Y(new_n8635_));
  MX2X1    g06199(.A(new_n8629_), .B(new_n8635_), .S0(new_n5094_), .Y(new_n8636_));
  INVX1    g06200(.A(new_n8636_), .Y(new_n8637_));
  MX2X1    g06201(.A(new_n8637_), .B(new_n8633_), .S0(new_n2766_), .Y(new_n8638_));
  AND2X1   g06202(.A(new_n7783_), .B(new_n4515_), .Y(new_n8639_));
  MX2X1    g06203(.A(new_n8635_), .B(new_n8628_), .S0(new_n2766_), .Y(new_n8640_));
  AOI21X1  g06204(.A0(new_n8640_), .A1(new_n8639_), .B0(new_n2953_), .Y(new_n8641_));
  OAI21X1  g06205(.A0(new_n8639_), .A1(new_n8638_), .B0(new_n8641_), .Y(new_n8642_));
  MX2X1    g06206(.A(new_n8637_), .B(new_n8633_), .S0(new_n2973_), .Y(new_n8643_));
  AND2X1   g06207(.A(new_n5033_), .B(new_n2980_), .Y(new_n8644_));
  MX2X1    g06208(.A(new_n8635_), .B(new_n8628_), .S0(new_n2973_), .Y(new_n8645_));
  AOI21X1  g06209(.A0(new_n8645_), .A1(new_n8644_), .B0(pi0299), .Y(new_n8646_));
  OAI21X1  g06210(.A0(new_n8644_), .A1(new_n8643_), .B0(new_n8646_), .Y(new_n8647_));
  AOI21X1  g06211(.A0(new_n8647_), .A1(new_n8642_), .B0(new_n5237_), .Y(new_n8648_));
  NOR2X1   g06212(.A(new_n8638_), .B(new_n2953_), .Y(new_n8649_));
  OAI21X1  g06213(.A0(new_n8643_), .A1(pi0299), .B0(new_n5237_), .Y(new_n8650_));
  NOR2X1   g06214(.A(new_n8650_), .B(new_n8649_), .Y(new_n8651_));
  OAI21X1  g06215(.A0(new_n8651_), .A1(new_n8648_), .B0(new_n6077_), .Y(new_n8652_));
  INVX1    g06216(.A(new_n7630_), .Y(new_n8653_));
  OR2X1    g06217(.A(new_n8610_), .B(new_n2785_), .Y(new_n8654_));
  MX2X1    g06218(.A(new_n8601_), .B(new_n3053_), .S0(new_n2784_), .Y(new_n8655_));
  AND2X1   g06219(.A(new_n8655_), .B(new_n8654_), .Y(new_n8656_));
  OAI22X1  g06220(.A0(new_n8656_), .A1(new_n6259_), .B0(new_n8606_), .B1(new_n5952_), .Y(new_n8657_));
  INVX1    g06221(.A(new_n8657_), .Y(new_n8658_));
  NOR2X1   g06222(.A(new_n8606_), .B(pi1093), .Y(new_n8659_));
  AOI21X1  g06223(.A0(new_n8617_), .A1(new_n2724_), .B0(new_n8659_), .Y(new_n8660_));
  OAI21X1  g06224(.A0(new_n8658_), .A1(new_n2724_), .B0(new_n8660_), .Y(new_n8661_));
  INVX1    g06225(.A(new_n8661_), .Y(new_n8662_));
  NOR4X1   g06226(.A(new_n7682_), .B(new_n6790_), .C(new_n5094_), .D(new_n2544_), .Y(new_n8663_));
  AOI22X1  g06227(.A0(new_n8663_), .A1(new_n8653_), .B0(new_n8662_), .B1(new_n5094_), .Y(new_n8664_));
  NOR3X1   g06228(.A(new_n8606_), .B(pi1093), .C(new_n2453_), .Y(new_n8665_));
  AOI21X1  g06229(.A0(new_n8655_), .A1(new_n8654_), .B0(pi0137), .Y(new_n8666_));
  AND2X1   g06230(.A(new_n8666_), .B(new_n2756_), .Y(new_n8667_));
  NOR4X1   g06231(.A(new_n8667_), .B(new_n8665_), .C(new_n8617_), .D(po1057), .Y(new_n8668_));
  OR2X1    g06232(.A(new_n8668_), .B(new_n8663_), .Y(new_n8669_));
  AOI21X1  g06233(.A0(new_n8630_), .A1(new_n6772_), .B0(new_n2723_), .Y(new_n8670_));
  AND2X1   g06234(.A(new_n8657_), .B(pi0137), .Y(new_n8671_));
  OR2X1    g06235(.A(new_n8666_), .B(new_n8665_), .Y(new_n8672_));
  OAI21X1  g06236(.A0(new_n8672_), .A1(new_n8671_), .B0(new_n5094_), .Y(new_n8673_));
  AOI21X1  g06237(.A0(new_n6259_), .A1(pi0137), .B0(new_n2785_), .Y(new_n8674_));
  OR4X1    g06238(.A(new_n8674_), .B(new_n7682_), .C(new_n6790_), .D(new_n2544_), .Y(new_n8675_));
  AOI21X1  g06239(.A0(new_n8675_), .A1(po1057), .B0(new_n2724_), .Y(new_n8676_));
  AOI22X1  g06240(.A0(new_n8676_), .A1(new_n8673_), .B0(new_n8670_), .B1(new_n8669_), .Y(new_n8677_));
  MX2X1    g06241(.A(new_n8677_), .B(new_n8664_), .S0(pi0210), .Y(new_n8678_));
  NOR4X1   g06242(.A(new_n8667_), .B(new_n8665_), .C(new_n8617_), .D(new_n2723_), .Y(new_n8679_));
  NOR3X1   g06243(.A(new_n8672_), .B(new_n8671_), .C(new_n2724_), .Y(new_n8680_));
  OR2X1    g06244(.A(new_n8680_), .B(new_n8679_), .Y(new_n8681_));
  INVX1    g06245(.A(new_n8639_), .Y(new_n8682_));
  AOI21X1  g06246(.A0(new_n8661_), .A1(pi0210), .B0(new_n8682_), .Y(new_n8683_));
  OAI21X1  g06247(.A0(new_n8681_), .A1(pi0210), .B0(new_n8683_), .Y(new_n8684_));
  AND2X1   g06248(.A(new_n8684_), .B(pi0299), .Y(new_n8685_));
  OAI21X1  g06249(.A0(new_n8678_), .A1(new_n8639_), .B0(new_n8685_), .Y(new_n8686_));
  MX2X1    g06250(.A(new_n8677_), .B(new_n8664_), .S0(pi0198), .Y(new_n8687_));
  MX2X1    g06251(.A(new_n8681_), .B(new_n8662_), .S0(pi0198), .Y(new_n8688_));
  AOI21X1  g06252(.A0(new_n8688_), .A1(new_n8644_), .B0(pi0299), .Y(new_n8689_));
  OAI21X1  g06253(.A0(new_n8687_), .A1(new_n8644_), .B0(new_n8689_), .Y(new_n8690_));
  AOI21X1  g06254(.A0(new_n8690_), .A1(new_n8686_), .B0(new_n5237_), .Y(new_n8691_));
  NOR2X1   g06255(.A(new_n8687_), .B(pi0299), .Y(new_n8692_));
  OAI21X1  g06256(.A0(new_n8678_), .A1(new_n2953_), .B0(new_n5237_), .Y(new_n8693_));
  OAI21X1  g06257(.A0(new_n8693_), .A1(new_n8692_), .B0(new_n6633_), .Y(new_n8694_));
  OR2X1    g06258(.A(new_n8694_), .B(new_n8691_), .Y(new_n8695_));
  AOI21X1  g06259(.A0(new_n8695_), .A1(new_n8652_), .B0(new_n7749_), .Y(po0234));
  OR4X1    g06260(.A(new_n2591_), .B(new_n2579_), .C(new_n2577_), .D(new_n2581_), .Y(new_n8697_));
  AND2X1   g06261(.A(new_n8697_), .B(new_n2474_), .Y(new_n8698_));
  NOR4X1   g06262(.A(new_n8698_), .B(new_n2598_), .C(new_n2477_), .D(pi0046), .Y(new_n8699_));
  NAND4X1  g06263(.A(new_n8699_), .B(new_n2483_), .C(new_n2482_), .D(new_n2481_), .Y(new_n8700_));
  NOR4X1   g06264(.A(new_n6789_), .B(new_n2593_), .C(new_n2591_), .D(new_n2474_), .Y(new_n8701_));
  OAI21X1  g06265(.A0(new_n8701_), .A1(new_n7734_), .B0(new_n7669_), .Y(new_n8702_));
  AOI21X1  g06266(.A0(new_n8700_), .A1(new_n7734_), .B0(new_n8702_), .Y(po0235));
  NOR3X1   g06267(.A(pi0468), .B(new_n5237_), .C(new_n5862_), .Y(po0236));
  INVX1    g06268(.A(pi0163), .Y(new_n8705_));
  OR2X1    g06269(.A(new_n7348_), .B(pi0163), .Y(new_n8706_));
  OAI22X1  g06270(.A0(new_n8706_), .A1(new_n7350_), .B0(new_n7351_), .B1(new_n8705_), .Y(new_n8707_));
  NOR2X1   g06271(.A(new_n8707_), .B(new_n5237_), .Y(new_n8708_));
  AOI21X1  g06272(.A0(new_n3026_), .A1(new_n3095_), .B0(new_n8708_), .Y(new_n8709_));
  INVX1    g06273(.A(pi0147), .Y(new_n8710_));
  NOR4X1   g06274(.A(pi0468), .B(pi0332), .C(new_n5237_), .D(new_n8710_), .Y(new_n8711_));
  AND2X1   g06275(.A(new_n8711_), .B(new_n6828_), .Y(new_n8712_));
  AOI21X1  g06276(.A0(new_n8708_), .A1(new_n6832_), .B0(new_n4991_), .Y(new_n8713_));
  OR4X1    g06277(.A(new_n8713_), .B(new_n8712_), .C(new_n8709_), .D(new_n3246_), .Y(new_n8714_));
  NOR2X1   g06278(.A(new_n7371_), .B(new_n6837_), .Y(new_n8715_));
  NOR4X1   g06279(.A(new_n7372_), .B(new_n8715_), .C(new_n5057_), .D(pi0184), .Y(new_n8716_));
  INVX1    g06280(.A(pi0184), .Y(new_n8717_));
  NOR3X1   g06281(.A(new_n7372_), .B(new_n8715_), .C(new_n5057_), .Y(new_n8718_));
  NOR3X1   g06282(.A(new_n8718_), .B(new_n5057_), .C(new_n8717_), .Y(new_n8719_));
  NOR3X1   g06283(.A(new_n8719_), .B(new_n8716_), .C(pi0299), .Y(new_n8720_));
  OR2X1    g06284(.A(new_n8720_), .B(new_n5237_), .Y(new_n8721_));
  AOI21X1  g06285(.A0(new_n8707_), .A1(pi0299), .B0(new_n8721_), .Y(new_n8722_));
  AOI21X1  g06286(.A0(new_n8722_), .A1(new_n6832_), .B0(new_n4991_), .Y(new_n8723_));
  NOR2X1   g06287(.A(new_n8723_), .B(pi0055), .Y(new_n8724_));
  MX2X1    g06288(.A(pi0187), .B(pi0147), .S0(pi0299), .Y(new_n8725_));
  AND2X1   g06289(.A(new_n8725_), .B(new_n5930_), .Y(new_n8726_));
  OAI21X1  g06290(.A0(new_n8726_), .A1(new_n6832_), .B0(pi0054), .Y(new_n8727_));
  AOI21X1  g06291(.A0(new_n8722_), .A1(new_n6832_), .B0(new_n8727_), .Y(new_n8728_));
  INVX1    g06292(.A(pi0187), .Y(new_n8729_));
  OAI21X1  g06293(.A0(new_n7490_), .A1(new_n8729_), .B0(pi0147), .Y(new_n8730_));
  AOI21X1  g06294(.A0(new_n7489_), .A1(new_n8729_), .B0(new_n8730_), .Y(new_n8731_));
  NOR4X1   g06295(.A(new_n6862_), .B(new_n4995_), .C(new_n8729_), .D(pi0147), .Y(new_n8732_));
  OAI21X1  g06296(.A0(new_n8732_), .A1(new_n8731_), .B0(pi0038), .Y(new_n8733_));
  INVX1    g06297(.A(pi0153), .Y(new_n8734_));
  OAI21X1  g06298(.A0(new_n7004_), .A1(pi0040), .B0(new_n2540_), .Y(new_n8735_));
  NOR3X1   g06299(.A(new_n7015_), .B(new_n4464_), .C(pi0040), .Y(new_n8736_));
  NOR2X1   g06300(.A(new_n8736_), .B(new_n8735_), .Y(new_n8737_));
  OR2X1    g06301(.A(new_n7049_), .B(new_n5057_), .Y(new_n8738_));
  OAI21X1  g06302(.A0(new_n8738_), .A1(new_n8737_), .B0(new_n8734_), .Y(new_n8739_));
  NOR2X1   g06303(.A(new_n7059_), .B(pi0040), .Y(new_n8740_));
  OAI21X1  g06304(.A0(new_n8740_), .A1(pi0095), .B0(pi0166), .Y(new_n8741_));
  AND2X1   g06305(.A(new_n2472_), .B(new_n2549_), .Y(new_n8742_));
  AOI21X1  g06306(.A0(new_n7783_), .A1(new_n8742_), .B0(new_n8734_), .Y(new_n8743_));
  OAI21X1  g06307(.A0(new_n8741_), .A1(new_n8738_), .B0(new_n8743_), .Y(new_n8744_));
  AND2X1   g06308(.A(new_n8744_), .B(pi0160), .Y(new_n8745_));
  NOR3X1   g06309(.A(new_n8736_), .B(new_n8735_), .C(pi0153), .Y(new_n8746_));
  INVX1    g06310(.A(pi0160), .Y(new_n8747_));
  AOI22X1  g06311(.A0(new_n7093_), .A1(new_n2899_), .B0(new_n6933_), .B1(new_n6930_), .Y(new_n8748_));
  INVX1    g06312(.A(new_n8748_), .Y(new_n8749_));
  OAI21X1  g06313(.A0(new_n8740_), .A1(pi0095), .B0(new_n8577_), .Y(new_n8750_));
  NAND3X1  g06314(.A(new_n8750_), .B(new_n8741_), .C(pi0153), .Y(new_n8751_));
  NAND4X1  g06315(.A(new_n8751_), .B(new_n8749_), .C(new_n5033_), .D(new_n8747_), .Y(new_n8752_));
  OAI21X1  g06316(.A0(new_n8752_), .A1(new_n8746_), .B0(pi0163), .Y(new_n8753_));
  AOI21X1  g06317(.A0(new_n8745_), .A1(new_n8739_), .B0(new_n8753_), .Y(new_n8754_));
  OAI21X1  g06318(.A0(new_n7108_), .A1(new_n7115_), .B0(new_n2549_), .Y(new_n8755_));
  AOI21X1  g06319(.A0(new_n8755_), .A1(new_n2540_), .B0(new_n8748_), .Y(new_n8756_));
  INVX1    g06320(.A(new_n8756_), .Y(new_n8757_));
  OAI21X1  g06321(.A0(new_n6985_), .A1(pi0040), .B0(new_n2456_), .Y(new_n8758_));
  AOI21X1  g06322(.A0(new_n8758_), .A1(new_n7033_), .B0(pi0095), .Y(new_n8759_));
  OAI21X1  g06323(.A0(new_n8759_), .A1(new_n8748_), .B0(pi0210), .Y(new_n8760_));
  AOI21X1  g06324(.A0(new_n8758_), .A1(new_n7050_), .B0(pi0095), .Y(new_n8761_));
  OR2X1    g06325(.A(new_n8761_), .B(new_n8748_), .Y(new_n8762_));
  AOI21X1  g06326(.A0(new_n8762_), .A1(new_n2766_), .B0(new_n7784_), .Y(new_n8763_));
  AOI21X1  g06327(.A0(new_n8763_), .A1(new_n8760_), .B0(pi0153), .Y(new_n8764_));
  OAI21X1  g06328(.A0(new_n8757_), .A1(new_n4464_), .B0(new_n8764_), .Y(new_n8765_));
  AOI21X1  g06329(.A0(new_n7041_), .A1(new_n7033_), .B0(pi0095), .Y(new_n8766_));
  OAI21X1  g06330(.A0(new_n8766_), .A1(new_n8748_), .B0(pi0210), .Y(new_n8767_));
  OAI21X1  g06331(.A0(new_n8748_), .A1(new_n7051_), .B0(new_n2766_), .Y(new_n8768_));
  AND2X1   g06332(.A(new_n5033_), .B(pi0166), .Y(new_n8769_));
  NAND3X1  g06333(.A(new_n8769_), .B(new_n8768_), .C(new_n8767_), .Y(new_n8770_));
  AOI21X1  g06334(.A0(new_n8749_), .A1(new_n7098_), .B0(pi0210), .Y(new_n8771_));
  AOI21X1  g06335(.A0(new_n8749_), .A1(new_n7095_), .B0(new_n2766_), .Y(new_n8772_));
  OR4X1    g06336(.A(new_n8772_), .B(new_n8771_), .C(new_n5057_), .D(pi0166), .Y(new_n8773_));
  AND2X1   g06337(.A(new_n8773_), .B(pi0153), .Y(new_n8774_));
  AOI21X1  g06338(.A0(new_n8774_), .A1(new_n8770_), .B0(pi0160), .Y(new_n8775_));
  INVX1    g06339(.A(new_n8769_), .Y(new_n8776_));
  NOR2X1   g06340(.A(new_n8776_), .B(new_n8755_), .Y(new_n8777_));
  NOR2X1   g06341(.A(new_n8761_), .B(new_n7049_), .Y(new_n8778_));
  NOR2X1   g06342(.A(new_n8778_), .B(pi0210), .Y(new_n8779_));
  OAI21X1  g06343(.A0(new_n8759_), .A1(new_n7049_), .B0(pi0210), .Y(new_n8780_));
  NAND2X1  g06344(.A(new_n8780_), .B(new_n7783_), .Y(new_n8781_));
  OAI21X1  g06345(.A0(new_n8781_), .A1(new_n8779_), .B0(new_n8734_), .Y(new_n8782_));
  NOR2X1   g06346(.A(new_n8782_), .B(new_n8777_), .Y(new_n8783_));
  AOI21X1  g06347(.A0(new_n7095_), .A1(new_n7093_), .B0(new_n2766_), .Y(new_n8784_));
  AOI21X1  g06348(.A0(new_n7098_), .A1(new_n7093_), .B0(pi0210), .Y(new_n8785_));
  NOR3X1   g06349(.A(new_n8785_), .B(new_n8784_), .C(new_n7784_), .Y(new_n8786_));
  AND2X1   g06350(.A(new_n7052_), .B(new_n2766_), .Y(new_n8787_));
  NOR2X1   g06351(.A(new_n8766_), .B(new_n7049_), .Y(new_n8788_));
  OAI21X1  g06352(.A0(new_n8788_), .A1(new_n2766_), .B0(new_n8769_), .Y(new_n8789_));
  OAI21X1  g06353(.A0(new_n8789_), .A1(new_n8787_), .B0(pi0153), .Y(new_n8790_));
  OAI21X1  g06354(.A0(new_n8790_), .A1(new_n8786_), .B0(pi0160), .Y(new_n8791_));
  OAI21X1  g06355(.A0(new_n8791_), .A1(new_n8783_), .B0(new_n8705_), .Y(new_n8792_));
  AOI21X1  g06356(.A0(new_n8775_), .A1(new_n8765_), .B0(new_n8792_), .Y(new_n8793_));
  AOI21X1  g06357(.A0(new_n8756_), .A1(new_n5057_), .B0(new_n2953_), .Y(new_n8794_));
  OAI21X1  g06358(.A0(new_n8793_), .A1(new_n8754_), .B0(new_n8794_), .Y(new_n8795_));
  AOI21X1  g06359(.A0(new_n7026_), .A1(new_n6977_), .B0(pi0040), .Y(new_n8796_));
  OAI21X1  g06360(.A0(new_n8796_), .A1(pi0095), .B0(new_n8749_), .Y(new_n8797_));
  OR2X1    g06361(.A(new_n8797_), .B(new_n5033_), .Y(new_n8798_));
  NOR2X1   g06362(.A(pi0299), .B(pi0175), .Y(new_n8799_));
  INVX1    g06363(.A(new_n8799_), .Y(new_n8800_));
  NOR3X1   g06364(.A(new_n7015_), .B(new_n7942_), .C(pi0040), .Y(new_n8801_));
  OAI21X1  g06365(.A0(new_n7093_), .A1(new_n5227_), .B0(new_n5033_), .Y(new_n8802_));
  AOI21X1  g06366(.A0(new_n8748_), .A1(new_n5227_), .B0(new_n8802_), .Y(new_n8803_));
  OAI21X1  g06367(.A0(new_n8801_), .A1(new_n8735_), .B0(new_n8803_), .Y(new_n8804_));
  AND2X1   g06368(.A(new_n5033_), .B(pi0189), .Y(new_n8805_));
  NAND2X1  g06369(.A(new_n8805_), .B(new_n8796_), .Y(new_n8806_));
  OAI21X1  g06370(.A0(new_n8761_), .A1(new_n7049_), .B0(new_n2973_), .Y(new_n8807_));
  OAI21X1  g06371(.A0(new_n8759_), .A1(new_n7049_), .B0(pi0198), .Y(new_n8808_));
  NAND3X1  g06372(.A(new_n8808_), .B(new_n8807_), .C(new_n7780_), .Y(new_n8809_));
  AND2X1   g06373(.A(new_n8717_), .B(pi0182), .Y(new_n8810_));
  AND2X1   g06374(.A(new_n8810_), .B(new_n8809_), .Y(new_n8811_));
  AOI22X1  g06375(.A0(new_n8811_), .A1(new_n8806_), .B0(new_n8804_), .B1(pi0184), .Y(new_n8812_));
  INVX1    g06376(.A(new_n7780_), .Y(new_n8813_));
  NOR3X1   g06377(.A(new_n8813_), .B(new_n7099_), .C(new_n7096_), .Y(new_n8814_));
  AND2X1   g06378(.A(new_n7052_), .B(new_n2973_), .Y(new_n8815_));
  OAI21X1  g06379(.A0(new_n8788_), .A1(new_n2973_), .B0(new_n8805_), .Y(new_n8816_));
  OAI21X1  g06380(.A0(new_n8816_), .A1(new_n8815_), .B0(pi0182), .Y(new_n8817_));
  NOR2X1   g06381(.A(new_n8748_), .B(new_n7051_), .Y(new_n8818_));
  NOR2X1   g06382(.A(new_n8818_), .B(pi0198), .Y(new_n8819_));
  OAI21X1  g06383(.A0(new_n8766_), .A1(new_n8748_), .B0(pi0198), .Y(new_n8820_));
  NAND2X1  g06384(.A(new_n8820_), .B(new_n8805_), .Y(new_n8821_));
  OAI21X1  g06385(.A0(new_n8821_), .A1(new_n8819_), .B0(new_n5227_), .Y(new_n8822_));
  OAI21X1  g06386(.A0(new_n8817_), .A1(new_n8814_), .B0(new_n8822_), .Y(new_n8823_));
  AND2X1   g06387(.A(new_n5227_), .B(pi0095), .Y(new_n8824_));
  NOR2X1   g06388(.A(new_n8748_), .B(new_n8813_), .Y(new_n8825_));
  OAI21X1  g06389(.A0(new_n8824_), .A1(new_n7100_), .B0(new_n8825_), .Y(new_n8826_));
  AOI21X1  g06390(.A0(new_n8826_), .A1(new_n8823_), .B0(pi0184), .Y(new_n8827_));
  AND2X1   g06391(.A(new_n2953_), .B(pi0175), .Y(new_n8828_));
  INVX1    g06392(.A(new_n8828_), .Y(new_n8829_));
  AND2X1   g06393(.A(new_n5033_), .B(pi0184), .Y(new_n8830_));
  AOI21X1  g06394(.A0(pi0189), .A1(new_n2540_), .B0(new_n2472_), .Y(new_n8831_));
  NOR3X1   g06395(.A(new_n8831_), .B(new_n7059_), .C(pi0040), .Y(new_n8832_));
  OAI21X1  g06396(.A0(new_n8832_), .A1(new_n8824_), .B0(new_n8830_), .Y(new_n8833_));
  AOI21X1  g06397(.A0(new_n8748_), .A1(new_n5227_), .B0(new_n8833_), .Y(new_n8834_));
  OR2X1    g06398(.A(new_n8834_), .B(new_n8829_), .Y(new_n8835_));
  OAI22X1  g06399(.A0(new_n8835_), .A1(new_n8827_), .B0(new_n8812_), .B1(new_n8800_), .Y(new_n8836_));
  OR2X1    g06400(.A(new_n8797_), .B(new_n7780_), .Y(new_n8837_));
  OAI21X1  g06401(.A0(new_n8759_), .A1(new_n8748_), .B0(pi0198), .Y(new_n8838_));
  AOI21X1  g06402(.A0(new_n8762_), .A1(new_n2973_), .B0(new_n8813_), .Y(new_n8839_));
  OR4X1    g06403(.A(pi0299), .B(pi0184), .C(pi0182), .D(pi0175), .Y(new_n8840_));
  AOI21X1  g06404(.A0(new_n8839_), .A1(new_n8838_), .B0(new_n8840_), .Y(new_n8841_));
  AOI22X1  g06405(.A0(new_n8841_), .A1(new_n8837_), .B0(new_n8836_), .B1(new_n8798_), .Y(new_n8842_));
  AOI21X1  g06406(.A0(new_n8842_), .A1(new_n8795_), .B0(new_n5237_), .Y(new_n8843_));
  NOR2X1   g06407(.A(new_n8797_), .B(pi0299), .Y(new_n8844_));
  OAI21X1  g06408(.A0(new_n8757_), .A1(new_n2953_), .B0(new_n5237_), .Y(new_n8845_));
  OAI21X1  g06409(.A0(new_n8845_), .A1(new_n8844_), .B0(new_n2959_), .Y(new_n8846_));
  NOR2X1   g06410(.A(new_n8742_), .B(new_n6886_), .Y(new_n8847_));
  NOR2X1   g06411(.A(new_n6885_), .B(pi0040), .Y(new_n8848_));
  NOR2X1   g06412(.A(new_n8848_), .B(pi0189), .Y(new_n8849_));
  OR2X1    g06413(.A(new_n6907_), .B(new_n2472_), .Y(new_n8850_));
  AND2X1   g06414(.A(new_n8850_), .B(new_n7025_), .Y(new_n8851_));
  AOI21X1  g06415(.A0(new_n6897_), .A1(new_n2607_), .B0(pi0040), .Y(new_n8852_));
  AOI22X1  g06416(.A0(new_n8852_), .A1(new_n6269_), .B0(new_n8742_), .B1(new_n5052_), .Y(new_n8853_));
  INVX1    g06417(.A(new_n8853_), .Y(new_n8854_));
  NOR4X1   g06418(.A(new_n8854_), .B(new_n8851_), .C(new_n5050_), .D(new_n7942_), .Y(new_n8855_));
  OAI21X1  g06419(.A0(new_n8855_), .A1(new_n8849_), .B0(pi0179), .Y(new_n8856_));
  OAI21X1  g06420(.A0(new_n6901_), .A1(new_n2472_), .B0(new_n7025_), .Y(new_n8857_));
  AOI21X1  g06421(.A0(new_n8857_), .A1(new_n8853_), .B0(pi0189), .Y(new_n8858_));
  MX2X1    g06422(.A(new_n8852_), .B(new_n8742_), .S0(new_n5052_), .Y(new_n8859_));
  INVX1    g06423(.A(new_n8859_), .Y(new_n8860_));
  AOI21X1  g06424(.A0(new_n5049_), .A1(new_n5048_), .B0(pi0179), .Y(new_n8861_));
  OAI21X1  g06425(.A0(new_n8860_), .A1(new_n7942_), .B0(new_n8861_), .Y(new_n8862_));
  OAI22X1  g06426(.A0(new_n8862_), .A1(new_n8858_), .B0(new_n8848_), .B1(new_n5051_), .Y(new_n8863_));
  INVX1    g06427(.A(new_n8863_), .Y(new_n8864_));
  AOI21X1  g06428(.A0(new_n8864_), .A1(new_n8856_), .B0(new_n6913_), .Y(new_n8865_));
  OAI21X1  g06429(.A0(new_n8865_), .A1(new_n8847_), .B0(new_n2953_), .Y(new_n8866_));
  INVX1    g06430(.A(new_n8866_), .Y(new_n8867_));
  NOR3X1   g06431(.A(new_n6893_), .B(new_n2607_), .C(pi0040), .Y(new_n8868_));
  OR2X1    g06432(.A(new_n8868_), .B(new_n2953_), .Y(new_n8869_));
  INVX1    g06433(.A(new_n8848_), .Y(new_n8870_));
  MX2X1    g06434(.A(new_n8860_), .B(new_n8870_), .S0(new_n5070_), .Y(new_n8871_));
  OAI21X1  g06435(.A0(new_n5070_), .A1(pi0166), .B0(new_n8871_), .Y(new_n8872_));
  NAND4X1  g06436(.A(new_n8857_), .B(new_n8853_), .C(new_n5071_), .D(new_n4464_), .Y(new_n8873_));
  AND2X1   g06437(.A(new_n8873_), .B(new_n6893_), .Y(new_n8874_));
  AOI21X1  g06438(.A0(new_n8874_), .A1(new_n8872_), .B0(new_n8869_), .Y(new_n8875_));
  INVX1    g06439(.A(pi0156), .Y(new_n8876_));
  AND2X1   g06440(.A(pi0232), .B(new_n8876_), .Y(new_n8877_));
  OAI21X1  g06441(.A0(new_n8875_), .A1(new_n8867_), .B0(new_n8877_), .Y(new_n8878_));
  NOR4X1   g06442(.A(new_n8854_), .B(new_n8851_), .C(new_n5070_), .D(new_n4464_), .Y(new_n8879_));
  AOI21X1  g06443(.A0(new_n5071_), .A1(pi0166), .B0(new_n8848_), .Y(new_n8880_));
  NOR3X1   g06444(.A(new_n8880_), .B(new_n8879_), .C(new_n6905_), .Y(new_n8881_));
  OAI21X1  g06445(.A0(new_n8881_), .A1(new_n8869_), .B0(new_n8866_), .Y(new_n8882_));
  AND2X1   g06446(.A(pi0232), .B(pi0156), .Y(new_n8883_));
  MX2X1    g06447(.A(new_n8860_), .B(new_n8870_), .S0(new_n5050_), .Y(new_n8884_));
  OAI21X1  g06448(.A0(new_n8742_), .A1(new_n6886_), .B0(new_n2953_), .Y(new_n8885_));
  AOI21X1  g06449(.A0(new_n8884_), .A1(new_n6886_), .B0(new_n8885_), .Y(new_n8886_));
  OAI21X1  g06450(.A0(new_n8871_), .A1(new_n6922_), .B0(new_n5237_), .Y(new_n8887_));
  OAI21X1  g06451(.A0(new_n8887_), .A1(new_n8886_), .B0(pi0039), .Y(new_n8888_));
  AOI21X1  g06452(.A0(new_n8883_), .A1(new_n8882_), .B0(new_n8888_), .Y(new_n8889_));
  AOI21X1  g06453(.A0(new_n8889_), .A1(new_n8878_), .B0(pi0038), .Y(new_n8890_));
  OAI21X1  g06454(.A0(new_n8846_), .A1(new_n8843_), .B0(new_n8890_), .Y(new_n8891_));
  AOI21X1  g06455(.A0(new_n8891_), .A1(new_n8733_), .B0(new_n3124_), .Y(new_n8892_));
  OAI21X1  g06456(.A0(new_n8726_), .A1(new_n2996_), .B0(new_n3026_), .Y(new_n8893_));
  NOR2X1   g06457(.A(pi0040), .B(pi0038), .Y(new_n8894_));
  INVX1    g06458(.A(new_n8894_), .Y(new_n8895_));
  NOR3X1   g06459(.A(new_n8895_), .B(new_n2607_), .C(new_n3156_), .Y(new_n8896_));
  OR2X1    g06460(.A(new_n8896_), .B(new_n8893_), .Y(new_n8897_));
  OAI22X1  g06461(.A0(new_n8897_), .A1(new_n3156_), .B0(new_n8722_), .B1(new_n3026_), .Y(new_n8898_));
  OAI21X1  g06462(.A0(new_n8898_), .A1(new_n8892_), .B0(new_n3105_), .Y(new_n8899_));
  NOR2X1   g06463(.A(new_n8722_), .B(new_n3095_), .Y(new_n8900_));
  OR2X1    g06464(.A(new_n8722_), .B(new_n3026_), .Y(new_n8901_));
  OAI21X1  g06465(.A0(new_n8742_), .A1(new_n2959_), .B0(new_n7320_), .Y(new_n8902_));
  AOI21X1  g06466(.A0(new_n6880_), .A1(new_n2607_), .B0(pi0040), .Y(new_n8903_));
  MX2X1    g06467(.A(pi0179), .B(pi0156), .S0(pi0299), .Y(new_n8904_));
  NAND3X1  g06468(.A(new_n8904_), .B(new_n5033_), .C(pi0232), .Y(new_n8905_));
  OAI21X1  g06469(.A0(new_n8905_), .A1(new_n2472_), .B0(new_n8903_), .Y(new_n8906_));
  AOI21X1  g06470(.A0(new_n8906_), .A1(new_n2959_), .B0(new_n8902_), .Y(new_n8907_));
  OAI21X1  g06471(.A0(new_n8907_), .A1(new_n8897_), .B0(new_n8901_), .Y(new_n8908_));
  AOI21X1  g06472(.A0(new_n8908_), .A1(new_n7185_), .B0(new_n8900_), .Y(new_n8909_));
  AOI21X1  g06473(.A0(new_n8909_), .A1(new_n8899_), .B0(pi0054), .Y(new_n8910_));
  OAI21X1  g06474(.A0(new_n8910_), .A1(new_n8728_), .B0(new_n4991_), .Y(new_n8911_));
  OR2X1    g06475(.A(new_n8713_), .B(new_n3128_), .Y(new_n8912_));
  OAI21X1  g06476(.A0(new_n8712_), .A1(new_n8709_), .B0(pi0054), .Y(new_n8913_));
  OAI21X1  g06477(.A0(new_n8707_), .A1(new_n5237_), .B0(pi0100), .Y(new_n8914_));
  AOI21X1  g06478(.A0(new_n6879_), .A1(new_n5057_), .B0(new_n6870_), .Y(new_n8915_));
  NAND3X1  g06479(.A(new_n8915_), .B(pi0232), .C(pi0163), .Y(new_n8916_));
  AOI21X1  g06480(.A0(new_n8916_), .A1(new_n8903_), .B0(pi0039), .Y(new_n8917_));
  OAI21X1  g06481(.A0(new_n8711_), .A1(new_n2996_), .B0(new_n3026_), .Y(new_n8918_));
  NOR2X1   g06482(.A(new_n8918_), .B(new_n8896_), .Y(new_n8919_));
  OAI21X1  g06483(.A0(new_n8917_), .A1(new_n8902_), .B0(new_n8919_), .Y(new_n8920_));
  AOI21X1  g06484(.A0(new_n8920_), .A1(new_n8914_), .B0(new_n5315_), .Y(new_n8921_));
  OAI21X1  g06485(.A0(new_n8918_), .A1(new_n8894_), .B0(new_n8914_), .Y(new_n8922_));
  OAI21X1  g06486(.A0(new_n8922_), .A1(new_n7180_), .B0(new_n7185_), .Y(new_n8923_));
  OAI21X1  g06487(.A0(new_n8708_), .A1(new_n3095_), .B0(new_n8923_), .Y(new_n8924_));
  OAI21X1  g06488(.A0(new_n8924_), .A1(new_n8921_), .B0(new_n3112_), .Y(new_n8925_));
  AOI21X1  g06489(.A0(new_n8925_), .A1(new_n8913_), .B0(pi0074), .Y(new_n8926_));
  OAI21X1  g06490(.A0(new_n8926_), .A1(new_n8912_), .B0(new_n3148_), .Y(new_n8927_));
  AOI21X1  g06491(.A0(new_n8911_), .A1(new_n8724_), .B0(new_n8927_), .Y(new_n8928_));
  NOR2X1   g06492(.A(new_n8708_), .B(new_n3095_), .Y(new_n8929_));
  AOI21X1  g06493(.A0(new_n8922_), .A1(new_n3095_), .B0(new_n8929_), .Y(new_n8930_));
  OAI21X1  g06494(.A0(new_n8930_), .A1(pi0054), .B0(new_n8913_), .Y(new_n8931_));
  AOI21X1  g06495(.A0(new_n8931_), .A1(new_n4991_), .B0(new_n8713_), .Y(new_n8932_));
  OAI21X1  g06496(.A0(new_n8932_), .A1(new_n3148_), .B0(new_n3246_), .Y(new_n8933_));
  OR2X1    g06497(.A(new_n8933_), .B(new_n7231_), .Y(new_n8934_));
  OAI21X1  g06498(.A0(new_n8934_), .A1(new_n8928_), .B0(new_n8714_), .Y(new_n8935_));
  NOR2X1   g06499(.A(new_n8935_), .B(pi0079), .Y(new_n8936_));
  INVX1    g06500(.A(new_n2545_), .Y(new_n8937_));
  NOR4X1   g06501(.A(new_n8937_), .B(pi0479), .C(new_n2540_), .D(pi0032), .Y(new_n8938_));
  OR4X1    g06502(.A(new_n8938_), .B(new_n7264_), .C(new_n5196_), .D(pi0040), .Y(new_n8939_));
  AND2X1   g06503(.A(new_n8939_), .B(new_n7783_), .Y(new_n8940_));
  NOR4X1   g06504(.A(new_n8938_), .B(new_n7288_), .C(new_n5196_), .D(pi0040), .Y(new_n8941_));
  OAI21X1  g06505(.A0(new_n8941_), .A1(new_n8776_), .B0(new_n8734_), .Y(new_n8942_));
  OAI21X1  g06506(.A0(new_n7264_), .A1(new_n7263_), .B0(new_n2766_), .Y(new_n8943_));
  NOR3X1   g06507(.A(new_n8938_), .B(new_n7261_), .C(pi0040), .Y(new_n8944_));
  AOI21X1  g06508(.A0(new_n8944_), .A1(new_n8943_), .B0(new_n7784_), .Y(new_n8945_));
  INVX1    g06509(.A(new_n7303_), .Y(new_n8946_));
  NOR4X1   g06510(.A(new_n8938_), .B(new_n8946_), .C(new_n7279_), .D(pi0040), .Y(new_n8947_));
  OAI21X1  g06511(.A0(new_n8947_), .A1(new_n8776_), .B0(pi0153), .Y(new_n8948_));
  OAI22X1  g06512(.A0(new_n8948_), .A1(new_n8945_), .B0(new_n8942_), .B1(new_n8940_), .Y(new_n8949_));
  OAI21X1  g06513(.A0(pi0468), .A1(pi0332), .B0(pi0040), .Y(new_n8950_));
  AND2X1   g06514(.A(new_n8950_), .B(pi0163), .Y(new_n8951_));
  AOI21X1  g06515(.A0(new_n8951_), .A1(new_n8949_), .B0(new_n8747_), .Y(new_n8952_));
  OAI21X1  g06516(.A0(new_n7262_), .A1(new_n8734_), .B0(new_n7535_), .Y(new_n8953_));
  AOI21X1  g06517(.A0(new_n7279_), .A1(pi0153), .B0(new_n8946_), .Y(new_n8954_));
  AND2X1   g06518(.A(pi0163), .B(new_n2549_), .Y(new_n8955_));
  OAI21X1  g06519(.A0(new_n8954_), .A1(new_n8776_), .B0(new_n8955_), .Y(new_n8956_));
  AOI21X1  g06520(.A0(new_n8953_), .A1(new_n7783_), .B0(new_n8956_), .Y(new_n8957_));
  NOR3X1   g06521(.A(new_n5057_), .B(new_n7272_), .C(new_n8734_), .Y(new_n8958_));
  OR4X1    g06522(.A(new_n7784_), .B(new_n7291_), .C(pi0095), .D(pi0032), .Y(new_n8959_));
  NAND3X1  g06523(.A(new_n8959_), .B(new_n8705_), .C(new_n2549_), .Y(new_n8960_));
  AOI21X1  g06524(.A0(new_n8958_), .A1(new_n7282_), .B0(new_n8960_), .Y(new_n8961_));
  NOR3X1   g06525(.A(new_n8961_), .B(new_n8957_), .C(pi0160), .Y(new_n8962_));
  NAND2X1  g06526(.A(new_n8938_), .B(new_n5033_), .Y(new_n8963_));
  AOI21X1  g06527(.A0(new_n8963_), .A1(new_n8961_), .B0(new_n2953_), .Y(new_n8964_));
  OAI21X1  g06528(.A0(new_n8962_), .A1(new_n8952_), .B0(new_n8964_), .Y(new_n8965_));
  NOR2X1   g06529(.A(new_n7264_), .B(new_n5220_), .Y(new_n8966_));
  OAI21X1  g06530(.A0(new_n7291_), .A1(new_n7272_), .B0(new_n8717_), .Y(new_n8967_));
  NAND2X1  g06531(.A(new_n8967_), .B(new_n7942_), .Y(new_n8968_));
  AOI21X1  g06532(.A0(new_n8966_), .A1(pi0184), .B0(new_n8968_), .Y(new_n8969_));
  AND2X1   g06533(.A(new_n8938_), .B(pi0182), .Y(new_n8970_));
  NOR3X1   g06534(.A(new_n7549_), .B(new_n7942_), .C(new_n8717_), .Y(new_n8971_));
  NOR3X1   g06535(.A(new_n8971_), .B(new_n8970_), .C(new_n8969_), .Y(new_n8972_));
  OAI21X1  g06536(.A0(new_n8972_), .A1(new_n5057_), .B0(new_n2549_), .Y(new_n8973_));
  INVX1    g06537(.A(new_n8970_), .Y(new_n8974_));
  NOR2X1   g06538(.A(new_n7282_), .B(new_n7942_), .Y(new_n8975_));
  OAI21X1  g06539(.A0(new_n7270_), .A1(pi0189), .B0(new_n7271_), .Y(new_n8976_));
  OAI21X1  g06540(.A0(new_n8976_), .A1(new_n8975_), .B0(new_n8974_), .Y(new_n8977_));
  AOI21X1  g06541(.A0(new_n8977_), .A1(new_n5033_), .B0(pi0184), .Y(new_n8978_));
  AND2X1   g06542(.A(pi0184), .B(new_n5227_), .Y(new_n8979_));
  OAI21X1  g06543(.A0(new_n7280_), .A1(new_n7942_), .B0(new_n8979_), .Y(new_n8980_));
  AOI21X1  g06544(.A0(new_n7780_), .A1(new_n7266_), .B0(new_n8980_), .Y(new_n8981_));
  OAI21X1  g06545(.A0(new_n8981_), .A1(new_n8978_), .B0(new_n2549_), .Y(new_n8982_));
  OAI21X1  g06546(.A0(new_n7265_), .A1(pi0198), .B0(new_n8944_), .Y(new_n8983_));
  NAND2X1  g06547(.A(new_n8983_), .B(new_n7780_), .Y(new_n8984_));
  OR4X1    g06548(.A(new_n8938_), .B(new_n7279_), .C(new_n5220_), .D(pi0040), .Y(new_n8985_));
  NAND3X1  g06549(.A(new_n8950_), .B(pi0184), .C(pi0182), .Y(new_n8986_));
  AOI21X1  g06550(.A0(new_n8985_), .A1(new_n8805_), .B0(new_n8986_), .Y(new_n8987_));
  AOI21X1  g06551(.A0(new_n8987_), .A1(new_n8984_), .B0(new_n8829_), .Y(new_n8988_));
  AOI22X1  g06552(.A0(new_n8988_), .A1(new_n8982_), .B0(new_n8973_), .B1(new_n8799_), .Y(new_n8989_));
  AOI21X1  g06553(.A0(new_n8989_), .A1(new_n8965_), .B0(pi0039), .Y(new_n8990_));
  NAND3X1  g06554(.A(new_n5033_), .B(new_n7271_), .C(new_n2545_), .Y(new_n8991_));
  AOI22X1  g06555(.A0(new_n6882_), .A1(new_n4464_), .B0(new_n5059_), .B1(pi0156), .Y(new_n8992_));
  NOR4X1   g06556(.A(new_n8992_), .B(new_n8991_), .C(new_n6905_), .D(new_n5070_), .Y(new_n8993_));
  NOR3X1   g06557(.A(new_n8993_), .B(new_n2953_), .C(pi0040), .Y(new_n8994_));
  AOI22X1  g06558(.A0(new_n6882_), .A1(new_n7942_), .B0(new_n5059_), .B1(pi0179), .Y(new_n8995_));
  NOR4X1   g06559(.A(new_n8995_), .B(new_n8991_), .C(new_n6913_), .D(new_n5050_), .Y(new_n8996_));
  OR2X1    g06560(.A(pi0299), .B(pi0040), .Y(new_n8997_));
  OAI21X1  g06561(.A0(new_n8997_), .A1(new_n8996_), .B0(pi0039), .Y(new_n8998_));
  OAI21X1  g06562(.A0(new_n8998_), .A1(new_n8994_), .B0(pi0232), .Y(new_n8999_));
  AOI21X1  g06563(.A0(new_n5237_), .A1(new_n2549_), .B0(pi0038), .Y(new_n9000_));
  OAI21X1  g06564(.A0(new_n8999_), .A1(new_n8990_), .B0(new_n9000_), .Y(new_n9001_));
  AOI21X1  g06565(.A0(new_n9001_), .A1(new_n8733_), .B0(new_n3124_), .Y(new_n9002_));
  OAI21X1  g06566(.A0(pi0040), .A1(pi0038), .B0(pi0087), .Y(new_n9003_));
  OAI22X1  g06567(.A0(new_n9003_), .A1(new_n8893_), .B0(new_n8722_), .B1(new_n3026_), .Y(new_n9004_));
  OAI21X1  g06568(.A0(new_n9004_), .A1(new_n9002_), .B0(new_n3105_), .Y(new_n9005_));
  NOR3X1   g06569(.A(new_n8905_), .B(new_n7188_), .C(new_n7272_), .Y(new_n9006_));
  AOI21X1  g06570(.A0(new_n9006_), .A1(new_n2545_), .B0(new_n8895_), .Y(new_n9007_));
  OAI21X1  g06571(.A0(new_n9007_), .A1(new_n8893_), .B0(new_n8901_), .Y(new_n9008_));
  AOI21X1  g06572(.A0(new_n9008_), .A1(new_n7185_), .B0(new_n8900_), .Y(new_n9009_));
  AOI21X1  g06573(.A0(new_n9009_), .A1(new_n9005_), .B0(pi0054), .Y(new_n9010_));
  OAI21X1  g06574(.A0(new_n9010_), .A1(new_n8728_), .B0(new_n4991_), .Y(new_n9011_));
  NOR4X1   g06575(.A(new_n7188_), .B(new_n5237_), .C(new_n8705_), .D(pi0092), .Y(new_n9012_));
  NAND4X1  g06576(.A(new_n9012_), .B(new_n5033_), .C(new_n7271_), .D(new_n2545_), .Y(new_n9013_));
  OR2X1    g06577(.A(new_n8918_), .B(pi0075), .Y(new_n9014_));
  AOI21X1  g06578(.A0(new_n9013_), .A1(new_n8894_), .B0(new_n9014_), .Y(new_n9015_));
  OAI21X1  g06579(.A0(new_n9015_), .A1(new_n8709_), .B0(new_n3112_), .Y(new_n9016_));
  AOI21X1  g06580(.A0(new_n9016_), .A1(new_n8913_), .B0(pi0074), .Y(new_n9017_));
  OAI21X1  g06581(.A0(new_n9017_), .A1(new_n8912_), .B0(new_n3148_), .Y(new_n9018_));
  AOI21X1  g06582(.A0(new_n9011_), .A1(new_n8724_), .B0(new_n9018_), .Y(new_n9019_));
  OAI21X1  g06583(.A0(new_n9019_), .A1(new_n8933_), .B0(new_n8714_), .Y(new_n9020_));
  OAI22X1  g06584(.A0(new_n9020_), .A1(new_n6816_), .B0(new_n7600_), .B1(pi0034), .Y(new_n9021_));
  AOI21X1  g06585(.A0(new_n6818_), .A1(new_n6817_), .B0(pi0079), .Y(new_n9022_));
  NOR2X1   g06586(.A(new_n9022_), .B(new_n8935_), .Y(new_n9023_));
  NOR3X1   g06587(.A(pi0954), .B(pi0034), .C(pi0033), .Y(new_n9024_));
  INVX1    g06588(.A(new_n9022_), .Y(new_n9025_));
  OAI21X1  g06589(.A0(new_n9025_), .A1(new_n9020_), .B0(new_n9024_), .Y(new_n9026_));
  OAI22X1  g06590(.A0(new_n9026_), .A1(new_n9023_), .B0(new_n9021_), .B1(new_n8936_), .Y(po0237));
  INVX1    g06591(.A(pi0588), .Y(new_n9028_));
  AND2X1   g06592(.A(pi1092), .B(pi0098), .Y(new_n9029_));
  AOI22X1  g06593(.A0(new_n9029_), .A1(pi1093), .B0(new_n2739_), .B1(new_n5928_), .Y(new_n9030_));
  AOI21X1  g06594(.A0(new_n9030_), .A1(new_n6630_), .B0(new_n9028_), .Y(new_n9031_));
  INVX1    g06595(.A(new_n9030_), .Y(new_n9032_));
  AND2X1   g06596(.A(new_n2739_), .B(new_n5928_), .Y(new_n9033_));
  NOR2X1   g06597(.A(new_n9033_), .B(new_n6309_), .Y(new_n9034_));
  INVX1    g06598(.A(new_n9034_), .Y(new_n9035_));
  NOR4X1   g06599(.A(new_n2756_), .B(new_n2755_), .C(new_n5903_), .D(new_n3095_), .Y(new_n9036_));
  INVX1    g06600(.A(new_n9036_), .Y(new_n9037_));
  NOR4X1   g06601(.A(new_n2756_), .B(new_n2755_), .C(new_n2722_), .D(new_n5903_), .Y(new_n9038_));
  NAND4X1  g06602(.A(new_n7834_), .B(new_n2475_), .C(new_n2681_), .D(new_n2474_), .Y(new_n9039_));
  OR4X1    g06603(.A(new_n9039_), .B(new_n5007_), .C(pi0110), .D(pi0047), .Y(new_n9040_));
  OR4X1    g06604(.A(new_n9040_), .B(new_n8252_), .C(new_n2579_), .D(pi0094), .Y(new_n9041_));
  NOR4X1   g06605(.A(new_n9041_), .B(new_n5908_), .C(pi0070), .D(new_n2516_), .Y(new_n9042_));
  NAND2X1  g06606(.A(pi0093), .B(pi0090), .Y(new_n9043_));
  NAND4X1  g06607(.A(new_n9043_), .B(new_n2532_), .C(new_n2492_), .D(new_n2726_), .Y(new_n9044_));
  NOR2X1   g06608(.A(new_n9044_), .B(new_n9041_), .Y(new_n9045_));
  AND2X1   g06609(.A(pi0950), .B(pi0824), .Y(new_n9046_));
  INVX1    g06610(.A(new_n9046_), .Y(new_n9047_));
  NOR2X1   g06611(.A(new_n9047_), .B(new_n5911_), .Y(new_n9048_));
  OAI21X1  g06612(.A0(new_n9045_), .A1(new_n9042_), .B0(new_n9048_), .Y(new_n9049_));
  AOI21X1  g06613(.A0(new_n9049_), .A1(new_n5903_), .B0(new_n2755_), .Y(new_n9050_));
  OR2X1    g06614(.A(new_n9050_), .B(new_n9038_), .Y(new_n9051_));
  OAI21X1  g06615(.A0(new_n9029_), .A1(new_n2722_), .B0(pi1093), .Y(new_n9052_));
  NOR2X1   g06616(.A(new_n9052_), .B(new_n3092_), .Y(new_n9053_));
  AND2X1   g06617(.A(new_n9053_), .B(new_n9051_), .Y(new_n9054_));
  AND2X1   g06618(.A(new_n9029_), .B(pi1093), .Y(new_n9055_));
  INVX1    g06619(.A(new_n9055_), .Y(new_n9056_));
  NAND4X1  g06620(.A(new_n9046_), .B(new_n3002_), .C(new_n2526_), .D(new_n2516_), .Y(new_n9057_));
  NOR4X1   g06621(.A(new_n9057_), .B(new_n9041_), .C(new_n5908_), .D(pi0070), .Y(new_n9058_));
  OAI21X1  g06622(.A0(new_n9058_), .A1(pi0098), .B0(pi1092), .Y(new_n9059_));
  INVX1    g06623(.A(new_n9059_), .Y(new_n9060_));
  NOR2X1   g06624(.A(new_n9052_), .B(new_n5999_), .Y(new_n9061_));
  OAI21X1  g06625(.A0(new_n9060_), .A1(new_n9038_), .B0(new_n9061_), .Y(new_n9062_));
  OAI21X1  g06626(.A0(new_n9056_), .A1(new_n3085_), .B0(new_n9062_), .Y(new_n9063_));
  OAI21X1  g06627(.A0(new_n9063_), .A1(new_n9054_), .B0(new_n3095_), .Y(new_n9064_));
  AOI21X1  g06628(.A0(new_n9064_), .A1(new_n9037_), .B0(new_n5928_), .Y(new_n9065_));
  OAI22X1  g06629(.A0(new_n9065_), .A1(new_n9035_), .B0(new_n9032_), .B1(new_n5893_), .Y(new_n9066_));
  MX2X1    g06630(.A(new_n9066_), .B(new_n9030_), .S0(pi0592), .Y(new_n9067_));
  NAND2X1  g06631(.A(new_n9067_), .B(new_n6550_), .Y(new_n9068_));
  NOR2X1   g06632(.A(new_n9030_), .B(pi1196), .Y(new_n9069_));
  NOR2X1   g06633(.A(new_n9069_), .B(new_n6550_), .Y(new_n9070_));
  INVX1    g06634(.A(new_n9070_), .Y(new_n9071_));
  INVX1    g06635(.A(pi0429), .Y(new_n9072_));
  INVX1    g06636(.A(pi0443), .Y(new_n9073_));
  MX2X1    g06637(.A(new_n9067_), .B(new_n9030_), .S0(new_n9073_), .Y(new_n9074_));
  INVX1    g06638(.A(new_n9074_), .Y(new_n9075_));
  MX2X1    g06639(.A(new_n9067_), .B(new_n9030_), .S0(pi0443), .Y(new_n9076_));
  INVX1    g06640(.A(new_n9076_), .Y(new_n9077_));
  MX2X1    g06641(.A(new_n9077_), .B(new_n9075_), .S0(new_n6598_), .Y(new_n9078_));
  AOI21X1  g06642(.A0(new_n9074_), .A1(pi0444), .B0(pi0436), .Y(new_n9079_));
  OAI21X1  g06643(.A0(new_n9077_), .A1(pi0444), .B0(new_n9079_), .Y(new_n9080_));
  AOI21X1  g06644(.A0(new_n9076_), .A1(pi0444), .B0(new_n6559_), .Y(new_n9081_));
  OAI21X1  g06645(.A0(new_n9075_), .A1(pi0444), .B0(new_n9081_), .Y(new_n9082_));
  AND2X1   g06646(.A(new_n9082_), .B(new_n9080_), .Y(new_n9083_));
  INVX1    g06647(.A(new_n9083_), .Y(new_n9084_));
  MX2X1    g06648(.A(new_n9084_), .B(new_n9078_), .S0(pi0435), .Y(new_n9085_));
  NAND2X1  g06649(.A(new_n9085_), .B(new_n9072_), .Y(new_n9086_));
  INVX1    g06650(.A(pi0435), .Y(new_n9087_));
  MX2X1    g06651(.A(new_n9084_), .B(new_n9078_), .S0(new_n9087_), .Y(new_n9088_));
  AOI21X1  g06652(.A0(new_n9088_), .A1(pi0429), .B0(new_n6564_), .Y(new_n9089_));
  AND2X1   g06653(.A(new_n9089_), .B(new_n9086_), .Y(new_n9090_));
  AND2X1   g06654(.A(new_n9088_), .B(new_n9072_), .Y(new_n9091_));
  AND2X1   g06655(.A(new_n9085_), .B(pi0429), .Y(new_n9092_));
  NOR3X1   g06656(.A(new_n9092_), .B(new_n9091_), .C(new_n6565_), .Y(new_n9093_));
  NOR3X1   g06657(.A(new_n9093_), .B(new_n9090_), .C(new_n6132_), .Y(new_n9094_));
  OAI21X1  g06658(.A0(new_n9094_), .A1(new_n9071_), .B0(new_n9068_), .Y(new_n9095_));
  MX2X1    g06659(.A(new_n9095_), .B(new_n9067_), .S0(pi0428), .Y(new_n9096_));
  MX2X1    g06660(.A(new_n9095_), .B(new_n9067_), .S0(new_n6528_), .Y(new_n9097_));
  MX2X1    g06661(.A(new_n9097_), .B(new_n9096_), .S0(new_n6527_), .Y(new_n9098_));
  MX2X1    g06662(.A(new_n9097_), .B(new_n9096_), .S0(pi0427), .Y(new_n9099_));
  MX2X1    g06663(.A(new_n9099_), .B(new_n9098_), .S0(pi0430), .Y(new_n9100_));
  MX2X1    g06664(.A(new_n9099_), .B(new_n9098_), .S0(new_n6582_), .Y(new_n9101_));
  MX2X1    g06665(.A(new_n9101_), .B(new_n9100_), .S0(pi0426), .Y(new_n9102_));
  MX2X1    g06666(.A(new_n9101_), .B(new_n9100_), .S0(new_n6585_), .Y(new_n9103_));
  MX2X1    g06667(.A(new_n9103_), .B(new_n9102_), .S0(pi0445), .Y(new_n9104_));
  NOR2X1   g06668(.A(new_n9104_), .B(new_n6522_), .Y(new_n9105_));
  MX2X1    g06669(.A(new_n9103_), .B(new_n9102_), .S0(new_n6589_), .Y(new_n9106_));
  OAI21X1  g06670(.A0(new_n9106_), .A1(pi0448), .B0(new_n6525_), .Y(new_n9107_));
  NOR2X1   g06671(.A(new_n9107_), .B(new_n9105_), .Y(new_n9108_));
  NOR2X1   g06672(.A(new_n9106_), .B(new_n6522_), .Y(new_n9109_));
  OAI21X1  g06673(.A0(new_n9104_), .A1(pi0448), .B0(new_n6623_), .Y(new_n9110_));
  OAI21X1  g06674(.A0(new_n9110_), .A1(new_n9109_), .B0(pi1199), .Y(new_n9111_));
  OR2X1    g06675(.A(new_n9095_), .B(pi1199), .Y(new_n9112_));
  AND2X1   g06676(.A(new_n9112_), .B(new_n6593_), .Y(new_n9113_));
  OAI21X1  g06677(.A0(new_n9111_), .A1(new_n9108_), .B0(new_n9113_), .Y(new_n9114_));
  OAI21X1  g06678(.A0(new_n9030_), .A1(new_n6074_), .B0(pi0590), .Y(new_n9115_));
  INVX1    g06679(.A(pi0354), .Y(new_n9116_));
  INVX1    g06680(.A(new_n9067_), .Y(new_n9117_));
  MX2X1    g06681(.A(new_n9117_), .B(new_n9032_), .S0(new_n6653_), .Y(new_n9118_));
  NOR2X1   g06682(.A(new_n9069_), .B(pi1198), .Y(new_n9119_));
  INVX1    g06683(.A(new_n9119_), .Y(new_n9120_));
  MX2X1    g06684(.A(new_n9117_), .B(new_n9032_), .S0(new_n6025_), .Y(new_n9121_));
  MX2X1    g06685(.A(new_n9067_), .B(new_n9030_), .S0(pi0455), .Y(new_n9122_));
  MX2X1    g06686(.A(new_n9067_), .B(new_n9030_), .S0(new_n6041_), .Y(new_n9123_));
  MX2X1    g06687(.A(new_n9123_), .B(new_n9122_), .S0(new_n6024_), .Y(new_n9124_));
  INVX1    g06688(.A(new_n9124_), .Y(new_n9125_));
  MX2X1    g06689(.A(new_n9125_), .B(new_n9121_), .S0(pi0355), .Y(new_n9126_));
  INVX1    g06690(.A(new_n9126_), .Y(new_n9127_));
  MX2X1    g06691(.A(new_n9125_), .B(new_n9121_), .S0(new_n6039_), .Y(new_n9128_));
  AOI21X1  g06692(.A0(new_n9128_), .A1(pi0458), .B0(new_n6031_), .Y(new_n9129_));
  OAI21X1  g06693(.A0(new_n9127_), .A1(pi0458), .B0(new_n9129_), .Y(new_n9130_));
  NAND2X1  g06694(.A(new_n9128_), .B(new_n6038_), .Y(new_n9131_));
  AOI21X1  g06695(.A0(new_n9126_), .A1(pi0458), .B0(new_n6051_), .Y(new_n9132_));
  AOI21X1  g06696(.A0(new_n9132_), .A1(new_n9131_), .B0(new_n6132_), .Y(new_n9133_));
  AND2X1   g06697(.A(new_n9133_), .B(new_n9130_), .Y(new_n9134_));
  OAI22X1  g06698(.A0(new_n9134_), .A1(new_n9120_), .B0(new_n9118_), .B1(new_n6055_), .Y(new_n9135_));
  MX2X1    g06699(.A(new_n9135_), .B(new_n9067_), .S0(new_n5892_), .Y(new_n9136_));
  OR2X1    g06700(.A(new_n9067_), .B(new_n6061_), .Y(new_n9137_));
  OAI22X1  g06701(.A0(new_n9137_), .A1(new_n6059_), .B0(new_n9136_), .B1(new_n6064_), .Y(new_n9138_));
  OAI22X1  g06702(.A0(new_n9137_), .A1(pi0351), .B0(new_n9136_), .B1(new_n6060_), .Y(new_n9139_));
  MX2X1    g06703(.A(new_n9139_), .B(new_n9138_), .S0(new_n5879_), .Y(new_n9140_));
  MX2X1    g06704(.A(new_n9139_), .B(new_n9138_), .S0(pi0461), .Y(new_n9141_));
  MX2X1    g06705(.A(new_n9141_), .B(new_n9140_), .S0(new_n5878_), .Y(new_n9142_));
  MX2X1    g06706(.A(new_n9141_), .B(new_n9140_), .S0(pi0357), .Y(new_n9143_));
  MX2X1    g06707(.A(new_n9143_), .B(new_n9142_), .S0(new_n5877_), .Y(new_n9144_));
  AND2X1   g06708(.A(new_n9144_), .B(new_n9116_), .Y(new_n9145_));
  AND2X1   g06709(.A(new_n9143_), .B(new_n5877_), .Y(new_n9146_));
  AOI21X1  g06710(.A0(new_n9142_), .A1(pi0356), .B0(new_n9146_), .Y(new_n9147_));
  OAI21X1  g06711(.A0(new_n9147_), .A1(new_n9116_), .B0(new_n5874_), .Y(new_n9148_));
  OR2X1    g06712(.A(new_n9148_), .B(new_n9145_), .Y(new_n9149_));
  AOI21X1  g06713(.A0(new_n9144_), .A1(pi0354), .B0(new_n5874_), .Y(new_n9150_));
  OAI21X1  g06714(.A0(new_n9147_), .A1(pi0354), .B0(new_n9150_), .Y(new_n9151_));
  AND2X1   g06715(.A(new_n9151_), .B(new_n6074_), .Y(new_n9152_));
  AOI21X1  g06716(.A0(new_n9152_), .A1(new_n9149_), .B0(new_n9115_), .Y(new_n9153_));
  OR2X1    g06717(.A(new_n6183_), .B(pi1197), .Y(new_n9154_));
  AOI21X1  g06718(.A0(new_n9030_), .A1(new_n6309_), .B0(new_n6378_), .Y(new_n9155_));
  INVX1    g06719(.A(pi0411), .Y(new_n9156_));
  INVX1    g06720(.A(new_n6191_), .Y(new_n9157_));
  AOI21X1  g06721(.A0(new_n9029_), .A1(new_n9156_), .B0(new_n9157_), .Y(new_n9158_));
  INVX1    g06722(.A(new_n9158_), .Y(new_n9159_));
  AOI21X1  g06723(.A0(new_n9050_), .A1(pi0411), .B0(new_n9159_), .Y(new_n9160_));
  INVX1    g06724(.A(new_n9029_), .Y(new_n9161_));
  OAI21X1  g06725(.A0(new_n9161_), .A1(new_n9156_), .B0(new_n9157_), .Y(new_n9162_));
  AOI21X1  g06726(.A0(new_n9050_), .A1(new_n9156_), .B0(new_n9162_), .Y(new_n9163_));
  NOR2X1   g06727(.A(new_n9163_), .B(new_n9160_), .Y(new_n9164_));
  OAI21X1  g06728(.A0(new_n9164_), .A1(new_n9038_), .B0(new_n9053_), .Y(new_n9165_));
  AOI21X1  g06729(.A0(new_n9060_), .A1(pi0411), .B0(new_n9159_), .Y(new_n9166_));
  AOI21X1  g06730(.A0(new_n9060_), .A1(new_n9156_), .B0(new_n9162_), .Y(new_n9167_));
  OAI22X1  g06731(.A0(new_n9167_), .A1(new_n9166_), .B0(new_n9056_), .B1(new_n2722_), .Y(new_n9168_));
  AOI22X1  g06732(.A0(new_n9168_), .A1(new_n9061_), .B0(new_n9055_), .B1(new_n3157_), .Y(new_n9169_));
  NAND2X1  g06733(.A(new_n9169_), .B(new_n9165_), .Y(new_n9170_));
  AOI21X1  g06734(.A0(new_n9170_), .A1(new_n3095_), .B0(new_n9036_), .Y(new_n9171_));
  OAI21X1  g06735(.A0(new_n9171_), .A1(new_n5928_), .B0(new_n9034_), .Y(new_n9172_));
  OAI22X1  g06736(.A0(new_n9033_), .A1(new_n9055_), .B0(new_n6132_), .B1(pi0592), .Y(new_n9173_));
  NAND2X1  g06737(.A(new_n9173_), .B(new_n6061_), .Y(new_n9174_));
  AOI21X1  g06738(.A0(new_n9172_), .A1(new_n9155_), .B0(new_n9174_), .Y(new_n9175_));
  NOR2X1   g06739(.A(new_n9062_), .B(new_n6210_), .Y(new_n9176_));
  MX2X1    g06740(.A(new_n9050_), .B(new_n9029_), .S0(new_n6210_), .Y(new_n9177_));
  AND2X1   g06741(.A(new_n9177_), .B(new_n9054_), .Y(new_n9178_));
  OR2X1    g06742(.A(new_n9178_), .B(new_n9176_), .Y(new_n9179_));
  OAI21X1  g06743(.A0(new_n9179_), .A1(new_n9170_), .B0(new_n9155_), .Y(new_n9180_));
  MX2X1    g06744(.A(new_n9059_), .B(new_n9161_), .S0(new_n6210_), .Y(new_n9181_));
  OAI22X1  g06745(.A0(new_n9181_), .A1(new_n9062_), .B0(new_n9056_), .B1(new_n3085_), .Y(new_n9182_));
  AOI21X1  g06746(.A0(new_n9030_), .A1(new_n6309_), .B0(new_n6454_), .Y(new_n9183_));
  OAI21X1  g06747(.A0(new_n9182_), .A1(new_n9178_), .B0(new_n9183_), .Y(new_n9184_));
  NAND2X1  g06748(.A(new_n9184_), .B(new_n9180_), .Y(new_n9185_));
  AND2X1   g06749(.A(pi0567), .B(new_n3095_), .Y(new_n9186_));
  NOR3X1   g06750(.A(new_n9033_), .B(new_n6216_), .C(new_n6309_), .Y(new_n9187_));
  OAI21X1  g06751(.A0(new_n9187_), .A1(new_n9030_), .B0(pi1199), .Y(new_n9188_));
  AOI21X1  g06752(.A0(new_n9186_), .A1(new_n9185_), .B0(new_n9188_), .Y(new_n9189_));
  NOR3X1   g06753(.A(new_n9189_), .B(new_n9175_), .C(new_n6183_), .Y(new_n9190_));
  AOI22X1  g06754(.A0(new_n9190_), .A1(new_n5889_), .B0(new_n9154_), .B1(new_n9117_), .Y(new_n9191_));
  NOR3X1   g06755(.A(new_n9067_), .B(new_n6700_), .C(new_n6055_), .Y(new_n9192_));
  OAI21X1  g06756(.A0(new_n9192_), .A1(new_n9190_), .B0(pi0333), .Y(new_n9193_));
  OAI21X1  g06757(.A0(new_n9191_), .A1(pi0333), .B0(new_n9193_), .Y(new_n9194_));
  AND2X1   g06758(.A(new_n9194_), .B(new_n6231_), .Y(new_n9195_));
  OAI21X1  g06759(.A0(new_n9192_), .A1(new_n9190_), .B0(new_n6172_), .Y(new_n9196_));
  OAI21X1  g06760(.A0(new_n9191_), .A1(new_n6172_), .B0(new_n9196_), .Y(new_n9197_));
  AOI21X1  g06761(.A0(new_n9197_), .A1(pi0391), .B0(new_n9195_), .Y(new_n9198_));
  OR2X1    g06762(.A(new_n9198_), .B(pi0392), .Y(new_n9199_));
  AND2X1   g06763(.A(new_n9197_), .B(new_n6231_), .Y(new_n9200_));
  AOI21X1  g06764(.A0(new_n9194_), .A1(pi0391), .B0(new_n9200_), .Y(new_n9201_));
  OAI21X1  g06765(.A0(new_n9201_), .A1(new_n6171_), .B0(new_n9199_), .Y(new_n9202_));
  MX2X1    g06766(.A(new_n9201_), .B(new_n9198_), .S0(pi0392), .Y(new_n9203_));
  OAI21X1  g06767(.A0(new_n9203_), .A1(new_n6170_), .B0(new_n6713_), .Y(new_n9204_));
  AOI21X1  g06768(.A0(new_n9202_), .A1(new_n6170_), .B0(new_n9204_), .Y(new_n9205_));
  OR2X1    g06769(.A(new_n9203_), .B(pi0393), .Y(new_n9206_));
  AOI21X1  g06770(.A0(new_n9202_), .A1(pi0393), .B0(new_n6713_), .Y(new_n9207_));
  AND2X1   g06771(.A(new_n9207_), .B(new_n9206_), .Y(new_n9208_));
  NOR3X1   g06772(.A(new_n9208_), .B(new_n9205_), .C(new_n6074_), .Y(new_n9209_));
  MX2X1    g06773(.A(new_n9066_), .B(new_n9030_), .S0(new_n6120_), .Y(new_n9210_));
  INVX1    g06774(.A(new_n9210_), .Y(new_n9211_));
  AOI21X1  g06775(.A0(new_n9030_), .A1(new_n6676_), .B0(new_n6061_), .Y(new_n9212_));
  OAI21X1  g06776(.A0(new_n9211_), .A1(new_n6676_), .B0(new_n9212_), .Y(new_n9213_));
  AOI22X1  g06777(.A0(new_n9032_), .A1(new_n5889_), .B0(new_n6090_), .B1(pi1196), .Y(new_n9214_));
  INVX1    g06778(.A(new_n9214_), .Y(new_n9215_));
  XOR2X1   g06779(.A(new_n6101_), .B(new_n6093_), .Y(new_n9216_));
  XOR2X1   g06780(.A(new_n9216_), .B(new_n6095_), .Y(new_n9217_));
  OAI21X1  g06781(.A0(new_n9217_), .A1(new_n9032_), .B0(pi1197), .Y(new_n9218_));
  AOI21X1  g06782(.A0(new_n9217_), .A1(new_n9210_), .B0(new_n9218_), .Y(new_n9219_));
  AOI21X1  g06783(.A0(new_n9210_), .A1(new_n6091_), .B0(pi1199), .Y(new_n9220_));
  OAI21X1  g06784(.A0(new_n9219_), .A1(new_n9215_), .B0(new_n9220_), .Y(new_n9221_));
  AND2X1   g06785(.A(new_n9221_), .B(new_n9213_), .Y(new_n9222_));
  OR2X1    g06786(.A(new_n9222_), .B(pi0374), .Y(new_n9223_));
  MX2X1    g06787(.A(new_n9222_), .B(new_n9210_), .S0(pi1198), .Y(new_n9224_));
  OAI21X1  g06788(.A0(new_n9224_), .A1(new_n6143_), .B0(new_n9223_), .Y(new_n9225_));
  XOR2X1   g06789(.A(new_n6351_), .B(pi0371), .Y(new_n9226_));
  XOR2X1   g06790(.A(new_n9226_), .B(new_n6081_), .Y(new_n9227_));
  INVX1    g06791(.A(new_n9227_), .Y(new_n9228_));
  MX2X1    g06792(.A(new_n9224_), .B(new_n9222_), .S0(pi0374), .Y(new_n9229_));
  OAI21X1  g06793(.A0(new_n9229_), .A1(new_n6082_), .B0(new_n9228_), .Y(new_n9230_));
  AOI21X1  g06794(.A0(new_n9225_), .A1(new_n6082_), .B0(new_n9230_), .Y(new_n9231_));
  AND2X1   g06795(.A(new_n9225_), .B(pi0369), .Y(new_n9232_));
  OAI21X1  g06796(.A0(new_n9229_), .A1(pi0369), .B0(new_n9227_), .Y(new_n9233_));
  OAI21X1  g06797(.A0(new_n9233_), .A1(new_n9232_), .B0(new_n6074_), .Y(new_n9234_));
  OAI21X1  g06798(.A0(new_n9234_), .A1(new_n9231_), .B0(new_n6168_), .Y(new_n9235_));
  OAI21X1  g06799(.A0(new_n9235_), .A1(new_n9209_), .B0(new_n9028_), .Y(new_n9236_));
  OAI21X1  g06800(.A0(new_n9236_), .A1(new_n9153_), .B0(new_n6077_), .Y(new_n9237_));
  AOI21X1  g06801(.A0(new_n9114_), .A1(new_n9031_), .B0(new_n9237_), .Y(new_n9238_));
  AND2X1   g06802(.A(new_n6256_), .B(new_n5938_), .Y(new_n9239_));
  AOI21X1  g06803(.A0(new_n9239_), .A1(new_n2722_), .B0(new_n9055_), .Y(new_n9240_));
  AOI21X1  g06804(.A0(new_n9240_), .A1(new_n5952_), .B0(new_n5983_), .Y(new_n9241_));
  OR2X1    g06805(.A(new_n9038_), .B(new_n3157_), .Y(new_n9242_));
  NOR3X1   g06806(.A(new_n9242_), .B(new_n9050_), .C(pi0087), .Y(new_n9243_));
  NOR3X1   g06807(.A(new_n9038_), .B(new_n3157_), .C(new_n3156_), .Y(new_n9244_));
  AOI21X1  g06808(.A0(new_n9244_), .A1(new_n9059_), .B0(new_n9243_), .Y(new_n9245_));
  OAI22X1  g06809(.A0(new_n9245_), .A1(new_n5952_), .B0(new_n9242_), .B1(new_n9241_), .Y(new_n9246_));
  AND2X1   g06810(.A(new_n5893_), .B(pi0567), .Y(new_n9247_));
  INVX1    g06811(.A(new_n9247_), .Y(new_n9248_));
  AND2X1   g06812(.A(new_n9239_), .B(new_n2722_), .Y(new_n9249_));
  NOR3X1   g06813(.A(new_n9055_), .B(new_n9249_), .C(new_n5924_), .Y(new_n9250_));
  OR2X1    g06814(.A(new_n9250_), .B(new_n9248_), .Y(new_n9251_));
  AOI21X1  g06815(.A0(new_n9246_), .A1(new_n3095_), .B0(new_n9251_), .Y(new_n9252_));
  OAI22X1  g06816(.A0(new_n9240_), .A1(new_n5893_), .B0(new_n2740_), .B1(pi0567), .Y(new_n9253_));
  NOR2X1   g06817(.A(new_n9253_), .B(new_n9252_), .Y(new_n9254_));
  MX2X1    g06818(.A(new_n9254_), .B(new_n9030_), .S0(pi0592), .Y(new_n9255_));
  INVX1    g06819(.A(new_n9255_), .Y(new_n9256_));
  MX2X1    g06820(.A(new_n9255_), .B(new_n9030_), .S0(new_n9073_), .Y(new_n9257_));
  INVX1    g06821(.A(new_n9257_), .Y(new_n9258_));
  MX2X1    g06822(.A(new_n9255_), .B(new_n9030_), .S0(pi0443), .Y(new_n9259_));
  INVX1    g06823(.A(new_n9259_), .Y(new_n9260_));
  MX2X1    g06824(.A(new_n9260_), .B(new_n9258_), .S0(new_n6598_), .Y(new_n9261_));
  NAND2X1  g06825(.A(new_n9259_), .B(new_n6552_), .Y(new_n9262_));
  AOI21X1  g06826(.A0(new_n9257_), .A1(pi0444), .B0(pi0436), .Y(new_n9263_));
  NAND2X1  g06827(.A(new_n9257_), .B(new_n6552_), .Y(new_n9264_));
  AOI21X1  g06828(.A0(new_n9259_), .A1(pi0444), .B0(new_n6559_), .Y(new_n9265_));
  AOI22X1  g06829(.A0(new_n9265_), .A1(new_n9264_), .B0(new_n9263_), .B1(new_n9262_), .Y(new_n9266_));
  INVX1    g06830(.A(new_n9266_), .Y(new_n9267_));
  MX2X1    g06831(.A(new_n9267_), .B(new_n9261_), .S0(pi0435), .Y(new_n9268_));
  INVX1    g06832(.A(new_n9268_), .Y(new_n9269_));
  MX2X1    g06833(.A(new_n9267_), .B(new_n9261_), .S0(new_n9087_), .Y(new_n9270_));
  AOI21X1  g06834(.A0(new_n9270_), .A1(pi0429), .B0(new_n6564_), .Y(new_n9271_));
  OAI21X1  g06835(.A0(new_n9269_), .A1(pi0429), .B0(new_n9271_), .Y(new_n9272_));
  AND2X1   g06836(.A(new_n9270_), .B(new_n9072_), .Y(new_n9273_));
  AND2X1   g06837(.A(new_n9268_), .B(pi0429), .Y(new_n9274_));
  NOR3X1   g06838(.A(new_n9274_), .B(new_n9273_), .C(new_n6565_), .Y(new_n9275_));
  NOR2X1   g06839(.A(new_n9275_), .B(new_n6132_), .Y(new_n9276_));
  AOI21X1  g06840(.A0(new_n9276_), .A1(new_n9272_), .B0(new_n9071_), .Y(new_n9277_));
  AOI21X1  g06841(.A0(new_n9255_), .A1(new_n6550_), .B0(new_n9277_), .Y(new_n9278_));
  MX2X1    g06842(.A(new_n9278_), .B(new_n9256_), .S0(new_n6528_), .Y(new_n9279_));
  MX2X1    g06843(.A(new_n9278_), .B(new_n9256_), .S0(pi0428), .Y(new_n9280_));
  MX2X1    g06844(.A(new_n9280_), .B(new_n9279_), .S0(new_n6527_), .Y(new_n9281_));
  MX2X1    g06845(.A(new_n9280_), .B(new_n9279_), .S0(pi0427), .Y(new_n9282_));
  MX2X1    g06846(.A(new_n9282_), .B(new_n9281_), .S0(pi0430), .Y(new_n9283_));
  MX2X1    g06847(.A(new_n9282_), .B(new_n9281_), .S0(new_n6582_), .Y(new_n9284_));
  MX2X1    g06848(.A(new_n9284_), .B(new_n9283_), .S0(pi0426), .Y(new_n9285_));
  MX2X1    g06849(.A(new_n9284_), .B(new_n9283_), .S0(new_n6585_), .Y(new_n9286_));
  MX2X1    g06850(.A(new_n9286_), .B(new_n9285_), .S0(pi0445), .Y(new_n9287_));
  OR2X1    g06851(.A(new_n9286_), .B(new_n6589_), .Y(new_n9288_));
  OAI21X1  g06852(.A0(new_n9285_), .A1(pi0445), .B0(new_n9288_), .Y(new_n9289_));
  OAI21X1  g06853(.A0(new_n9289_), .A1(pi0448), .B0(new_n6623_), .Y(new_n9290_));
  AOI21X1  g06854(.A0(new_n9287_), .A1(pi0448), .B0(new_n9290_), .Y(new_n9291_));
  AND2X1   g06855(.A(new_n9287_), .B(new_n6522_), .Y(new_n9292_));
  OAI21X1  g06856(.A0(new_n9289_), .A1(new_n6522_), .B0(new_n6525_), .Y(new_n9293_));
  OAI21X1  g06857(.A0(new_n9293_), .A1(new_n9292_), .B0(pi1199), .Y(new_n9294_));
  AOI21X1  g06858(.A0(new_n9278_), .A1(new_n6061_), .B0(new_n6630_), .Y(new_n9295_));
  OAI21X1  g06859(.A0(new_n9294_), .A1(new_n9291_), .B0(new_n9295_), .Y(new_n9296_));
  MX2X1    g06860(.A(new_n9256_), .B(new_n9032_), .S0(new_n6653_), .Y(new_n9297_));
  MX2X1    g06861(.A(new_n9256_), .B(new_n9032_), .S0(new_n6025_), .Y(new_n9298_));
  MX2X1    g06862(.A(new_n9255_), .B(new_n9030_), .S0(pi0455), .Y(new_n9299_));
  MX2X1    g06863(.A(new_n9255_), .B(new_n9030_), .S0(new_n6041_), .Y(new_n9300_));
  MX2X1    g06864(.A(new_n9300_), .B(new_n9299_), .S0(new_n6024_), .Y(new_n9301_));
  INVX1    g06865(.A(new_n9301_), .Y(new_n9302_));
  MX2X1    g06866(.A(new_n9302_), .B(new_n9298_), .S0(new_n6039_), .Y(new_n9303_));
  NAND2X1  g06867(.A(new_n9303_), .B(new_n6038_), .Y(new_n9304_));
  MX2X1    g06868(.A(new_n9302_), .B(new_n9298_), .S0(pi0355), .Y(new_n9305_));
  AOI21X1  g06869(.A0(new_n9305_), .A1(pi0458), .B0(new_n6051_), .Y(new_n9306_));
  NAND2X1  g06870(.A(new_n9306_), .B(new_n9304_), .Y(new_n9307_));
  NAND2X1  g06871(.A(new_n9305_), .B(new_n6038_), .Y(new_n9308_));
  AOI21X1  g06872(.A0(new_n9303_), .A1(pi0458), .B0(new_n6031_), .Y(new_n9309_));
  AOI21X1  g06873(.A0(new_n9309_), .A1(new_n9308_), .B0(new_n6132_), .Y(new_n9310_));
  AND2X1   g06874(.A(new_n9310_), .B(new_n9307_), .Y(new_n9311_));
  OAI22X1  g06875(.A0(new_n9311_), .A1(new_n9120_), .B0(new_n9297_), .B1(new_n6055_), .Y(new_n9312_));
  MX2X1    g06876(.A(new_n9312_), .B(new_n9255_), .S0(new_n5892_), .Y(new_n9313_));
  INVX1    g06877(.A(new_n9313_), .Y(new_n9314_));
  NOR2X1   g06878(.A(new_n9255_), .B(new_n6061_), .Y(new_n9315_));
  AOI22X1  g06879(.A0(new_n9315_), .A1(pi0351), .B0(new_n9314_), .B1(new_n6336_), .Y(new_n9316_));
  AOI22X1  g06880(.A0(new_n9315_), .A1(new_n6059_), .B0(new_n9314_), .B1(new_n6251_), .Y(new_n9317_));
  MX2X1    g06881(.A(new_n9317_), .B(new_n9316_), .S0(new_n5879_), .Y(new_n9318_));
  MX2X1    g06882(.A(new_n9317_), .B(new_n9316_), .S0(pi0461), .Y(new_n9319_));
  MX2X1    g06883(.A(new_n9319_), .B(new_n9318_), .S0(new_n5878_), .Y(new_n9320_));
  MX2X1    g06884(.A(new_n9319_), .B(new_n9318_), .S0(pi0357), .Y(new_n9321_));
  MX2X1    g06885(.A(new_n9321_), .B(new_n9320_), .S0(new_n5877_), .Y(new_n9322_));
  INVX1    g06886(.A(new_n5874_), .Y(new_n9323_));
  OR2X1    g06887(.A(new_n9321_), .B(pi0356), .Y(new_n9324_));
  OAI21X1  g06888(.A0(new_n9320_), .A1(new_n5877_), .B0(new_n9324_), .Y(new_n9325_));
  AOI21X1  g06889(.A0(new_n9325_), .A1(pi0354), .B0(new_n9323_), .Y(new_n9326_));
  OAI21X1  g06890(.A0(new_n9322_), .A1(pi0354), .B0(new_n9326_), .Y(new_n9327_));
  NAND2X1  g06891(.A(new_n9325_), .B(new_n9116_), .Y(new_n9328_));
  OR2X1    g06892(.A(new_n9322_), .B(new_n9116_), .Y(new_n9329_));
  AND2X1   g06893(.A(new_n9329_), .B(new_n9323_), .Y(new_n9330_));
  AOI21X1  g06894(.A0(new_n9330_), .A1(new_n9328_), .B0(pi0591), .Y(new_n9331_));
  AOI21X1  g06895(.A0(new_n9331_), .A1(new_n9327_), .B0(new_n9115_), .Y(new_n9332_));
  MX2X1    g06896(.A(new_n9254_), .B(new_n9030_), .S0(new_n6120_), .Y(new_n9333_));
  MX2X1    g06897(.A(new_n9333_), .B(new_n9030_), .S0(pi0367), .Y(new_n9334_));
  MX2X1    g06898(.A(new_n9333_), .B(new_n9030_), .S0(new_n6095_), .Y(new_n9335_));
  MX2X1    g06899(.A(new_n9335_), .B(new_n9334_), .S0(new_n6093_), .Y(new_n9336_));
  OR2X1    g06900(.A(new_n9336_), .B(new_n6096_), .Y(new_n9337_));
  MX2X1    g06901(.A(new_n9335_), .B(new_n9334_), .S0(new_n6094_), .Y(new_n9338_));
  INVX1    g06902(.A(new_n9338_), .Y(new_n9339_));
  AOI21X1  g06903(.A0(new_n9339_), .A1(new_n6096_), .B0(new_n6100_), .Y(new_n9340_));
  NOR2X1   g06904(.A(new_n9336_), .B(new_n6097_), .Y(new_n9341_));
  OAI21X1  g06905(.A0(new_n9338_), .A1(new_n6096_), .B0(new_n6100_), .Y(new_n9342_));
  OAI21X1  g06906(.A0(new_n9342_), .A1(new_n9341_), .B0(pi1197), .Y(new_n9343_));
  AOI21X1  g06907(.A0(new_n9340_), .A1(new_n9337_), .B0(new_n9343_), .Y(new_n9344_));
  AOI21X1  g06908(.A0(new_n9333_), .A1(new_n6091_), .B0(pi1199), .Y(new_n9345_));
  OAI21X1  g06909(.A0(new_n9344_), .A1(new_n9215_), .B0(new_n9345_), .Y(new_n9346_));
  INVX1    g06910(.A(new_n9333_), .Y(new_n9347_));
  MX2X1    g06911(.A(new_n9347_), .B(new_n9032_), .S0(new_n6676_), .Y(new_n9348_));
  NAND2X1  g06912(.A(new_n9348_), .B(pi1199), .Y(new_n9349_));
  AND2X1   g06913(.A(new_n9349_), .B(new_n9346_), .Y(new_n9350_));
  AOI22X1  g06914(.A0(new_n9348_), .A1(new_n6138_), .B0(new_n9347_), .B1(pi1198), .Y(new_n9351_));
  OAI21X1  g06915(.A0(new_n9346_), .A1(pi1198), .B0(new_n9351_), .Y(new_n9352_));
  NAND2X1  g06916(.A(new_n9352_), .B(pi0374), .Y(new_n9353_));
  OAI21X1  g06917(.A0(new_n9350_), .A1(pi0374), .B0(new_n9353_), .Y(new_n9354_));
  AOI21X1  g06918(.A0(new_n9349_), .A1(new_n9346_), .B0(new_n6143_), .Y(new_n9355_));
  AOI21X1  g06919(.A0(new_n9352_), .A1(new_n6143_), .B0(new_n9355_), .Y(new_n9356_));
  OAI21X1  g06920(.A0(new_n9356_), .A1(pi0369), .B0(new_n9227_), .Y(new_n9357_));
  AOI21X1  g06921(.A0(new_n9354_), .A1(pi0369), .B0(new_n9357_), .Y(new_n9358_));
  OAI21X1  g06922(.A0(new_n9356_), .A1(new_n6082_), .B0(new_n9228_), .Y(new_n9359_));
  AOI21X1  g06923(.A0(new_n9354_), .A1(new_n6082_), .B0(new_n9359_), .Y(new_n9360_));
  NOR3X1   g06924(.A(new_n9360_), .B(new_n9358_), .C(pi0591), .Y(new_n9361_));
  XOR2X1   g06925(.A(pi0404), .B(pi0397), .Y(new_n9362_));
  XOR2X1   g06926(.A(new_n9362_), .B(pi0411), .Y(new_n9363_));
  XOR2X1   g06927(.A(new_n9363_), .B(new_n6184_), .Y(new_n9364_));
  OR2X1    g06928(.A(new_n9364_), .B(new_n5939_), .Y(new_n9365_));
  AND2X1   g06929(.A(new_n9365_), .B(new_n9161_), .Y(new_n9366_));
  INVX1    g06930(.A(pi0412), .Y(new_n9367_));
  AOI21X1  g06931(.A0(new_n9364_), .A1(new_n5938_), .B0(new_n9029_), .Y(new_n9368_));
  OR2X1    g06932(.A(new_n9368_), .B(new_n9367_), .Y(new_n9369_));
  AND2X1   g06933(.A(new_n9369_), .B(new_n6189_), .Y(new_n9370_));
  OAI21X1  g06934(.A0(new_n9366_), .A1(pi0412), .B0(new_n9370_), .Y(new_n9371_));
  INVX1    g06935(.A(new_n9368_), .Y(new_n9372_));
  AOI21X1  g06936(.A0(new_n9372_), .A1(new_n9367_), .B0(new_n6189_), .Y(new_n9373_));
  OAI21X1  g06937(.A0(new_n9366_), .A1(new_n9367_), .B0(new_n9373_), .Y(new_n9374_));
  NAND3X1  g06938(.A(new_n9374_), .B(new_n9371_), .C(new_n5952_), .Y(new_n9375_));
  AOI21X1  g06939(.A0(new_n9375_), .A1(new_n9161_), .B0(new_n5983_), .Y(new_n9376_));
  NOR2X1   g06940(.A(new_n9376_), .B(new_n9038_), .Y(new_n9377_));
  MX2X1    g06941(.A(new_n9377_), .B(new_n2740_), .S0(new_n5928_), .Y(new_n9378_));
  NOR2X1   g06942(.A(new_n9378_), .B(new_n9034_), .Y(new_n9379_));
  INVX1    g06943(.A(new_n9379_), .Y(new_n9380_));
  NOR3X1   g06944(.A(new_n9038_), .B(new_n3157_), .C(pi0087), .Y(new_n9381_));
  INVX1    g06945(.A(new_n9375_), .Y(new_n9382_));
  NOR3X1   g06946(.A(new_n9163_), .B(new_n9160_), .C(new_n5952_), .Y(new_n9383_));
  OAI21X1  g06947(.A0(new_n9383_), .A1(new_n9382_), .B0(new_n5982_), .Y(new_n9384_));
  NAND2X1  g06948(.A(new_n9384_), .B(new_n9381_), .Y(new_n9385_));
  NOR3X1   g06949(.A(new_n9167_), .B(new_n9166_), .C(new_n5952_), .Y(new_n9386_));
  OAI21X1  g06950(.A0(new_n9386_), .A1(new_n9382_), .B0(new_n5982_), .Y(new_n9387_));
  AOI22X1  g06951(.A0(new_n9387_), .A1(new_n9244_), .B0(new_n9377_), .B1(new_n3157_), .Y(new_n9388_));
  AND2X1   g06952(.A(new_n9388_), .B(new_n9385_), .Y(new_n9389_));
  AOI21X1  g06953(.A0(new_n9377_), .A1(pi0075), .B0(new_n9248_), .Y(new_n9390_));
  OAI21X1  g06954(.A0(new_n9389_), .A1(pi0075), .B0(new_n9390_), .Y(new_n9391_));
  AOI21X1  g06955(.A0(new_n9391_), .A1(new_n9380_), .B0(new_n6378_), .Y(new_n9392_));
  OAI21X1  g06956(.A0(new_n9392_), .A1(new_n9069_), .B0(new_n6061_), .Y(new_n9393_));
  NOR4X1   g06957(.A(new_n2755_), .B(new_n5096_), .C(new_n5251_), .D(pi0122), .Y(new_n9394_));
  NOR2X1   g06958(.A(new_n6210_), .B(new_n5939_), .Y(new_n9395_));
  NOR3X1   g06959(.A(new_n9395_), .B(new_n9029_), .C(pi0122), .Y(new_n9396_));
  NOR2X1   g06960(.A(new_n9396_), .B(new_n9052_), .Y(new_n9397_));
  OAI21X1  g06961(.A0(new_n9394_), .A1(new_n9029_), .B0(new_n9397_), .Y(new_n9398_));
  MX2X1    g06962(.A(new_n9398_), .B(new_n2740_), .S0(new_n5928_), .Y(new_n9399_));
  OAI21X1  g06963(.A0(new_n9377_), .A1(new_n5928_), .B0(new_n9399_), .Y(new_n9400_));
  AND2X1   g06964(.A(new_n9400_), .B(new_n9035_), .Y(new_n9401_));
  INVX1    g06965(.A(new_n9401_), .Y(new_n9402_));
  NOR3X1   g06966(.A(new_n9397_), .B(new_n9376_), .C(new_n3157_), .Y(new_n9403_));
  NOR3X1   g06967(.A(new_n9242_), .B(new_n9177_), .C(pi0087), .Y(new_n9404_));
  AOI21X1  g06968(.A0(new_n9050_), .A1(new_n9156_), .B0(new_n6191_), .Y(new_n9405_));
  OAI21X1  g06969(.A0(new_n9405_), .A1(new_n9160_), .B0(new_n9404_), .Y(new_n9406_));
  OR2X1    g06970(.A(new_n9059_), .B(new_n6210_), .Y(new_n9407_));
  AND2X1   g06971(.A(new_n9244_), .B(new_n9407_), .Y(new_n9408_));
  OAI21X1  g06972(.A0(new_n9167_), .A1(new_n9166_), .B0(new_n9408_), .Y(new_n9409_));
  AOI21X1  g06973(.A0(new_n9395_), .A1(new_n5952_), .B0(new_n9382_), .Y(new_n9410_));
  INVX1    g06974(.A(new_n9410_), .Y(new_n9411_));
  AOI21X1  g06975(.A0(new_n9409_), .A1(new_n9406_), .B0(new_n9411_), .Y(new_n9412_));
  OAI21X1  g06976(.A0(new_n9412_), .A1(new_n9403_), .B0(new_n3095_), .Y(new_n9413_));
  OAI21X1  g06977(.A0(new_n3138_), .A1(pi0075), .B0(new_n9398_), .Y(new_n9414_));
  OR2X1    g06978(.A(new_n9414_), .B(new_n9376_), .Y(new_n9415_));
  NAND3X1  g06979(.A(new_n9415_), .B(new_n9413_), .C(new_n9247_), .Y(new_n9416_));
  AND2X1   g06980(.A(new_n9416_), .B(new_n9402_), .Y(new_n9417_));
  NOR2X1   g06981(.A(new_n9399_), .B(new_n9034_), .Y(new_n9418_));
  AOI21X1  g06982(.A0(new_n9244_), .A1(new_n9181_), .B0(new_n9404_), .Y(new_n9419_));
  OAI22X1  g06983(.A0(new_n9419_), .A1(new_n5952_), .B0(new_n9397_), .B1(new_n3157_), .Y(new_n9420_));
  AND2X1   g06984(.A(new_n9414_), .B(new_n9247_), .Y(new_n9421_));
  INVX1    g06985(.A(new_n9421_), .Y(new_n9422_));
  AOI21X1  g06986(.A0(new_n9420_), .A1(new_n3095_), .B0(new_n9422_), .Y(new_n9423_));
  OAI21X1  g06987(.A0(new_n9423_), .A1(new_n9418_), .B0(new_n6453_), .Y(new_n9424_));
  OAI21X1  g06988(.A0(new_n9417_), .A1(new_n6378_), .B0(new_n9424_), .Y(new_n9425_));
  AOI22X1  g06989(.A0(new_n9425_), .A1(pi1199), .B0(new_n9032_), .B1(pi0592), .Y(new_n9426_));
  AND2X1   g06990(.A(new_n9426_), .B(new_n9393_), .Y(new_n9427_));
  INVX1    g06991(.A(new_n9427_), .Y(new_n9428_));
  MX2X1    g06992(.A(new_n9428_), .B(new_n9256_), .S0(new_n9154_), .Y(new_n9429_));
  MX2X1    g06993(.A(new_n9427_), .B(new_n9255_), .S0(new_n6183_), .Y(new_n9430_));
  INVX1    g06994(.A(new_n9430_), .Y(new_n9431_));
  MX2X1    g06995(.A(new_n9431_), .B(new_n9429_), .S0(pi0333), .Y(new_n9432_));
  MX2X1    g06996(.A(new_n9431_), .B(new_n9429_), .S0(new_n6172_), .Y(new_n9433_));
  MX2X1    g06997(.A(new_n9433_), .B(new_n9432_), .S0(pi0391), .Y(new_n9434_));
  MX2X1    g06998(.A(new_n9433_), .B(new_n9432_), .S0(new_n6231_), .Y(new_n9435_));
  MX2X1    g06999(.A(new_n9435_), .B(new_n9434_), .S0(pi0392), .Y(new_n9436_));
  MX2X1    g07000(.A(new_n9435_), .B(new_n9434_), .S0(new_n6171_), .Y(new_n9437_));
  MX2X1    g07001(.A(new_n9437_), .B(new_n9436_), .S0(pi0393), .Y(new_n9438_));
  NOR2X1   g07002(.A(new_n9438_), .B(new_n6375_), .Y(new_n9439_));
  MX2X1    g07003(.A(new_n9437_), .B(new_n9436_), .S0(new_n6170_), .Y(new_n9440_));
  OAI21X1  g07004(.A0(new_n9440_), .A1(new_n6713_), .B0(pi0591), .Y(new_n9441_));
  OAI21X1  g07005(.A0(new_n9441_), .A1(new_n9439_), .B0(new_n6168_), .Y(new_n9442_));
  OAI21X1  g07006(.A0(new_n9442_), .A1(new_n9361_), .B0(new_n9028_), .Y(new_n9443_));
  OAI21X1  g07007(.A0(new_n9443_), .A1(new_n9332_), .B0(new_n6633_), .Y(new_n9444_));
  AOI21X1  g07008(.A0(new_n9296_), .A1(new_n9031_), .B0(new_n9444_), .Y(new_n9445_));
  OR4X1    g07009(.A(new_n9445_), .B(new_n9238_), .C(po1038), .D(pi0080), .Y(new_n9446_));
  AND2X1   g07010(.A(new_n9030_), .B(new_n6673_), .Y(new_n9447_));
  OAI21X1  g07011(.A0(new_n9378_), .A1(new_n6378_), .B0(new_n9173_), .Y(new_n9448_));
  INVX1    g07012(.A(new_n9448_), .Y(new_n9449_));
  OAI22X1  g07013(.A0(new_n9399_), .A1(new_n6454_), .B0(new_n9030_), .B1(new_n6120_), .Y(new_n9450_));
  AOI21X1  g07014(.A0(new_n9400_), .A1(new_n6377_), .B0(new_n9450_), .Y(new_n9451_));
  MX2X1    g07015(.A(new_n9451_), .B(new_n9449_), .S0(new_n6061_), .Y(new_n9452_));
  MX2X1    g07016(.A(new_n9452_), .B(new_n9447_), .S0(new_n9154_), .Y(new_n9453_));
  MX2X1    g07017(.A(new_n9452_), .B(new_n9447_), .S0(new_n6183_), .Y(new_n9454_));
  MX2X1    g07018(.A(new_n9454_), .B(new_n9453_), .S0(pi0333), .Y(new_n9455_));
  XOR2X1   g07019(.A(new_n6376_), .B(pi0392), .Y(new_n9456_));
  OR2X1    g07020(.A(new_n9453_), .B(pi0333), .Y(new_n9457_));
  OAI21X1  g07021(.A0(new_n9454_), .A1(new_n6172_), .B0(new_n9457_), .Y(new_n9458_));
  AOI21X1  g07022(.A0(new_n9458_), .A1(new_n6231_), .B0(new_n9456_), .Y(new_n9459_));
  OAI21X1  g07023(.A0(new_n9455_), .A1(new_n6231_), .B0(new_n9459_), .Y(new_n9460_));
  NAND2X1  g07024(.A(new_n9458_), .B(pi0391), .Y(new_n9461_));
  OR2X1    g07025(.A(new_n9455_), .B(pi0391), .Y(new_n9462_));
  AND2X1   g07026(.A(new_n9462_), .B(new_n9456_), .Y(new_n9463_));
  AOI21X1  g07027(.A0(new_n9463_), .A1(new_n9461_), .B0(new_n6074_), .Y(new_n9464_));
  NAND2X1  g07028(.A(new_n6687_), .B(new_n6673_), .Y(new_n9465_));
  OAI21X1  g07029(.A0(new_n6678_), .A1(new_n6638_), .B0(new_n6055_), .Y(new_n9466_));
  AND2X1   g07030(.A(new_n9466_), .B(new_n6702_), .Y(new_n9467_));
  AOI21X1  g07031(.A0(new_n9467_), .A1(new_n9465_), .B0(new_n9032_), .Y(new_n9468_));
  OAI21X1  g07032(.A0(new_n9468_), .A1(pi0591), .B0(new_n6168_), .Y(new_n9469_));
  AOI21X1  g07033(.A0(new_n9464_), .A1(new_n9460_), .B0(new_n9469_), .Y(new_n9470_));
  INVX1    g07034(.A(new_n9447_), .Y(new_n9471_));
  OR4X1    g07035(.A(new_n9032_), .B(new_n6674_), .C(new_n6656_), .D(new_n6064_), .Y(new_n9472_));
  AND2X1   g07036(.A(new_n9472_), .B(new_n9471_), .Y(new_n9473_));
  NOR4X1   g07037(.A(new_n9032_), .B(new_n6674_), .C(new_n6656_), .D(new_n6060_), .Y(new_n9474_));
  NOR2X1   g07038(.A(new_n9474_), .B(new_n9447_), .Y(new_n9475_));
  MX2X1    g07039(.A(new_n9475_), .B(new_n9473_), .S0(pi0461), .Y(new_n9476_));
  MX2X1    g07040(.A(new_n9475_), .B(new_n9473_), .S0(new_n5879_), .Y(new_n9477_));
  MX2X1    g07041(.A(new_n9477_), .B(new_n9476_), .S0(pi0357), .Y(new_n9478_));
  MX2X1    g07042(.A(new_n9477_), .B(new_n9476_), .S0(new_n5878_), .Y(new_n9479_));
  MX2X1    g07043(.A(new_n9479_), .B(new_n9478_), .S0(pi0356), .Y(new_n9480_));
  INVX1    g07044(.A(new_n9480_), .Y(new_n9481_));
  MX2X1    g07045(.A(new_n9479_), .B(new_n9478_), .S0(new_n5877_), .Y(new_n9482_));
  AOI21X1  g07046(.A0(new_n9482_), .A1(new_n9116_), .B0(new_n9323_), .Y(new_n9483_));
  OAI21X1  g07047(.A0(new_n9481_), .A1(new_n9116_), .B0(new_n9483_), .Y(new_n9484_));
  NAND2X1  g07048(.A(new_n9482_), .B(pi0354), .Y(new_n9485_));
  AOI21X1  g07049(.A0(new_n9480_), .A1(new_n9116_), .B0(new_n5874_), .Y(new_n9486_));
  AOI21X1  g07050(.A0(new_n9486_), .A1(new_n9485_), .B0(pi0591), .Y(new_n9487_));
  AOI21X1  g07051(.A0(new_n9487_), .A1(new_n9484_), .B0(new_n9115_), .Y(new_n9488_));
  OR2X1    g07052(.A(new_n9488_), .B(pi0588), .Y(new_n9489_));
  AND2X1   g07053(.A(new_n6550_), .B(pi0592), .Y(new_n9490_));
  OAI21X1  g07054(.A0(new_n6726_), .A1(new_n6550_), .B0(new_n6310_), .Y(new_n9491_));
  OAI21X1  g07055(.A0(new_n9491_), .A1(new_n9490_), .B0(new_n9030_), .Y(new_n9492_));
  MX2X1    g07056(.A(new_n9492_), .B(new_n9471_), .S0(new_n6528_), .Y(new_n9493_));
  INVX1    g07057(.A(new_n9493_), .Y(new_n9494_));
  MX2X1    g07058(.A(new_n9492_), .B(new_n9471_), .S0(pi0428), .Y(new_n9495_));
  INVX1    g07059(.A(new_n9495_), .Y(new_n9496_));
  MX2X1    g07060(.A(new_n9496_), .B(new_n9494_), .S0(new_n6527_), .Y(new_n9497_));
  MX2X1    g07061(.A(new_n9496_), .B(new_n9494_), .S0(pi0427), .Y(new_n9498_));
  MX2X1    g07062(.A(new_n9498_), .B(new_n9497_), .S0(new_n6582_), .Y(new_n9499_));
  MX2X1    g07063(.A(new_n9498_), .B(new_n9497_), .S0(pi0430), .Y(new_n9500_));
  MX2X1    g07064(.A(new_n9500_), .B(new_n9499_), .S0(new_n6585_), .Y(new_n9501_));
  OR2X1    g07065(.A(new_n9501_), .B(pi0445), .Y(new_n9502_));
  MX2X1    g07066(.A(new_n9500_), .B(new_n9499_), .S0(pi0426), .Y(new_n9503_));
  OAI21X1  g07067(.A0(new_n9503_), .A1(new_n6589_), .B0(new_n9502_), .Y(new_n9504_));
  MX2X1    g07068(.A(new_n9503_), .B(new_n9501_), .S0(pi0445), .Y(new_n9505_));
  OAI21X1  g07069(.A0(new_n9505_), .A1(pi0448), .B0(new_n6525_), .Y(new_n9506_));
  AOI21X1  g07070(.A0(new_n9504_), .A1(pi0448), .B0(new_n9506_), .Y(new_n9507_));
  OAI21X1  g07071(.A0(new_n9505_), .A1(new_n6522_), .B0(new_n6623_), .Y(new_n9508_));
  AOI21X1  g07072(.A0(new_n9504_), .A1(new_n6522_), .B0(new_n9508_), .Y(new_n9509_));
  OR2X1    g07073(.A(new_n9509_), .B(new_n6061_), .Y(new_n9510_));
  AOI21X1  g07074(.A0(new_n9492_), .A1(new_n6061_), .B0(new_n6630_), .Y(new_n9511_));
  OAI21X1  g07075(.A0(new_n9510_), .A1(new_n9507_), .B0(new_n9511_), .Y(new_n9512_));
  AOI21X1  g07076(.A0(new_n9512_), .A1(new_n9031_), .B0(new_n6077_), .Y(new_n9513_));
  OAI21X1  g07077(.A0(new_n9489_), .A1(new_n9470_), .B0(new_n9513_), .Y(new_n9514_));
  OR2X1    g07078(.A(new_n6520_), .B(pi0080), .Y(new_n9515_));
  AOI21X1  g07079(.A0(new_n9030_), .A1(new_n6077_), .B0(new_n9515_), .Y(new_n9516_));
  AOI21X1  g07080(.A0(new_n9516_), .A1(new_n9514_), .B0(pi0217), .Y(new_n9517_));
  OAI21X1  g07081(.A0(new_n9030_), .A1(pi0080), .B0(pi0217), .Y(new_n9518_));
  NAND2X1  g07082(.A(new_n9518_), .B(new_n6748_), .Y(new_n9519_));
  AOI21X1  g07083(.A0(new_n9517_), .A1(new_n9446_), .B0(new_n9519_), .Y(po0238));
  OR4X1    g07084(.A(new_n8454_), .B(po1038), .C(new_n3131_), .D(new_n2461_), .Y(new_n9521_));
  NAND3X1  g07085(.A(new_n2510_), .B(new_n7734_), .C(pi0081), .Y(new_n9522_));
  INVX1    g07086(.A(pi0068), .Y(new_n9523_));
  OR2X1    g07087(.A(new_n2468_), .B(pi0036), .Y(new_n9524_));
  OR4X1    g07088(.A(new_n8265_), .B(new_n9524_), .C(pi0081), .D(new_n9523_), .Y(new_n9525_));
  OR4X1    g07089(.A(new_n9525_), .B(new_n6782_), .C(new_n2647_), .D(pi0064), .Y(new_n9526_));
  AOI21X1  g07090(.A0(new_n9526_), .A1(new_n9522_), .B0(new_n9521_), .Y(po0239));
  AND2X1   g07091(.A(pi0314), .B(pi0069), .Y(new_n9528_));
  INVX1    g07092(.A(pi0066), .Y(new_n9529_));
  NOR4X1   g07093(.A(new_n2470_), .B(new_n2464_), .C(pi0073), .D(new_n9529_), .Y(new_n9530_));
  AOI21X1  g07094(.A0(new_n9528_), .A1(new_n2612_), .B0(new_n9530_), .Y(new_n9531_));
  NOR4X1   g07095(.A(new_n9531_), .B(new_n8325_), .C(new_n8324_), .D(new_n2463_), .Y(po0240));
  INVX1    g07096(.A(new_n2617_), .Y(new_n9533_));
  NOR3X1   g07097(.A(new_n8325_), .B(new_n2484_), .C(new_n2478_), .Y(new_n9534_));
  OR4X1    g07098(.A(new_n6775_), .B(pi0069), .C(pi0068), .D(pi0067), .Y(new_n9535_));
  OR4X1    g07099(.A(new_n9535_), .B(new_n2621_), .C(new_n2468_), .D(pi0036), .Y(new_n9536_));
  NAND2X1  g07100(.A(new_n9536_), .B(new_n2614_), .Y(new_n9537_));
  AND2X1   g07101(.A(new_n9537_), .B(new_n9534_), .Y(new_n9538_));
  AOI21X1  g07102(.A0(new_n9538_), .A1(new_n9533_), .B0(pi0314), .Y(new_n9539_));
  NOR4X1   g07103(.A(new_n9535_), .B(new_n2621_), .C(new_n9524_), .D(new_n2463_), .Y(new_n9540_));
  AOI21X1  g07104(.A0(new_n9540_), .A1(new_n9534_), .B0(new_n7734_), .Y(new_n9541_));
  NOR3X1   g07105(.A(new_n9541_), .B(new_n9539_), .C(new_n7670_), .Y(po0241));
  NAND2X1  g07106(.A(new_n8505_), .B(new_n3130_), .Y(new_n9543_));
  AND2X1   g07107(.A(pi0299), .B(pi0211), .Y(new_n9544_));
  AND2X1   g07108(.A(pi0299), .B(pi0219), .Y(new_n9545_));
  NOR3X1   g07109(.A(new_n9545_), .B(new_n9544_), .C(new_n8131_), .Y(new_n9546_));
  INVX1    g07110(.A(new_n9546_), .Y(new_n9547_));
  NOR3X1   g07111(.A(new_n9547_), .B(new_n9543_), .C(po1038), .Y(po0242));
  NOR3X1   g07112(.A(new_n8325_), .B(new_n2463_), .C(pi0069), .Y(new_n9549_));
  NOR3X1   g07113(.A(new_n8544_), .B(new_n2469_), .C(new_n2465_), .Y(new_n9550_));
  NOR2X1   g07114(.A(new_n8326_), .B(pi0314), .Y(new_n9551_));
  AOI22X1  g07115(.A0(new_n9551_), .A1(new_n9550_), .B0(new_n9549_), .B1(new_n5154_), .Y(new_n9552_));
  NOR2X1   g07116(.A(new_n9552_), .B(new_n8324_), .Y(po0243));
  AOI22X1  g07117(.A0(new_n8519_), .A1(new_n5962_), .B0(new_n8516_), .B1(new_n5960_), .Y(new_n9554_));
  NOR2X1   g07118(.A(new_n9554_), .B(new_n8245_), .Y(po0244));
  NOR3X1   g07119(.A(new_n8325_), .B(new_n2664_), .C(new_n2478_), .Y(new_n9556_));
  NOR4X1   g07120(.A(new_n7749_), .B(new_n8284_), .C(new_n2484_), .D(new_n7734_), .Y(new_n9557_));
  AND2X1   g07121(.A(new_n9557_), .B(new_n9556_), .Y(po0245));
  AOI21X1  g07122(.A0(new_n8277_), .A1(new_n5938_), .B0(pi1093), .Y(new_n9559_));
  NOR4X1   g07123(.A(pi0110), .B(pi0091), .C(pi0058), .D(pi0047), .Y(new_n9560_));
  NOR4X1   g07124(.A(new_n9039_), .B(new_n8275_), .C(new_n8252_), .D(pi0094), .Y(new_n9561_));
  NAND4X1  g07125(.A(new_n9561_), .B(new_n9560_), .C(new_n7667_), .D(new_n5938_), .Y(new_n9562_));
  AND2X1   g07126(.A(new_n9562_), .B(pi1093), .Y(new_n9563_));
  OR4X1    g07127(.A(new_n9563_), .B(new_n9559_), .C(new_n7607_), .D(new_n3131_), .Y(new_n9564_));
  AND2X1   g07128(.A(new_n5938_), .B(new_n2486_), .Y(new_n9565_));
  NAND4X1  g07129(.A(new_n9565_), .B(new_n3130_), .C(new_n3002_), .D(new_n2756_), .Y(new_n9566_));
  NOR3X1   g07130(.A(new_n9566_), .B(new_n8561_), .C(new_n2682_), .Y(new_n9567_));
  OAI21X1  g07131(.A0(new_n9567_), .A1(new_n6077_), .B0(new_n6520_), .Y(new_n9568_));
  AOI21X1  g07132(.A0(new_n9564_), .A1(new_n6077_), .B0(new_n9568_), .Y(po0246));
  NAND4X1  g07133(.A(new_n7680_), .B(new_n6786_), .C(new_n6871_), .D(new_n2460_), .Y(new_n9570_));
  NOR3X1   g07134(.A(new_n9570_), .B(new_n5908_), .C(new_n2726_), .Y(new_n9571_));
  AND2X1   g07135(.A(new_n6520_), .B(new_n3135_), .Y(new_n9572_));
  INVX1    g07136(.A(new_n9572_), .Y(new_n9573_));
  NOR4X1   g07137(.A(new_n9573_), .B(new_n5843_), .C(new_n3003_), .D(pi0092), .Y(new_n9574_));
  OAI21X1  g07138(.A0(new_n9571_), .A1(pi0070), .B0(new_n9574_), .Y(new_n9575_));
  AOI21X1  g07139(.A0(new_n6805_), .A1(pi0070), .B0(new_n9575_), .Y(po0247));
  OAI21X1  g07140(.A0(new_n7268_), .A1(pi1050), .B0(new_n2701_), .Y(new_n9577_));
  NAND2X1  g07141(.A(new_n9577_), .B(new_n8470_), .Y(new_n9578_));
  NOR3X1   g07142(.A(new_n9578_), .B(new_n5898_), .C(new_n2702_), .Y(po0248));
  INVX1    g07143(.A(new_n7686_), .Y(new_n9580_));
  INVX1    g07144(.A(new_n5942_), .Y(new_n9581_));
  OAI22X1  g07145(.A0(new_n7662_), .A1(new_n7657_), .B0(new_n9581_), .B1(pi0058), .Y(new_n9582_));
  AND2X1   g07146(.A(new_n7667_), .B(new_n2778_), .Y(new_n9583_));
  OR4X1    g07147(.A(new_n8314_), .B(new_n2778_), .C(new_n2744_), .D(new_n5787_), .Y(new_n9584_));
  OAI21X1  g07148(.A0(new_n9584_), .A1(new_n9581_), .B0(new_n2959_), .Y(new_n9585_));
  AOI21X1  g07149(.A0(new_n9583_), .A1(new_n9582_), .B0(new_n9585_), .Y(new_n9586_));
  NOR4X1   g07150(.A(new_n9586_), .B(new_n9580_), .C(new_n5965_), .D(pi0038), .Y(po0249));
  NAND4X1  g07151(.A(new_n3137_), .B(new_n3098_), .C(pi1050), .D(new_n7734_), .Y(new_n9588_));
  OR4X1    g07152(.A(new_n9588_), .B(new_n3003_), .C(new_n2555_), .D(new_n3100_), .Y(new_n9589_));
  INVX1    g07153(.A(new_n8244_), .Y(new_n9590_));
  NOR4X1   g07154(.A(new_n2953_), .B(new_n2437_), .C(new_n2438_), .D(pi0215), .Y(new_n9591_));
  NOR4X1   g07155(.A(pi0299), .B(new_n2961_), .C(pi0223), .D(new_n2960_), .Y(new_n9592_));
  AOI22X1  g07156(.A0(new_n9592_), .A1(new_n5962_), .B0(new_n9591_), .B1(new_n5960_), .Y(new_n9593_));
  OR4X1    g07157(.A(new_n9593_), .B(new_n9590_), .C(new_n3139_), .D(pi0100), .Y(new_n9594_));
  AOI21X1  g07158(.A0(new_n9594_), .A1(new_n9589_), .B0(new_n9573_), .Y(po0250));
  OR4X1    g07159(.A(new_n3003_), .B(new_n2709_), .C(pi1050), .D(pi0070), .Y(new_n9596_));
  AND2X1   g07160(.A(new_n9572_), .B(new_n3230_), .Y(new_n9597_));
  INVX1    g07161(.A(new_n5011_), .Y(new_n9598_));
  NOR4X1   g07162(.A(new_n8314_), .B(new_n9598_), .C(new_n2726_), .D(new_n2531_), .Y(new_n9599_));
  OAI21X1  g07163(.A0(new_n9599_), .A1(pi0092), .B0(new_n9597_), .Y(new_n9600_));
  AOI21X1  g07164(.A0(new_n9596_), .A1(pi0092), .B0(new_n9600_), .Y(po0251));
  NAND4X1  g07165(.A(new_n8300_), .B(new_n6806_), .C(new_n2491_), .D(new_n2726_), .Y(new_n9602_));
  INVX1    g07166(.A(new_n9602_), .Y(new_n9603_));
  AOI21X1  g07167(.A0(new_n9603_), .A1(new_n2723_), .B0(new_n2756_), .Y(new_n9604_));
  NOR4X1   g07168(.A(new_n2498_), .B(pi0841), .C(pi0060), .D(pi0053), .Y(new_n9605_));
  AOI21X1  g07169(.A0(new_n8298_), .A1(new_n9605_), .B0(new_n2594_), .Y(new_n9606_));
  NAND4X1  g07170(.A(new_n7667_), .B(new_n2505_), .C(pi0252), .D(new_n2502_), .Y(new_n9607_));
  OAI22X1  g07171(.A0(new_n9607_), .A1(new_n9606_), .B0(new_n9604_), .B1(new_n2785_), .Y(new_n9608_));
  AND2X1   g07172(.A(new_n9608_), .B(new_n6773_), .Y(new_n9609_));
  OAI22X1  g07173(.A0(new_n9609_), .A1(new_n9603_), .B0(new_n9608_), .B1(new_n3053_), .Y(new_n9610_));
  OAI21X1  g07174(.A0(new_n9603_), .A1(new_n6763_), .B0(new_n7668_), .Y(new_n9611_));
  AOI21X1  g07175(.A0(new_n9610_), .A1(new_n6763_), .B0(new_n9611_), .Y(po0252));
  OR4X1    g07176(.A(new_n8531_), .B(new_n5257_), .C(new_n5058_), .D(new_n3285_), .Y(new_n9613_));
  NOR4X1   g07177(.A(new_n8534_), .B(new_n8533_), .C(new_n5074_), .D(pi0216), .Y(new_n9614_));
  OAI21X1  g07178(.A0(new_n5256_), .A1(new_n5249_), .B0(new_n9614_), .Y(new_n9615_));
  AND2X1   g07179(.A(new_n9615_), .B(pi0039), .Y(new_n9616_));
  NOR4X1   g07180(.A(new_n8557_), .B(new_n2458_), .C(new_n2540_), .D(pi0032), .Y(new_n9617_));
  NAND4X1  g07181(.A(new_n7667_), .B(new_n2491_), .C(new_n2726_), .D(new_n2445_), .Y(new_n9618_));
  OAI21X1  g07182(.A0(new_n9618_), .A1(new_n9570_), .B0(new_n2959_), .Y(new_n9619_));
  OAI21X1  g07183(.A0(new_n9619_), .A1(new_n9617_), .B0(new_n7689_), .Y(new_n9620_));
  AOI21X1  g07184(.A0(new_n9616_), .A1(new_n9613_), .B0(new_n9620_), .Y(po0253));
  NAND4X1  g07185(.A(new_n7774_), .B(new_n2457_), .C(pi0095), .D(new_n2456_), .Y(new_n9622_));
  NOR3X1   g07186(.A(po0840), .B(new_n2897_), .C(new_n2454_), .Y(new_n9623_));
  AND2X1   g07187(.A(new_n6773_), .B(pi0479), .Y(new_n9624_));
  NAND4X1  g07188(.A(new_n2715_), .B(pi0096), .C(new_n5134_), .D(new_n2518_), .Y(new_n9625_));
  NOR4X1   g07189(.A(new_n9625_), .B(new_n9624_), .C(new_n2727_), .D(new_n2710_), .Y(new_n9626_));
  OAI21X1  g07190(.A0(new_n9626_), .A1(new_n9623_), .B0(new_n2540_), .Y(new_n9627_));
  AOI21X1  g07191(.A0(new_n9627_), .A1(new_n9622_), .B0(new_n7749_), .Y(po0254));
  INVX1    g07192(.A(pi0593), .Y(new_n9629_));
  OR4X1    g07193(.A(new_n8536_), .B(new_n5257_), .C(new_n9629_), .D(new_n2959_), .Y(new_n9630_));
  AOI21X1  g07194(.A0(new_n9624_), .A1(new_n5019_), .B0(po0740), .Y(new_n9631_));
  OR4X1    g07195(.A(new_n9631_), .B(new_n8582_), .C(new_n7673_), .D(pi0096), .Y(new_n9632_));
  AOI21X1  g07196(.A0(new_n9632_), .A1(new_n9630_), .B0(new_n7690_), .Y(po0255));
  MX2X1    g07197(.A(new_n8577_), .B(new_n3074_), .S0(pi0092), .Y(new_n9634_));
  NAND4X1  g07198(.A(new_n9572_), .B(new_n3230_), .C(pi1050), .D(pi0314), .Y(new_n9635_));
  NOR2X1   g07199(.A(new_n9635_), .B(new_n9634_), .Y(po0256));
  AND2X1   g07200(.A(pi0099), .B(new_n2548_), .Y(new_n9637_));
  OR2X1    g07201(.A(new_n9637_), .B(new_n6291_), .Y(new_n9638_));
  AOI21X1  g07202(.A0(new_n9637_), .A1(new_n2724_), .B0(new_n7761_), .Y(new_n9639_));
  INVX1    g07203(.A(new_n9637_), .Y(new_n9640_));
  NOR2X1   g07204(.A(new_n9640_), .B(new_n7776_), .Y(new_n9641_));
  AOI21X1  g07205(.A0(new_n8200_), .A1(new_n5089_), .B0(new_n9641_), .Y(new_n9642_));
  OAI21X1  g07206(.A0(new_n9642_), .A1(new_n7874_), .B0(new_n9639_), .Y(new_n9643_));
  AOI21X1  g07207(.A0(new_n9643_), .A1(new_n9638_), .B0(pi0039), .Y(new_n9644_));
  NOR4X1   g07208(.A(new_n7784_), .B(new_n4613_), .C(new_n6900_), .D(pi0072), .Y(new_n9645_));
  NOR3X1   g07209(.A(pi0299), .B(new_n7008_), .C(pi0072), .Y(new_n9646_));
  AND2X1   g07210(.A(new_n9646_), .B(new_n7781_), .Y(new_n9647_));
  AOI21X1  g07211(.A0(new_n9645_), .A1(pi0299), .B0(new_n9647_), .Y(new_n9648_));
  OR2X1    g07212(.A(new_n9648_), .B(new_n5237_), .Y(new_n9649_));
  AND2X1   g07213(.A(new_n9649_), .B(pi0039), .Y(new_n9650_));
  OR2X1    g07214(.A(new_n9650_), .B(new_n5788_), .Y(new_n9651_));
  AOI21X1  g07215(.A0(new_n9640_), .A1(new_n2959_), .B0(new_n9650_), .Y(new_n9652_));
  AOI21X1  g07216(.A0(new_n9652_), .A1(new_n5788_), .B0(new_n3095_), .Y(new_n9653_));
  OAI21X1  g07217(.A0(new_n9651_), .A1(new_n9644_), .B0(new_n9653_), .Y(new_n9654_));
  AOI21X1  g07218(.A0(pi0072), .A1(pi0041), .B0(new_n7770_), .Y(new_n9655_));
  INVX1    g07219(.A(new_n9655_), .Y(new_n9656_));
  NOR2X1   g07220(.A(new_n9656_), .B(new_n7819_), .Y(new_n9657_));
  NOR3X1   g07221(.A(new_n9657_), .B(new_n8083_), .C(new_n2724_), .Y(new_n9658_));
  INVX1    g07222(.A(new_n7823_), .Y(new_n9659_));
  AOI21X1  g07223(.A0(new_n9655_), .A1(new_n9659_), .B0(new_n8084_), .Y(new_n9660_));
  OAI21X1  g07224(.A0(new_n9660_), .A1(new_n9658_), .B0(pi0228), .Y(new_n9661_));
  NOR4X1   g07225(.A(new_n7853_), .B(new_n7903_), .C(pi0101), .D(pi0044), .Y(new_n9662_));
  NOR2X1   g07226(.A(new_n9662_), .B(pi0228), .Y(new_n9663_));
  OAI21X1  g07227(.A0(new_n9656_), .A1(new_n7859_), .B0(new_n9663_), .Y(new_n9664_));
  AND2X1   g07228(.A(new_n9664_), .B(new_n2959_), .Y(new_n9665_));
  OR2X1    g07229(.A(new_n9648_), .B(new_n7892_), .Y(new_n9666_));
  AOI21X1  g07230(.A0(new_n8218_), .A1(pi0287), .B0(new_n9666_), .Y(new_n9667_));
  OR2X1    g07231(.A(new_n9667_), .B(new_n5792_), .Y(new_n9668_));
  AOI21X1  g07232(.A0(new_n9665_), .A1(new_n9661_), .B0(new_n9668_), .Y(new_n9669_));
  INVX1    g07233(.A(new_n9639_), .Y(new_n9670_));
  OAI22X1  g07234(.A0(new_n9640_), .A1(new_n7872_), .B0(new_n7767_), .B1(new_n7903_), .Y(new_n9671_));
  AND2X1   g07235(.A(new_n9671_), .B(new_n7873_), .Y(new_n9672_));
  OAI21X1  g07236(.A0(new_n9672_), .A1(new_n9670_), .B0(new_n9638_), .Y(new_n9673_));
  AOI21X1  g07237(.A0(new_n9673_), .A1(new_n2959_), .B0(new_n9650_), .Y(new_n9674_));
  INVX1    g07238(.A(new_n9652_), .Y(new_n9675_));
  AOI21X1  g07239(.A0(new_n9675_), .A1(pi0038), .B0(pi0087), .Y(new_n9676_));
  OAI21X1  g07240(.A0(new_n9674_), .A1(new_n5086_), .B0(new_n9676_), .Y(new_n9677_));
  NOR3X1   g07241(.A(new_n7765_), .B(new_n7903_), .C(new_n3013_), .Y(new_n9678_));
  AOI21X1  g07242(.A0(new_n7870_), .A1(pi0228), .B0(new_n9640_), .Y(new_n9679_));
  OR4X1    g07243(.A(new_n9679_), .B(new_n9678_), .C(new_n3066_), .D(pi0100), .Y(new_n9680_));
  AOI21X1  g07244(.A0(new_n9675_), .A1(new_n3138_), .B0(new_n3156_), .Y(new_n9681_));
  AOI21X1  g07245(.A0(new_n9681_), .A1(new_n9680_), .B0(pi0075), .Y(new_n9682_));
  OAI21X1  g07246(.A0(new_n9677_), .A1(new_n9669_), .B0(new_n9682_), .Y(new_n9683_));
  AOI21X1  g07247(.A0(new_n9683_), .A1(new_n9654_), .B0(new_n6309_), .Y(new_n9684_));
  OAI21X1  g07248(.A0(new_n9652_), .A1(new_n5893_), .B0(new_n6520_), .Y(new_n9685_));
  AOI21X1  g07249(.A0(new_n9645_), .A1(pi0232), .B0(new_n2959_), .Y(new_n9686_));
  OAI22X1  g07250(.A0(new_n9637_), .A1(pi0039), .B0(new_n5118_), .B1(pi0057), .Y(new_n9687_));
  OAI22X1  g07251(.A0(new_n9687_), .A1(new_n9686_), .B0(new_n9685_), .B1(new_n9684_), .Y(po0257));
  INVX1    g07252(.A(new_n5929_), .Y(new_n9689_));
  OR2X1    g07253(.A(new_n7611_), .B(new_n5930_), .Y(new_n9690_));
  AND2X1   g07254(.A(new_n9690_), .B(pi0129), .Y(new_n9691_));
  AOI21X1  g07255(.A0(po1057), .A1(new_n5088_), .B0(new_n5098_), .Y(new_n9692_));
  NOR2X1   g07256(.A(new_n9692_), .B(new_n5083_), .Y(new_n9693_));
  NAND2X1  g07257(.A(new_n7611_), .B(pi0129), .Y(new_n9694_));
  AOI21X1  g07258(.A0(new_n9694_), .A1(new_n7613_), .B0(new_n9693_), .Y(new_n9695_));
  OAI21X1  g07259(.A0(new_n9691_), .A1(new_n9689_), .B0(new_n9695_), .Y(new_n9696_));
  NOR4X1   g07260(.A(new_n7188_), .B(new_n3026_), .C(pi0075), .D(pi0038), .Y(new_n9697_));
  NOR4X1   g07261(.A(new_n6812_), .B(new_n6810_), .C(new_n6773_), .D(pi0024), .Y(new_n9698_));
  AOI21X1  g07262(.A0(new_n9697_), .A1(new_n9696_), .B0(new_n9698_), .Y(new_n9699_));
  NOR3X1   g07263(.A(new_n9699_), .B(new_n8306_), .C(new_n3074_), .Y(po0258));
  AND2X1   g07264(.A(pi0101), .B(new_n2548_), .Y(new_n9701_));
  OR2X1    g07265(.A(new_n9701_), .B(new_n6291_), .Y(new_n9702_));
  AOI21X1  g07266(.A0(new_n9701_), .A1(new_n2724_), .B0(new_n7761_), .Y(new_n9703_));
  OAI21X1  g07267(.A0(new_n5093_), .A1(new_n5090_), .B0(new_n2723_), .Y(new_n9704_));
  OR2X1    g07268(.A(new_n7775_), .B(pi0044), .Y(new_n9705_));
  AOI22X1  g07269(.A0(new_n9705_), .A1(new_n9701_), .B0(new_n7766_), .B1(new_n5932_), .Y(new_n9706_));
  OAI21X1  g07270(.A0(new_n9706_), .A1(new_n9704_), .B0(new_n9703_), .Y(new_n9707_));
  AOI21X1  g07271(.A0(new_n9707_), .A1(new_n9702_), .B0(pi0039), .Y(new_n9708_));
  INVX1    g07272(.A(new_n3215_), .Y(new_n9709_));
  NOR4X1   g07273(.A(new_n5057_), .B(new_n9709_), .C(new_n6900_), .D(pi0072), .Y(new_n9710_));
  NAND4X1  g07274(.A(new_n7780_), .B(pi0174), .C(new_n7548_), .D(new_n2548_), .Y(new_n9711_));
  AOI21X1  g07275(.A0(new_n9711_), .A1(new_n2953_), .B0(new_n5237_), .Y(new_n9712_));
  OAI21X1  g07276(.A0(new_n9710_), .A1(new_n2953_), .B0(new_n9712_), .Y(new_n9713_));
  AND2X1   g07277(.A(new_n9713_), .B(pi0039), .Y(new_n9714_));
  OR2X1    g07278(.A(new_n9714_), .B(new_n5788_), .Y(new_n9715_));
  AOI21X1  g07279(.A0(pi0101), .A1(new_n2548_), .B0(pi0039), .Y(new_n9716_));
  AOI21X1  g07280(.A0(new_n9713_), .A1(pi0039), .B0(new_n9716_), .Y(new_n9717_));
  AOI21X1  g07281(.A0(new_n9717_), .A1(new_n5788_), .B0(new_n3095_), .Y(new_n9718_));
  OAI21X1  g07282(.A0(new_n9715_), .A1(new_n9708_), .B0(new_n9718_), .Y(new_n9719_));
  OAI21X1  g07283(.A0(new_n7809_), .A1(pi0101), .B0(new_n2723_), .Y(new_n9720_));
  AOI21X1  g07284(.A0(new_n7818_), .A1(pi0101), .B0(new_n9720_), .Y(new_n9721_));
  OR2X1    g07285(.A(new_n7826_), .B(new_n2723_), .Y(new_n9722_));
  AOI21X1  g07286(.A0(new_n7822_), .A1(pi0101), .B0(new_n9722_), .Y(new_n9723_));
  OAI21X1  g07287(.A0(new_n9723_), .A1(new_n9721_), .B0(pi0228), .Y(new_n9724_));
  NAND2X1  g07288(.A(new_n7858_), .B(pi0101), .Y(new_n9725_));
  NAND3X1  g07289(.A(new_n9725_), .B(new_n7855_), .C(new_n3013_), .Y(new_n9726_));
  AND2X1   g07290(.A(new_n9726_), .B(new_n2959_), .Y(new_n9727_));
  NOR3X1   g07291(.A(new_n5057_), .B(new_n9709_), .C(new_n6900_), .Y(new_n9728_));
  AOI21X1  g07292(.A0(new_n9728_), .A1(new_n8219_), .B0(new_n2953_), .Y(new_n9729_));
  NOR4X1   g07293(.A(new_n8220_), .B(new_n8813_), .C(new_n7008_), .D(pi0144), .Y(new_n9730_));
  OAI21X1  g07294(.A0(new_n9730_), .A1(pi0299), .B0(new_n7891_), .Y(new_n9731_));
  OAI21X1  g07295(.A0(new_n9731_), .A1(new_n9729_), .B0(new_n3277_), .Y(new_n9732_));
  AOI21X1  g07296(.A0(new_n9727_), .A1(new_n9724_), .B0(new_n9732_), .Y(new_n9733_));
  INVX1    g07297(.A(new_n9703_), .Y(new_n9734_));
  OAI21X1  g07298(.A0(new_n8223_), .A1(pi0044), .B0(new_n9701_), .Y(new_n9735_));
  AOI21X1  g07299(.A0(new_n9735_), .A1(new_n7767_), .B0(new_n9704_), .Y(new_n9736_));
  OAI21X1  g07300(.A0(new_n9736_), .A1(new_n9734_), .B0(new_n9702_), .Y(new_n9737_));
  AOI21X1  g07301(.A0(new_n9737_), .A1(new_n2959_), .B0(new_n9714_), .Y(new_n9738_));
  OR2X1    g07302(.A(new_n9717_), .B(new_n2996_), .Y(new_n9739_));
  AND2X1   g07303(.A(new_n9739_), .B(new_n3156_), .Y(new_n9740_));
  OAI21X1  g07304(.A0(new_n9738_), .A1(new_n5086_), .B0(new_n9740_), .Y(new_n9741_));
  OR2X1    g07305(.A(new_n8231_), .B(pi0101), .Y(new_n9742_));
  OAI21X1  g07306(.A0(new_n8230_), .A1(new_n7869_), .B0(new_n9701_), .Y(new_n9743_));
  NAND3X1  g07307(.A(new_n9743_), .B(new_n9742_), .C(new_n2959_), .Y(new_n9744_));
  AOI21X1  g07308(.A0(new_n9713_), .A1(pi0039), .B0(new_n3156_), .Y(new_n9745_));
  AOI21X1  g07309(.A0(new_n9745_), .A1(new_n9744_), .B0(pi0075), .Y(new_n9746_));
  OAI21X1  g07310(.A0(new_n9741_), .A1(new_n9733_), .B0(new_n9746_), .Y(new_n9747_));
  AOI21X1  g07311(.A0(new_n9747_), .A1(new_n9719_), .B0(new_n6309_), .Y(new_n9748_));
  OAI21X1  g07312(.A0(new_n9717_), .A1(new_n5893_), .B0(new_n6520_), .Y(new_n9749_));
  AOI21X1  g07313(.A0(new_n9710_), .A1(pi0232), .B0(new_n2959_), .Y(new_n9750_));
  OR2X1    g07314(.A(new_n9716_), .B(new_n6520_), .Y(new_n9751_));
  OAI22X1  g07315(.A0(new_n9751_), .A1(new_n9750_), .B0(new_n9749_), .B1(new_n9748_), .Y(po0259));
  INVX1    g07316(.A(new_n2669_), .Y(new_n9753_));
  INVX1    g07317(.A(new_n6871_), .Y(new_n9754_));
  NOR4X1   g07318(.A(new_n9521_), .B(new_n9754_), .C(new_n9753_), .D(new_n2472_), .Y(po0260));
  OAI21X1  g07319(.A0(new_n9556_), .A1(pi0109), .B0(new_n5137_), .Y(new_n9756_));
  NOR3X1   g07320(.A(new_n7749_), .B(new_n8284_), .C(new_n5007_), .Y(new_n9757_));
  NOR3X1   g07321(.A(new_n2818_), .B(new_n2480_), .C(new_n2481_), .Y(new_n9758_));
  OAI21X1  g07322(.A0(new_n9758_), .A1(new_n7734_), .B0(new_n9757_), .Y(new_n9759_));
  AOI21X1  g07323(.A0(new_n9756_), .A1(new_n7734_), .B0(new_n9759_), .Y(po0261));
  OAI21X1  g07324(.A0(new_n6763_), .A1(new_n6633_), .B0(new_n7608_), .Y(new_n9761_));
  NAND3X1  g07325(.A(new_n9761_), .B(new_n7843_), .C(new_n7667_), .Y(new_n9762_));
  NOR3X1   g07326(.A(new_n8284_), .B(new_n5939_), .C(pi0047), .Y(new_n9763_));
  OAI21X1  g07327(.A0(new_n9561_), .A1(pi0110), .B0(new_n9763_), .Y(new_n9764_));
  OR4X1    g07328(.A(new_n9764_), .B(new_n2566_), .C(pi0091), .D(pi0058), .Y(new_n9765_));
  INVX1    g07329(.A(new_n5970_), .Y(new_n9766_));
  INVX1    g07330(.A(new_n7607_), .Y(new_n9767_));
  NAND2X1  g07331(.A(new_n9562_), .B(po1057), .Y(new_n9768_));
  NAND3X1  g07332(.A(new_n9768_), .B(new_n9767_), .C(new_n9766_), .Y(new_n9769_));
  AOI21X1  g07333(.A0(new_n9765_), .A1(new_n5094_), .B0(new_n9769_), .Y(new_n9770_));
  NOR3X1   g07334(.A(new_n9765_), .B(new_n7607_), .C(new_n9766_), .Y(new_n9771_));
  OAI21X1  g07335(.A0(new_n9771_), .A1(new_n9770_), .B0(new_n6633_), .Y(new_n9772_));
  AOI21X1  g07336(.A0(new_n9772_), .A1(new_n9762_), .B0(new_n7749_), .Y(po0262));
  NOR3X1   g07337(.A(new_n8443_), .B(new_n8438_), .C(new_n5787_), .Y(new_n9774_));
  NAND2X1  g07338(.A(new_n8443_), .B(new_n2493_), .Y(new_n9775_));
  NAND2X1  g07339(.A(new_n9775_), .B(new_n2500_), .Y(new_n9776_));
  NOR3X1   g07340(.A(new_n9776_), .B(new_n2506_), .C(pi0024), .Y(new_n9777_));
  OAI21X1  g07341(.A0(new_n9777_), .A1(new_n9774_), .B0(pi0841), .Y(new_n9778_));
  NAND3X1  g07342(.A(new_n8430_), .B(new_n2726_), .C(new_n5787_), .Y(new_n9779_));
  AOI21X1  g07343(.A0(new_n9779_), .A1(new_n9778_), .B0(new_n7670_), .Y(po0264));
  NOR3X1   g07344(.A(new_n8490_), .B(new_n7670_), .C(pi0999), .Y(po0265));
  AND2X1   g07345(.A(new_n2583_), .B(pi0108), .Y(new_n9782_));
  AOI21X1  g07346(.A0(new_n5905_), .A1(new_n2880_), .B0(pi0108), .Y(new_n9783_));
  OR4X1    g07347(.A(new_n9783_), .B(new_n9782_), .C(new_n2504_), .D(new_n7842_), .Y(new_n9784_));
  OAI21X1  g07348(.A0(new_n5906_), .A1(new_n2506_), .B0(pi0314), .Y(new_n9785_));
  NOR3X1   g07349(.A(new_n7736_), .B(new_n5908_), .C(pi0070), .Y(new_n9786_));
  NAND2X1  g07350(.A(new_n9786_), .B(new_n9785_), .Y(new_n9787_));
  AOI21X1  g07351(.A0(new_n9784_), .A1(new_n7734_), .B0(new_n9787_), .Y(new_n9788_));
  NAND4X1  g07352(.A(new_n7735_), .B(new_n5907_), .C(pi0252), .D(new_n5134_), .Y(new_n9789_));
  OAI21X1  g07353(.A0(new_n9789_), .A1(new_n9784_), .B0(new_n2516_), .Y(new_n9790_));
  NOR3X1   g07354(.A(new_n5911_), .B(new_n3157_), .C(new_n2869_), .Y(new_n9791_));
  OAI21X1  g07355(.A0(new_n9790_), .A1(new_n9788_), .B0(new_n9791_), .Y(new_n9792_));
  NAND3X1  g07356(.A(new_n6756_), .B(new_n5104_), .C(new_n3095_), .Y(new_n9793_));
  AOI21X1  g07357(.A0(new_n9792_), .A1(new_n3156_), .B0(new_n9793_), .Y(po0266));
  OR4X1    g07358(.A(new_n8489_), .B(new_n2586_), .C(new_n2581_), .D(pi0050), .Y(new_n9795_));
  NOR3X1   g07359(.A(new_n9795_), .B(new_n7670_), .C(new_n7734_), .Y(po0267));
  NAND4X1  g07360(.A(new_n9560_), .B(pi0111), .C(new_n2481_), .D(new_n2648_), .Y(new_n9797_));
  OR2X1    g07361(.A(new_n9797_), .B(new_n2478_), .Y(new_n9798_));
  NOR4X1   g07362(.A(new_n9798_), .B(new_n8326_), .C(new_n2647_), .D(pi0068), .Y(new_n9799_));
  NOR3X1   g07363(.A(new_n7609_), .B(new_n5970_), .C(new_n5094_), .Y(new_n9800_));
  AOI22X1  g07364(.A0(new_n9800_), .A1(new_n7843_), .B0(new_n9799_), .B1(pi0314), .Y(new_n9801_));
  NOR2X1   g07365(.A(new_n9801_), .B(new_n7670_), .Y(po0268));
  AND2X1   g07366(.A(new_n9799_), .B(new_n7734_), .Y(new_n9803_));
  AOI22X1  g07367(.A0(new_n9803_), .A1(new_n6972_), .B0(new_n7774_), .B1(pi0072), .Y(new_n9804_));
  NOR3X1   g07368(.A(new_n9804_), .B(new_n7749_), .C(new_n7666_), .Y(po0269));
  NAND2X1  g07369(.A(new_n5860_), .B(pi0124), .Y(po0270));
  INVX1    g07370(.A(pi0113), .Y(new_n9807_));
  NOR3X1   g07371(.A(new_n9807_), .B(pi0072), .C(pi0039), .Y(new_n9808_));
  OAI21X1  g07372(.A0(new_n7823_), .A1(new_n2723_), .B0(new_n7770_), .Y(new_n9809_));
  NOR2X1   g07373(.A(new_n9809_), .B(new_n7820_), .Y(new_n9810_));
  OAI21X1  g07374(.A0(new_n7902_), .A1(new_n2548_), .B0(pi0113), .Y(new_n9811_));
  NOR2X1   g07375(.A(new_n9811_), .B(new_n9810_), .Y(new_n9812_));
  OAI21X1  g07376(.A0(new_n8085_), .A1(pi0113), .B0(pi0228), .Y(new_n9813_));
  NAND2X1  g07377(.A(new_n7929_), .B(pi0113), .Y(new_n9814_));
  AOI21X1  g07378(.A0(new_n9662_), .A1(new_n9807_), .B0(pi0228), .Y(new_n9815_));
  AOI21X1  g07379(.A0(new_n9815_), .A1(new_n9814_), .B0(pi0039), .Y(new_n9816_));
  OAI21X1  g07380(.A0(new_n9813_), .A1(new_n9812_), .B0(new_n9816_), .Y(new_n9817_));
  AND2X1   g07381(.A(pi0113), .B(new_n2548_), .Y(new_n9818_));
  INVX1    g07382(.A(new_n9818_), .Y(new_n9819_));
  AND2X1   g07383(.A(new_n6291_), .B(new_n2723_), .Y(new_n9820_));
  INVX1    g07384(.A(new_n9820_), .Y(new_n9821_));
  OR4X1    g07385(.A(new_n7869_), .B(new_n5972_), .C(new_n7903_), .D(pi0101), .Y(new_n9822_));
  AOI21X1  g07386(.A0(new_n9822_), .A1(new_n5093_), .B0(new_n9821_), .Y(new_n9823_));
  OR2X1    g07387(.A(new_n9823_), .B(new_n9819_), .Y(new_n9824_));
  NAND3X1  g07388(.A(new_n6291_), .B(new_n5093_), .C(new_n2723_), .Y(new_n9825_));
  OR4X1    g07389(.A(new_n9825_), .B(new_n7767_), .C(new_n7903_), .D(pi0113), .Y(new_n9826_));
  AOI21X1  g07390(.A0(new_n9826_), .A1(new_n9824_), .B0(pi0039), .Y(new_n9827_));
  OAI22X1  g07391(.A0(new_n9827_), .A1(new_n5086_), .B0(new_n9808_), .B1(new_n2996_), .Y(new_n9828_));
  AOI21X1  g07392(.A0(new_n9817_), .A1(new_n3277_), .B0(new_n9828_), .Y(new_n9829_));
  NOR3X1   g07393(.A(new_n7869_), .B(new_n5090_), .C(new_n3013_), .Y(new_n9830_));
  NOR2X1   g07394(.A(new_n9819_), .B(new_n9830_), .Y(new_n9831_));
  AOI21X1  g07395(.A0(new_n9678_), .A1(new_n9807_), .B0(new_n9831_), .Y(new_n9832_));
  AOI21X1  g07396(.A0(new_n9808_), .A1(new_n5792_), .B0(new_n3156_), .Y(new_n9833_));
  OAI21X1  g07397(.A0(new_n9832_), .A1(new_n3138_), .B0(new_n9833_), .Y(new_n9834_));
  OAI21X1  g07398(.A0(new_n9829_), .A1(pi0087), .B0(new_n9834_), .Y(new_n9835_));
  OR4X1    g07399(.A(new_n7775_), .B(new_n7903_), .C(pi0101), .D(pi0044), .Y(new_n9836_));
  AOI21X1  g07400(.A0(new_n9836_), .A1(new_n5093_), .B0(new_n9821_), .Y(new_n9837_));
  OAI22X1  g07401(.A0(new_n9837_), .A1(new_n9819_), .B0(new_n9826_), .B1(new_n7764_), .Y(new_n9838_));
  NAND2X1  g07402(.A(new_n9838_), .B(new_n3091_), .Y(new_n9839_));
  AOI21X1  g07403(.A0(new_n9808_), .A1(new_n5788_), .B0(new_n3095_), .Y(new_n9840_));
  AOI22X1  g07404(.A0(new_n9840_), .A1(new_n9839_), .B0(new_n9835_), .B1(new_n3095_), .Y(new_n9841_));
  MX2X1    g07405(.A(new_n9841_), .B(new_n9808_), .S0(new_n8306_), .Y(po0271));
  NOR3X1   g07406(.A(new_n7907_), .B(pi0072), .C(pi0039), .Y(new_n9843_));
  OAI21X1  g07407(.A0(new_n8120_), .A1(new_n7907_), .B0(new_n8367_), .Y(new_n9844_));
  AND2X1   g07408(.A(pi0114), .B(new_n2548_), .Y(new_n9845_));
  INVX1    g07409(.A(new_n9845_), .Y(new_n9846_));
  AOI21X1  g07410(.A0(new_n9846_), .A1(new_n8368_), .B0(new_n3092_), .Y(new_n9847_));
  OAI21X1  g07411(.A0(new_n9844_), .A1(new_n7995_), .B0(new_n9847_), .Y(new_n9848_));
  AOI21X1  g07412(.A0(new_n9843_), .A1(new_n5788_), .B0(new_n3095_), .Y(new_n9849_));
  MX2X1    g07413(.A(new_n8088_), .B(new_n8079_), .S0(pi0114), .Y(new_n9850_));
  OAI21X1  g07414(.A0(new_n9845_), .A1(new_n7898_), .B0(new_n2959_), .Y(new_n9851_));
  AOI21X1  g07415(.A0(new_n9850_), .A1(new_n7898_), .B0(new_n9851_), .Y(new_n9852_));
  NOR3X1   g07416(.A(new_n7964_), .B(new_n7962_), .C(pi0114), .Y(new_n9853_));
  OAI21X1  g07417(.A0(new_n7968_), .A1(new_n7907_), .B0(new_n8367_), .Y(new_n9854_));
  AOI21X1  g07418(.A0(new_n9846_), .A1(new_n8368_), .B0(pi0039), .Y(new_n9855_));
  OAI21X1  g07419(.A0(new_n9854_), .A1(new_n9853_), .B0(new_n9855_), .Y(new_n9856_));
  OAI21X1  g07420(.A0(new_n9843_), .A1(new_n2996_), .B0(new_n3156_), .Y(new_n9857_));
  AOI21X1  g07421(.A0(new_n9856_), .A1(new_n5085_), .B0(new_n9857_), .Y(new_n9858_));
  OAI21X1  g07422(.A0(new_n9852_), .A1(new_n5792_), .B0(new_n9858_), .Y(new_n9859_));
  NOR4X1   g07423(.A(new_n7869_), .B(new_n7909_), .C(new_n5090_), .D(new_n3013_), .Y(new_n9860_));
  AOI21X1  g07424(.A0(new_n9860_), .A1(new_n7898_), .B0(new_n9846_), .Y(new_n9861_));
  OR4X1    g07425(.A(new_n9861_), .B(new_n7985_), .C(pi0100), .D(pi0038), .Y(new_n9862_));
  NOR2X1   g07426(.A(new_n9843_), .B(new_n3277_), .Y(new_n9863_));
  NOR2X1   g07427(.A(new_n9863_), .B(new_n8340_), .Y(new_n9864_));
  AOI21X1  g07428(.A0(new_n9864_), .A1(new_n9862_), .B0(pi0075), .Y(new_n9865_));
  AOI22X1  g07429(.A0(new_n9865_), .A1(new_n9859_), .B0(new_n9849_), .B1(new_n9848_), .Y(new_n9866_));
  MX2X1    g07430(.A(new_n9866_), .B(new_n9843_), .S0(new_n8306_), .Y(po0272));
  NOR3X1   g07431(.A(new_n7898_), .B(pi0072), .C(pi0039), .Y(new_n9868_));
  NOR4X1   g07432(.A(pi0114), .B(pi0052), .C(pi0043), .D(pi0042), .Y(new_n9869_));
  NOR4X1   g07433(.A(new_n9869_), .B(new_n7964_), .C(new_n7764_), .D(pi0115), .Y(new_n9870_));
  OAI21X1  g07434(.A0(new_n8120_), .A1(new_n7898_), .B0(new_n9820_), .Y(new_n9871_));
  OR2X1    g07435(.A(new_n7898_), .B(pi0072), .Y(new_n9872_));
  AOI21X1  g07436(.A0(new_n9872_), .A1(new_n9821_), .B0(new_n3092_), .Y(new_n9873_));
  OAI21X1  g07437(.A0(new_n9871_), .A1(new_n9870_), .B0(new_n9873_), .Y(new_n9874_));
  AOI21X1  g07438(.A0(new_n9868_), .A1(new_n5788_), .B0(new_n3095_), .Y(new_n9875_));
  OAI21X1  g07439(.A0(new_n8087_), .A1(pi0115), .B0(new_n2959_), .Y(new_n9876_));
  AOI21X1  g07440(.A0(new_n8079_), .A1(pi0115), .B0(new_n9876_), .Y(new_n9877_));
  NOR3X1   g07441(.A(new_n9869_), .B(new_n7964_), .C(pi0115), .Y(new_n9878_));
  OAI21X1  g07442(.A0(new_n7968_), .A1(new_n7898_), .B0(new_n9820_), .Y(new_n9879_));
  AOI21X1  g07443(.A0(new_n9872_), .A1(new_n9821_), .B0(pi0039), .Y(new_n9880_));
  OAI21X1  g07444(.A0(new_n9879_), .A1(new_n9878_), .B0(new_n9880_), .Y(new_n9881_));
  OAI21X1  g07445(.A0(new_n9868_), .A1(new_n2996_), .B0(new_n3156_), .Y(new_n9882_));
  AOI21X1  g07446(.A0(new_n9881_), .A1(new_n5085_), .B0(new_n9882_), .Y(new_n9883_));
  OAI21X1  g07447(.A0(new_n9877_), .A1(new_n5792_), .B0(new_n9883_), .Y(new_n9884_));
  OAI21X1  g07448(.A0(new_n9872_), .A1(new_n9860_), .B0(new_n3277_), .Y(new_n9885_));
  NOR2X1   g07449(.A(new_n9868_), .B(new_n3277_), .Y(new_n9886_));
  NOR2X1   g07450(.A(new_n9886_), .B(new_n8340_), .Y(new_n9887_));
  OAI21X1  g07451(.A0(new_n9885_), .A1(new_n7984_), .B0(new_n9887_), .Y(new_n9888_));
  AND2X1   g07452(.A(new_n9888_), .B(new_n3095_), .Y(new_n9889_));
  AOI22X1  g07453(.A0(new_n9889_), .A1(new_n9884_), .B0(new_n9875_), .B1(new_n9874_), .Y(new_n9890_));
  MX2X1    g07454(.A(new_n9890_), .B(new_n9868_), .S0(new_n8306_), .Y(po0273));
  AND2X1   g07455(.A(pi0116), .B(new_n2548_), .Y(new_n9892_));
  AND2X1   g07456(.A(new_n9892_), .B(new_n2959_), .Y(new_n9893_));
  AND2X1   g07457(.A(new_n7919_), .B(pi0116), .Y(new_n9894_));
  OR2X1    g07458(.A(new_n9894_), .B(new_n2723_), .Y(new_n9895_));
  OAI21X1  g07459(.A0(new_n7905_), .A1(new_n2724_), .B0(pi0116), .Y(new_n9896_));
  NAND2X1  g07460(.A(new_n9896_), .B(new_n7911_), .Y(new_n9897_));
  OAI21X1  g07461(.A0(new_n8347_), .A1(new_n2723_), .B0(pi0228), .Y(new_n9898_));
  AOI21X1  g07462(.A0(new_n9897_), .A1(new_n9895_), .B0(new_n9898_), .Y(new_n9899_));
  OR2X1    g07463(.A(new_n7932_), .B(pi0228), .Y(new_n9900_));
  AOI21X1  g07464(.A0(new_n7930_), .A1(pi0116), .B0(new_n9900_), .Y(new_n9901_));
  NOR3X1   g07465(.A(new_n9901_), .B(new_n9899_), .C(pi0039), .Y(new_n9902_));
  INVX1    g07466(.A(new_n9892_), .Y(new_n9903_));
  AOI21X1  g07467(.A0(new_n6291_), .A1(new_n2723_), .B0(new_n9903_), .Y(new_n9904_));
  OAI21X1  g07468(.A0(new_n9822_), .A1(pi0113), .B0(new_n9892_), .Y(new_n9905_));
  AOI21X1  g07469(.A0(new_n9905_), .A1(new_n7964_), .B0(new_n9825_), .Y(new_n9906_));
  OAI21X1  g07470(.A0(new_n9906_), .A1(new_n9904_), .B0(new_n2959_), .Y(new_n9907_));
  AOI21X1  g07471(.A0(new_n9892_), .A1(new_n2959_), .B0(new_n2996_), .Y(new_n9908_));
  OR2X1    g07472(.A(new_n9908_), .B(pi0087), .Y(new_n9909_));
  AOI21X1  g07473(.A0(new_n9907_), .A1(new_n5085_), .B0(new_n9909_), .Y(new_n9910_));
  OAI21X1  g07474(.A0(new_n9902_), .A1(new_n5792_), .B0(new_n9910_), .Y(new_n9911_));
  AOI21X1  g07475(.A0(new_n9830_), .A1(new_n9807_), .B0(new_n9903_), .Y(new_n9912_));
  NOR3X1   g07476(.A(new_n9912_), .B(new_n7983_), .C(pi0038), .Y(new_n9913_));
  OAI21X1  g07477(.A0(new_n9913_), .A1(new_n9908_), .B0(new_n3026_), .Y(new_n9914_));
  AOI21X1  g07478(.A0(new_n9892_), .A1(new_n2959_), .B0(new_n3026_), .Y(new_n9915_));
  NOR2X1   g07479(.A(new_n9915_), .B(new_n8340_), .Y(new_n9916_));
  AOI21X1  g07480(.A0(new_n9916_), .A1(new_n9914_), .B0(pi0075), .Y(new_n9917_));
  AOI22X1  g07481(.A0(new_n9892_), .A1(new_n7996_), .B0(new_n7963_), .B1(new_n5932_), .Y(new_n9918_));
  OAI22X1  g07482(.A0(new_n9918_), .A1(new_n9825_), .B0(new_n9903_), .B1(new_n9820_), .Y(new_n9919_));
  NAND2X1  g07483(.A(new_n9919_), .B(new_n3091_), .Y(new_n9920_));
  AOI21X1  g07484(.A0(new_n9893_), .A1(new_n5788_), .B0(new_n3095_), .Y(new_n9921_));
  AOI22X1  g07485(.A0(new_n9921_), .A1(new_n9920_), .B0(new_n9917_), .B1(new_n9911_), .Y(new_n9922_));
  MX2X1    g07486(.A(new_n9922_), .B(new_n9893_), .S0(new_n8306_), .Y(po0274));
  OAI22X1  g07487(.A0(new_n5832_), .A1(new_n3408_), .B0(new_n3407_), .B1(pi0100), .Y(new_n9924_));
  AOI21X1  g07488(.A0(new_n9924_), .A1(new_n2996_), .B0(pi0087), .Y(new_n9925_));
  OAI21X1  g07489(.A0(new_n9925_), .A1(new_n5106_), .B0(new_n3100_), .Y(new_n9926_));
  AND2X1   g07490(.A(new_n5794_), .B(new_n3112_), .Y(new_n9927_));
  NAND3X1  g07491(.A(new_n9927_), .B(new_n9926_), .C(new_n4991_), .Y(new_n9928_));
  AOI21X1  g07492(.A0(new_n9928_), .A1(new_n3128_), .B0(new_n5822_), .Y(new_n9929_));
  OAI21X1  g07493(.A0(new_n9929_), .A1(pi0056), .B0(new_n4990_), .Y(new_n9930_));
  OR2X1    g07494(.A(new_n5113_), .B(pi0057), .Y(new_n9931_));
  AOI21X1  g07495(.A0(new_n9930_), .A1(new_n3245_), .B0(new_n9931_), .Y(po0275));
  INVX1    g07496(.A(new_n7369_), .Y(new_n9933_));
  NAND2X1  g07497(.A(new_n5033_), .B(pi0163), .Y(new_n9934_));
  AOI21X1  g07498(.A0(new_n9934_), .A1(new_n8707_), .B0(pi0150), .Y(new_n9935_));
  INVX1    g07499(.A(pi0150), .Y(new_n9936_));
  NOR4X1   g07500(.A(new_n8706_), .B(new_n7350_), .C(new_n5057_), .D(new_n9936_), .Y(new_n9937_));
  NOR2X1   g07501(.A(new_n9937_), .B(new_n9935_), .Y(new_n9938_));
  NOR2X1   g07502(.A(new_n9938_), .B(new_n5237_), .Y(new_n9939_));
  AOI21X1  g07503(.A0(new_n9939_), .A1(new_n6832_), .B0(new_n4991_), .Y(new_n9940_));
  INVX1    g07504(.A(pi0165), .Y(new_n9941_));
  OAI22X1  g07505(.A0(new_n6855_), .A1(new_n9941_), .B0(pi0054), .B1(pi0038), .Y(new_n9942_));
  OR2X1    g07506(.A(new_n9942_), .B(new_n6832_), .Y(new_n9943_));
  AOI21X1  g07507(.A0(new_n9939_), .A1(new_n6832_), .B0(pi0074), .Y(new_n9944_));
  AOI21X1  g07508(.A0(new_n9944_), .A1(new_n9943_), .B0(new_n9940_), .Y(new_n9945_));
  OAI21X1  g07509(.A0(new_n9945_), .A1(new_n3148_), .B0(new_n3246_), .Y(new_n9946_));
  AND2X1   g07510(.A(new_n9946_), .B(new_n9933_), .Y(new_n9947_));
  NOR3X1   g07511(.A(new_n9937_), .B(new_n9935_), .C(new_n2953_), .Y(new_n9948_));
  OR2X1    g07512(.A(new_n8718_), .B(pi0184), .Y(new_n9949_));
  OAI21X1  g07513(.A0(new_n9949_), .A1(pi0185), .B0(new_n5033_), .Y(new_n9950_));
  AOI21X1  g07514(.A0(new_n9949_), .A1(pi0185), .B0(new_n9950_), .Y(new_n9951_));
  OAI21X1  g07515(.A0(new_n9951_), .A1(pi0299), .B0(pi0232), .Y(new_n9952_));
  NOR3X1   g07516(.A(new_n9952_), .B(new_n9948_), .C(new_n6828_), .Y(new_n9953_));
  OR2X1    g07517(.A(new_n9953_), .B(new_n4991_), .Y(new_n9954_));
  AND2X1   g07518(.A(new_n9954_), .B(new_n3128_), .Y(new_n9955_));
  MX2X1    g07519(.A(pi0143), .B(pi0165), .S0(pi0299), .Y(new_n9956_));
  AND2X1   g07520(.A(new_n9956_), .B(new_n5930_), .Y(new_n9957_));
  OAI21X1  g07521(.A0(new_n9957_), .A1(new_n6832_), .B0(pi0054), .Y(new_n9958_));
  NOR2X1   g07522(.A(new_n9958_), .B(new_n9953_), .Y(new_n9959_));
  INVX1    g07523(.A(pi0143), .Y(new_n9960_));
  OAI21X1  g07524(.A0(new_n7490_), .A1(new_n9960_), .B0(pi0165), .Y(new_n9961_));
  AOI21X1  g07525(.A0(new_n7489_), .A1(new_n9960_), .B0(new_n9961_), .Y(new_n9962_));
  NAND3X1  g07526(.A(new_n7486_), .B(new_n9941_), .C(pi0143), .Y(new_n9963_));
  NAND2X1  g07527(.A(new_n9963_), .B(pi0038), .Y(new_n9964_));
  OAI21X1  g07528(.A0(new_n9964_), .A1(new_n9962_), .B0(new_n3123_), .Y(new_n9965_));
  INVX1    g07529(.A(new_n7078_), .Y(new_n9966_));
  OR2X1    g07530(.A(pi0168), .B(new_n3325_), .Y(new_n9967_));
  NOR2X1   g07531(.A(new_n9967_), .B(new_n7136_), .Y(new_n9968_));
  AND2X1   g07532(.A(new_n7133_), .B(new_n4351_), .Y(new_n9969_));
  OR2X1    g07533(.A(new_n9969_), .B(pi0151), .Y(new_n9970_));
  AOI21X1  g07534(.A0(new_n7130_), .A1(pi0168), .B0(new_n9970_), .Y(new_n9971_));
  OAI22X1  g07535(.A0(new_n9971_), .A1(new_n9968_), .B0(new_n9966_), .B1(new_n5033_), .Y(new_n9972_));
  NOR2X1   g07536(.A(new_n7078_), .B(new_n5033_), .Y(new_n9973_));
  INVX1    g07537(.A(new_n9973_), .Y(new_n9974_));
  OAI21X1  g07538(.A0(new_n7114_), .A1(new_n5057_), .B0(new_n9974_), .Y(new_n9975_));
  AND2X1   g07539(.A(pi0168), .B(pi0151), .Y(new_n9976_));
  AOI21X1  g07540(.A0(new_n9976_), .A1(new_n9975_), .B0(new_n9936_), .Y(new_n9977_));
  NAND3X1  g07541(.A(new_n9974_), .B(new_n7017_), .C(pi0168), .Y(new_n9978_));
  NOR3X1   g07542(.A(new_n9973_), .B(new_n7161_), .C(pi0168), .Y(new_n9979_));
  NOR2X1   g07543(.A(new_n9979_), .B(new_n3325_), .Y(new_n9980_));
  AND2X1   g07544(.A(new_n5033_), .B(pi0168), .Y(new_n9981_));
  INVX1    g07545(.A(new_n9981_), .Y(new_n9982_));
  AND2X1   g07546(.A(new_n9982_), .B(new_n7078_), .Y(new_n9983_));
  OAI21X1  g07547(.A0(new_n7399_), .A1(new_n4351_), .B0(new_n3325_), .Y(new_n9984_));
  OAI21X1  g07548(.A0(new_n9984_), .A1(new_n9983_), .B0(new_n9936_), .Y(new_n9985_));
  AOI21X1  g07549(.A0(new_n9980_), .A1(new_n9978_), .B0(new_n9985_), .Y(new_n9986_));
  OR2X1    g07550(.A(new_n9986_), .B(new_n2953_), .Y(new_n9987_));
  AOI21X1  g07551(.A0(new_n9977_), .A1(new_n9972_), .B0(new_n9987_), .Y(new_n9988_));
  INVX1    g07552(.A(pi0173), .Y(new_n9989_));
  AND2X1   g07553(.A(new_n7078_), .B(new_n5057_), .Y(new_n9990_));
  OAI21X1  g07554(.A0(new_n9990_), .A1(new_n7055_), .B0(new_n9989_), .Y(new_n9991_));
  NOR2X1   g07555(.A(new_n9973_), .B(new_n9989_), .Y(new_n9992_));
  OAI21X1  g07556(.A0(new_n6978_), .A1(new_n5057_), .B0(new_n9992_), .Y(new_n9993_));
  AND2X1   g07557(.A(new_n9993_), .B(pi0185), .Y(new_n9994_));
  NOR3X1   g07558(.A(new_n9973_), .B(new_n7018_), .C(new_n9989_), .Y(new_n9995_));
  INVX1    g07559(.A(pi0185), .Y(new_n9996_));
  AOI21X1  g07560(.A0(new_n7078_), .A1(new_n5057_), .B0(new_n7061_), .Y(new_n9997_));
  OAI21X1  g07561(.A0(new_n9997_), .A1(pi0173), .B0(new_n9996_), .Y(new_n9998_));
  OAI21X1  g07562(.A0(new_n9998_), .A1(new_n9995_), .B0(pi0190), .Y(new_n9999_));
  AOI21X1  g07563(.A0(new_n9994_), .A1(new_n9991_), .B0(new_n9999_), .Y(new_n10000_));
  AOI21X1  g07564(.A0(new_n7075_), .A1(new_n9989_), .B0(new_n5057_), .Y(new_n10001_));
  OAI21X1  g07565(.A0(new_n7419_), .A1(new_n9989_), .B0(new_n10001_), .Y(new_n10002_));
  AOI21X1  g07566(.A0(new_n7078_), .A1(new_n5057_), .B0(new_n9996_), .Y(new_n10003_));
  INVX1    g07567(.A(pi0190), .Y(new_n10004_));
  NOR3X1   g07568(.A(new_n9973_), .B(new_n7161_), .C(new_n9989_), .Y(new_n10005_));
  OAI21X1  g07569(.A0(new_n9966_), .A1(pi0173), .B0(new_n9996_), .Y(new_n10006_));
  OAI21X1  g07570(.A0(new_n10006_), .A1(new_n10005_), .B0(new_n10004_), .Y(new_n10007_));
  AOI21X1  g07571(.A0(new_n10003_), .A1(new_n10002_), .B0(new_n10007_), .Y(new_n10008_));
  OR2X1    g07572(.A(new_n10008_), .B(pi0299), .Y(new_n10009_));
  OAI21X1  g07573(.A0(new_n10009_), .A1(new_n10000_), .B0(pi0232), .Y(new_n10010_));
  AOI21X1  g07574(.A0(new_n7078_), .A1(new_n5237_), .B0(pi0039), .Y(new_n10011_));
  OAI21X1  g07575(.A0(new_n10010_), .A1(new_n9988_), .B0(new_n10011_), .Y(new_n10012_));
  AOI22X1  g07576(.A0(new_n6901_), .A1(pi0157), .B0(new_n6907_), .B1(pi0168), .Y(new_n10013_));
  NOR4X1   g07577(.A(new_n10013_), .B(new_n6905_), .C(new_n5070_), .D(new_n5057_), .Y(new_n10014_));
  MX2X1    g07578(.A(new_n10014_), .B(pi0178), .S0(new_n2953_), .Y(new_n10015_));
  AOI21X1  g07579(.A0(new_n7465_), .A1(pi0178), .B0(pi0190), .Y(new_n10016_));
  OAI22X1  g07580(.A0(new_n10016_), .A1(pi0299), .B0(new_n10015_), .B1(new_n6870_), .Y(new_n10017_));
  OAI21X1  g07581(.A0(new_n6869_), .A1(new_n5051_), .B0(new_n6886_), .Y(new_n10018_));
  NOR3X1   g07582(.A(new_n10018_), .B(new_n6890_), .C(pi0178), .Y(new_n10019_));
  INVX1    g07583(.A(pi0178), .Y(new_n10020_));
  NOR3X1   g07584(.A(new_n10018_), .B(new_n6923_), .C(new_n10020_), .Y(new_n10021_));
  OAI21X1  g07585(.A0(new_n6886_), .A1(new_n6870_), .B0(new_n2953_), .Y(new_n10022_));
  OR4X1    g07586(.A(new_n10022_), .B(new_n10021_), .C(new_n10019_), .D(new_n10004_), .Y(new_n10023_));
  NAND3X1  g07587(.A(new_n10023_), .B(new_n10017_), .C(pi0232), .Y(new_n10024_));
  AOI21X1  g07588(.A0(new_n6869_), .A1(new_n5237_), .B0(new_n2959_), .Y(new_n10025_));
  AOI21X1  g07589(.A0(new_n10025_), .A1(new_n10024_), .B0(pi0038), .Y(new_n10026_));
  AOI21X1  g07590(.A0(new_n10026_), .A1(new_n10012_), .B0(new_n9965_), .Y(new_n10027_));
  OAI21X1  g07591(.A0(new_n9952_), .A1(new_n9948_), .B0(pi0100), .Y(new_n10028_));
  OAI21X1  g07592(.A0(new_n9957_), .A1(new_n2996_), .B0(new_n7329_), .Y(new_n10029_));
  OAI21X1  g07593(.A0(new_n10029_), .A1(new_n7229_), .B0(new_n10028_), .Y(new_n10030_));
  OAI21X1  g07594(.A0(new_n10030_), .A1(new_n10027_), .B0(new_n3105_), .Y(new_n10031_));
  OR2X1    g07595(.A(new_n9952_), .B(new_n9948_), .Y(new_n10032_));
  AND2X1   g07596(.A(new_n10032_), .B(pi0075), .Y(new_n10033_));
  OAI21X1  g07597(.A0(new_n9957_), .A1(new_n2996_), .B0(new_n3026_), .Y(new_n10034_));
  MX2X1    g07598(.A(pi0178), .B(pi0157), .S0(pi0299), .Y(new_n10035_));
  AND2X1   g07599(.A(new_n10035_), .B(new_n5930_), .Y(new_n10036_));
  AOI21X1  g07600(.A0(new_n10036_), .A1(new_n7502_), .B0(new_n7230_), .Y(new_n10037_));
  OAI21X1  g07601(.A0(new_n10037_), .A1(new_n10034_), .B0(new_n10028_), .Y(new_n10038_));
  AOI21X1  g07602(.A0(new_n10038_), .A1(new_n7185_), .B0(new_n10033_), .Y(new_n10039_));
  AOI21X1  g07603(.A0(new_n10039_), .A1(new_n10031_), .B0(pi0054), .Y(new_n10040_));
  OAI21X1  g07604(.A0(new_n10040_), .A1(new_n9959_), .B0(new_n4991_), .Y(new_n10041_));
  OR2X1    g07605(.A(new_n9940_), .B(new_n3128_), .Y(new_n10042_));
  INVX1    g07606(.A(new_n9944_), .Y(new_n10043_));
  NOR4X1   g07607(.A(pi0468), .B(pi0332), .C(new_n5237_), .D(new_n9936_), .Y(new_n10044_));
  NOR4X1   g07608(.A(new_n6878_), .B(new_n7188_), .C(pi0095), .D(pi0092), .Y(new_n10045_));
  AND2X1   g07609(.A(new_n10045_), .B(new_n10044_), .Y(new_n10046_));
  NAND3X1  g07610(.A(new_n6869_), .B(new_n3112_), .C(new_n2996_), .Y(new_n10047_));
  OAI21X1  g07611(.A0(new_n10047_), .A1(new_n10046_), .B0(new_n9942_), .Y(new_n10048_));
  AOI21X1  g07612(.A0(new_n10048_), .A1(new_n6828_), .B0(new_n10043_), .Y(new_n10049_));
  OAI21X1  g07613(.A0(new_n10049_), .A1(new_n10042_), .B0(new_n3148_), .Y(new_n10050_));
  AOI21X1  g07614(.A0(new_n10041_), .A1(new_n9955_), .B0(new_n10050_), .Y(new_n10051_));
  NOR2X1   g07615(.A(new_n9939_), .B(new_n6828_), .Y(new_n10052_));
  NOR4X1   g07616(.A(new_n6832_), .B(new_n5057_), .C(new_n5237_), .D(new_n9941_), .Y(new_n10053_));
  OR4X1    g07617(.A(new_n10053_), .B(new_n10052_), .C(new_n9940_), .D(new_n3246_), .Y(new_n10054_));
  OAI21X1  g07618(.A0(new_n10051_), .A1(new_n9947_), .B0(new_n10054_), .Y(new_n10055_));
  NOR2X1   g07619(.A(new_n10055_), .B(new_n6817_), .Y(new_n10056_));
  NOR4X1   g07620(.A(pi0954), .B(pi0079), .C(pi0034), .D(pi0033), .Y(new_n10057_));
  INVX1    g07621(.A(new_n10057_), .Y(new_n10058_));
  OAI21X1  g07622(.A0(new_n5256_), .A1(new_n5249_), .B0(new_n6269_), .Y(new_n10059_));
  INVX1    g07623(.A(pi0157), .Y(new_n10060_));
  AOI21X1  g07624(.A0(new_n7241_), .A1(new_n10060_), .B0(new_n4351_), .Y(new_n10061_));
  OR2X1    g07625(.A(pi0168), .B(pi0157), .Y(new_n10062_));
  OAI22X1  g07626(.A0(new_n10062_), .A1(new_n7235_), .B0(new_n7237_), .B1(new_n10060_), .Y(new_n10063_));
  OAI21X1  g07627(.A0(new_n10063_), .A1(new_n10061_), .B0(new_n10059_), .Y(new_n10064_));
  INVX1    g07628(.A(new_n9592_), .Y(new_n10065_));
  AND2X1   g07629(.A(new_n7239_), .B(pi1091), .Y(new_n10066_));
  NAND4X1  g07630(.A(new_n10066_), .B(new_n5051_), .C(new_n5033_), .D(new_n10020_), .Y(new_n10067_));
  AOI21X1  g07631(.A0(new_n10067_), .A1(new_n10059_), .B0(new_n10004_), .Y(new_n10068_));
  NAND3X1  g07632(.A(new_n5261_), .B(new_n5051_), .C(new_n5033_), .Y(new_n10069_));
  NAND3X1  g07633(.A(new_n10059_), .B(new_n10069_), .C(pi0178), .Y(new_n10070_));
  OAI21X1  g07634(.A0(new_n5256_), .A1(new_n5249_), .B0(new_n8518_), .Y(new_n10071_));
  AOI21X1  g07635(.A0(new_n10071_), .A1(new_n10020_), .B0(pi0190), .Y(new_n10072_));
  AOI21X1  g07636(.A0(new_n10072_), .A1(new_n10070_), .B0(new_n10068_), .Y(new_n10073_));
  OAI21X1  g07637(.A0(new_n10073_), .A1(new_n10065_), .B0(pi0232), .Y(new_n10074_));
  AOI21X1  g07638(.A0(new_n10064_), .A1(new_n9591_), .B0(new_n10074_), .Y(new_n10075_));
  NOR3X1   g07639(.A(new_n6913_), .B(new_n5797_), .C(new_n5257_), .Y(new_n10076_));
  OAI21X1  g07640(.A0(new_n6906_), .A1(new_n6269_), .B0(new_n9591_), .Y(new_n10077_));
  OAI21X1  g07641(.A0(new_n10077_), .A1(new_n5257_), .B0(new_n5237_), .Y(new_n10078_));
  OAI21X1  g07642(.A0(new_n10078_), .A1(new_n10076_), .B0(pi0039), .Y(new_n10079_));
  NOR2X1   g07643(.A(new_n7282_), .B(new_n4351_), .Y(new_n10080_));
  OAI21X1  g07644(.A0(new_n7270_), .A1(pi0168), .B0(new_n3325_), .Y(new_n10081_));
  OAI22X1  g07645(.A0(new_n10081_), .A1(new_n10080_), .B0(new_n9967_), .B1(new_n7291_), .Y(new_n10082_));
  AOI21X1  g07646(.A0(new_n10082_), .A1(new_n7273_), .B0(new_n9936_), .Y(new_n10083_));
  OAI21X1  g07647(.A0(new_n7262_), .A1(pi0151), .B0(new_n7535_), .Y(new_n10084_));
  AOI21X1  g07648(.A0(new_n7279_), .A1(new_n3325_), .B0(new_n8946_), .Y(new_n10085_));
  OAI21X1  g07649(.A0(new_n10085_), .A1(new_n9982_), .B0(new_n9936_), .Y(new_n10086_));
  AOI21X1  g07650(.A0(new_n10084_), .A1(new_n4351_), .B0(new_n10086_), .Y(new_n10087_));
  AOI21X1  g07651(.A0(new_n8943_), .A1(new_n7262_), .B0(new_n5033_), .Y(new_n10088_));
  NOR2X1   g07652(.A(new_n10088_), .B(new_n2953_), .Y(new_n10089_));
  OAI21X1  g07653(.A0(new_n10087_), .A1(new_n10083_), .B0(new_n10089_), .Y(new_n10090_));
  NOR2X1   g07654(.A(new_n7291_), .B(new_n7666_), .Y(new_n10091_));
  INVX1    g07655(.A(new_n10091_), .Y(new_n10092_));
  NAND4X1  g07656(.A(new_n7269_), .B(new_n7267_), .C(new_n5189_), .D(new_n9989_), .Y(new_n10093_));
  OAI21X1  g07657(.A0(new_n10092_), .A1(new_n9989_), .B0(new_n10093_), .Y(new_n10094_));
  NOR3X1   g07658(.A(pi0468), .B(pi0332), .C(pi0190), .Y(new_n10095_));
  NAND4X1  g07659(.A(new_n7282_), .B(new_n7273_), .C(pi0190), .D(new_n9989_), .Y(new_n10096_));
  NAND2X1  g07660(.A(new_n10096_), .B(pi0185), .Y(new_n10097_));
  AOI21X1  g07661(.A0(new_n10095_), .A1(new_n10094_), .B0(new_n10097_), .Y(new_n10098_));
  OAI21X1  g07662(.A0(new_n7262_), .A1(pi0173), .B0(new_n8966_), .Y(new_n10099_));
  NOR3X1   g07663(.A(new_n7288_), .B(new_n5220_), .C(new_n9989_), .Y(new_n10100_));
  NOR3X1   g07664(.A(new_n10100_), .B(new_n7280_), .C(new_n10004_), .Y(new_n10101_));
  OR2X1    g07665(.A(new_n10101_), .B(pi0185), .Y(new_n10102_));
  AOI21X1  g07666(.A0(new_n10099_), .A1(new_n10004_), .B0(new_n10102_), .Y(new_n10103_));
  AOI21X1  g07667(.A0(new_n7266_), .A1(new_n5057_), .B0(pi0299), .Y(new_n10104_));
  OAI21X1  g07668(.A0(new_n10103_), .A1(new_n10098_), .B0(new_n10104_), .Y(new_n10105_));
  AOI21X1  g07669(.A0(new_n10105_), .A1(new_n10090_), .B0(new_n5237_), .Y(new_n10106_));
  NOR2X1   g07670(.A(new_n7265_), .B(new_n5019_), .Y(new_n10107_));
  OR2X1    g07671(.A(new_n7261_), .B(pi0232), .Y(new_n10108_));
  OAI21X1  g07672(.A0(new_n10108_), .A1(new_n10107_), .B0(new_n2959_), .Y(new_n10109_));
  OAI22X1  g07673(.A0(new_n10109_), .A1(new_n10106_), .B0(new_n10079_), .B1(new_n10075_), .Y(new_n10110_));
  AOI21X1  g07674(.A0(new_n10110_), .A1(new_n2996_), .B0(new_n9965_), .Y(new_n10111_));
  NAND2X1  g07675(.A(new_n10029_), .B(new_n10028_), .Y(new_n10112_));
  OAI21X1  g07676(.A0(new_n10112_), .A1(new_n10111_), .B0(new_n3105_), .Y(new_n10113_));
  NOR4X1   g07677(.A(new_n10036_), .B(new_n3066_), .C(new_n3074_), .D(pi0087), .Y(new_n10114_));
  OAI21X1  g07678(.A0(new_n10114_), .A1(new_n10034_), .B0(new_n10028_), .Y(new_n10115_));
  AOI21X1  g07679(.A0(new_n10115_), .A1(new_n7185_), .B0(new_n10033_), .Y(new_n10116_));
  AOI21X1  g07680(.A0(new_n10116_), .A1(new_n10113_), .B0(pi0054), .Y(new_n10117_));
  OAI21X1  g07681(.A0(new_n10117_), .A1(new_n9959_), .B0(new_n4991_), .Y(new_n10118_));
  AND2X1   g07682(.A(new_n9944_), .B(new_n9943_), .Y(new_n10119_));
  NOR4X1   g07683(.A(new_n5057_), .B(new_n5237_), .C(new_n9941_), .D(new_n3112_), .Y(new_n10120_));
  NOR3X1   g07684(.A(pi0087), .B(pi0039), .C(pi0038), .Y(new_n10121_));
  NAND3X1  g07685(.A(new_n6828_), .B(new_n10121_), .C(new_n3100_), .Y(new_n10122_));
  OR4X1    g07686(.A(new_n10122_), .B(new_n10120_), .C(new_n10044_), .D(new_n3074_), .Y(new_n10123_));
  AOI21X1  g07687(.A0(new_n10123_), .A1(new_n10119_), .B0(new_n10042_), .Y(new_n10124_));
  OR2X1    g07688(.A(new_n10124_), .B(new_n5324_), .Y(new_n10125_));
  AOI21X1  g07689(.A0(new_n10118_), .A1(new_n9955_), .B0(new_n10125_), .Y(new_n10126_));
  OAI21X1  g07690(.A0(new_n10126_), .A1(new_n9946_), .B0(new_n10054_), .Y(new_n10127_));
  OAI21X1  g07691(.A0(new_n10127_), .A1(pi0118), .B0(new_n10058_), .Y(new_n10128_));
  NOR3X1   g07692(.A(new_n10055_), .B(new_n6818_), .C(pi0118), .Y(new_n10129_));
  NOR2X1   g07693(.A(new_n6818_), .B(pi0118), .Y(new_n10130_));
  OAI21X1  g07694(.A0(new_n10130_), .A1(new_n10127_), .B0(new_n10057_), .Y(new_n10131_));
  OAI22X1  g07695(.A0(new_n10131_), .A1(new_n10129_), .B0(new_n10128_), .B1(new_n10056_), .Y(po0276));
  NAND2X1  g07696(.A(pi0228), .B(pi0128), .Y(new_n10133_));
  INVX1    g07697(.A(pi0128), .Y(new_n10134_));
  NAND3X1  g07698(.A(new_n5962_), .B(new_n4780_), .C(new_n2971_), .Y(new_n10135_));
  NOR2X1   g07699(.A(pi0221), .B(pi0216), .Y(new_n10136_));
  INVX1    g07700(.A(new_n10136_), .Y(new_n10137_));
  NAND3X1  g07701(.A(new_n5960_), .B(new_n4898_), .C(new_n10137_), .Y(new_n10138_));
  AOI21X1  g07702(.A0(new_n10138_), .A1(new_n10135_), .B0(new_n2959_), .Y(new_n10139_));
  OR2X1    g07703(.A(new_n7662_), .B(new_n8560_), .Y(new_n10140_));
  AOI21X1  g07704(.A0(new_n10140_), .A1(new_n8698_), .B0(new_n2598_), .Y(new_n10141_));
  NOR4X1   g07705(.A(new_n5250_), .B(new_n2588_), .C(pi0108), .D(pi0046), .Y(new_n10142_));
  OAI21X1  g07706(.A0(new_n10141_), .A1(pi0097), .B0(new_n10142_), .Y(new_n10143_));
  MX2X1    g07707(.A(new_n5228_), .B(new_n5131_), .S0(pi0299), .Y(new_n10144_));
  NAND2X1  g07708(.A(new_n10144_), .B(new_n5930_), .Y(new_n10145_));
  AOI22X1  g07709(.A0(new_n10145_), .A1(pi0109), .B0(new_n8699_), .B1(new_n5250_), .Y(new_n10146_));
  MX2X1    g07710(.A(new_n5203_), .B(new_n5175_), .S0(new_n10145_), .Y(new_n10147_));
  AOI21X1  g07711(.A0(new_n10146_), .A1(new_n10143_), .B0(new_n10147_), .Y(new_n10148_));
  AOI21X1  g07712(.A0(new_n3255_), .A1(pi0091), .B0(new_n2744_), .Y(new_n10149_));
  OAI21X1  g07713(.A0(new_n10148_), .A1(pi0091), .B0(new_n10149_), .Y(new_n10150_));
  NAND4X1  g07714(.A(new_n3002_), .B(new_n2532_), .C(new_n2526_), .D(new_n2959_), .Y(new_n10151_));
  AOI21X1  g07715(.A0(new_n10150_), .A1(new_n2561_), .B0(new_n10151_), .Y(new_n10152_));
  OAI21X1  g07716(.A0(new_n10152_), .A1(new_n10139_), .B0(new_n2996_), .Y(new_n10153_));
  MX2X1    g07717(.A(new_n10153_), .B(new_n10134_), .S0(pi0228), .Y(new_n10154_));
  OAI21X1  g07718(.A0(new_n3632_), .A1(new_n3066_), .B0(new_n10133_), .Y(new_n10155_));
  AOI21X1  g07719(.A0(new_n10155_), .A1(pi0100), .B0(pi0087), .Y(new_n10156_));
  OAI21X1  g07720(.A0(new_n10154_), .A1(pi0100), .B0(new_n10156_), .Y(new_n10157_));
  AOI21X1  g07721(.A0(new_n10133_), .A1(pi0087), .B0(pi0075), .Y(new_n10158_));
  AOI22X1  g07722(.A0(new_n10121_), .A1(new_n5836_), .B0(pi0228), .B1(pi0128), .Y(new_n10159_));
  OAI21X1  g07723(.A0(new_n10159_), .A1(new_n3095_), .B0(new_n3100_), .Y(new_n10160_));
  AOI21X1  g07724(.A0(new_n10158_), .A1(new_n10157_), .B0(new_n10160_), .Y(new_n10161_));
  NAND2X1  g07725(.A(new_n10133_), .B(pi0092), .Y(new_n10162_));
  OAI21X1  g07726(.A0(new_n10162_), .A1(new_n5844_), .B0(new_n9572_), .Y(new_n10163_));
  OAI22X1  g07727(.A0(new_n10163_), .A1(new_n10161_), .B0(new_n10133_), .B1(new_n9572_), .Y(po0277));
  INVX1    g07728(.A(pi0818), .Y(new_n10165_));
  OR2X1    g07729(.A(pi0080), .B(pi0031), .Y(new_n10166_));
  NOR2X1   g07730(.A(new_n10166_), .B(new_n10165_), .Y(new_n10167_));
  INVX1    g07731(.A(new_n10167_), .Y(new_n10168_));
  AOI21X1  g07732(.A0(new_n9249_), .A1(new_n6309_), .B0(new_n6077_), .Y(new_n10169_));
  NOR2X1   g07733(.A(new_n5893_), .B(pi0120), .Y(new_n10170_));
  NAND2X1  g07734(.A(new_n10170_), .B(new_n2756_), .Y(new_n10171_));
  AND2X1   g07735(.A(new_n10171_), .B(new_n10169_), .Y(new_n10172_));
  AND2X1   g07736(.A(new_n5933_), .B(new_n3630_), .Y(new_n10173_));
  INVX1    g07737(.A(pi0120), .Y(new_n10174_));
  AOI21X1  g07738(.A0(new_n9239_), .A1(new_n2722_), .B0(new_n10174_), .Y(new_n10175_));
  INVX1    g07739(.A(new_n10175_), .Y(new_n10176_));
  OAI21X1  g07740(.A0(new_n10176_), .A1(new_n5975_), .B0(new_n10173_), .Y(new_n10177_));
  AND2X1   g07741(.A(pi1093), .B(new_n10174_), .Y(new_n10178_));
  OAI21X1  g07742(.A0(new_n10178_), .A1(new_n5976_), .B0(new_n10177_), .Y(new_n10179_));
  AND2X1   g07743(.A(new_n6291_), .B(new_n3065_), .Y(new_n10180_));
  NAND4X1  g07744(.A(new_n2783_), .B(new_n2722_), .C(pi0824), .D(new_n5952_), .Y(new_n10181_));
  AND2X1   g07745(.A(new_n10181_), .B(new_n10178_), .Y(new_n10182_));
  OAI21X1  g07746(.A0(new_n10182_), .A1(new_n10175_), .B0(pi0100), .Y(new_n10183_));
  AOI21X1  g07747(.A0(new_n10180_), .A1(new_n10179_), .B0(new_n10183_), .Y(new_n10184_));
  NAND3X1  g07748(.A(new_n5919_), .B(new_n5913_), .C(new_n2756_), .Y(new_n10185_));
  OAI21X1  g07749(.A0(new_n10185_), .A1(new_n10174_), .B0(new_n2959_), .Y(new_n10186_));
  NOR4X1   g07750(.A(new_n5939_), .B(new_n5911_), .C(new_n5910_), .D(pi0829), .Y(new_n10187_));
  OR2X1    g07751(.A(new_n10187_), .B(pi0122), .Y(new_n10188_));
  AOI21X1  g07752(.A0(new_n7805_), .A1(new_n5949_), .B0(new_n10188_), .Y(new_n10189_));
  OAI21X1  g07753(.A0(new_n5912_), .A1(new_n5952_), .B0(new_n8273_), .Y(new_n10190_));
  OAI21X1  g07754(.A0(new_n10190_), .A1(new_n10189_), .B0(new_n2781_), .Y(new_n10191_));
  NOR3X1   g07755(.A(new_n5939_), .B(new_n5911_), .C(new_n5910_), .Y(new_n10192_));
  OR4X1    g07756(.A(new_n10192_), .B(new_n9394_), .C(new_n2756_), .D(pi1091), .Y(new_n10193_));
  NAND2X1  g07757(.A(new_n10193_), .B(new_n10191_), .Y(new_n10194_));
  NOR2X1   g07758(.A(new_n10182_), .B(new_n10175_), .Y(new_n10195_));
  INVX1    g07759(.A(new_n10195_), .Y(new_n10196_));
  INVX1    g07760(.A(new_n10182_), .Y(new_n10197_));
  NOR3X1   g07761(.A(new_n5959_), .B(new_n2755_), .C(new_n2722_), .Y(new_n10198_));
  OAI22X1  g07762(.A0(new_n10198_), .A1(new_n10197_), .B0(new_n10176_), .B1(new_n10066_), .Y(new_n10199_));
  MX2X1    g07763(.A(new_n10199_), .B(new_n10196_), .S0(new_n6270_), .Y(new_n10200_));
  NAND2X1  g07764(.A(new_n10200_), .B(new_n5070_), .Y(new_n10201_));
  MX2X1    g07765(.A(new_n10199_), .B(new_n10196_), .S0(new_n5052_), .Y(new_n10202_));
  AOI21X1  g07766(.A0(new_n10202_), .A1(new_n5071_), .B0(new_n6284_), .Y(new_n10203_));
  OAI21X1  g07767(.A0(new_n10196_), .A1(new_n6283_), .B0(pi0299), .Y(new_n10204_));
  AOI21X1  g07768(.A0(new_n10203_), .A1(new_n10201_), .B0(new_n10204_), .Y(new_n10205_));
  NAND2X1  g07769(.A(new_n10200_), .B(new_n5050_), .Y(new_n10206_));
  AOI21X1  g07770(.A0(new_n10202_), .A1(new_n5051_), .B0(new_n6278_), .Y(new_n10207_));
  OAI21X1  g07771(.A0(new_n10196_), .A1(new_n6277_), .B0(new_n2953_), .Y(new_n10208_));
  AOI21X1  g07772(.A0(new_n10207_), .A1(new_n10206_), .B0(new_n10208_), .Y(new_n10209_));
  OR2X1    g07773(.A(new_n10209_), .B(new_n2959_), .Y(new_n10210_));
  OAI22X1  g07774(.A0(new_n10210_), .A1(new_n10205_), .B0(new_n10194_), .B1(new_n10186_), .Y(new_n10211_));
  INVX1    g07775(.A(new_n9249_), .Y(new_n10212_));
  NOR2X1   g07776(.A(pi1093), .B(pi0120), .Y(new_n10213_));
  AOI21X1  g07777(.A0(new_n10213_), .A1(pi0038), .B0(pi0100), .Y(new_n10214_));
  OAI21X1  g07778(.A0(new_n10212_), .A1(new_n2996_), .B0(new_n10214_), .Y(new_n10215_));
  AOI21X1  g07779(.A0(new_n10211_), .A1(new_n2996_), .B0(new_n10215_), .Y(new_n10216_));
  OAI21X1  g07780(.A0(new_n10216_), .A1(new_n10184_), .B0(new_n3156_), .Y(new_n10217_));
  INVX1    g07781(.A(new_n10213_), .Y(new_n10218_));
  NOR3X1   g07782(.A(new_n9394_), .B(new_n2756_), .C(pi1091), .Y(new_n10219_));
  INVX1    g07783(.A(new_n10219_), .Y(new_n10220_));
  OAI21X1  g07784(.A0(new_n10220_), .A1(new_n6301_), .B0(new_n5988_), .Y(new_n10221_));
  NAND4X1  g07785(.A(new_n6256_), .B(new_n5938_), .C(new_n3157_), .D(new_n2722_), .Y(new_n10222_));
  AND2X1   g07786(.A(new_n10222_), .B(pi0087), .Y(new_n10223_));
  NAND4X1  g07787(.A(new_n10223_), .B(new_n10221_), .C(new_n10218_), .D(new_n5989_), .Y(new_n10224_));
  AOI21X1  g07788(.A0(new_n10224_), .A1(new_n10217_), .B0(pi0075), .Y(new_n10225_));
  OR4X1    g07789(.A(new_n10182_), .B(new_n10175_), .C(new_n6855_), .D(new_n9689_), .Y(new_n10226_));
  AND2X1   g07790(.A(new_n5933_), .B(new_n5932_), .Y(new_n10227_));
  OR2X1    g07791(.A(new_n10197_), .B(new_n10227_), .Y(new_n10228_));
  AOI21X1  g07792(.A0(new_n6256_), .A1(new_n5938_), .B0(pi1091), .Y(new_n10229_));
  OAI21X1  g07793(.A0(new_n10229_), .A1(new_n6253_), .B0(pi0120), .Y(new_n10230_));
  NAND3X1  g07794(.A(new_n10230_), .B(new_n10228_), .C(new_n9766_), .Y(new_n10231_));
  AOI21X1  g07795(.A0(new_n10231_), .A1(new_n10226_), .B0(new_n3092_), .Y(new_n10232_));
  OAI21X1  g07796(.A0(new_n10196_), .A1(new_n3091_), .B0(pi0075), .Y(new_n10233_));
  OAI21X1  g07797(.A0(new_n10233_), .A1(new_n10232_), .B0(new_n5893_), .Y(new_n10234_));
  OAI21X1  g07798(.A0(new_n10234_), .A1(new_n10225_), .B0(new_n10172_), .Y(new_n10235_));
  NAND2X1  g07799(.A(new_n10218_), .B(new_n5989_), .Y(new_n10236_));
  INVX1    g07800(.A(new_n10214_), .Y(new_n10237_));
  OAI21X1  g07801(.A0(new_n10192_), .A1(new_n5983_), .B0(new_n10191_), .Y(new_n10238_));
  OR4X1    g07802(.A(new_n5069_), .B(new_n5065_), .C(new_n6269_), .D(new_n2756_), .Y(new_n10239_));
  AOI21X1  g07803(.A0(new_n5071_), .A1(new_n5052_), .B0(new_n6284_), .Y(new_n10240_));
  AND2X1   g07804(.A(new_n10240_), .B(new_n10239_), .Y(new_n10241_));
  OAI21X1  g07805(.A0(pi1093), .A1(pi0120), .B0(pi0299), .Y(new_n10242_));
  AOI21X1  g07806(.A0(new_n10241_), .A1(new_n10066_), .B0(new_n10242_), .Y(new_n10243_));
  NOR3X1   g07807(.A(new_n6269_), .B(new_n5051_), .C(new_n2756_), .Y(new_n10244_));
  OAI21X1  g07808(.A0(new_n5053_), .A1(new_n5050_), .B0(new_n6277_), .Y(new_n10245_));
  NOR4X1   g07809(.A(new_n10245_), .B(new_n10244_), .C(new_n7240_), .D(new_n2722_), .Y(new_n10246_));
  OR2X1    g07810(.A(new_n10213_), .B(pi0299), .Y(new_n10247_));
  OAI21X1  g07811(.A0(new_n10247_), .A1(new_n10246_), .B0(pi0039), .Y(new_n10248_));
  OAI22X1  g07812(.A0(new_n10248_), .A1(new_n10243_), .B0(new_n10238_), .B1(new_n10186_), .Y(new_n10249_));
  AOI21X1  g07813(.A0(new_n10249_), .A1(new_n2996_), .B0(new_n10237_), .Y(new_n10250_));
  MX2X1    g07814(.A(new_n10173_), .B(new_n5975_), .S0(pi0120), .Y(new_n10251_));
  OAI21X1  g07815(.A0(pi1093), .A1(pi0120), .B0(pi0100), .Y(new_n10252_));
  AOI21X1  g07816(.A0(new_n10251_), .A1(new_n10180_), .B0(new_n10252_), .Y(new_n10253_));
  OAI21X1  g07817(.A0(new_n10253_), .A1(new_n10250_), .B0(new_n3156_), .Y(new_n10254_));
  AOI21X1  g07818(.A0(new_n10254_), .A1(new_n10236_), .B0(pi0075), .Y(new_n10255_));
  OAI21X1  g07819(.A0(new_n10213_), .A1(new_n5936_), .B0(new_n5893_), .Y(new_n10256_));
  AOI21X1  g07820(.A0(new_n10170_), .A1(new_n2756_), .B0(new_n6633_), .Y(new_n10257_));
  OAI21X1  g07821(.A0(new_n10256_), .A1(new_n10255_), .B0(new_n10257_), .Y(new_n10258_));
  AOI21X1  g07822(.A0(new_n10258_), .A1(new_n10235_), .B0(new_n10168_), .Y(new_n10259_));
  NOR3X1   g07823(.A(new_n10182_), .B(new_n10175_), .C(new_n6077_), .Y(new_n10260_));
  OR2X1    g07824(.A(new_n10260_), .B(new_n10174_), .Y(new_n10261_));
  OR4X1    g07825(.A(new_n10260_), .B(new_n10213_), .C(new_n10166_), .D(new_n10165_), .Y(new_n10262_));
  AND2X1   g07826(.A(new_n10262_), .B(po1038), .Y(new_n10263_));
  AOI21X1  g07827(.A0(new_n10263_), .A1(new_n10261_), .B0(new_n6748_), .Y(new_n10264_));
  INVX1    g07828(.A(new_n6748_), .Y(new_n10265_));
  NAND3X1  g07829(.A(pi1092), .B(pi0982), .C(pi0951), .Y(new_n10266_));
  NOR2X1   g07830(.A(new_n10266_), .B(new_n2756_), .Y(new_n10267_));
  NOR2X1   g07831(.A(new_n10267_), .B(pi0120), .Y(new_n10268_));
  NOR2X1   g07832(.A(new_n10268_), .B(new_n10260_), .Y(new_n10269_));
  INVX1    g07833(.A(new_n10269_), .Y(new_n10270_));
  AOI21X1  g07834(.A0(new_n10270_), .A1(new_n10263_), .B0(new_n10265_), .Y(new_n10271_));
  OAI22X1  g07835(.A0(new_n10271_), .A1(new_n10264_), .B0(new_n10259_), .B1(po1038), .Y(new_n10272_));
  INVX1    g07836(.A(new_n10172_), .Y(new_n10273_));
  NAND4X1  g07837(.A(new_n5933_), .B(new_n5932_), .C(pi1093), .D(pi0120), .Y(new_n10274_));
  NOR3X1   g07838(.A(new_n10266_), .B(new_n2756_), .C(pi1091), .Y(new_n10275_));
  NOR2X1   g07839(.A(new_n10275_), .B(pi0120), .Y(new_n10276_));
  INVX1    g07840(.A(new_n10276_), .Y(new_n10277_));
  NOR3X1   g07841(.A(new_n10266_), .B(new_n2756_), .C(new_n2722_), .Y(new_n10278_));
  INVX1    g07842(.A(new_n10278_), .Y(new_n10279_));
  OR4X1    g07843(.A(pi0122), .B(pi0096), .C(pi0093), .D(pi0072), .Y(new_n10280_));
  OR4X1    g07844(.A(new_n10280_), .B(new_n2738_), .C(pi0090), .D(pi0024), .Y(new_n10281_));
  OR4X1    g07845(.A(new_n10281_), .B(new_n7666_), .C(new_n5193_), .D(new_n3053_), .Y(new_n10282_));
  NOR3X1   g07846(.A(new_n10282_), .B(new_n5094_), .C(new_n2829_), .Y(new_n10283_));
  AOI21X1  g07847(.A0(new_n10283_), .A1(new_n2550_), .B0(new_n10279_), .Y(new_n10284_));
  OR2X1    g07848(.A(new_n10284_), .B(new_n10277_), .Y(new_n10285_));
  AOI21X1  g07849(.A0(new_n10285_), .A1(new_n10274_), .B0(new_n5970_), .Y(new_n10286_));
  INVX1    g07850(.A(new_n10268_), .Y(new_n10287_));
  OAI21X1  g07851(.A0(new_n10287_), .A1(new_n9766_), .B0(new_n3091_), .Y(new_n10288_));
  AOI21X1  g07852(.A0(new_n10287_), .A1(new_n3092_), .B0(new_n3095_), .Y(new_n10289_));
  OAI21X1  g07853(.A0(new_n10288_), .A1(new_n10286_), .B0(new_n10289_), .Y(new_n10290_));
  OR4X1    g07854(.A(new_n3003_), .B(new_n2709_), .C(new_n5096_), .D(pi0070), .Y(new_n10291_));
  OR4X1    g07855(.A(new_n5094_), .B(new_n2829_), .C(new_n5258_), .D(pi0122), .Y(new_n10292_));
  OAI21X1  g07856(.A0(new_n10292_), .A1(new_n10291_), .B0(new_n10278_), .Y(new_n10293_));
  AOI22X1  g07857(.A0(new_n10293_), .A1(new_n10276_), .B0(new_n5975_), .B1(pi0120), .Y(new_n10294_));
  NAND2X1  g07858(.A(new_n6291_), .B(new_n2959_), .Y(new_n10295_));
  OAI21X1  g07859(.A0(new_n10295_), .A1(new_n10294_), .B0(pi0100), .Y(new_n10296_));
  NOR2X1   g07860(.A(new_n10287_), .B(new_n10180_), .Y(new_n10297_));
  AOI21X1  g07861(.A0(new_n10296_), .A1(new_n2996_), .B0(new_n10297_), .Y(new_n10298_));
  AOI21X1  g07862(.A0(new_n10268_), .A1(new_n6278_), .B0(pi0299), .Y(new_n10299_));
  OR2X1    g07863(.A(new_n10268_), .B(new_n6393_), .Y(new_n10300_));
  NOR2X1   g07864(.A(new_n10268_), .B(new_n6391_), .Y(new_n10301_));
  AOI21X1  g07865(.A0(new_n10301_), .A1(new_n5050_), .B0(new_n6278_), .Y(new_n10302_));
  OAI21X1  g07866(.A0(new_n10300_), .A1(new_n5050_), .B0(new_n10302_), .Y(new_n10303_));
  AOI21X1  g07867(.A0(new_n10268_), .A1(new_n6284_), .B0(new_n2953_), .Y(new_n10304_));
  AOI21X1  g07868(.A0(new_n10301_), .A1(new_n5070_), .B0(new_n6284_), .Y(new_n10305_));
  OAI21X1  g07869(.A0(new_n10300_), .A1(new_n5070_), .B0(new_n10305_), .Y(new_n10306_));
  AOI22X1  g07870(.A0(new_n10306_), .A1(new_n10304_), .B0(new_n10303_), .B1(new_n10299_), .Y(new_n10307_));
  INVX1    g07871(.A(new_n5937_), .Y(new_n10308_));
  INVX1    g07872(.A(new_n10267_), .Y(new_n10309_));
  OR4X1    g07873(.A(new_n2582_), .B(new_n2579_), .C(new_n5903_), .D(pi0088), .Y(new_n10310_));
  AOI21X1  g07874(.A0(new_n10310_), .A1(new_n2880_), .B0(new_n2748_), .Y(new_n10311_));
  AOI21X1  g07875(.A0(new_n10311_), .A1(new_n2743_), .B0(new_n5943_), .Y(new_n10312_));
  OAI21X1  g07876(.A0(new_n10312_), .A1(new_n2520_), .B0(new_n5899_), .Y(new_n10313_));
  AOI21X1  g07877(.A0(new_n10313_), .A1(new_n5897_), .B0(pi0051), .Y(new_n10314_));
  OAI21X1  g07878(.A0(new_n10314_), .A1(new_n2869_), .B0(new_n2526_), .Y(new_n10315_));
  NAND4X1  g07879(.A(new_n10315_), .B(new_n7806_), .C(pi0950), .D(new_n2548_), .Y(new_n10316_));
  NOR3X1   g07880(.A(new_n10266_), .B(new_n5258_), .C(pi0122), .Y(new_n10317_));
  OR4X1    g07881(.A(new_n10310_), .B(new_n6954_), .C(pi0090), .D(pi0058), .Y(new_n10318_));
  OR4X1    g07882(.A(new_n10318_), .B(new_n5012_), .C(pi0070), .D(pi0035), .Y(new_n10319_));
  OR4X1    g07883(.A(new_n3256_), .B(new_n2869_), .C(new_n5096_), .D(pi0096), .Y(new_n10320_));
  AOI21X1  g07884(.A0(new_n10319_), .A1(new_n5901_), .B0(new_n10320_), .Y(new_n10321_));
  AOI21X1  g07885(.A0(new_n10321_), .A1(pi0824), .B0(new_n10266_), .Y(new_n10322_));
  NAND2X1  g07886(.A(new_n10322_), .B(new_n5258_), .Y(new_n10323_));
  AND2X1   g07887(.A(pi1092), .B(pi0829), .Y(new_n10324_));
  NAND4X1  g07888(.A(new_n10324_), .B(pi0982), .C(pi0951), .D(pi0122), .Y(new_n10325_));
  OAI21X1  g07889(.A0(new_n10325_), .A1(new_n10321_), .B0(new_n10323_), .Y(new_n10326_));
  AOI21X1  g07890(.A0(new_n10317_), .A1(new_n10316_), .B0(new_n10326_), .Y(new_n10327_));
  OAI22X1  g07891(.A0(new_n10327_), .A1(new_n10308_), .B0(new_n10309_), .B1(new_n8273_), .Y(new_n10328_));
  AND2X1   g07892(.A(new_n10328_), .B(pi1091), .Y(new_n10329_));
  INVX1    g07893(.A(new_n10275_), .Y(new_n10330_));
  AOI21X1  g07894(.A0(new_n10321_), .A1(pi0824), .B0(new_n10330_), .Y(new_n10331_));
  NOR3X1   g07895(.A(new_n10331_), .B(new_n10329_), .C(pi0120), .Y(new_n10332_));
  INVX1    g07896(.A(new_n10185_), .Y(new_n10333_));
  OR2X1    g07897(.A(new_n10238_), .B(new_n10333_), .Y(new_n10334_));
  OAI21X1  g07898(.A0(new_n10334_), .A1(new_n10174_), .B0(new_n2959_), .Y(new_n10335_));
  OAI22X1  g07899(.A0(new_n10335_), .A1(new_n10332_), .B0(new_n10307_), .B1(new_n2959_), .Y(new_n10336_));
  AOI21X1  g07900(.A0(new_n10336_), .A1(new_n3277_), .B0(new_n10298_), .Y(new_n10337_));
  AOI21X1  g07901(.A0(new_n10268_), .A1(new_n3157_), .B0(new_n3156_), .Y(new_n10338_));
  OAI22X1  g07902(.A0(new_n2780_), .A1(pi0833), .B0(pi0829), .B1(pi0824), .Y(new_n10339_));
  OAI21X1  g07903(.A0(new_n10339_), .A1(new_n10291_), .B0(new_n10278_), .Y(new_n10340_));
  OAI21X1  g07904(.A0(new_n10291_), .A1(new_n5251_), .B0(new_n10275_), .Y(new_n10341_));
  AOI21X1  g07905(.A0(new_n10341_), .A1(new_n10340_), .B0(pi0120), .Y(new_n10342_));
  MX2X1    g07906(.A(new_n5986_), .B(new_n5981_), .S0(new_n5982_), .Y(new_n10343_));
  OAI21X1  g07907(.A0(new_n10343_), .A1(new_n10174_), .B0(new_n3085_), .Y(new_n10344_));
  OAI21X1  g07908(.A0(new_n10344_), .A1(new_n10342_), .B0(new_n10338_), .Y(new_n10345_));
  AND2X1   g07909(.A(new_n10345_), .B(new_n3095_), .Y(new_n10346_));
  OAI21X1  g07910(.A0(new_n10337_), .A1(pi0087), .B0(new_n10346_), .Y(new_n10347_));
  AOI21X1  g07911(.A0(new_n10347_), .A1(new_n10290_), .B0(new_n6309_), .Y(new_n10348_));
  NOR2X1   g07912(.A(new_n10176_), .B(new_n5975_), .Y(new_n10349_));
  NOR4X1   g07913(.A(new_n10266_), .B(new_n9394_), .C(new_n2756_), .D(pi1091), .Y(new_n10350_));
  INVX1    g07914(.A(new_n10350_), .Y(new_n10351_));
  AOI21X1  g07915(.A0(new_n10351_), .A1(new_n10293_), .B0(pi0120), .Y(new_n10352_));
  OAI21X1  g07916(.A0(new_n10352_), .A1(new_n10349_), .B0(new_n6291_), .Y(new_n10353_));
  NOR2X1   g07917(.A(new_n10268_), .B(new_n10195_), .Y(new_n10354_));
  AOI21X1  g07918(.A0(new_n10354_), .A1(new_n7761_), .B0(new_n3066_), .Y(new_n10355_));
  OAI21X1  g07919(.A0(new_n10354_), .A1(new_n3065_), .B0(pi0100), .Y(new_n10356_));
  AOI21X1  g07920(.A0(new_n10355_), .A1(new_n10353_), .B0(new_n10356_), .Y(new_n10357_));
  NAND4X1  g07921(.A(new_n10193_), .B(new_n10191_), .C(new_n10185_), .D(pi0120), .Y(new_n10358_));
  AND2X1   g07922(.A(new_n10322_), .B(new_n10219_), .Y(new_n10359_));
  OR2X1    g07923(.A(new_n10359_), .B(pi0120), .Y(new_n10360_));
  OAI21X1  g07924(.A0(new_n10360_), .A1(new_n10329_), .B0(new_n10358_), .Y(new_n10361_));
  AOI21X1  g07925(.A0(new_n10278_), .A1(new_n5959_), .B0(new_n10350_), .Y(new_n10362_));
  OAI22X1  g07926(.A0(new_n10362_), .A1(pi0120), .B0(new_n10176_), .B1(new_n10066_), .Y(new_n10363_));
  NOR3X1   g07927(.A(new_n10268_), .B(new_n10195_), .C(new_n6269_), .Y(new_n10364_));
  AOI21X1  g07928(.A0(new_n10363_), .A1(new_n6269_), .B0(new_n10364_), .Y(new_n10365_));
  OR2X1    g07929(.A(new_n10365_), .B(new_n5051_), .Y(new_n10366_));
  MX2X1    g07930(.A(new_n10363_), .B(new_n10354_), .S0(new_n5052_), .Y(new_n10367_));
  AOI21X1  g07931(.A0(new_n10367_), .A1(new_n5051_), .B0(new_n6278_), .Y(new_n10368_));
  OAI21X1  g07932(.A0(new_n10196_), .A1(new_n6277_), .B0(new_n10299_), .Y(new_n10369_));
  AOI21X1  g07933(.A0(new_n10368_), .A1(new_n10366_), .B0(new_n10369_), .Y(new_n10370_));
  OR2X1    g07934(.A(new_n10365_), .B(new_n5071_), .Y(new_n10371_));
  AOI21X1  g07935(.A0(new_n10367_), .A1(new_n5071_), .B0(new_n6284_), .Y(new_n10372_));
  OAI21X1  g07936(.A0(new_n6283_), .A1(new_n10212_), .B0(new_n10304_), .Y(new_n10373_));
  AOI21X1  g07937(.A0(new_n10372_), .A1(new_n10371_), .B0(new_n10373_), .Y(new_n10374_));
  NOR3X1   g07938(.A(new_n10374_), .B(new_n10370_), .C(new_n2959_), .Y(new_n10375_));
  AOI21X1  g07939(.A0(new_n10361_), .A1(new_n2959_), .B0(new_n10375_), .Y(new_n10376_));
  OR2X1    g07940(.A(new_n10376_), .B(pi0038), .Y(new_n10377_));
  OAI21X1  g07941(.A0(new_n10268_), .A1(new_n10195_), .B0(pi0038), .Y(new_n10378_));
  AND2X1   g07942(.A(new_n10378_), .B(new_n3026_), .Y(new_n10379_));
  AOI21X1  g07943(.A0(new_n10379_), .A1(new_n10377_), .B0(new_n10357_), .Y(new_n10380_));
  NAND2X1  g07944(.A(new_n10351_), .B(new_n10340_), .Y(new_n10381_));
  AOI22X1  g07945(.A0(new_n10381_), .A1(new_n10342_), .B0(new_n10344_), .B1(new_n10221_), .Y(new_n10382_));
  NAND2X1  g07946(.A(new_n10338_), .B(new_n10222_), .Y(new_n10383_));
  OAI22X1  g07947(.A0(new_n10383_), .A1(new_n10382_), .B0(new_n10380_), .B1(pi0087), .Y(new_n10384_));
  OAI21X1  g07948(.A0(new_n10268_), .A1(new_n10195_), .B0(new_n5970_), .Y(new_n10385_));
  OAI21X1  g07949(.A0(new_n10350_), .A1(new_n10284_), .B0(new_n10174_), .Y(new_n10386_));
  NAND3X1  g07950(.A(new_n10386_), .B(new_n10230_), .C(new_n9766_), .Y(new_n10387_));
  AOI21X1  g07951(.A0(new_n10387_), .A1(new_n10385_), .B0(new_n3092_), .Y(new_n10388_));
  OAI21X1  g07952(.A0(new_n10354_), .A1(new_n3091_), .B0(pi0075), .Y(new_n10389_));
  OAI21X1  g07953(.A0(new_n10389_), .A1(new_n10388_), .B0(new_n5893_), .Y(new_n10390_));
  AOI21X1  g07954(.A0(new_n10384_), .A1(new_n3095_), .B0(new_n10390_), .Y(new_n10391_));
  OAI22X1  g07955(.A0(new_n10391_), .A1(new_n10273_), .B0(new_n10348_), .B1(new_n6633_), .Y(new_n10392_));
  OAI21X1  g07956(.A0(new_n10266_), .A1(new_n2756_), .B0(new_n10170_), .Y(new_n10393_));
  AND2X1   g07957(.A(new_n10393_), .B(new_n10271_), .Y(new_n10394_));
  OAI21X1  g07958(.A0(new_n10194_), .A1(new_n10333_), .B0(new_n2959_), .Y(new_n10395_));
  NOR2X1   g07959(.A(new_n10229_), .B(new_n6272_), .Y(new_n10396_));
  MX2X1    g07960(.A(new_n10396_), .B(new_n9249_), .S0(new_n6270_), .Y(new_n10397_));
  MX2X1    g07961(.A(new_n10396_), .B(new_n9249_), .S0(new_n5052_), .Y(new_n10398_));
  INVX1    g07962(.A(new_n10398_), .Y(new_n10399_));
  AOI21X1  g07963(.A0(new_n10399_), .A1(new_n5051_), .B0(new_n6278_), .Y(new_n10400_));
  OAI21X1  g07964(.A0(new_n10397_), .A1(new_n5051_), .B0(new_n10400_), .Y(new_n10401_));
  AOI21X1  g07965(.A0(new_n6278_), .A1(new_n9249_), .B0(pi0299), .Y(new_n10402_));
  AOI21X1  g07966(.A0(new_n10399_), .A1(new_n5071_), .B0(new_n6284_), .Y(new_n10403_));
  OAI21X1  g07967(.A0(new_n10397_), .A1(new_n5071_), .B0(new_n10403_), .Y(new_n10404_));
  AOI21X1  g07968(.A0(new_n6284_), .A1(new_n9249_), .B0(new_n2953_), .Y(new_n10405_));
  AOI22X1  g07969(.A0(new_n10405_), .A1(new_n10404_), .B0(new_n10402_), .B1(new_n10401_), .Y(new_n10406_));
  OAI21X1  g07970(.A0(new_n10406_), .A1(new_n2959_), .B0(new_n2996_), .Y(new_n10407_));
  INVX1    g07971(.A(new_n10407_), .Y(new_n10408_));
  AOI21X1  g07972(.A0(new_n9249_), .A1(pi0038), .B0(pi0100), .Y(new_n10409_));
  INVX1    g07973(.A(new_n10409_), .Y(new_n10410_));
  AOI21X1  g07974(.A0(new_n10408_), .A1(new_n10395_), .B0(new_n10410_), .Y(new_n10411_));
  AOI21X1  g07975(.A0(new_n10212_), .A1(new_n5978_), .B0(new_n10411_), .Y(new_n10412_));
  NOR2X1   g07976(.A(new_n10412_), .B(pi0087), .Y(new_n10413_));
  AOI21X1  g07977(.A0(new_n10223_), .A1(new_n10221_), .B0(new_n10413_), .Y(new_n10414_));
  NOR3X1   g07978(.A(new_n10229_), .B(new_n6253_), .C(new_n6252_), .Y(new_n10415_));
  AOI21X1  g07979(.A0(new_n9249_), .A1(new_n6252_), .B0(new_n3095_), .Y(new_n10416_));
  INVX1    g07980(.A(new_n10416_), .Y(new_n10417_));
  OAI22X1  g07981(.A0(new_n10417_), .A1(new_n10415_), .B0(new_n10414_), .B1(pi0075), .Y(new_n10418_));
  NAND2X1  g07982(.A(new_n10418_), .B(new_n10169_), .Y(new_n10419_));
  AOI21X1  g07983(.A0(new_n10334_), .A1(new_n2959_), .B0(new_n5966_), .Y(new_n10420_));
  OAI21X1  g07984(.A0(new_n10420_), .A1(pi0100), .B0(new_n5979_), .Y(new_n10421_));
  AOI21X1  g07985(.A0(new_n10421_), .A1(new_n3156_), .B0(new_n5989_), .Y(new_n10422_));
  OAI21X1  g07986(.A0(new_n10422_), .A1(pi0075), .B0(new_n5936_), .Y(new_n10423_));
  NOR2X1   g07987(.A(new_n10170_), .B(new_n6633_), .Y(new_n10424_));
  NOR2X1   g07988(.A(new_n10260_), .B(new_n5893_), .Y(new_n10425_));
  AOI21X1  g07989(.A0(new_n10424_), .A1(new_n10423_), .B0(new_n10425_), .Y(new_n10426_));
  NAND2X1  g07990(.A(new_n10426_), .B(new_n10419_), .Y(new_n10427_));
  AND2X1   g07991(.A(new_n10264_), .B(pi0120), .Y(new_n10428_));
  AOI22X1  g07992(.A0(new_n10428_), .A1(new_n10427_), .B0(new_n10394_), .B1(new_n10392_), .Y(new_n10429_));
  OAI21X1  g07993(.A0(new_n10429_), .A1(new_n10167_), .B0(new_n10272_), .Y(po0278));
  OR4X1    g07994(.A(pi0136), .B(pi0135), .C(pi0134), .D(pi0130), .Y(new_n10431_));
  NOR4X1   g07995(.A(new_n10431_), .B(pi0132), .C(pi0126), .D(pi0121), .Y(new_n10432_));
  INVX1    g07996(.A(new_n10432_), .Y(new_n10433_));
  NOR2X1   g07997(.A(pi0133), .B(pi0125), .Y(new_n10434_));
  XOR2X1   g07998(.A(new_n10434_), .B(pi0121), .Y(new_n10435_));
  AND2X1   g07999(.A(new_n10435_), .B(new_n10433_), .Y(new_n10436_));
  NOR4X1   g08000(.A(pi0084), .B(pi0071), .C(pi0068), .D(pi0067), .Y(new_n10437_));
  INVX1    g08001(.A(new_n10437_), .Y(new_n10438_));
  OR4X1    g08002(.A(new_n10438_), .B(new_n10436_), .C(pi0087), .D(pi0051), .Y(new_n10439_));
  AND2X1   g08003(.A(new_n10437_), .B(new_n2516_), .Y(new_n10440_));
  NOR4X1   g08004(.A(pi0468), .B(pi0332), .C(pi0146), .D(new_n2516_), .Y(new_n10441_));
  NOR2X1   g08005(.A(new_n10441_), .B(new_n4613_), .Y(new_n10442_));
  AND2X1   g08006(.A(pi0146), .B(pi0051), .Y(new_n10443_));
  NOR4X1   g08007(.A(new_n10443_), .B(new_n10442_), .C(new_n10440_), .D(new_n5057_), .Y(new_n10444_));
  AOI21X1  g08008(.A0(new_n9934_), .A1(pi0087), .B0(new_n5237_), .Y(new_n10445_));
  OAI21X1  g08009(.A0(new_n10444_), .A1(pi0087), .B0(new_n10445_), .Y(new_n10446_));
  NAND3X1  g08010(.A(new_n10446_), .B(new_n10439_), .C(po1038), .Y(new_n10447_));
  NOR4X1   g08011(.A(pi0468), .B(pi0332), .C(pi0142), .D(new_n2516_), .Y(new_n10448_));
  NOR2X1   g08012(.A(new_n10448_), .B(new_n7548_), .Y(new_n10449_));
  INVX1    g08013(.A(new_n10449_), .Y(new_n10450_));
  NOR2X1   g08014(.A(new_n10440_), .B(new_n5057_), .Y(new_n10451_));
  INVX1    g08015(.A(new_n10451_), .Y(new_n10452_));
  AOI21X1  g08016(.A0(pi0142), .A1(pi0051), .B0(new_n10452_), .Y(new_n10453_));
  AOI21X1  g08017(.A0(new_n10453_), .A1(new_n10450_), .B0(pi0299), .Y(new_n10454_));
  OAI21X1  g08018(.A0(new_n10444_), .A1(new_n2953_), .B0(pi0232), .Y(new_n10455_));
  NOR2X1   g08019(.A(new_n10455_), .B(new_n10454_), .Y(new_n10456_));
  INVX1    g08020(.A(new_n10456_), .Y(new_n10457_));
  AOI21X1  g08021(.A0(new_n10457_), .A1(pi0038), .B0(pi0100), .Y(new_n10458_));
  INVX1    g08022(.A(new_n10440_), .Y(new_n10459_));
  AOI21X1  g08023(.A0(new_n10459_), .A1(pi0038), .B0(pi0100), .Y(new_n10460_));
  INVX1    g08024(.A(pi0179), .Y(new_n10461_));
  INVX1    g08025(.A(new_n10448_), .Y(new_n10462_));
  NAND4X1  g08026(.A(new_n7660_), .B(new_n2615_), .C(new_n2614_), .D(new_n7658_), .Y(new_n10463_));
  NOR4X1   g08027(.A(new_n10463_), .B(new_n2621_), .C(new_n8560_), .D(new_n9524_), .Y(new_n10464_));
  INVX1    g08028(.A(new_n10464_), .Y(new_n10465_));
  NAND3X1  g08029(.A(new_n5907_), .B(new_n2526_), .C(new_n5134_), .Y(new_n10466_));
  OR4X1    g08030(.A(new_n10466_), .B(new_n6954_), .C(new_n2498_), .D(pi0058), .Y(new_n10467_));
  NOR4X1   g08031(.A(new_n10467_), .B(new_n10465_), .C(new_n7666_), .D(new_n2548_), .Y(new_n10468_));
  INVX1    g08032(.A(new_n10468_), .Y(new_n10469_));
  AOI21X1  g08033(.A0(new_n10466_), .A1(new_n10437_), .B0(pi0051), .Y(new_n10470_));
  OR4X1    g08034(.A(new_n10463_), .B(new_n2621_), .C(new_n2468_), .D(pi0036), .Y(new_n10471_));
  NOR4X1   g08035(.A(new_n10471_), .B(new_n2476_), .C(new_n2581_), .D(pi0050), .Y(new_n10472_));
  AOI21X1  g08036(.A0(new_n10464_), .A1(pi0086), .B0(new_n10472_), .Y(new_n10473_));
  INVX1    g08037(.A(new_n6768_), .Y(new_n10474_));
  NOR4X1   g08038(.A(new_n10474_), .B(new_n7842_), .C(new_n2474_), .D(pi0024), .Y(new_n10475_));
  AOI21X1  g08039(.A0(new_n10475_), .A1(new_n10464_), .B0(new_n10438_), .Y(new_n10476_));
  OAI21X1  g08040(.A0(new_n10473_), .A1(new_n8307_), .B0(new_n10476_), .Y(new_n10477_));
  AND2X1   g08041(.A(new_n10477_), .B(new_n10470_), .Y(new_n10478_));
  AND2X1   g08042(.A(new_n10478_), .B(new_n3002_), .Y(new_n10479_));
  NOR3X1   g08043(.A(new_n10466_), .B(new_n7734_), .C(pi0024), .Y(new_n10480_));
  NAND3X1  g08044(.A(new_n10480_), .B(new_n10472_), .C(new_n6769_), .Y(new_n10481_));
  NOR2X1   g08045(.A(new_n10481_), .B(new_n3256_), .Y(new_n10482_));
  NOR2X1   g08046(.A(new_n10482_), .B(new_n10459_), .Y(new_n10483_));
  INVX1    g08047(.A(new_n10483_), .Y(new_n10484_));
  NOR2X1   g08048(.A(new_n10484_), .B(new_n10479_), .Y(new_n10485_));
  MX2X1    g08049(.A(new_n10485_), .B(new_n10440_), .S0(new_n5033_), .Y(new_n10486_));
  NAND2X1  g08050(.A(new_n10486_), .B(new_n10469_), .Y(new_n10487_));
  NOR4X1   g08051(.A(new_n10482_), .B(new_n10479_), .C(new_n10468_), .D(new_n10459_), .Y(new_n10488_));
  NOR2X1   g08052(.A(new_n10488_), .B(new_n5033_), .Y(new_n10489_));
  AND2X1   g08053(.A(new_n5033_), .B(pi0051), .Y(new_n10490_));
  AND2X1   g08054(.A(new_n8218_), .B(pi0072), .Y(new_n10491_));
  OR2X1    g08055(.A(new_n10491_), .B(new_n10490_), .Y(new_n10492_));
  AND2X1   g08056(.A(new_n10492_), .B(new_n5033_), .Y(new_n10493_));
  NOR2X1   g08057(.A(new_n10493_), .B(new_n10489_), .Y(new_n10494_));
  INVX1    g08058(.A(new_n10494_), .Y(new_n10495_));
  MX2X1    g08059(.A(new_n10495_), .B(new_n10487_), .S0(pi0144), .Y(new_n10496_));
  AOI21X1  g08060(.A0(new_n10496_), .A1(new_n10462_), .B0(new_n5225_), .Y(new_n10497_));
  OR4X1    g08061(.A(new_n10466_), .B(new_n7734_), .C(pi0051), .D(pi0024), .Y(new_n10498_));
  NOR4X1   g08062(.A(new_n10498_), .B(new_n8541_), .C(new_n2586_), .D(new_n2581_), .Y(new_n10499_));
  AND2X1   g08063(.A(new_n5033_), .B(new_n3002_), .Y(new_n10500_));
  AND2X1   g08064(.A(new_n10500_), .B(new_n10499_), .Y(new_n10501_));
  OR4X1    g08065(.A(new_n10501_), .B(new_n10493_), .C(new_n10489_), .D(new_n2972_), .Y(new_n10502_));
  OAI21X1  g08066(.A0(new_n10499_), .A1(pi0072), .B0(new_n5190_), .Y(new_n10503_));
  MX2X1    g08067(.A(new_n10503_), .B(new_n10488_), .S0(new_n5057_), .Y(new_n10504_));
  AOI21X1  g08068(.A0(new_n10504_), .A1(new_n2972_), .B0(pi0144), .Y(new_n10505_));
  NOR2X1   g08069(.A(new_n10485_), .B(new_n5033_), .Y(new_n10506_));
  NOR4X1   g08070(.A(new_n10506_), .B(new_n10482_), .C(new_n10468_), .D(new_n10451_), .Y(new_n10507_));
  OAI21X1  g08071(.A0(new_n10507_), .A1(new_n10450_), .B0(new_n5225_), .Y(new_n10508_));
  AOI21X1  g08072(.A0(new_n10505_), .A1(new_n10502_), .B0(new_n10508_), .Y(new_n10509_));
  NOR3X1   g08073(.A(new_n10509_), .B(new_n10497_), .C(new_n10461_), .Y(new_n10510_));
  INVX1    g08074(.A(new_n10489_), .Y(new_n10511_));
  INVX1    g08075(.A(new_n8701_), .Y(new_n10512_));
  MX2X1    g08076(.A(new_n10512_), .B(new_n8700_), .S0(pi0024), .Y(new_n10513_));
  MX2X1    g08077(.A(new_n10513_), .B(new_n8700_), .S0(pi0314), .Y(new_n10514_));
  NAND4X1  g08078(.A(new_n5907_), .B(new_n3002_), .C(new_n2526_), .D(new_n5134_), .Y(new_n10515_));
  OAI21X1  g08079(.A0(new_n10515_), .A1(new_n10514_), .B0(new_n2516_), .Y(new_n10516_));
  OAI21X1  g08080(.A0(new_n10516_), .A1(new_n10491_), .B0(new_n5033_), .Y(new_n10517_));
  NAND3X1  g08081(.A(new_n10517_), .B(new_n10511_), .C(pi0142), .Y(new_n10518_));
  AND2X1   g08082(.A(new_n10488_), .B(new_n5057_), .Y(new_n10519_));
  OAI21X1  g08083(.A0(new_n10514_), .A1(new_n2487_), .B0(new_n2548_), .Y(new_n10520_));
  AOI21X1  g08084(.A0(new_n10520_), .A1(new_n5190_), .B0(new_n5057_), .Y(new_n10521_));
  OAI21X1  g08085(.A0(new_n10521_), .A1(new_n10519_), .B0(new_n2972_), .Y(new_n10522_));
  NAND3X1  g08086(.A(new_n10522_), .B(new_n10518_), .C(new_n7548_), .Y(new_n10523_));
  INVX1    g08087(.A(new_n10488_), .Y(new_n10524_));
  AOI21X1  g08088(.A0(new_n10524_), .A1(new_n10449_), .B0(pi0180), .Y(new_n10525_));
  NOR2X1   g08089(.A(new_n10513_), .B(new_n2487_), .Y(new_n10526_));
  OAI21X1  g08090(.A0(new_n10526_), .A1(pi0072), .B0(new_n5190_), .Y(new_n10527_));
  AOI21X1  g08091(.A0(new_n10527_), .A1(new_n5033_), .B0(new_n10519_), .Y(new_n10528_));
  NOR2X1   g08092(.A(new_n10528_), .B(pi0142), .Y(new_n10529_));
  INVX1    g08093(.A(new_n10500_), .Y(new_n10530_));
  NOR3X1   g08094(.A(new_n10513_), .B(new_n10530_), .C(new_n2487_), .Y(new_n10531_));
  NOR4X1   g08095(.A(new_n10531_), .B(new_n10493_), .C(new_n10489_), .D(new_n2972_), .Y(new_n10532_));
  NOR3X1   g08096(.A(new_n10532_), .B(new_n10529_), .C(pi0144), .Y(new_n10533_));
  NOR3X1   g08097(.A(new_n10479_), .B(new_n10468_), .C(new_n10459_), .Y(new_n10534_));
  NOR3X1   g08098(.A(pi0468), .B(pi0332), .C(pi0051), .Y(new_n10535_));
  INVX1    g08099(.A(new_n10535_), .Y(new_n10536_));
  NOR2X1   g08100(.A(new_n10536_), .B(new_n10534_), .Y(new_n10537_));
  NOR2X1   g08101(.A(new_n10537_), .B(new_n10489_), .Y(new_n10538_));
  INVX1    g08102(.A(new_n10479_), .Y(new_n10539_));
  AOI21X1  g08103(.A0(new_n10539_), .A1(new_n10440_), .B0(new_n5057_), .Y(new_n10540_));
  NOR4X1   g08104(.A(new_n10437_), .B(pi0468), .C(pi0332), .D(pi0051), .Y(new_n10541_));
  OAI22X1  g08105(.A0(new_n10541_), .A1(new_n10500_), .B0(new_n10478_), .B1(new_n3256_), .Y(new_n10542_));
  INVX1    g08106(.A(new_n10542_), .Y(new_n10543_));
  MX2X1    g08107(.A(new_n10543_), .B(new_n10540_), .S0(new_n2972_), .Y(new_n10544_));
  OR2X1    g08108(.A(new_n10544_), .B(new_n10486_), .Y(new_n10545_));
  AOI21X1  g08109(.A0(new_n10545_), .A1(new_n10538_), .B0(new_n7548_), .Y(new_n10546_));
  OR2X1    g08110(.A(new_n10546_), .B(new_n5225_), .Y(new_n10547_));
  OAI21X1  g08111(.A0(new_n10547_), .A1(new_n10533_), .B0(new_n10461_), .Y(new_n10548_));
  AOI21X1  g08112(.A0(new_n10525_), .A1(new_n10523_), .B0(new_n10548_), .Y(new_n10549_));
  OAI21X1  g08113(.A0(new_n10549_), .A1(new_n10510_), .B0(new_n2953_), .Y(new_n10550_));
  INVX1    g08114(.A(new_n7107_), .Y(new_n10551_));
  NOR2X1   g08115(.A(new_n10441_), .B(pi0161), .Y(new_n10552_));
  NAND3X1  g08116(.A(new_n10486_), .B(new_n10469_), .C(pi0146), .Y(new_n10553_));
  AOI21X1  g08117(.A0(new_n10469_), .A1(new_n10437_), .B0(new_n10536_), .Y(new_n10554_));
  NOR3X1   g08118(.A(new_n10554_), .B(new_n10489_), .C(pi0146), .Y(new_n10555_));
  NOR2X1   g08119(.A(new_n10555_), .B(new_n4613_), .Y(new_n10556_));
  AOI22X1  g08120(.A0(new_n10556_), .A1(new_n10553_), .B0(new_n10552_), .B1(new_n10495_), .Y(new_n10557_));
  OR4X1    g08121(.A(new_n10501_), .B(new_n10493_), .C(new_n10489_), .D(new_n2800_), .Y(new_n10558_));
  AOI21X1  g08122(.A0(new_n10504_), .A1(new_n2800_), .B0(pi0161), .Y(new_n10559_));
  INVX1    g08123(.A(new_n10490_), .Y(new_n10560_));
  NOR3X1   g08124(.A(new_n10536_), .B(new_n10468_), .C(new_n10438_), .Y(new_n10561_));
  OAI21X1  g08125(.A0(new_n10481_), .A1(new_n3256_), .B0(new_n10561_), .Y(new_n10562_));
  AOI22X1  g08126(.A0(new_n10562_), .A1(new_n10560_), .B0(new_n10459_), .B1(pi0146), .Y(new_n10563_));
  NOR3X1   g08127(.A(new_n10563_), .B(new_n10519_), .C(new_n4613_), .Y(new_n10564_));
  AOI21X1  g08128(.A0(new_n10559_), .A1(new_n10558_), .B0(new_n10564_), .Y(new_n10565_));
  OAI22X1  g08129(.A0(new_n10565_), .A1(new_n7140_), .B0(new_n10557_), .B1(new_n10551_), .Y(new_n10566_));
  OAI21X1  g08130(.A0(new_n10521_), .A1(new_n10519_), .B0(new_n2800_), .Y(new_n10567_));
  NAND3X1  g08131(.A(new_n10517_), .B(new_n10511_), .C(pi0146), .Y(new_n10568_));
  NAND3X1  g08132(.A(new_n10568_), .B(new_n10567_), .C(new_n7139_), .Y(new_n10569_));
  OR4X1    g08133(.A(new_n10531_), .B(new_n10493_), .C(new_n10489_), .D(new_n2800_), .Y(new_n10570_));
  AND2X1   g08134(.A(new_n10570_), .B(new_n7107_), .Y(new_n10571_));
  OAI21X1  g08135(.A0(new_n10528_), .A1(pi0146), .B0(new_n10571_), .Y(new_n10572_));
  NAND3X1  g08136(.A(new_n10572_), .B(new_n10569_), .C(new_n4613_), .Y(new_n10573_));
  MX2X1    g08137(.A(new_n10543_), .B(new_n10540_), .S0(new_n2800_), .Y(new_n10574_));
  OAI21X1  g08138(.A0(new_n10574_), .A1(new_n10486_), .B0(new_n10538_), .Y(new_n10575_));
  NAND2X1  g08139(.A(new_n10575_), .B(new_n7107_), .Y(new_n10576_));
  OR4X1    g08140(.A(new_n10488_), .B(new_n10441_), .C(new_n2953_), .D(pi0158), .Y(new_n10577_));
  AND2X1   g08141(.A(new_n10577_), .B(pi0161), .Y(new_n10578_));
  AOI21X1  g08142(.A0(new_n10578_), .A1(new_n10576_), .B0(pi0156), .Y(new_n10579_));
  AOI22X1  g08143(.A0(new_n10579_), .A1(new_n10573_), .B0(new_n10566_), .B1(pi0156), .Y(new_n10580_));
  AOI21X1  g08144(.A0(new_n10580_), .A1(new_n10550_), .B0(new_n7300_), .Y(new_n10581_));
  NOR4X1   g08145(.A(new_n10467_), .B(new_n10471_), .C(new_n3256_), .D(new_n8560_), .Y(new_n10582_));
  NOR2X1   g08146(.A(new_n10582_), .B(new_n10459_), .Y(new_n10583_));
  INVX1    g08147(.A(new_n10583_), .Y(new_n10584_));
  AOI21X1  g08148(.A0(new_n10584_), .A1(new_n5057_), .B0(new_n5046_), .Y(new_n10585_));
  INVX1    g08149(.A(new_n10585_), .Y(new_n10586_));
  AND2X1   g08150(.A(new_n2964_), .B(pi0222), .Y(new_n10587_));
  NOR2X1   g08151(.A(new_n5911_), .B(new_n2555_), .Y(new_n10588_));
  NOR2X1   g08152(.A(new_n10588_), .B(pi0051), .Y(new_n10589_));
  MX2X1    g08153(.A(new_n10589_), .B(new_n10583_), .S0(new_n5057_), .Y(new_n10590_));
  OAI21X1  g08154(.A0(new_n10590_), .A1(new_n2972_), .B0(new_n10587_), .Y(new_n10591_));
  AOI21X1  g08155(.A0(new_n10586_), .A1(new_n2972_), .B0(new_n10591_), .Y(new_n10592_));
  OR2X1    g08156(.A(new_n10592_), .B(new_n6886_), .Y(new_n10593_));
  NOR3X1   g08157(.A(pi0468), .B(pi0332), .C(pi0287), .Y(new_n10594_));
  AOI21X1  g08158(.A0(new_n10594_), .A1(new_n2516_), .B0(new_n10590_), .Y(new_n10595_));
  NAND3X1  g08159(.A(new_n10595_), .B(new_n10462_), .C(pi0224), .Y(new_n10596_));
  OAI22X1  g08160(.A0(new_n10448_), .A1(new_n10440_), .B0(pi0223), .B1(new_n2960_), .Y(new_n10597_));
  OAI21X1  g08161(.A0(pi0223), .A1(new_n2960_), .B0(new_n10541_), .Y(new_n10598_));
  NAND3X1  g08162(.A(new_n10598_), .B(new_n10597_), .C(new_n7548_), .Y(new_n10599_));
  AOI21X1  g08163(.A0(new_n10596_), .A1(new_n10593_), .B0(new_n10599_), .Y(new_n10600_));
  INVX1    g08164(.A(new_n10541_), .Y(new_n10601_));
  INVX1    g08165(.A(new_n10594_), .Y(new_n10602_));
  NOR2X1   g08166(.A(new_n10583_), .B(pi0051), .Y(new_n10603_));
  INVX1    g08167(.A(new_n10603_), .Y(new_n10604_));
  AOI22X1  g08168(.A0(new_n10604_), .A1(new_n7862_), .B0(new_n10602_), .B1(new_n10601_), .Y(new_n10605_));
  OR2X1    g08169(.A(new_n10605_), .B(new_n10453_), .Y(new_n10606_));
  AND2X1   g08170(.A(new_n10606_), .B(new_n6886_), .Y(new_n10607_));
  AND2X1   g08171(.A(new_n10597_), .B(pi0144), .Y(new_n10608_));
  MX2X1    g08172(.A(new_n10583_), .B(new_n5033_), .S0(pi0051), .Y(new_n10609_));
  INVX1    g08173(.A(new_n10609_), .Y(new_n10610_));
  OAI21X1  g08174(.A0(new_n2972_), .A1(new_n2516_), .B0(new_n10587_), .Y(new_n10611_));
  OAI21X1  g08175(.A0(new_n10611_), .A1(new_n10610_), .B0(new_n10608_), .Y(new_n10612_));
  AOI21X1  g08176(.A0(new_n10607_), .A1(new_n10437_), .B0(new_n10612_), .Y(new_n10613_));
  OR2X1    g08177(.A(new_n10613_), .B(new_n5226_), .Y(new_n10614_));
  AND2X1   g08178(.A(new_n10612_), .B(new_n5226_), .Y(new_n10615_));
  OAI21X1  g08179(.A0(new_n10599_), .A1(new_n10592_), .B0(new_n10615_), .Y(new_n10616_));
  AND2X1   g08180(.A(new_n10616_), .B(new_n2953_), .Y(new_n10617_));
  OAI21X1  g08181(.A0(new_n10614_), .A1(new_n10600_), .B0(new_n10617_), .Y(new_n10618_));
  OAI21X1  g08182(.A0(new_n10583_), .A1(new_n10441_), .B0(pi0161), .Y(new_n10619_));
  NOR2X1   g08183(.A(new_n10585_), .B(pi0146), .Y(new_n10620_));
  OAI21X1  g08184(.A0(new_n10590_), .A1(new_n2800_), .B0(new_n4613_), .Y(new_n10621_));
  OAI21X1  g08185(.A0(new_n10621_), .A1(new_n10620_), .B0(new_n10619_), .Y(new_n10622_));
  AND2X1   g08186(.A(new_n10622_), .B(new_n5241_), .Y(new_n10623_));
  AOI21X1  g08187(.A0(new_n10602_), .A1(new_n10582_), .B0(new_n10459_), .Y(new_n10624_));
  INVX1    g08188(.A(new_n10624_), .Y(new_n10625_));
  AOI22X1  g08189(.A0(new_n10625_), .A1(new_n10442_), .B0(new_n10595_), .B1(new_n10552_), .Y(new_n10626_));
  OAI22X1  g08190(.A0(new_n10626_), .A1(new_n2438_), .B0(new_n10623_), .B1(new_n6893_), .Y(new_n10627_));
  OAI21X1  g08191(.A0(new_n10444_), .A1(new_n10440_), .B0(new_n5242_), .Y(new_n10628_));
  AND2X1   g08192(.A(new_n10628_), .B(new_n7457_), .Y(new_n10629_));
  NAND2X1  g08193(.A(new_n10628_), .B(new_n7429_), .Y(new_n10630_));
  OAI21X1  g08194(.A0(new_n10630_), .A1(new_n10623_), .B0(pi0232), .Y(new_n10631_));
  AOI21X1  g08195(.A0(new_n10629_), .A1(new_n10627_), .B0(new_n10631_), .Y(new_n10632_));
  MX2X1    g08196(.A(new_n10587_), .B(new_n5241_), .S0(pi0299), .Y(new_n10633_));
  NAND3X1  g08197(.A(new_n10437_), .B(new_n5237_), .C(new_n2516_), .Y(new_n10634_));
  AOI21X1  g08198(.A0(new_n10633_), .A1(new_n10582_), .B0(new_n10634_), .Y(new_n10635_));
  OR2X1    g08199(.A(new_n10635_), .B(new_n2959_), .Y(new_n10636_));
  AOI21X1  g08200(.A0(new_n10632_), .A1(new_n10618_), .B0(new_n10636_), .Y(new_n10637_));
  NOR3X1   g08201(.A(new_n10488_), .B(pi0232), .C(pi0039), .Y(new_n10638_));
  NOR3X1   g08202(.A(new_n10638_), .B(new_n10637_), .C(new_n10581_), .Y(new_n10639_));
  OAI22X1  g08203(.A0(new_n10639_), .A1(pi0038), .B0(new_n10460_), .B1(new_n10458_), .Y(new_n10640_));
  INVX1    g08204(.A(new_n5821_), .Y(new_n10641_));
  AOI21X1  g08205(.A0(new_n10440_), .A1(pi0100), .B0(new_n10641_), .Y(new_n10642_));
  INVX1    g08206(.A(new_n10642_), .Y(new_n10643_));
  AOI21X1  g08207(.A0(new_n10456_), .A1(pi0100), .B0(new_n10643_), .Y(new_n10644_));
  AND2X1   g08208(.A(new_n3125_), .B(new_n3156_), .Y(new_n10645_));
  OAI21X1  g08209(.A0(new_n10438_), .A1(pi0051), .B0(new_n10645_), .Y(new_n10646_));
  MX2X1    g08210(.A(new_n8717_), .B(new_n8705_), .S0(pi0299), .Y(new_n10647_));
  OR4X1    g08211(.A(new_n10647_), .B(pi0468), .C(pi0332), .D(new_n5237_), .Y(new_n10648_));
  AOI22X1  g08212(.A0(new_n10648_), .A1(pi0087), .B0(new_n10435_), .B1(new_n10433_), .Y(new_n10649_));
  OAI21X1  g08213(.A0(new_n10646_), .A1(new_n10456_), .B0(new_n10649_), .Y(new_n10650_));
  AOI21X1  g08214(.A0(new_n10644_), .A1(new_n10640_), .B0(new_n10650_), .Y(new_n10651_));
  INVX1    g08215(.A(new_n10443_), .Y(new_n10652_));
  AND2X1   g08216(.A(new_n10516_), .B(new_n5033_), .Y(new_n10653_));
  AOI21X1  g08217(.A0(new_n10653_), .A1(new_n10652_), .B0(new_n4613_), .Y(new_n10654_));
  OR4X1    g08218(.A(new_n10485_), .B(pi0468), .C(pi0332), .D(pi0146), .Y(new_n10655_));
  INVX1    g08219(.A(new_n10481_), .Y(new_n10656_));
  OR4X1    g08220(.A(new_n10656_), .B(new_n10477_), .C(new_n10466_), .D(new_n10438_), .Y(new_n10657_));
  AOI21X1  g08221(.A0(new_n10657_), .A1(new_n10470_), .B0(new_n3256_), .Y(new_n10658_));
  AOI21X1  g08222(.A0(new_n10601_), .A1(new_n10530_), .B0(new_n10658_), .Y(new_n10659_));
  AOI21X1  g08223(.A0(new_n10659_), .A1(pi0146), .B0(pi0161), .Y(new_n10660_));
  AND2X1   g08224(.A(new_n10660_), .B(new_n10655_), .Y(new_n10661_));
  OAI21X1  g08225(.A0(new_n10661_), .A1(new_n10654_), .B0(new_n7107_), .Y(new_n10662_));
  INVX1    g08226(.A(new_n10442_), .Y(new_n10663_));
  OAI22X1  g08227(.A0(new_n10574_), .A1(pi0161), .B0(new_n10531_), .B1(new_n10663_), .Y(new_n10664_));
  AOI21X1  g08228(.A0(new_n10664_), .A1(new_n7139_), .B0(new_n5237_), .Y(new_n10665_));
  AOI21X1  g08229(.A0(new_n10665_), .A1(new_n10662_), .B0(new_n8876_), .Y(new_n10666_));
  NAND2X1  g08230(.A(pi0142), .B(pi0051), .Y(new_n10667_));
  AND2X1   g08231(.A(new_n10653_), .B(new_n10667_), .Y(new_n10668_));
  OR4X1    g08232(.A(new_n10485_), .B(pi0468), .C(pi0332), .D(pi0142), .Y(new_n10669_));
  AOI21X1  g08233(.A0(new_n10659_), .A1(pi0142), .B0(pi0144), .Y(new_n10670_));
  AOI21X1  g08234(.A0(new_n10670_), .A1(new_n10669_), .B0(new_n5225_), .Y(new_n10671_));
  OAI21X1  g08235(.A0(new_n10668_), .A1(new_n7548_), .B0(new_n10671_), .Y(new_n10672_));
  NOR2X1   g08236(.A(new_n10531_), .B(new_n10450_), .Y(new_n10673_));
  OAI21X1  g08237(.A0(new_n10544_), .A1(pi0144), .B0(new_n5225_), .Y(new_n10674_));
  NOR2X1   g08238(.A(new_n10674_), .B(new_n10673_), .Y(new_n10675_));
  NOR2X1   g08239(.A(new_n10675_), .B(new_n10461_), .Y(new_n10676_));
  OR2X1    g08240(.A(new_n10501_), .B(new_n10450_), .Y(new_n10677_));
  AOI21X1  g08241(.A0(new_n10481_), .A1(new_n10437_), .B0(pi0051), .Y(new_n10678_));
  OAI22X1  g08242(.A0(new_n10678_), .A1(new_n3256_), .B0(new_n10541_), .B1(new_n10500_), .Y(new_n10679_));
  OR2X1    g08243(.A(new_n10679_), .B(new_n2972_), .Y(new_n10680_));
  OR4X1    g08244(.A(new_n10483_), .B(pi0468), .C(pi0332), .D(pi0142), .Y(new_n10681_));
  NAND3X1  g08245(.A(new_n10681_), .B(new_n10680_), .C(new_n7548_), .Y(new_n10682_));
  NAND3X1  g08246(.A(new_n10682_), .B(new_n10677_), .C(pi0180), .Y(new_n10683_));
  AND2X1   g08247(.A(new_n10453_), .B(new_n10450_), .Y(new_n10684_));
  AOI21X1  g08248(.A0(new_n10684_), .A1(new_n5225_), .B0(pi0179), .Y(new_n10685_));
  AOI22X1  g08249(.A0(new_n10685_), .A1(new_n10683_), .B0(new_n10676_), .B1(new_n10672_), .Y(new_n10686_));
  OAI21X1  g08250(.A0(new_n10686_), .A1(pi0299), .B0(new_n2959_), .Y(new_n10687_));
  OAI21X1  g08251(.A0(new_n3003_), .A1(new_n2555_), .B0(pi0142), .Y(new_n10688_));
  NOR2X1   g08252(.A(new_n10588_), .B(pi0142), .Y(new_n10689_));
  NAND4X1  g08253(.A(new_n10594_), .B(pi0224), .C(new_n2964_), .D(pi0222), .Y(new_n10690_));
  NOR2X1   g08254(.A(new_n10690_), .B(new_n10689_), .Y(new_n10691_));
  AOI21X1  g08255(.A0(new_n10691_), .A1(new_n10688_), .B0(new_n10450_), .Y(new_n10692_));
  OR2X1    g08256(.A(new_n10453_), .B(pi0144), .Y(new_n10693_));
  OAI21X1  g08257(.A0(new_n10693_), .A1(new_n10607_), .B0(pi0181), .Y(new_n10694_));
  AOI21X1  g08258(.A0(new_n10684_), .A1(new_n5226_), .B0(pi0299), .Y(new_n10695_));
  OAI21X1  g08259(.A0(new_n10694_), .A1(new_n10692_), .B0(new_n10695_), .Y(new_n10696_));
  NOR4X1   g08260(.A(new_n5057_), .B(new_n3003_), .C(new_n2555_), .D(pi0287), .Y(new_n10697_));
  INVX1    g08261(.A(new_n10605_), .Y(new_n10698_));
  AOI21X1  g08262(.A0(new_n10698_), .A1(new_n10552_), .B0(new_n6905_), .Y(new_n10699_));
  OAI21X1  g08263(.A0(new_n10697_), .A1(new_n10663_), .B0(new_n10699_), .Y(new_n10700_));
  AOI21X1  g08264(.A0(new_n10444_), .A1(new_n6905_), .B0(new_n7458_), .Y(new_n10701_));
  NOR3X1   g08265(.A(new_n10444_), .B(new_n2953_), .C(pi0159), .Y(new_n10702_));
  OR2X1    g08266(.A(new_n10702_), .B(new_n7892_), .Y(new_n10703_));
  AOI21X1  g08267(.A0(new_n10701_), .A1(new_n10700_), .B0(new_n10703_), .Y(new_n10704_));
  AOI21X1  g08268(.A0(new_n10704_), .A1(new_n10696_), .B0(pi0038), .Y(new_n10705_));
  OAI21X1  g08269(.A0(new_n10687_), .A1(new_n10666_), .B0(new_n10705_), .Y(new_n10706_));
  INVX1    g08270(.A(new_n10458_), .Y(new_n10707_));
  INVX1    g08271(.A(new_n10501_), .Y(new_n10708_));
  NOR2X1   g08272(.A(new_n10679_), .B(new_n2800_), .Y(new_n10709_));
  NOR3X1   g08273(.A(new_n10483_), .B(new_n5057_), .C(pi0146), .Y(new_n10710_));
  NOR3X1   g08274(.A(new_n10710_), .B(new_n10709_), .C(pi0161), .Y(new_n10711_));
  AOI21X1  g08275(.A0(new_n10708_), .A1(new_n10442_), .B0(new_n10711_), .Y(new_n10712_));
  NOR3X1   g08276(.A(new_n10444_), .B(new_n2953_), .C(pi0158), .Y(new_n10713_));
  NOR2X1   g08277(.A(new_n10713_), .B(new_n5237_), .Y(new_n10714_));
  OAI21X1  g08278(.A0(new_n10712_), .A1(new_n10551_), .B0(new_n10714_), .Y(new_n10715_));
  NOR3X1   g08279(.A(pi0156), .B(pi0039), .C(pi0038), .Y(new_n10716_));
  AOI21X1  g08280(.A0(new_n10716_), .A1(new_n10715_), .B0(new_n10707_), .Y(new_n10717_));
  OAI21X1  g08281(.A0(new_n10457_), .A1(new_n3026_), .B0(new_n5821_), .Y(new_n10718_));
  AOI21X1  g08282(.A0(new_n10717_), .A1(new_n10706_), .B0(new_n10718_), .Y(new_n10719_));
  INVX1    g08283(.A(new_n10645_), .Y(new_n10720_));
  NAND2X1  g08284(.A(new_n10648_), .B(pi0087), .Y(new_n10721_));
  AND2X1   g08285(.A(new_n10721_), .B(new_n10436_), .Y(new_n10722_));
  OAI21X1  g08286(.A0(new_n10720_), .A1(new_n10456_), .B0(new_n10722_), .Y(new_n10723_));
  OAI21X1  g08287(.A0(new_n10723_), .A1(new_n10719_), .B0(new_n6520_), .Y(new_n10724_));
  OAI21X1  g08288(.A0(new_n10724_), .A1(new_n10651_), .B0(new_n10447_), .Y(po0279));
  OAI21X1  g08289(.A0(new_n10418_), .A1(new_n6309_), .B0(new_n10169_), .Y(new_n10726_));
  OAI21X1  g08290(.A0(new_n10423_), .A1(new_n6309_), .B0(new_n6077_), .Y(new_n10727_));
  NAND3X1  g08291(.A(new_n10727_), .B(new_n10726_), .C(new_n6520_), .Y(new_n10728_));
  OAI21X1  g08292(.A0(new_n6746_), .A1(new_n10212_), .B0(new_n10728_), .Y(po0280));
  NAND4X1  g08293(.A(new_n6882_), .B(new_n5241_), .C(new_n8515_), .D(new_n2482_), .Y(new_n10730_));
  NOR4X1   g08294(.A(new_n8240_), .B(new_n7609_), .C(new_n5094_), .D(new_n2482_), .Y(new_n10731_));
  OAI21X1  g08295(.A0(new_n10731_), .A1(pi0039), .B0(po1038), .Y(new_n10732_));
  AOI21X1  g08296(.A0(new_n10730_), .A1(pi0039), .B0(new_n10732_), .Y(new_n10733_));
  NOR4X1   g08297(.A(new_n3125_), .B(pi0100), .C(pi0087), .D(pi0038), .Y(new_n10734_));
  NOR2X1   g08298(.A(new_n10730_), .B(new_n2953_), .Y(new_n10735_));
  NAND3X1  g08299(.A(new_n2953_), .B(new_n2964_), .C(pi0222), .Y(new_n10736_));
  NOR4X1   g08300(.A(new_n6883_), .B(new_n10736_), .C(new_n5058_), .D(pi0110), .Y(new_n10737_));
  NOR3X1   g08301(.A(new_n10737_), .B(new_n10735_), .C(new_n2959_), .Y(new_n10738_));
  NOR3X1   g08302(.A(new_n7842_), .B(new_n2480_), .C(pi0109), .Y(new_n10739_));
  INVX1    g08303(.A(new_n5158_), .Y(new_n10740_));
  INVX1    g08304(.A(new_n2464_), .Y(new_n10741_));
  NOR2X1   g08305(.A(new_n2651_), .B(pi0036), .Y(new_n10742_));
  OAI21X1  g08306(.A0(new_n5150_), .A1(pi0111), .B0(new_n10742_), .Y(new_n10743_));
  OAI21X1  g08307(.A0(new_n2612_), .A1(new_n7658_), .B0(new_n2659_), .Y(new_n10744_));
  AOI21X1  g08308(.A0(new_n10743_), .A1(new_n10741_), .B0(new_n10744_), .Y(new_n10745_));
  OAI21X1  g08309(.A0(new_n10745_), .A1(pi0083), .B0(new_n9533_), .Y(new_n10746_));
  AOI21X1  g08310(.A0(new_n10746_), .A1(new_n2663_), .B0(new_n10740_), .Y(new_n10747_));
  OAI21X1  g08311(.A0(new_n10747_), .A1(pi0081), .B0(new_n8542_), .Y(new_n10748_));
  AOI21X1  g08312(.A0(new_n10748_), .A1(new_n2701_), .B0(new_n2485_), .Y(new_n10749_));
  NOR2X1   g08313(.A(new_n10739_), .B(new_n2701_), .Y(new_n10750_));
  NOR2X1   g08314(.A(new_n10750_), .B(new_n6971_), .Y(new_n10751_));
  NOR4X1   g08315(.A(new_n2485_), .B(pi0093), .C(pi0090), .D(new_n2548_), .Y(new_n10752_));
  AOI22X1  g08316(.A0(new_n10752_), .A1(new_n10739_), .B0(new_n10751_), .B1(new_n10749_), .Y(new_n10753_));
  OAI21X1  g08317(.A0(new_n10753_), .A1(new_n7666_), .B0(new_n2482_), .Y(new_n10754_));
  NOR2X1   g08318(.A(new_n2702_), .B(pi0093), .Y(new_n10755_));
  AOI21X1  g08319(.A0(new_n10749_), .A1(new_n10755_), .B0(pi0072), .Y(new_n10756_));
  OR2X1    g08320(.A(new_n9800_), .B(new_n5191_), .Y(new_n10757_));
  OAI21X1  g08321(.A0(new_n10757_), .A1(new_n10756_), .B0(new_n2959_), .Y(new_n10758_));
  AOI21X1  g08322(.A0(new_n10754_), .A1(new_n9800_), .B0(new_n10758_), .Y(new_n10759_));
  OAI21X1  g08323(.A0(new_n10759_), .A1(new_n10738_), .B0(new_n10734_), .Y(new_n10760_));
  INVX1    g08324(.A(new_n10734_), .Y(new_n10761_));
  AOI21X1  g08325(.A0(new_n9800_), .A1(pi0110), .B0(pi0039), .Y(new_n10762_));
  OAI21X1  g08326(.A0(new_n10762_), .A1(new_n10738_), .B0(new_n10761_), .Y(new_n10763_));
  AND2X1   g08327(.A(new_n10763_), .B(new_n6520_), .Y(new_n10764_));
  AOI21X1  g08328(.A0(new_n10764_), .A1(new_n10760_), .B0(new_n10733_), .Y(po0281));
  INVX1    g08329(.A(pi0125), .Y(new_n10766_));
  XOR2X1   g08330(.A(pi0133), .B(pi0125), .Y(new_n10767_));
  AOI21X1  g08331(.A0(new_n10432_), .A1(new_n10766_), .B0(new_n10767_), .Y(new_n10768_));
  INVX1    g08332(.A(new_n10768_), .Y(new_n10769_));
  AOI22X1  g08333(.A0(new_n10541_), .A1(new_n6900_), .B0(new_n10490_), .B1(pi0172), .Y(new_n10770_));
  INVX1    g08334(.A(new_n10770_), .Y(new_n10771_));
  AOI22X1  g08335(.A0(new_n10771_), .A1(pi0232), .B0(new_n10769_), .B1(new_n10440_), .Y(new_n10772_));
  NOR4X1   g08336(.A(pi0468), .B(pi0332), .C(new_n5237_), .D(new_n3156_), .Y(new_n10773_));
  AOI21X1  g08337(.A0(new_n10773_), .A1(pi0162), .B0(new_n6520_), .Y(new_n10774_));
  OAI21X1  g08338(.A0(new_n10772_), .A1(pi0087), .B0(new_n10774_), .Y(new_n10775_));
  INVX1    g08339(.A(new_n10491_), .Y(new_n10776_));
  NOR3X1   g08340(.A(pi0468), .B(pi0332), .C(pi0152), .Y(new_n10777_));
  AOI21X1  g08341(.A0(new_n10554_), .A1(new_n6900_), .B0(pi0197), .Y(new_n10778_));
  OAI21X1  g08342(.A0(new_n10777_), .A1(new_n10776_), .B0(new_n10778_), .Y(new_n10779_));
  INVX1    g08343(.A(new_n10482_), .Y(new_n10780_));
  AND2X1   g08344(.A(new_n10491_), .B(new_n5057_), .Y(new_n10781_));
  INVX1    g08345(.A(new_n10781_), .Y(new_n10782_));
  AOI22X1  g08346(.A0(new_n10782_), .A1(new_n10536_), .B0(new_n10561_), .B1(new_n10780_), .Y(new_n10783_));
  OR2X1    g08347(.A(new_n7347_), .B(pi0152), .Y(new_n10784_));
  OR2X1    g08348(.A(new_n10784_), .B(new_n10783_), .Y(new_n10785_));
  AOI22X1  g08349(.A0(new_n10785_), .A1(new_n10779_), .B0(new_n10490_), .B1(pi0172), .Y(new_n10786_));
  AOI21X1  g08350(.A0(new_n8218_), .A1(pi0072), .B0(new_n5033_), .Y(new_n10787_));
  AOI21X1  g08351(.A0(new_n10503_), .A1(new_n5033_), .B0(new_n10787_), .Y(new_n10788_));
  NOR3X1   g08352(.A(new_n10501_), .B(new_n10491_), .C(new_n10490_), .Y(new_n10789_));
  AND2X1   g08353(.A(pi0197), .B(pi0152), .Y(new_n10790_));
  OAI21X1  g08354(.A0(new_n10789_), .A1(new_n3601_), .B0(new_n10790_), .Y(new_n10791_));
  AOI21X1  g08355(.A0(new_n10788_), .A1(new_n3601_), .B0(new_n10791_), .Y(new_n10792_));
  OAI21X1  g08356(.A0(new_n10792_), .A1(new_n10786_), .B0(new_n7477_), .Y(new_n10793_));
  NOR2X1   g08357(.A(new_n10787_), .B(new_n10521_), .Y(new_n10794_));
  NOR2X1   g08358(.A(new_n10516_), .B(new_n10491_), .Y(new_n10795_));
  NOR2X1   g08359(.A(new_n10787_), .B(new_n10795_), .Y(new_n10796_));
  INVX1    g08360(.A(new_n10796_), .Y(new_n10797_));
  OAI21X1  g08361(.A0(new_n10797_), .A1(new_n3601_), .B0(pi0152), .Y(new_n10798_));
  AOI21X1  g08362(.A0(new_n10794_), .A1(new_n3601_), .B0(new_n10798_), .Y(new_n10799_));
  AOI22X1  g08363(.A0(new_n10782_), .A1(new_n10536_), .B0(new_n10488_), .B1(new_n5033_), .Y(new_n10800_));
  AOI21X1  g08364(.A0(new_n10490_), .A1(pi0172), .B0(pi0152), .Y(new_n10801_));
  INVX1    g08365(.A(new_n10801_), .Y(new_n10802_));
  OAI21X1  g08366(.A0(new_n10802_), .A1(new_n10800_), .B0(pi0197), .Y(new_n10803_));
  AOI21X1  g08367(.A0(new_n10527_), .A1(new_n5033_), .B0(new_n10787_), .Y(new_n10804_));
  INVX1    g08368(.A(new_n10804_), .Y(new_n10805_));
  NOR2X1   g08369(.A(new_n10781_), .B(new_n10537_), .Y(new_n10806_));
  INVX1    g08370(.A(new_n10806_), .Y(new_n10807_));
  AOI21X1  g08371(.A0(new_n10807_), .A1(new_n6900_), .B0(pi0172), .Y(new_n10808_));
  OAI21X1  g08372(.A0(new_n10805_), .A1(new_n6900_), .B0(new_n10808_), .Y(new_n10809_));
  OAI21X1  g08373(.A0(new_n10531_), .A1(new_n10492_), .B0(pi0152), .Y(new_n10810_));
  INVX1    g08374(.A(new_n10561_), .Y(new_n10811_));
  NOR4X1   g08375(.A(new_n10811_), .B(new_n10479_), .C(new_n10468_), .D(new_n10459_), .Y(new_n10812_));
  NOR2X1   g08376(.A(new_n10812_), .B(new_n10787_), .Y(new_n10813_));
  AOI21X1  g08377(.A0(new_n10813_), .A1(new_n6900_), .B0(new_n3601_), .Y(new_n10814_));
  AOI21X1  g08378(.A0(new_n10814_), .A1(new_n10810_), .B0(pi0197), .Y(new_n10815_));
  AOI21X1  g08379(.A0(new_n10815_), .A1(new_n10809_), .B0(new_n7482_), .Y(new_n10816_));
  OAI21X1  g08380(.A0(new_n10803_), .A1(new_n10799_), .B0(new_n10816_), .Y(new_n10817_));
  AOI21X1  g08381(.A0(new_n10817_), .A1(new_n10793_), .B0(new_n2953_), .Y(new_n10818_));
  NAND2X1  g08382(.A(new_n10788_), .B(pi0145), .Y(new_n10819_));
  AOI21X1  g08383(.A0(new_n10491_), .A1(new_n5224_), .B0(new_n7008_), .Y(new_n10820_));
  NAND2X1  g08384(.A(new_n10783_), .B(pi0145), .Y(new_n10821_));
  AOI21X1  g08385(.A0(new_n10491_), .A1(new_n5057_), .B0(new_n10554_), .Y(new_n10822_));
  INVX1    g08386(.A(new_n10822_), .Y(new_n10823_));
  AOI21X1  g08387(.A0(new_n10823_), .A1(new_n5224_), .B0(pi0174), .Y(new_n10824_));
  AOI22X1  g08388(.A0(new_n10824_), .A1(new_n10821_), .B0(new_n10820_), .B1(new_n10819_), .Y(new_n10825_));
  MX2X1    g08389(.A(new_n10560_), .B(new_n5224_), .S0(new_n10501_), .Y(new_n10826_));
  AOI21X1  g08390(.A0(new_n10826_), .A1(new_n10776_), .B0(new_n7008_), .Y(new_n10827_));
  AOI21X1  g08391(.A0(new_n10780_), .A1(new_n10560_), .B0(new_n5224_), .Y(new_n10828_));
  OAI21X1  g08392(.A0(new_n10828_), .A1(new_n10811_), .B0(new_n7008_), .Y(new_n10829_));
  OAI21X1  g08393(.A0(new_n10829_), .A1(new_n10787_), .B0(pi0193), .Y(new_n10830_));
  OAI22X1  g08394(.A0(new_n10830_), .A1(new_n10827_), .B0(new_n10825_), .B1(pi0193), .Y(new_n10831_));
  NAND2X1  g08395(.A(new_n10831_), .B(new_n7464_), .Y(new_n10832_));
  OAI21X1  g08396(.A0(new_n10805_), .A1(pi0145), .B0(new_n7083_), .Y(new_n10833_));
  AOI21X1  g08397(.A0(new_n10794_), .A1(pi0145), .B0(new_n10833_), .Y(new_n10834_));
  NOR3X1   g08398(.A(new_n10787_), .B(new_n10795_), .C(new_n5224_), .Y(new_n10835_));
  NOR2X1   g08399(.A(new_n10531_), .B(new_n10492_), .Y(new_n10836_));
  OAI21X1  g08400(.A0(new_n10836_), .A1(pi0145), .B0(pi0193), .Y(new_n10837_));
  OAI21X1  g08401(.A0(new_n10837_), .A1(new_n10835_), .B0(pi0174), .Y(new_n10838_));
  NAND2X1  g08402(.A(new_n10813_), .B(pi0193), .Y(new_n10839_));
  OAI21X1  g08403(.A0(new_n10781_), .A1(new_n10537_), .B0(new_n7083_), .Y(new_n10840_));
  NAND3X1  g08404(.A(new_n10840_), .B(new_n10839_), .C(new_n5224_), .Y(new_n10841_));
  NOR4X1   g08405(.A(pi0468), .B(pi0332), .C(new_n7083_), .D(new_n2516_), .Y(new_n10842_));
  NOR3X1   g08406(.A(new_n10842_), .B(new_n10800_), .C(new_n5224_), .Y(new_n10843_));
  NOR2X1   g08407(.A(new_n10843_), .B(pi0174), .Y(new_n10844_));
  AOI21X1  g08408(.A0(new_n10844_), .A1(new_n10841_), .B0(new_n7565_), .Y(new_n10845_));
  OAI21X1  g08409(.A0(new_n10838_), .A1(new_n10834_), .B0(new_n10845_), .Y(new_n10846_));
  AOI21X1  g08410(.A0(new_n10846_), .A1(new_n10832_), .B0(pi0038), .Y(new_n10847_));
  OAI21X1  g08411(.A0(new_n10847_), .A1(new_n10818_), .B0(new_n7299_), .Y(new_n10848_));
  MX2X1    g08412(.A(new_n6283_), .B(new_n6277_), .S0(new_n2953_), .Y(new_n10849_));
  AOI21X1  g08413(.A0(new_n10849_), .A1(new_n3630_), .B0(pi0232), .Y(new_n10850_));
  NOR2X1   g08414(.A(new_n10850_), .B(new_n2959_), .Y(new_n10851_));
  MX2X1    g08415(.A(new_n10583_), .B(new_n3074_), .S0(new_n5057_), .Y(new_n10852_));
  MX2X1    g08416(.A(new_n10589_), .B(new_n3074_), .S0(new_n5057_), .Y(new_n10853_));
  MX2X1    g08417(.A(new_n10853_), .B(new_n10852_), .S0(new_n6900_), .Y(new_n10854_));
  AND2X1   g08418(.A(new_n3601_), .B(pi0051), .Y(new_n10855_));
  OAI21X1  g08419(.A0(new_n10855_), .A1(new_n10854_), .B0(new_n2438_), .Y(new_n10856_));
  OAI22X1  g08420(.A0(new_n10856_), .A1(new_n5242_), .B0(new_n10771_), .B1(new_n6283_), .Y(new_n10857_));
  AND2X1   g08421(.A(new_n10857_), .B(new_n7139_), .Y(new_n10858_));
  INVX1    g08422(.A(new_n10587_), .Y(new_n10859_));
  NOR3X1   g08423(.A(new_n10602_), .B(new_n5911_), .C(new_n2555_), .Y(new_n10860_));
  NOR2X1   g08424(.A(new_n10860_), .B(new_n10490_), .Y(new_n10861_));
  AOI21X1  g08425(.A0(new_n10861_), .A1(pi0224), .B0(new_n10859_), .Y(new_n10862_));
  INVX1    g08426(.A(new_n10862_), .Y(new_n10863_));
  AND2X1   g08427(.A(new_n10853_), .B(new_n6277_), .Y(new_n10864_));
  OAI21X1  g08428(.A0(new_n10864_), .A1(new_n10863_), .B0(new_n10560_), .Y(new_n10865_));
  AND2X1   g08429(.A(new_n10865_), .B(pi0174), .Y(new_n10866_));
  AOI21X1  g08430(.A0(new_n10594_), .A1(new_n10582_), .B0(new_n2961_), .Y(new_n10867_));
  OR2X1    g08431(.A(new_n10867_), .B(new_n10859_), .Y(new_n10868_));
  AOI22X1  g08432(.A0(new_n10868_), .A1(new_n10452_), .B0(new_n10852_), .B1(new_n6277_), .Y(new_n10869_));
  INVX1    g08433(.A(new_n10869_), .Y(new_n10870_));
  OAI21X1  g08434(.A0(new_n10870_), .A1(pi0174), .B0(pi0193), .Y(new_n10871_));
  OR2X1    g08435(.A(new_n10871_), .B(new_n10866_), .Y(new_n10872_));
  MX2X1    g08436(.A(new_n10604_), .B(new_n3074_), .S0(new_n5057_), .Y(new_n10873_));
  NAND2X1  g08437(.A(new_n10873_), .B(new_n2961_), .Y(new_n10874_));
  AOI21X1  g08438(.A0(new_n10698_), .A1(pi0224), .B0(new_n10859_), .Y(new_n10875_));
  AOI22X1  g08439(.A0(new_n10875_), .A1(new_n10874_), .B0(new_n10541_), .B1(new_n10859_), .Y(new_n10876_));
  AOI21X1  g08440(.A0(new_n10690_), .A1(new_n6278_), .B0(new_n3074_), .Y(new_n10877_));
  AOI21X1  g08441(.A0(new_n10877_), .A1(pi0174), .B0(pi0193), .Y(new_n10878_));
  OAI21X1  g08442(.A0(new_n10876_), .A1(pi0174), .B0(new_n10878_), .Y(new_n10879_));
  AND2X1   g08443(.A(new_n10879_), .B(pi0180), .Y(new_n10880_));
  AOI21X1  g08444(.A0(new_n10452_), .A1(new_n6278_), .B0(new_n10873_), .Y(new_n10881_));
  NOR3X1   g08445(.A(new_n6278_), .B(new_n3003_), .C(new_n2555_), .Y(new_n10882_));
  INVX1    g08446(.A(new_n10882_), .Y(new_n10883_));
  OAI22X1  g08447(.A0(new_n10883_), .A1(new_n7008_), .B0(new_n10560_), .B1(new_n7083_), .Y(new_n10884_));
  AOI21X1  g08448(.A0(new_n10881_), .A1(new_n7008_), .B0(new_n10884_), .Y(new_n10885_));
  OAI21X1  g08449(.A0(new_n10885_), .A1(pi0180), .B0(new_n2953_), .Y(new_n10886_));
  AOI21X1  g08450(.A0(new_n10880_), .A1(new_n10872_), .B0(new_n10886_), .Y(new_n10887_));
  INVX1    g08451(.A(new_n10861_), .Y(new_n10888_));
  AOI21X1  g08452(.A0(new_n10594_), .A1(new_n10582_), .B0(new_n10451_), .Y(new_n10889_));
  AOI21X1  g08453(.A0(new_n10889_), .A1(new_n6900_), .B0(new_n3601_), .Y(new_n10890_));
  OAI21X1  g08454(.A0(new_n10888_), .A1(new_n6900_), .B0(new_n10890_), .Y(new_n10891_));
  OR2X1    g08455(.A(new_n10697_), .B(new_n6900_), .Y(new_n10892_));
  AOI21X1  g08456(.A0(new_n10698_), .A1(new_n6900_), .B0(pi0172), .Y(new_n10893_));
  AOI21X1  g08457(.A0(new_n10893_), .A1(new_n10892_), .B0(new_n2438_), .Y(new_n10894_));
  AOI21X1  g08458(.A0(new_n10894_), .A1(new_n10891_), .B0(new_n5242_), .Y(new_n10895_));
  OAI21X1  g08459(.A0(new_n10770_), .A1(new_n5241_), .B0(new_n7107_), .Y(new_n10896_));
  AOI21X1  g08460(.A0(new_n10895_), .A1(new_n10856_), .B0(new_n10896_), .Y(new_n10897_));
  NOR3X1   g08461(.A(new_n10897_), .B(new_n10887_), .C(new_n10858_), .Y(new_n10898_));
  OAI21X1  g08462(.A0(new_n10898_), .A1(new_n5237_), .B0(new_n10851_), .Y(new_n10899_));
  AOI21X1  g08463(.A0(new_n10776_), .A1(new_n5237_), .B0(pi0039), .Y(new_n10900_));
  NOR2X1   g08464(.A(new_n10900_), .B(pi0038), .Y(new_n10901_));
  NAND2X1  g08465(.A(new_n10901_), .B(new_n10899_), .Y(new_n10902_));
  AND2X1   g08466(.A(new_n10770_), .B(pi0299), .Y(new_n10903_));
  AND2X1   g08467(.A(new_n10541_), .B(new_n7008_), .Y(new_n10904_));
  OR2X1    g08468(.A(new_n10842_), .B(pi0299), .Y(new_n10905_));
  OAI21X1  g08469(.A0(new_n10905_), .A1(new_n10904_), .B0(pi0232), .Y(new_n10906_));
  NOR2X1   g08470(.A(new_n10906_), .B(new_n10903_), .Y(new_n10907_));
  INVX1    g08471(.A(new_n10907_), .Y(new_n10908_));
  AOI21X1  g08472(.A0(new_n10908_), .A1(pi0038), .B0(pi0100), .Y(new_n10909_));
  NAND3X1  g08473(.A(new_n10909_), .B(new_n10902_), .C(new_n10848_), .Y(new_n10910_));
  AOI21X1  g08474(.A0(new_n10907_), .A1(pi0100), .B0(new_n10641_), .Y(new_n10911_));
  MX2X1    g08475(.A(new_n7349_), .B(new_n7398_), .S0(new_n2953_), .Y(new_n10912_));
  OAI21X1  g08476(.A0(new_n10912_), .A1(new_n6855_), .B0(pi0087), .Y(new_n10913_));
  AND2X1   g08477(.A(new_n10913_), .B(new_n10768_), .Y(new_n10914_));
  OAI21X1  g08478(.A0(new_n10907_), .A1(new_n10720_), .B0(new_n10914_), .Y(new_n10915_));
  AOI21X1  g08479(.A0(new_n10911_), .A1(new_n10910_), .B0(new_n10915_), .Y(new_n10916_));
  NOR3X1   g08480(.A(new_n10514_), .B(new_n10530_), .C(new_n2487_), .Y(new_n10917_));
  NOR3X1   g08481(.A(new_n10917_), .B(new_n10506_), .C(pi0145), .Y(new_n10918_));
  OR2X1    g08482(.A(new_n10531_), .B(new_n10506_), .Y(new_n10919_));
  OAI21X1  g08483(.A0(new_n10919_), .A1(new_n5224_), .B0(new_n7008_), .Y(new_n10920_));
  OR2X1    g08484(.A(new_n10659_), .B(new_n10506_), .Y(new_n10921_));
  AOI21X1  g08485(.A0(new_n10482_), .A1(new_n5057_), .B0(new_n10459_), .Y(new_n10922_));
  INVX1    g08486(.A(new_n10922_), .Y(new_n10923_));
  NOR2X1   g08487(.A(new_n10923_), .B(new_n10479_), .Y(new_n10924_));
  INVX1    g08488(.A(new_n10924_), .Y(new_n10925_));
  AOI21X1  g08489(.A0(new_n10484_), .A1(new_n5224_), .B0(new_n10925_), .Y(new_n10926_));
  AOI21X1  g08490(.A0(new_n10926_), .A1(new_n3002_), .B0(new_n7008_), .Y(new_n10927_));
  AOI21X1  g08491(.A0(new_n10927_), .A1(new_n10921_), .B0(new_n7083_), .Y(new_n10928_));
  OAI21X1  g08492(.A0(new_n10920_), .A1(new_n10918_), .B0(new_n10928_), .Y(new_n10929_));
  NOR3X1   g08493(.A(new_n10653_), .B(new_n10506_), .C(pi0145), .Y(new_n10930_));
  NOR4X1   g08494(.A(new_n10531_), .B(new_n10506_), .C(new_n5224_), .D(pi0051), .Y(new_n10931_));
  OR2X1    g08495(.A(new_n10931_), .B(pi0174), .Y(new_n10932_));
  OR2X1    g08496(.A(new_n10926_), .B(new_n7008_), .Y(new_n10933_));
  AND2X1   g08497(.A(new_n10933_), .B(new_n7083_), .Y(new_n10934_));
  OAI21X1  g08498(.A0(new_n10932_), .A1(new_n10930_), .B0(new_n10934_), .Y(new_n10935_));
  NAND3X1  g08499(.A(new_n10935_), .B(new_n10929_), .C(new_n7464_), .Y(new_n10936_));
  MX2X1    g08500(.A(new_n10485_), .B(new_n2516_), .S0(new_n5033_), .Y(new_n10937_));
  NOR4X1   g08501(.A(new_n10530_), .B(new_n10498_), .C(new_n9795_), .D(pi0145), .Y(new_n10938_));
  OAI22X1  g08502(.A0(new_n10938_), .A1(pi0174), .B0(new_n10438_), .B1(new_n5224_), .Y(new_n10939_));
  AOI21X1  g08503(.A0(new_n10479_), .A1(new_n5057_), .B0(new_n10484_), .Y(new_n10940_));
  AOI22X1  g08504(.A0(new_n10940_), .A1(pi0174), .B0(new_n10939_), .B1(new_n10937_), .Y(new_n10941_));
  AND2X1   g08505(.A(pi0174), .B(new_n5224_), .Y(new_n10942_));
  AOI22X1  g08506(.A0(new_n10942_), .A1(new_n10679_), .B0(new_n10601_), .B1(pi0145), .Y(new_n10943_));
  OAI21X1  g08507(.A0(new_n10938_), .A1(pi0174), .B0(new_n10943_), .Y(new_n10944_));
  NOR2X1   g08508(.A(new_n10506_), .B(new_n7083_), .Y(new_n10945_));
  AOI21X1  g08509(.A0(new_n10945_), .A1(new_n10944_), .B0(new_n7565_), .Y(new_n10946_));
  OAI21X1  g08510(.A0(new_n10941_), .A1(pi0193), .B0(new_n10946_), .Y(new_n10947_));
  AOI21X1  g08511(.A0(new_n10947_), .A1(new_n10936_), .B0(pi0038), .Y(new_n10948_));
  NOR2X1   g08512(.A(new_n10917_), .B(new_n10506_), .Y(new_n10949_));
  AOI21X1  g08513(.A0(new_n10921_), .A1(pi0152), .B0(new_n3601_), .Y(new_n10950_));
  OAI21X1  g08514(.A0(new_n10949_), .A1(pi0152), .B0(new_n10950_), .Y(new_n10951_));
  AND2X1   g08515(.A(new_n10653_), .B(new_n6900_), .Y(new_n10952_));
  OAI21X1  g08516(.A0(new_n10777_), .A1(new_n10485_), .B0(new_n3601_), .Y(new_n10953_));
  OAI21X1  g08517(.A0(new_n10953_), .A1(new_n10952_), .B0(new_n10951_), .Y(new_n10954_));
  AND2X1   g08518(.A(new_n10919_), .B(new_n6900_), .Y(new_n10955_));
  OAI21X1  g08519(.A0(new_n10485_), .A1(new_n5033_), .B0(new_n10542_), .Y(new_n10956_));
  NOR2X1   g08520(.A(new_n10956_), .B(new_n3601_), .Y(new_n10957_));
  OAI21X1  g08521(.A0(new_n10925_), .A1(pi0172), .B0(pi0152), .Y(new_n10958_));
  AOI21X1  g08522(.A0(new_n10490_), .A1(new_n3601_), .B0(new_n7347_), .Y(new_n10959_));
  OAI21X1  g08523(.A0(new_n10958_), .A1(new_n10957_), .B0(new_n10959_), .Y(new_n10960_));
  AND2X1   g08524(.A(new_n7477_), .B(pi0299), .Y(new_n10961_));
  OAI21X1  g08525(.A0(new_n10960_), .A1(new_n10955_), .B0(new_n10961_), .Y(new_n10962_));
  AOI21X1  g08526(.A0(new_n10954_), .A1(new_n7347_), .B0(new_n10962_), .Y(new_n10963_));
  OR4X1    g08527(.A(new_n10501_), .B(new_n10506_), .C(new_n10490_), .D(pi0152), .Y(new_n10964_));
  AOI21X1  g08528(.A0(new_n10940_), .A1(pi0152), .B0(pi0172), .Y(new_n10965_));
  AND2X1   g08529(.A(new_n10965_), .B(new_n10964_), .Y(new_n10966_));
  NOR3X1   g08530(.A(new_n10501_), .B(new_n10506_), .C(pi0152), .Y(new_n10967_));
  INVX1    g08531(.A(new_n10679_), .Y(new_n10968_));
  NOR3X1   g08532(.A(new_n10968_), .B(new_n10506_), .C(new_n6900_), .Y(new_n10969_));
  NOR3X1   g08533(.A(new_n10969_), .B(new_n10967_), .C(new_n3601_), .Y(new_n10970_));
  NOR3X1   g08534(.A(new_n10970_), .B(new_n10966_), .C(pi0197), .Y(new_n10971_));
  OAI22X1  g08535(.A0(new_n10601_), .A1(new_n6900_), .B0(new_n10485_), .B1(new_n5033_), .Y(new_n10972_));
  OAI21X1  g08536(.A0(new_n10601_), .A1(pi0152), .B0(new_n3601_), .Y(new_n10973_));
  OAI21X1  g08537(.A0(new_n10973_), .A1(new_n10486_), .B0(pi0197), .Y(new_n10974_));
  AOI21X1  g08538(.A0(new_n10972_), .A1(pi0172), .B0(new_n10974_), .Y(new_n10975_));
  NOR4X1   g08539(.A(new_n10975_), .B(new_n10971_), .C(new_n7482_), .D(new_n2953_), .Y(new_n10976_));
  OR2X1    g08540(.A(new_n10976_), .B(new_n10963_), .Y(new_n10977_));
  OAI21X1  g08541(.A0(new_n10977_), .A1(new_n10948_), .B0(new_n7299_), .Y(new_n10978_));
  NOR2X1   g08542(.A(new_n10909_), .B(new_n10460_), .Y(new_n10979_));
  OAI21X1  g08543(.A0(new_n10771_), .A1(new_n10440_), .B0(new_n6905_), .Y(new_n10980_));
  NOR2X1   g08544(.A(new_n10589_), .B(new_n5057_), .Y(new_n10981_));
  INVX1    g08545(.A(new_n10981_), .Y(new_n10982_));
  OAI22X1  g08546(.A0(new_n10777_), .A1(new_n10583_), .B0(new_n10982_), .B1(pi0152), .Y(new_n10983_));
  OAI21X1  g08547(.A0(new_n10610_), .A1(new_n6900_), .B0(pi0172), .Y(new_n10984_));
  AOI21X1  g08548(.A0(new_n10585_), .A1(new_n6900_), .B0(new_n10984_), .Y(new_n10985_));
  OR2X1    g08549(.A(new_n10985_), .B(new_n6905_), .Y(new_n10986_));
  AOI21X1  g08550(.A0(new_n10983_), .A1(new_n3601_), .B0(new_n10986_), .Y(new_n10987_));
  OAI21X1  g08551(.A0(new_n10560_), .A1(new_n3601_), .B0(pi0152), .Y(new_n10988_));
  OAI21X1  g08552(.A0(new_n10988_), .A1(new_n10624_), .B0(new_n6893_), .Y(new_n10989_));
  AOI21X1  g08553(.A0(new_n10801_), .A1(new_n10595_), .B0(new_n10989_), .Y(new_n10990_));
  OAI22X1  g08554(.A0(new_n10990_), .A1(new_n10551_), .B0(new_n10987_), .B1(new_n7140_), .Y(new_n10991_));
  OAI21X1  g08555(.A0(pi0468), .A1(pi0332), .B0(pi0051), .Y(new_n10992_));
  AOI21X1  g08556(.A0(new_n10438_), .A1(new_n5057_), .B0(new_n6886_), .Y(new_n10993_));
  AOI22X1  g08557(.A0(new_n10993_), .A1(new_n10992_), .B0(new_n10585_), .B1(new_n6886_), .Y(new_n10994_));
  AOI21X1  g08558(.A0(new_n10582_), .A1(new_n6886_), .B0(new_n10459_), .Y(new_n10995_));
  OAI21X1  g08559(.A0(new_n10995_), .A1(new_n10490_), .B0(pi0174), .Y(new_n10996_));
  AND2X1   g08560(.A(new_n10996_), .B(new_n5225_), .Y(new_n10997_));
  OAI21X1  g08561(.A0(new_n10994_), .A1(pi0174), .B0(new_n10997_), .Y(new_n10998_));
  INVX1    g08562(.A(new_n7944_), .Y(new_n10999_));
  AOI21X1  g08563(.A0(new_n10584_), .A1(new_n5057_), .B0(new_n6913_), .Y(new_n11000_));
  AOI22X1  g08564(.A0(new_n11000_), .A1(new_n10999_), .B0(new_n10993_), .B1(new_n10992_), .Y(new_n11001_));
  NOR2X1   g08565(.A(new_n10624_), .B(pi0051), .Y(new_n11002_));
  NOR2X1   g08566(.A(new_n11002_), .B(new_n5057_), .Y(new_n11003_));
  OR2X1    g08567(.A(new_n11003_), .B(new_n10995_), .Y(new_n11004_));
  AOI21X1  g08568(.A0(new_n11004_), .A1(pi0174), .B0(new_n5225_), .Y(new_n11005_));
  OAI21X1  g08569(.A0(new_n11001_), .A1(pi0174), .B0(new_n11005_), .Y(new_n11006_));
  NAND3X1  g08570(.A(new_n11006_), .B(new_n10998_), .C(pi0193), .Y(new_n11007_));
  AOI22X1  g08571(.A0(new_n10993_), .A1(new_n2516_), .B0(new_n10590_), .B1(new_n6886_), .Y(new_n11008_));
  OR4X1    g08572(.A(pi0468), .B(pi0332), .C(pi0287), .D(pi0051), .Y(new_n11009_));
  OR2X1    g08573(.A(new_n11009_), .B(new_n5225_), .Y(new_n11010_));
  NAND3X1  g08574(.A(new_n11010_), .B(new_n11008_), .C(new_n7008_), .Y(new_n11011_));
  NAND2X1  g08575(.A(new_n10624_), .B(pi0180), .Y(new_n11012_));
  NOR2X1   g08576(.A(new_n10995_), .B(new_n7008_), .Y(new_n11013_));
  AOI21X1  g08577(.A0(new_n11013_), .A1(new_n11012_), .B0(pi0193), .Y(new_n11014_));
  AOI21X1  g08578(.A0(new_n11014_), .A1(new_n11011_), .B0(pi0299), .Y(new_n11015_));
  AOI22X1  g08579(.A0(new_n11015_), .A1(new_n11007_), .B0(new_n10991_), .B1(new_n10980_), .Y(new_n11016_));
  AOI21X1  g08580(.A0(new_n10582_), .A1(new_n6893_), .B0(new_n10459_), .Y(new_n11017_));
  MX2X1    g08581(.A(new_n11017_), .B(new_n10995_), .S0(new_n2953_), .Y(new_n11018_));
  NOR2X1   g08582(.A(new_n11018_), .B(pi0232), .Y(new_n11019_));
  NOR2X1   g08583(.A(new_n11019_), .B(new_n2959_), .Y(new_n11020_));
  OAI21X1  g08584(.A0(new_n11016_), .A1(new_n5237_), .B0(new_n11020_), .Y(new_n11021_));
  OAI21X1  g08585(.A0(new_n10485_), .A1(pi0232), .B0(new_n2959_), .Y(new_n11022_));
  AND2X1   g08586(.A(new_n11022_), .B(new_n2996_), .Y(new_n11023_));
  AOI21X1  g08587(.A0(new_n11023_), .A1(new_n11021_), .B0(new_n10979_), .Y(new_n11024_));
  OAI21X1  g08588(.A0(new_n10908_), .A1(new_n3026_), .B0(new_n10642_), .Y(new_n11025_));
  AOI21X1  g08589(.A0(new_n11024_), .A1(new_n10978_), .B0(new_n11025_), .Y(new_n11026_));
  AND2X1   g08590(.A(new_n10913_), .B(new_n10769_), .Y(new_n11027_));
  OAI21X1  g08591(.A0(new_n10907_), .A1(new_n10646_), .B0(new_n11027_), .Y(new_n11028_));
  OAI21X1  g08592(.A0(new_n11028_), .A1(new_n11026_), .B0(new_n6520_), .Y(new_n11029_));
  OAI21X1  g08593(.A0(new_n11029_), .A1(new_n10916_), .B0(new_n10775_), .Y(po0282));
  OAI21X1  g08594(.A0(new_n10797_), .A1(new_n8734_), .B0(pi0157), .Y(new_n11031_));
  AOI21X1  g08595(.A0(new_n10794_), .A1(new_n8734_), .B0(new_n11031_), .Y(new_n11032_));
  OAI21X1  g08596(.A0(new_n10789_), .A1(new_n8734_), .B0(new_n10060_), .Y(new_n11033_));
  AOI21X1  g08597(.A0(new_n10788_), .A1(new_n8734_), .B0(new_n11033_), .Y(new_n11034_));
  OAI21X1  g08598(.A0(new_n11034_), .A1(new_n11032_), .B0(pi0166), .Y(new_n11035_));
  AND2X1   g08599(.A(new_n10800_), .B(pi0157), .Y(new_n11036_));
  AND2X1   g08600(.A(new_n10783_), .B(new_n10060_), .Y(new_n11037_));
  NOR4X1   g08601(.A(pi0468), .B(pi0332), .C(new_n8734_), .D(new_n2516_), .Y(new_n11038_));
  OR4X1    g08602(.A(new_n11038_), .B(new_n11037_), .C(new_n11036_), .D(pi0166), .Y(new_n11039_));
  AOI21X1  g08603(.A0(new_n11039_), .A1(new_n11035_), .B0(new_n7458_), .Y(new_n11040_));
  AND2X1   g08604(.A(new_n10800_), .B(new_n7942_), .Y(new_n11041_));
  NOR3X1   g08605(.A(new_n10787_), .B(new_n10521_), .C(new_n7942_), .Y(new_n11042_));
  OAI21X1  g08606(.A0(new_n11042_), .A1(new_n11041_), .B0(pi0178), .Y(new_n11043_));
  OR2X1    g08607(.A(new_n10783_), .B(pi0189), .Y(new_n11044_));
  OR2X1    g08608(.A(new_n10788_), .B(new_n7942_), .Y(new_n11045_));
  NAND3X1  g08609(.A(new_n11045_), .B(new_n11044_), .C(new_n10020_), .Y(new_n11046_));
  AOI21X1  g08610(.A0(new_n11046_), .A1(new_n11043_), .B0(new_n5226_), .Y(new_n11047_));
  OAI21X1  g08611(.A0(new_n10806_), .A1(pi0189), .B0(pi0178), .Y(new_n11048_));
  AOI21X1  g08612(.A0(new_n10804_), .A1(pi0189), .B0(new_n11048_), .Y(new_n11049_));
  OAI21X1  g08613(.A0(new_n10776_), .A1(new_n7942_), .B0(new_n10020_), .Y(new_n11050_));
  OR2X1    g08614(.A(new_n10822_), .B(pi0189), .Y(new_n11051_));
  NOR2X1   g08615(.A(new_n11050_), .B(new_n10490_), .Y(new_n11052_));
  AOI21X1  g08616(.A0(new_n11052_), .A1(new_n11051_), .B0(pi0181), .Y(new_n11053_));
  OAI21X1  g08617(.A0(new_n11050_), .A1(new_n10823_), .B0(new_n11053_), .Y(new_n11054_));
  OAI21X1  g08618(.A0(new_n11054_), .A1(new_n11049_), .B0(new_n8799_), .Y(new_n11055_));
  OAI21X1  g08619(.A0(new_n10531_), .A1(new_n10492_), .B0(pi0166), .Y(new_n11056_));
  AOI21X1  g08620(.A0(new_n10813_), .A1(new_n4464_), .B0(new_n8734_), .Y(new_n11057_));
  NAND2X1  g08621(.A(new_n10804_), .B(pi0166), .Y(new_n11058_));
  AOI21X1  g08622(.A0(new_n10807_), .A1(new_n4464_), .B0(pi0153), .Y(new_n11059_));
  AOI22X1  g08623(.A0(new_n11059_), .A1(new_n11058_), .B0(new_n11057_), .B1(new_n11056_), .Y(new_n11060_));
  OR2X1    g08624(.A(new_n11038_), .B(pi0157), .Y(new_n11061_));
  AOI21X1  g08625(.A0(new_n10491_), .A1(pi0166), .B0(new_n11061_), .Y(new_n11062_));
  OAI21X1  g08626(.A0(new_n10822_), .A1(pi0166), .B0(new_n11062_), .Y(new_n11063_));
  OAI21X1  g08627(.A0(new_n11060_), .A1(new_n10060_), .B0(new_n11063_), .Y(new_n11064_));
  NAND2X1  g08628(.A(new_n10937_), .B(new_n7942_), .Y(new_n11065_));
  AND2X1   g08629(.A(new_n11065_), .B(new_n10796_), .Y(new_n11066_));
  OR2X1    g08630(.A(new_n11041_), .B(new_n10020_), .Y(new_n11067_));
  OR4X1    g08631(.A(new_n10501_), .B(new_n10491_), .C(new_n10490_), .D(new_n7942_), .Y(new_n11068_));
  OAI21X1  g08632(.A0(new_n11044_), .A1(new_n10490_), .B0(new_n11068_), .Y(new_n11069_));
  AOI21X1  g08633(.A0(new_n11069_), .A1(new_n10020_), .B0(new_n5226_), .Y(new_n11070_));
  OAI21X1  g08634(.A0(new_n11067_), .A1(new_n11066_), .B0(new_n11070_), .Y(new_n11071_));
  AOI21X1  g08635(.A0(new_n10813_), .A1(new_n7942_), .B0(new_n10020_), .Y(new_n11072_));
  OAI21X1  g08636(.A0(new_n10836_), .A1(new_n7942_), .B0(new_n11072_), .Y(new_n11073_));
  AOI21X1  g08637(.A0(new_n11073_), .A1(new_n11053_), .B0(new_n8829_), .Y(new_n11074_));
  AOI22X1  g08638(.A0(new_n11074_), .A1(new_n11071_), .B0(new_n11064_), .B1(new_n7429_), .Y(new_n11075_));
  OAI21X1  g08639(.A0(new_n11055_), .A1(new_n11047_), .B0(new_n11075_), .Y(new_n11076_));
  OAI21X1  g08640(.A0(new_n11076_), .A1(new_n11040_), .B0(pi0232), .Y(new_n11077_));
  INVX1    g08641(.A(new_n10851_), .Y(new_n11078_));
  NOR3X1   g08642(.A(new_n10431_), .B(pi0132), .C(pi0126), .Y(new_n11079_));
  INVX1    g08643(.A(pi0126), .Y(new_n11080_));
  NOR3X1   g08644(.A(pi0133), .B(pi0125), .C(pi0121), .Y(new_n11081_));
  XOR2X1   g08645(.A(new_n11081_), .B(new_n11080_), .Y(new_n11082_));
  NOR2X1   g08646(.A(new_n11082_), .B(new_n11079_), .Y(new_n11083_));
  AND2X1   g08647(.A(new_n10881_), .B(new_n7942_), .Y(new_n11084_));
  OAI21X1  g08648(.A0(new_n10883_), .A1(new_n7942_), .B0(new_n5227_), .Y(new_n11085_));
  NOR3X1   g08649(.A(new_n11085_), .B(new_n11084_), .C(new_n10490_), .Y(new_n11086_));
  OAI21X1  g08650(.A0(new_n10870_), .A1(pi0189), .B0(pi0182), .Y(new_n11087_));
  AOI21X1  g08651(.A0(new_n10865_), .A1(pi0189), .B0(new_n11087_), .Y(new_n11088_));
  OAI21X1  g08652(.A0(new_n11088_), .A1(new_n11086_), .B0(new_n8828_), .Y(new_n11089_));
  INVX1    g08653(.A(new_n10697_), .Y(new_n11090_));
  AOI21X1  g08654(.A0(new_n10605_), .A1(new_n4464_), .B0(pi0153), .Y(new_n11091_));
  OAI21X1  g08655(.A0(new_n11090_), .A1(new_n4464_), .B0(new_n11091_), .Y(new_n11092_));
  OAI21X1  g08656(.A0(new_n10860_), .A1(new_n10490_), .B0(pi0166), .Y(new_n11093_));
  INVX1    g08657(.A(new_n10889_), .Y(new_n11094_));
  AOI21X1  g08658(.A0(new_n11094_), .A1(new_n4464_), .B0(new_n8734_), .Y(new_n11095_));
  AOI21X1  g08659(.A0(new_n11095_), .A1(new_n11093_), .B0(new_n8747_), .Y(new_n11096_));
  AOI21X1  g08660(.A0(new_n11096_), .A1(new_n11092_), .B0(new_n2438_), .Y(new_n11097_));
  INVX1    g08661(.A(new_n10852_), .Y(new_n11098_));
  INVX1    g08662(.A(new_n10853_), .Y(new_n11099_));
  MX2X1    g08663(.A(new_n11099_), .B(new_n11098_), .S0(new_n4464_), .Y(new_n11100_));
  OR2X1    g08664(.A(pi0153), .B(new_n2516_), .Y(new_n11101_));
  AOI21X1  g08665(.A0(new_n11101_), .A1(new_n11100_), .B0(pi0216), .Y(new_n11102_));
  OR4X1    g08666(.A(new_n11102_), .B(new_n11097_), .C(new_n2437_), .D(pi0215), .Y(new_n11103_));
  NOR2X1   g08667(.A(new_n10541_), .B(pi0051), .Y(new_n11104_));
  INVX1    g08668(.A(new_n11104_), .Y(new_n11105_));
  AOI21X1  g08669(.A0(new_n10438_), .A1(new_n7784_), .B0(pi0051), .Y(new_n11106_));
  OR2X1    g08670(.A(new_n11106_), .B(new_n11038_), .Y(new_n11107_));
  AND2X1   g08671(.A(new_n11107_), .B(new_n11105_), .Y(new_n11108_));
  OAI21X1  g08672(.A0(new_n2438_), .A1(pi0160), .B0(new_n5241_), .Y(new_n11109_));
  AOI21X1  g08673(.A0(new_n11109_), .A1(new_n11108_), .B0(new_n2953_), .Y(new_n11110_));
  OR2X1    g08674(.A(new_n11085_), .B(new_n11084_), .Y(new_n11111_));
  AOI21X1  g08675(.A0(new_n10877_), .A1(pi0189), .B0(new_n5227_), .Y(new_n11112_));
  OAI21X1  g08676(.A0(new_n10876_), .A1(pi0189), .B0(new_n11112_), .Y(new_n11113_));
  AOI21X1  g08677(.A0(new_n11113_), .A1(new_n11111_), .B0(new_n8800_), .Y(new_n11114_));
  AOI21X1  g08678(.A0(new_n11110_), .A1(new_n11103_), .B0(new_n11114_), .Y(new_n11115_));
  AOI21X1  g08679(.A0(new_n11115_), .A1(new_n11089_), .B0(new_n5237_), .Y(new_n11116_));
  OAI21X1  g08680(.A0(new_n11116_), .A1(new_n11078_), .B0(new_n11083_), .Y(new_n11117_));
  AOI21X1  g08681(.A0(new_n11077_), .A1(new_n10900_), .B0(new_n11117_), .Y(new_n11118_));
  INVX1    g08682(.A(new_n10485_), .Y(new_n11119_));
  AOI22X1  g08683(.A0(new_n10653_), .A1(new_n7942_), .B0(new_n11119_), .B1(new_n8813_), .Y(new_n11120_));
  NOR2X1   g08684(.A(new_n11120_), .B(pi0178), .Y(new_n11121_));
  AND2X1   g08685(.A(new_n10940_), .B(pi0189), .Y(new_n11122_));
  AOI21X1  g08686(.A0(new_n10937_), .A1(new_n7942_), .B0(new_n10020_), .Y(new_n11123_));
  NOR3X1   g08687(.A(new_n10501_), .B(new_n10506_), .C(pi0189), .Y(new_n11124_));
  NOR2X1   g08688(.A(new_n11124_), .B(new_n10020_), .Y(new_n11125_));
  NOR2X1   g08689(.A(new_n11125_), .B(new_n11123_), .Y(new_n11126_));
  OAI21X1  g08690(.A0(new_n11126_), .A1(new_n11122_), .B0(new_n5226_), .Y(new_n11127_));
  AOI21X1  g08691(.A0(new_n10924_), .A1(pi0189), .B0(pi0178), .Y(new_n11128_));
  OAI21X1  g08692(.A0(new_n11065_), .A1(new_n10531_), .B0(new_n11128_), .Y(new_n11129_));
  NAND2X1  g08693(.A(new_n10486_), .B(pi0189), .Y(new_n11130_));
  AOI21X1  g08694(.A0(new_n11130_), .A1(new_n11123_), .B0(new_n5226_), .Y(new_n11131_));
  AOI21X1  g08695(.A0(new_n11131_), .A1(new_n11129_), .B0(new_n8800_), .Y(new_n11132_));
  OAI21X1  g08696(.A0(new_n11127_), .A1(new_n11121_), .B0(new_n11132_), .Y(new_n11133_));
  OAI21X1  g08697(.A0(new_n10917_), .A1(new_n10506_), .B0(new_n4464_), .Y(new_n11134_));
  AOI21X1  g08698(.A0(new_n10921_), .A1(pi0166), .B0(new_n8734_), .Y(new_n11135_));
  NAND3X1  g08699(.A(new_n10516_), .B(new_n5033_), .C(new_n4464_), .Y(new_n11136_));
  AOI21X1  g08700(.A0(new_n11119_), .A1(new_n7784_), .B0(pi0153), .Y(new_n11137_));
  AOI22X1  g08701(.A0(new_n11137_), .A1(new_n11136_), .B0(new_n11135_), .B1(new_n11134_), .Y(new_n11138_));
  INVX1    g08702(.A(new_n7429_), .Y(new_n11139_));
  OAI21X1  g08703(.A0(new_n10501_), .A1(new_n10506_), .B0(new_n4464_), .Y(new_n11140_));
  OAI22X1  g08704(.A0(new_n10940_), .A1(new_n4464_), .B0(new_n7784_), .B1(new_n2516_), .Y(new_n11141_));
  NOR2X1   g08705(.A(new_n10968_), .B(new_n10506_), .Y(new_n11142_));
  NAND2X1  g08706(.A(pi0166), .B(pi0153), .Y(new_n11143_));
  OAI21X1  g08707(.A0(new_n11143_), .A1(new_n11142_), .B0(pi0157), .Y(new_n11144_));
  AOI21X1  g08708(.A0(new_n11141_), .A1(new_n8734_), .B0(new_n11144_), .Y(new_n11145_));
  AOI21X1  g08709(.A0(new_n11145_), .A1(new_n11140_), .B0(new_n11139_), .Y(new_n11146_));
  OAI21X1  g08710(.A0(new_n11138_), .A1(pi0157), .B0(new_n11146_), .Y(new_n11147_));
  OAI21X1  g08711(.A0(new_n10921_), .A1(new_n7942_), .B0(new_n10020_), .Y(new_n11148_));
  AOI21X1  g08712(.A0(new_n10949_), .A1(new_n7942_), .B0(new_n11148_), .Y(new_n11149_));
  NOR3X1   g08713(.A(new_n10968_), .B(new_n10506_), .C(new_n7942_), .Y(new_n11150_));
  NOR3X1   g08714(.A(new_n11150_), .B(new_n11124_), .C(new_n10020_), .Y(new_n11151_));
  OR2X1    g08715(.A(new_n11151_), .B(pi0181), .Y(new_n11152_));
  AOI21X1  g08716(.A0(new_n10542_), .A1(pi0189), .B0(pi0178), .Y(new_n11153_));
  OAI21X1  g08717(.A0(new_n10531_), .A1(pi0189), .B0(new_n11153_), .Y(new_n11154_));
  NOR2X1   g08718(.A(new_n10437_), .B(pi0051), .Y(new_n11155_));
  INVX1    g08719(.A(new_n11155_), .Y(new_n11156_));
  NOR4X1   g08720(.A(new_n11156_), .B(new_n5057_), .C(new_n7942_), .D(new_n10020_), .Y(new_n11157_));
  NOR3X1   g08721(.A(new_n11157_), .B(new_n10506_), .C(new_n5226_), .Y(new_n11158_));
  AOI21X1  g08722(.A0(new_n11158_), .A1(new_n11154_), .B0(new_n8829_), .Y(new_n11159_));
  OAI21X1  g08723(.A0(new_n11152_), .A1(new_n11149_), .B0(new_n11159_), .Y(new_n11160_));
  AND2X1   g08724(.A(new_n10919_), .B(new_n4464_), .Y(new_n11161_));
  NAND3X1  g08725(.A(new_n10956_), .B(pi0166), .C(pi0153), .Y(new_n11162_));
  OAI22X1  g08726(.A0(new_n10924_), .A1(new_n4464_), .B0(new_n7784_), .B1(new_n2516_), .Y(new_n11163_));
  AOI21X1  g08727(.A0(new_n11163_), .A1(new_n8734_), .B0(pi0157), .Y(new_n11164_));
  NAND2X1  g08728(.A(new_n11164_), .B(new_n11162_), .Y(new_n11165_));
  OAI22X1  g08729(.A0(new_n10601_), .A1(new_n4464_), .B0(new_n10485_), .B1(new_n5033_), .Y(new_n11166_));
  NAND2X1  g08730(.A(new_n11166_), .B(pi0153), .Y(new_n11167_));
  NOR3X1   g08731(.A(new_n11108_), .B(new_n10486_), .C(pi0153), .Y(new_n11168_));
  NOR2X1   g08732(.A(new_n11168_), .B(new_n10060_), .Y(new_n11169_));
  AOI21X1  g08733(.A0(new_n11169_), .A1(new_n11167_), .B0(new_n7458_), .Y(new_n11170_));
  OAI21X1  g08734(.A0(new_n11165_), .A1(new_n11161_), .B0(new_n11170_), .Y(new_n11171_));
  NAND4X1  g08735(.A(new_n11171_), .B(new_n11160_), .C(new_n11147_), .D(new_n11133_), .Y(new_n11172_));
  AOI21X1  g08736(.A0(new_n11172_), .A1(pi0232), .B0(new_n11022_), .Y(new_n11173_));
  INVX1    g08737(.A(new_n11020_), .Y(new_n11174_));
  INVX1    g08738(.A(new_n11083_), .Y(new_n11175_));
  MX2X1    g08739(.A(new_n10625_), .B(new_n10595_), .S0(new_n4464_), .Y(new_n11176_));
  NOR2X1   g08740(.A(new_n11038_), .B(new_n8747_), .Y(new_n11177_));
  AND2X1   g08741(.A(new_n11177_), .B(new_n11176_), .Y(new_n11178_));
  OAI22X1  g08742(.A0(new_n10982_), .A1(pi0166), .B0(new_n10583_), .B1(new_n7783_), .Y(new_n11179_));
  OAI21X1  g08743(.A0(new_n10610_), .A1(new_n4464_), .B0(pi0153), .Y(new_n11180_));
  AOI21X1  g08744(.A0(new_n10585_), .A1(new_n4464_), .B0(new_n11180_), .Y(new_n11181_));
  AOI21X1  g08745(.A0(new_n11179_), .A1(new_n8734_), .B0(new_n11181_), .Y(new_n11182_));
  OAI21X1  g08746(.A0(new_n11182_), .A1(pi0160), .B0(new_n6893_), .Y(new_n11183_));
  AOI21X1  g08747(.A0(new_n11107_), .A1(new_n6905_), .B0(new_n2953_), .Y(new_n11184_));
  OAI21X1  g08748(.A0(new_n11183_), .A1(new_n11178_), .B0(new_n11184_), .Y(new_n11185_));
  INVX1    g08749(.A(new_n11008_), .Y(new_n11186_));
  NOR2X1   g08750(.A(new_n10995_), .B(new_n7942_), .Y(new_n11187_));
  OAI21X1  g08751(.A0(new_n10625_), .A1(new_n5227_), .B0(new_n11187_), .Y(new_n11188_));
  OAI21X1  g08752(.A0(new_n11009_), .A1(new_n5227_), .B0(new_n7942_), .Y(new_n11189_));
  OAI21X1  g08753(.A0(new_n11189_), .A1(new_n11186_), .B0(new_n11188_), .Y(new_n11190_));
  NOR2X1   g08754(.A(new_n10994_), .B(pi0189), .Y(new_n11191_));
  OAI21X1  g08755(.A0(new_n10995_), .A1(new_n10490_), .B0(pi0189), .Y(new_n11192_));
  NAND2X1  g08756(.A(new_n11192_), .B(new_n5227_), .Y(new_n11193_));
  AOI21X1  g08757(.A0(new_n11004_), .A1(pi0189), .B0(new_n5227_), .Y(new_n11194_));
  OAI21X1  g08758(.A0(new_n11001_), .A1(pi0189), .B0(new_n11194_), .Y(new_n11195_));
  OAI21X1  g08759(.A0(new_n11193_), .A1(new_n11191_), .B0(new_n11195_), .Y(new_n11196_));
  AOI22X1  g08760(.A0(new_n11196_), .A1(new_n8828_), .B0(new_n11190_), .B1(new_n8799_), .Y(new_n11197_));
  AOI21X1  g08761(.A0(new_n11197_), .A1(new_n11185_), .B0(new_n5237_), .Y(new_n11198_));
  OAI21X1  g08762(.A0(new_n11198_), .A1(new_n11174_), .B0(new_n11175_), .Y(new_n11199_));
  OAI21X1  g08763(.A0(new_n11199_), .A1(new_n11173_), .B0(new_n3277_), .Y(new_n11200_));
  AOI21X1  g08764(.A0(new_n11107_), .A1(new_n11105_), .B0(new_n2953_), .Y(new_n11201_));
  AND2X1   g08765(.A(new_n10541_), .B(new_n7942_), .Y(new_n11202_));
  INVX1    g08766(.A(pi0175), .Y(new_n11203_));
  OAI21X1  g08767(.A0(new_n10560_), .A1(new_n11203_), .B0(new_n2953_), .Y(new_n11204_));
  OAI21X1  g08768(.A0(new_n11204_), .A1(new_n11202_), .B0(pi0232), .Y(new_n11205_));
  NOR2X1   g08769(.A(new_n11205_), .B(new_n11201_), .Y(new_n11206_));
  AND2X1   g08770(.A(new_n10440_), .B(new_n5792_), .Y(new_n11207_));
  INVX1    g08771(.A(new_n11207_), .Y(new_n11208_));
  OAI21X1  g08772(.A0(new_n11208_), .A1(new_n11083_), .B0(new_n5821_), .Y(new_n11209_));
  AOI21X1  g08773(.A0(new_n11206_), .A1(new_n5792_), .B0(new_n11209_), .Y(new_n11210_));
  OAI21X1  g08774(.A0(new_n11200_), .A1(new_n11118_), .B0(new_n11210_), .Y(new_n11211_));
  MX2X1    g08775(.A(pi0185), .B(pi0150), .S0(pi0299), .Y(new_n11212_));
  AND2X1   g08776(.A(new_n11212_), .B(new_n5930_), .Y(new_n11213_));
  OAI22X1  g08777(.A0(new_n11213_), .A1(new_n3156_), .B0(new_n11206_), .B1(new_n10720_), .Y(new_n11214_));
  AND2X1   g08778(.A(new_n10440_), .B(new_n3156_), .Y(new_n11215_));
  OAI21X1  g08779(.A0(new_n11082_), .A1(new_n11079_), .B0(new_n11215_), .Y(new_n11216_));
  AOI21X1  g08780(.A0(new_n11216_), .A1(new_n11214_), .B0(po1038), .Y(new_n11217_));
  AOI21X1  g08781(.A0(new_n11105_), .A1(pi0232), .B0(new_n11175_), .Y(new_n11218_));
  OAI22X1  g08782(.A0(new_n11106_), .A1(new_n11038_), .B0(new_n10440_), .B1(pi0232), .Y(new_n11219_));
  OAI21X1  g08783(.A0(new_n11219_), .A1(new_n11218_), .B0(new_n3156_), .Y(new_n11220_));
  OR2X1    g08784(.A(new_n10044_), .B(new_n3156_), .Y(new_n11221_));
  AND2X1   g08785(.A(new_n11221_), .B(po1038), .Y(new_n11222_));
  AOI22X1  g08786(.A0(new_n11222_), .A1(new_n11220_), .B0(new_n11217_), .B1(new_n11211_), .Y(po0283));
  NOR4X1   g08787(.A(new_n3242_), .B(new_n3003_), .C(new_n2555_), .D(new_n5095_), .Y(new_n11224_));
  AOI21X1  g08788(.A0(new_n4995_), .A1(pi0129), .B0(new_n2996_), .Y(new_n11225_));
  INVX1    g08789(.A(new_n2870_), .Y(new_n11226_));
  NOR2X1   g08790(.A(new_n5011_), .B(new_n2531_), .Y(new_n11227_));
  OR2X1    g08791(.A(new_n11227_), .B(new_n2515_), .Y(new_n11228_));
  OR2X1    g08792(.A(pi0102), .B(pi0081), .Y(new_n11229_));
  OR2X1    g08793(.A(new_n11229_), .B(new_n2673_), .Y(new_n11230_));
  AOI21X1  g08794(.A0(new_n11230_), .A1(new_n2604_), .B0(new_n2577_), .Y(new_n11231_));
  OAI21X1  g08795(.A0(new_n11231_), .A1(new_n2685_), .B0(new_n2601_), .Y(new_n11232_));
  AOI21X1  g08796(.A0(new_n11232_), .A1(new_n2687_), .B0(new_n2745_), .Y(new_n11233_));
  OR2X1    g08797(.A(new_n11233_), .B(new_n2599_), .Y(new_n11234_));
  AOI21X1  g08798(.A0(new_n11234_), .A1(new_n2474_), .B0(new_n2598_), .Y(new_n11235_));
  OAI21X1  g08799(.A0(new_n11235_), .A1(pi0097), .B0(new_n2589_), .Y(new_n11236_));
  AOI21X1  g08800(.A0(new_n11236_), .A1(new_n2576_), .B0(new_n2585_), .Y(new_n11237_));
  OAI21X1  g08801(.A0(new_n11237_), .A1(new_n2697_), .B0(new_n2575_), .Y(new_n11238_));
  AOI21X1  g08802(.A0(new_n11238_), .A1(new_n2573_), .B0(new_n2572_), .Y(new_n11239_));
  NAND2X1  g08803(.A(new_n11239_), .B(po0740), .Y(new_n11240_));
  OAI21X1  g08804(.A0(new_n11235_), .A1(new_n2596_), .B0(new_n2589_), .Y(new_n11241_));
  AOI21X1  g08805(.A0(new_n11241_), .A1(new_n2576_), .B0(new_n2585_), .Y(new_n11242_));
  OAI21X1  g08806(.A0(new_n11242_), .A1(new_n2697_), .B0(new_n2575_), .Y(new_n11243_));
  AOI21X1  g08807(.A0(new_n11243_), .A1(new_n2573_), .B0(new_n2572_), .Y(new_n11244_));
  NOR4X1   g08808(.A(new_n5970_), .B(new_n5094_), .C(new_n3053_), .D(new_n7846_), .Y(new_n11245_));
  INVX1    g08809(.A(new_n11245_), .Y(new_n11246_));
  AOI21X1  g08810(.A0(new_n11244_), .A1(new_n5922_), .B0(new_n11246_), .Y(new_n11247_));
  INVX1    g08811(.A(pi0127), .Y(new_n11248_));
  NAND2X1  g08812(.A(new_n11239_), .B(new_n11248_), .Y(new_n11249_));
  AOI21X1  g08813(.A0(new_n11244_), .A1(pi0127), .B0(new_n11245_), .Y(new_n11250_));
  AOI22X1  g08814(.A0(new_n11250_), .A1(new_n11249_), .B0(new_n11247_), .B1(new_n11240_), .Y(new_n11251_));
  OAI21X1  g08815(.A0(new_n11251_), .A1(new_n2565_), .B0(new_n2857_), .Y(new_n11252_));
  AOI21X1  g08816(.A0(new_n11252_), .A1(new_n2541_), .B0(new_n11228_), .Y(new_n11253_));
  OAI21X1  g08817(.A0(new_n11253_), .A1(pi0070), .B0(new_n11226_), .Y(new_n11254_));
  AOI21X1  g08818(.A0(new_n11254_), .A1(new_n2516_), .B0(new_n2557_), .Y(new_n11255_));
  OAI21X1  g08819(.A0(new_n11255_), .A1(new_n3194_), .B0(new_n2552_), .Y(new_n11256_));
  AOI21X1  g08820(.A0(new_n11256_), .A1(new_n2715_), .B0(new_n3202_), .Y(new_n11257_));
  NOR3X1   g08821(.A(new_n2716_), .B(new_n5095_), .C(pi0039), .Y(new_n11258_));
  OAI21X1  g08822(.A0(new_n11257_), .A1(pi0095), .B0(new_n11258_), .Y(new_n11259_));
  AOI21X1  g08823(.A0(new_n6761_), .A1(pi0039), .B0(pi0038), .Y(new_n11260_));
  AOI21X1  g08824(.A0(new_n11260_), .A1(new_n11259_), .B0(new_n11225_), .Y(new_n11261_));
  OAI21X1  g08825(.A0(new_n10121_), .A1(new_n3085_), .B0(new_n6761_), .Y(new_n11262_));
  AOI21X1  g08826(.A0(new_n11262_), .A1(new_n3124_), .B0(pi0075), .Y(new_n11263_));
  OAI21X1  g08827(.A0(new_n11261_), .A1(new_n3124_), .B0(new_n11263_), .Y(new_n11264_));
  NAND3X1  g08828(.A(new_n5789_), .B(pi0129), .C(pi0075), .Y(new_n11265_));
  AND2X1   g08829(.A(new_n11265_), .B(new_n3100_), .Y(new_n11266_));
  OAI21X1  g08830(.A0(pi0129), .A1(new_n3100_), .B0(new_n9927_), .Y(new_n11267_));
  AOI21X1  g08831(.A0(new_n11266_), .A1(new_n11264_), .B0(new_n11267_), .Y(new_n11268_));
  NAND3X1  g08832(.A(new_n3105_), .B(new_n3091_), .C(pi0054), .Y(new_n11269_));
  OAI21X1  g08833(.A0(new_n11269_), .A1(new_n6762_), .B0(new_n4991_), .Y(new_n11270_));
  NAND3X1  g08834(.A(new_n5789_), .B(new_n5319_), .C(pi0129), .Y(new_n11271_));
  AOI21X1  g08835(.A0(new_n11271_), .A1(pi0074), .B0(pi0055), .Y(new_n11272_));
  OAI21X1  g08836(.A0(new_n11270_), .A1(new_n11268_), .B0(new_n11272_), .Y(new_n11273_));
  NOR2X1   g08837(.A(new_n3125_), .B(new_n3128_), .Y(new_n11274_));
  NAND3X1  g08838(.A(new_n11274_), .B(new_n5789_), .C(pi0129), .Y(new_n11275_));
  AOI21X1  g08839(.A0(new_n11275_), .A1(new_n11273_), .B0(pi0056), .Y(new_n11276_));
  XOR2X1   g08840(.A(pi0062), .B(pi0056), .Y(new_n11277_));
  OAI22X1  g08841(.A0(new_n11277_), .A1(new_n11276_), .B0(new_n11224_), .B1(new_n3148_), .Y(new_n11278_));
  AOI21X1  g08842(.A0(new_n11224_), .A1(new_n3148_), .B0(new_n3246_), .Y(new_n11279_));
  OR2X1    g08843(.A(new_n11279_), .B(new_n4982_), .Y(new_n11280_));
  AOI21X1  g08844(.A0(new_n11278_), .A1(new_n3246_), .B0(new_n11280_), .Y(po0284));
  INVX1    g08845(.A(new_n5112_), .Y(new_n11282_));
  NOR2X1   g08846(.A(new_n5822_), .B(new_n4993_), .Y(new_n11283_));
  AOI21X1  g08847(.A0(new_n3407_), .A1(new_n2996_), .B0(new_n4998_), .Y(new_n11284_));
  NOR4X1   g08848(.A(new_n5098_), .B(new_n5086_), .C(new_n3074_), .D(pi0039), .Y(new_n11285_));
  OR2X1    g08849(.A(new_n11285_), .B(pi0087), .Y(new_n11286_));
  OAI21X1  g08850(.A0(new_n11286_), .A1(new_n11284_), .B0(new_n5105_), .Y(new_n11287_));
  NOR3X1   g08851(.A(new_n7851_), .B(new_n5970_), .C(new_n5094_), .Y(new_n11288_));
  OAI21X1  g08852(.A0(new_n11288_), .A1(pi0129), .B0(new_n6811_), .Y(new_n11289_));
  AOI21X1  g08853(.A0(new_n11288_), .A1(po0740), .B0(new_n11289_), .Y(new_n11290_));
  AOI21X1  g08854(.A0(new_n11290_), .A1(new_n3630_), .B0(new_n5107_), .Y(new_n11291_));
  OAI21X1  g08855(.A0(new_n5817_), .A1(new_n3112_), .B0(new_n5794_), .Y(new_n11292_));
  AOI21X1  g08856(.A0(new_n11291_), .A1(new_n11287_), .B0(new_n11292_), .Y(new_n11293_));
  OAI21X1  g08857(.A0(new_n11293_), .A1(new_n6755_), .B0(new_n11283_), .Y(new_n11294_));
  AOI21X1  g08858(.A0(new_n11294_), .A1(new_n3143_), .B0(new_n4989_), .Y(new_n11295_));
  OAI21X1  g08859(.A0(new_n11295_), .A1(pi0062), .B0(new_n11282_), .Y(new_n11296_));
  AOI21X1  g08860(.A0(new_n11296_), .A1(new_n3246_), .B0(new_n4985_), .Y(po0286));
  OR2X1    g08861(.A(new_n11018_), .B(pi0051), .Y(new_n11298_));
  AOI21X1  g08862(.A0(new_n11298_), .A1(new_n5237_), .B0(new_n9590_), .Y(new_n11299_));
  AND2X1   g08863(.A(new_n2953_), .B(pi0191), .Y(new_n11300_));
  AND2X1   g08864(.A(new_n11008_), .B(new_n2516_), .Y(new_n11301_));
  OAI21X1  g08865(.A0(new_n10602_), .A1(new_n7398_), .B0(new_n11301_), .Y(new_n11302_));
  NAND2X1  g08866(.A(new_n11302_), .B(new_n11300_), .Y(new_n11303_));
  NOR3X1   g08867(.A(new_n10594_), .B(new_n10590_), .C(pi0051), .Y(new_n11304_));
  NOR2X1   g08868(.A(new_n11002_), .B(pi0169), .Y(new_n11305_));
  NOR3X1   g08869(.A(new_n11305_), .B(new_n6905_), .C(new_n7349_), .Y(new_n11306_));
  OAI21X1  g08870(.A0(new_n11304_), .A1(new_n4210_), .B0(new_n11306_), .Y(new_n11307_));
  AND2X1   g08871(.A(new_n5033_), .B(pi0169), .Y(new_n11308_));
  OAI21X1  g08872(.A0(new_n3003_), .A1(new_n2555_), .B0(new_n11308_), .Y(new_n11309_));
  INVX1    g08873(.A(new_n11308_), .Y(new_n11310_));
  OR4X1    g08874(.A(new_n2437_), .B(new_n2438_), .C(pi0215), .D(pi0162), .Y(new_n11311_));
  AOI21X1  g08875(.A0(new_n11310_), .A1(new_n10604_), .B0(new_n11311_), .Y(new_n11312_));
  NOR3X1   g08876(.A(new_n10437_), .B(new_n6893_), .C(pi0051), .Y(new_n11313_));
  INVX1    g08877(.A(new_n11313_), .Y(new_n11314_));
  OAI21X1  g08878(.A0(new_n11314_), .A1(new_n11308_), .B0(pi0299), .Y(new_n11315_));
  AOI21X1  g08879(.A0(new_n11312_), .A1(new_n11309_), .B0(new_n11315_), .Y(new_n11316_));
  NOR2X1   g08880(.A(pi0299), .B(pi0191), .Y(new_n11317_));
  INVX1    g08881(.A(new_n11003_), .Y(new_n11318_));
  NOR2X1   g08882(.A(new_n10995_), .B(pi0051), .Y(new_n11319_));
  OAI21X1  g08883(.A0(new_n11318_), .A1(new_n7398_), .B0(new_n11319_), .Y(new_n11320_));
  AOI22X1  g08884(.A0(new_n11320_), .A1(new_n11317_), .B0(new_n11316_), .B1(new_n11307_), .Y(new_n11321_));
  AND2X1   g08885(.A(new_n11321_), .B(new_n11303_), .Y(new_n11322_));
  OAI21X1  g08886(.A0(new_n11322_), .A1(new_n5237_), .B0(new_n11299_), .Y(new_n11323_));
  OR4X1    g08887(.A(new_n6845_), .B(pi0468), .C(pi0332), .D(new_n5237_), .Y(new_n11324_));
  NAND3X1  g08888(.A(new_n11324_), .B(new_n11155_), .C(new_n9590_), .Y(new_n11325_));
  AND2X1   g08889(.A(new_n11325_), .B(new_n3026_), .Y(new_n11326_));
  AOI21X1  g08890(.A0(new_n11324_), .A1(new_n11155_), .B0(new_n11104_), .Y(new_n11327_));
  AOI21X1  g08891(.A0(new_n11327_), .A1(pi0100), .B0(new_n10641_), .Y(new_n11328_));
  OAI21X1  g08892(.A0(new_n10459_), .A1(new_n3026_), .B0(new_n11328_), .Y(new_n11329_));
  AOI21X1  g08893(.A0(new_n11326_), .A1(new_n11323_), .B0(new_n11329_), .Y(new_n11330_));
  INVX1    g08894(.A(new_n11327_), .Y(new_n11331_));
  AOI22X1  g08895(.A0(new_n11331_), .A1(new_n10645_), .B0(new_n7496_), .B1(pi0087), .Y(new_n11332_));
  INVX1    g08896(.A(pi0130), .Y(new_n11333_));
  INVX1    g08897(.A(pi0132), .Y(new_n11334_));
  NOR4X1   g08898(.A(pi0133), .B(pi0126), .C(pi0125), .D(pi0121), .Y(new_n11335_));
  AOI21X1  g08899(.A0(new_n11335_), .A1(new_n11334_), .B0(new_n11333_), .Y(new_n11336_));
  INVX1    g08900(.A(new_n11335_), .Y(new_n11337_));
  NOR3X1   g08901(.A(new_n11337_), .B(pi0132), .C(pi0130), .Y(new_n11338_));
  OAI21X1  g08902(.A0(new_n11338_), .A1(new_n11336_), .B0(new_n10431_), .Y(new_n11339_));
  OAI21X1  g08903(.A0(new_n11332_), .A1(new_n11215_), .B0(new_n11339_), .Y(new_n11340_));
  AND2X1   g08904(.A(new_n10889_), .B(new_n10992_), .Y(new_n11341_));
  MX2X1    g08905(.A(new_n10589_), .B(new_n10583_), .S0(new_n5033_), .Y(new_n11342_));
  MX2X1    g08906(.A(new_n11342_), .B(new_n11341_), .S0(pi0224), .Y(new_n11343_));
  MX2X1    g08907(.A(new_n11343_), .B(new_n11104_), .S0(new_n10859_), .Y(new_n11344_));
  MX2X1    g08908(.A(new_n11342_), .B(new_n11104_), .S0(new_n6278_), .Y(new_n11345_));
  INVX1    g08909(.A(new_n11345_), .Y(new_n11346_));
  OAI21X1  g08910(.A0(new_n11346_), .A1(pi0140), .B0(new_n11300_), .Y(new_n11347_));
  AOI21X1  g08911(.A0(new_n11344_), .A1(pi0140), .B0(new_n11347_), .Y(new_n11348_));
  NOR2X1   g08912(.A(new_n10583_), .B(new_n5057_), .Y(new_n11349_));
  NOR2X1   g08913(.A(new_n11308_), .B(new_n10589_), .Y(new_n11350_));
  AOI21X1  g08914(.A0(new_n11349_), .A1(pi0169), .B0(new_n11350_), .Y(new_n11351_));
  NOR3X1   g08915(.A(new_n10860_), .B(pi0169), .C(pi0051), .Y(new_n11352_));
  NAND3X1  g08916(.A(new_n10889_), .B(new_n10992_), .C(pi0169), .Y(new_n11353_));
  NAND3X1  g08917(.A(new_n11353_), .B(pi0216), .C(pi0162), .Y(new_n11354_));
  OAI22X1  g08918(.A0(new_n11354_), .A1(new_n11352_), .B0(new_n11351_), .B1(pi0216), .Y(new_n11355_));
  AND2X1   g08919(.A(new_n10541_), .B(pi0169), .Y(new_n11356_));
  OR2X1    g08920(.A(new_n11356_), .B(pi0051), .Y(new_n11357_));
  OAI21X1  g08921(.A0(new_n2438_), .A1(pi0162), .B0(new_n5241_), .Y(new_n11358_));
  AOI22X1  g08922(.A0(new_n11358_), .A1(new_n11357_), .B0(new_n11355_), .B1(new_n5241_), .Y(new_n11359_));
  AOI21X1  g08923(.A0(new_n10862_), .A1(new_n10588_), .B0(pi0051), .Y(new_n11360_));
  AND2X1   g08924(.A(new_n11360_), .B(pi0140), .Y(new_n11361_));
  AOI21X1  g08925(.A0(new_n10588_), .A1(new_n6277_), .B0(pi0051), .Y(new_n11362_));
  INVX1    g08926(.A(new_n11362_), .Y(new_n11363_));
  OAI21X1  g08927(.A0(new_n11363_), .A1(pi0140), .B0(new_n11317_), .Y(new_n11364_));
  OAI22X1  g08928(.A0(new_n11364_), .A1(new_n11361_), .B0(new_n11359_), .B1(new_n2953_), .Y(new_n11365_));
  OAI21X1  g08929(.A0(new_n11365_), .A1(new_n11348_), .B0(pi0232), .Y(new_n11366_));
  AOI21X1  g08930(.A0(new_n10849_), .A1(new_n10588_), .B0(pi0051), .Y(new_n11367_));
  OAI21X1  g08931(.A0(new_n11367_), .A1(pi0232), .B0(pi0039), .Y(new_n11368_));
  INVX1    g08932(.A(new_n11368_), .Y(new_n11369_));
  INVX1    g08933(.A(new_n10795_), .Y(new_n11370_));
  AOI21X1  g08934(.A0(new_n11370_), .A1(new_n5237_), .B0(pi0039), .Y(new_n11371_));
  MX2X1    g08935(.A(new_n11370_), .B(new_n10524_), .S0(new_n5033_), .Y(new_n11372_));
  AOI21X1  g08936(.A0(new_n10795_), .A1(new_n6845_), .B0(new_n5237_), .Y(new_n11373_));
  OAI21X1  g08937(.A0(new_n11372_), .A1(new_n6845_), .B0(new_n11373_), .Y(new_n11374_));
  AOI22X1  g08938(.A0(new_n11374_), .A1(new_n11371_), .B0(new_n11369_), .B1(new_n11366_), .Y(new_n11375_));
  AOI21X1  g08939(.A0(new_n11331_), .A1(pi0038), .B0(pi0100), .Y(new_n11376_));
  OAI21X1  g08940(.A0(new_n11375_), .A1(pi0038), .B0(new_n11376_), .Y(new_n11377_));
  AND2X1   g08941(.A(new_n11377_), .B(new_n11328_), .Y(new_n11378_));
  OR2X1    g08942(.A(new_n11338_), .B(new_n11336_), .Y(new_n11379_));
  NAND3X1  g08943(.A(new_n11379_), .B(new_n11332_), .C(new_n10431_), .Y(new_n11380_));
  OAI22X1  g08944(.A0(new_n11380_), .A1(new_n11378_), .B0(new_n11340_), .B1(new_n11330_), .Y(new_n11381_));
  NOR4X1   g08945(.A(new_n11356_), .B(new_n11339_), .C(pi0087), .D(pi0051), .Y(new_n11382_));
  NOR4X1   g08946(.A(pi0468), .B(pi0332), .C(new_n5237_), .D(new_n4210_), .Y(new_n11383_));
  NOR4X1   g08947(.A(new_n11383_), .B(new_n10437_), .C(pi0087), .D(pi0051), .Y(new_n11384_));
  OAI22X1  g08948(.A0(new_n7355_), .A1(new_n3156_), .B0(new_n5118_), .B1(pi0057), .Y(new_n11385_));
  NOR3X1   g08949(.A(new_n11385_), .B(new_n11384_), .C(new_n11382_), .Y(new_n11386_));
  AOI21X1  g08950(.A0(new_n11381_), .A1(new_n6520_), .B0(new_n11386_), .Y(po0287));
  OAI21X1  g08951(.A0(new_n5813_), .A1(new_n3026_), .B0(new_n3156_), .Y(new_n11388_));
  AOI21X1  g08952(.A0(new_n10153_), .A1(new_n3026_), .B0(new_n11388_), .Y(new_n11389_));
  OAI21X1  g08953(.A0(new_n11389_), .A1(pi0075), .B0(new_n5791_), .Y(new_n11390_));
  NAND3X1  g08954(.A(new_n8435_), .B(new_n5794_), .C(new_n3112_), .Y(new_n11391_));
  AOI21X1  g08955(.A0(new_n11390_), .A1(new_n3100_), .B0(new_n11391_), .Y(po0288));
  AOI22X1  g08956(.A0(new_n10560_), .A1(new_n9982_), .B0(new_n3325_), .B1(pi0051), .Y(new_n11393_));
  AND2X1   g08957(.A(new_n11393_), .B(new_n10451_), .Y(new_n11394_));
  OR2X1    g08958(.A(new_n10431_), .B(pi0132), .Y(new_n11395_));
  XOR2X1   g08959(.A(new_n11335_), .B(pi0132), .Y(new_n11396_));
  AND2X1   g08960(.A(new_n11396_), .B(new_n11395_), .Y(new_n11397_));
  INVX1    g08961(.A(new_n11397_), .Y(new_n11398_));
  AOI22X1  g08962(.A0(new_n11398_), .A1(new_n10440_), .B0(new_n11394_), .B1(pi0232), .Y(new_n11399_));
  AOI21X1  g08963(.A0(new_n10773_), .A1(pi0164), .B0(new_n6520_), .Y(new_n11400_));
  OAI21X1  g08964(.A0(new_n11399_), .A1(pi0087), .B0(new_n11400_), .Y(new_n11401_));
  NOR3X1   g08965(.A(new_n10516_), .B(new_n10491_), .C(new_n3325_), .Y(new_n11402_));
  AOI21X1  g08966(.A0(new_n10520_), .A1(new_n5190_), .B0(pi0151), .Y(new_n11403_));
  NOR3X1   g08967(.A(new_n11403_), .B(new_n11402_), .C(pi0168), .Y(new_n11404_));
  OAI21X1  g08968(.A0(pi0151), .A1(new_n2516_), .B0(pi0168), .Y(new_n11405_));
  OAI21X1  g08969(.A0(new_n11405_), .A1(new_n10488_), .B0(new_n5033_), .Y(new_n11406_));
  OR2X1    g08970(.A(new_n11406_), .B(new_n11404_), .Y(new_n11407_));
  AOI21X1  g08971(.A0(new_n10527_), .A1(new_n5057_), .B0(new_n8747_), .Y(new_n11408_));
  NOR2X1   g08972(.A(new_n10531_), .B(new_n10493_), .Y(new_n11409_));
  OAI21X1  g08973(.A0(new_n10527_), .A1(new_n5033_), .B0(new_n11409_), .Y(new_n11410_));
  OR2X1    g08974(.A(new_n10812_), .B(new_n4351_), .Y(new_n11411_));
  AOI21X1  g08975(.A0(new_n10527_), .A1(new_n5057_), .B0(new_n11411_), .Y(new_n11412_));
  OR2X1    g08976(.A(new_n11412_), .B(new_n3325_), .Y(new_n11413_));
  AOI21X1  g08977(.A0(new_n11410_), .A1(new_n4351_), .B0(new_n11413_), .Y(new_n11414_));
  NOR2X1   g08978(.A(new_n10527_), .B(new_n9981_), .Y(new_n11415_));
  NOR3X1   g08979(.A(new_n10536_), .B(new_n10534_), .C(new_n4351_), .Y(new_n11416_));
  OR2X1    g08980(.A(new_n11416_), .B(pi0151), .Y(new_n11417_));
  OAI21X1  g08981(.A0(new_n11417_), .A1(new_n11415_), .B0(new_n8747_), .Y(new_n11418_));
  OAI21X1  g08982(.A0(new_n11418_), .A1(new_n11414_), .B0(pi0299), .Y(new_n11419_));
  AOI21X1  g08983(.A0(new_n11408_), .A1(new_n11407_), .B0(new_n11419_), .Y(new_n11420_));
  OR2X1    g08984(.A(pi0299), .B(pi0190), .Y(new_n11421_));
  INVX1    g08985(.A(new_n10527_), .Y(new_n11422_));
  OAI21X1  g08986(.A0(new_n11422_), .A1(new_n5033_), .B0(pi0182), .Y(new_n11423_));
  AOI21X1  g08987(.A0(new_n11422_), .A1(new_n5227_), .B0(pi0173), .Y(new_n11424_));
  OAI21X1  g08988(.A0(new_n11423_), .A1(new_n10521_), .B0(new_n11424_), .Y(new_n11425_));
  MX2X1    g08989(.A(new_n10527_), .B(new_n10795_), .S0(new_n5033_), .Y(new_n11426_));
  AOI21X1  g08990(.A0(new_n11410_), .A1(new_n5227_), .B0(new_n9989_), .Y(new_n11427_));
  OAI21X1  g08991(.A0(new_n11426_), .A1(new_n5227_), .B0(new_n11427_), .Y(new_n11428_));
  AOI21X1  g08992(.A0(new_n11428_), .A1(new_n11425_), .B0(new_n11421_), .Y(new_n11429_));
  NOR2X1   g08993(.A(new_n10527_), .B(new_n5033_), .Y(new_n11430_));
  OR4X1    g08994(.A(new_n10481_), .B(new_n7272_), .C(new_n2458_), .D(new_n5227_), .Y(new_n11431_));
  OAI21X1  g08995(.A0(pi0173), .A1(new_n2516_), .B0(new_n5033_), .Y(new_n11432_));
  AOI21X1  g08996(.A0(new_n11431_), .A1(new_n10534_), .B0(new_n11432_), .Y(new_n11433_));
  NOR4X1   g08997(.A(new_n11433_), .B(new_n11430_), .C(pi0299), .D(new_n10004_), .Y(new_n11434_));
  OR4X1    g08998(.A(new_n11434_), .B(new_n11429_), .C(new_n11420_), .D(new_n5237_), .Y(new_n11435_));
  OR2X1    g08999(.A(new_n10527_), .B(pi0232), .Y(new_n11436_));
  AOI21X1  g09000(.A0(new_n11436_), .A1(new_n11435_), .B0(pi0039), .Y(new_n11437_));
  AOI21X1  g09001(.A0(new_n10605_), .A1(pi0168), .B0(pi0151), .Y(new_n11438_));
  OAI21X1  g09002(.A0(new_n11090_), .A1(pi0168), .B0(new_n11438_), .Y(new_n11439_));
  OAI21X1  g09003(.A0(new_n10860_), .A1(new_n10490_), .B0(new_n4351_), .Y(new_n11440_));
  AOI21X1  g09004(.A0(new_n11094_), .A1(pi0168), .B0(new_n3325_), .Y(new_n11441_));
  AOI21X1  g09005(.A0(new_n11441_), .A1(new_n11440_), .B0(new_n7129_), .Y(new_n11442_));
  AOI21X1  g09006(.A0(new_n11442_), .A1(new_n11439_), .B0(new_n2438_), .Y(new_n11443_));
  OR2X1    g09007(.A(pi0151), .B(new_n2516_), .Y(new_n11444_));
  MX2X1    g09008(.A(new_n11099_), .B(new_n11098_), .S0(pi0168), .Y(new_n11445_));
  AOI21X1  g09009(.A0(new_n11445_), .A1(new_n11444_), .B0(pi0216), .Y(new_n11446_));
  NOR3X1   g09010(.A(new_n11446_), .B(new_n11443_), .C(new_n5242_), .Y(new_n11447_));
  INVX1    g09011(.A(new_n11394_), .Y(new_n11448_));
  AOI21X1  g09012(.A0(pi0216), .A1(new_n7129_), .B0(new_n5242_), .Y(new_n11449_));
  OAI21X1  g09013(.A0(new_n11449_), .A1(new_n11448_), .B0(pi0299), .Y(new_n11450_));
  AND2X1   g09014(.A(new_n2953_), .B(pi0190), .Y(new_n11451_));
  OR2X1    g09015(.A(new_n10873_), .B(pi0183), .Y(new_n11452_));
  AND2X1   g09016(.A(new_n11452_), .B(new_n9989_), .Y(new_n11453_));
  OAI21X1  g09017(.A0(new_n10876_), .A1(new_n6928_), .B0(new_n11453_), .Y(new_n11454_));
  NAND3X1  g09018(.A(new_n10452_), .B(new_n6278_), .C(new_n6928_), .Y(new_n11455_));
  OAI21X1  g09019(.A0(new_n11098_), .A1(new_n6278_), .B0(new_n6928_), .Y(new_n11456_));
  NAND3X1  g09020(.A(new_n11456_), .B(new_n10870_), .C(pi0173), .Y(new_n11457_));
  NAND3X1  g09021(.A(new_n11457_), .B(new_n11455_), .C(new_n11454_), .Y(new_n11458_));
  NOR3X1   g09022(.A(new_n10882_), .B(new_n10490_), .C(pi0183), .Y(new_n11459_));
  NOR2X1   g09023(.A(new_n11459_), .B(new_n9989_), .Y(new_n11460_));
  OAI21X1  g09024(.A0(new_n10865_), .A1(new_n6928_), .B0(new_n11460_), .Y(new_n11461_));
  AOI21X1  g09025(.A0(new_n6278_), .A1(new_n6928_), .B0(pi0173), .Y(new_n11462_));
  AOI21X1  g09026(.A0(new_n11462_), .A1(new_n10877_), .B0(new_n11421_), .Y(new_n11463_));
  AOI22X1  g09027(.A0(new_n11463_), .A1(new_n11461_), .B0(new_n11458_), .B1(new_n11451_), .Y(new_n11464_));
  OAI21X1  g09028(.A0(new_n11450_), .A1(new_n11447_), .B0(new_n11464_), .Y(new_n11465_));
  AOI21X1  g09029(.A0(new_n11465_), .A1(pi0232), .B0(new_n11078_), .Y(new_n11466_));
  OAI21X1  g09030(.A0(new_n11466_), .A1(new_n11437_), .B0(new_n3277_), .Y(new_n11467_));
  NOR4X1   g09031(.A(pi0468), .B(pi0332), .C(new_n9989_), .D(new_n2516_), .Y(new_n11468_));
  OR2X1    g09032(.A(new_n11468_), .B(pi0299), .Y(new_n11469_));
  AOI21X1  g09033(.A0(new_n10541_), .A1(pi0190), .B0(new_n11469_), .Y(new_n11470_));
  AOI21X1  g09034(.A0(new_n11393_), .A1(new_n10451_), .B0(new_n2953_), .Y(new_n11471_));
  OR4X1    g09035(.A(new_n11471_), .B(new_n11470_), .C(new_n3277_), .D(new_n5237_), .Y(new_n11472_));
  AND2X1   g09036(.A(new_n11472_), .B(new_n5821_), .Y(new_n11473_));
  NOR3X1   g09037(.A(new_n11471_), .B(new_n11470_), .C(new_n5237_), .Y(new_n11474_));
  AOI21X1  g09038(.A0(new_n6850_), .A1(pi0087), .B0(new_n11398_), .Y(new_n11475_));
  OAI21X1  g09039(.A0(new_n11474_), .A1(new_n10720_), .B0(new_n11475_), .Y(new_n11476_));
  AOI21X1  g09040(.A0(new_n11473_), .A1(new_n11467_), .B0(new_n11476_), .Y(new_n11477_));
  AND2X1   g09041(.A(new_n11471_), .B(new_n10459_), .Y(new_n11478_));
  OAI21X1  g09042(.A0(new_n10609_), .A1(pi0168), .B0(pi0151), .Y(new_n11479_));
  AOI21X1  g09043(.A0(new_n10586_), .A1(pi0168), .B0(new_n11479_), .Y(new_n11480_));
  OAI21X1  g09044(.A0(new_n10583_), .A1(new_n9981_), .B0(new_n3325_), .Y(new_n11481_));
  AOI21X1  g09045(.A0(new_n10981_), .A1(pi0168), .B0(new_n11481_), .Y(new_n11482_));
  NOR3X1   g09046(.A(new_n11482_), .B(new_n11480_), .C(pi0149), .Y(new_n11483_));
  AOI21X1  g09047(.A0(new_n11444_), .A1(new_n10888_), .B0(new_n10590_), .Y(new_n11484_));
  NOR2X1   g09048(.A(new_n11484_), .B(new_n4351_), .Y(new_n11485_));
  OAI21X1  g09049(.A0(new_n11393_), .A1(new_n10624_), .B0(new_n4351_), .Y(new_n11486_));
  NAND2X1  g09050(.A(new_n11486_), .B(pi0149), .Y(new_n11487_));
  OAI21X1  g09051(.A0(new_n11487_), .A1(new_n11485_), .B0(new_n6893_), .Y(new_n11488_));
  OAI22X1  g09052(.A0(new_n11488_), .A1(new_n11483_), .B0(new_n11478_), .B1(new_n9591_), .Y(new_n11489_));
  NOR2X1   g09053(.A(new_n10994_), .B(pi0183), .Y(new_n11490_));
  OAI21X1  g09054(.A0(new_n11001_), .A1(new_n6928_), .B0(pi0173), .Y(new_n11491_));
  OAI21X1  g09055(.A0(new_n11009_), .A1(new_n6928_), .B0(new_n9989_), .Y(new_n11492_));
  OAI22X1  g09056(.A0(new_n11492_), .A1(new_n11186_), .B0(new_n11491_), .B1(new_n11490_), .Y(new_n11493_));
  OR4X1    g09057(.A(new_n11468_), .B(new_n10995_), .C(pi0299), .D(pi0190), .Y(new_n11494_));
  AOI21X1  g09058(.A0(new_n10624_), .A1(pi0183), .B0(new_n11494_), .Y(new_n11495_));
  AOI21X1  g09059(.A0(new_n11493_), .A1(new_n11451_), .B0(new_n11495_), .Y(new_n11496_));
  AOI21X1  g09060(.A0(new_n11496_), .A1(new_n11489_), .B0(new_n5237_), .Y(new_n11497_));
  OAI21X1  g09061(.A0(new_n11497_), .A1(new_n11019_), .B0(pi0039), .Y(new_n11498_));
  OAI21X1  g09062(.A0(new_n10483_), .A1(pi0151), .B0(new_n4351_), .Y(new_n11499_));
  AOI21X1  g09063(.A0(new_n10968_), .A1(pi0151), .B0(new_n11499_), .Y(new_n11500_));
  AOI21X1  g09064(.A0(new_n10490_), .A1(new_n3325_), .B0(new_n4351_), .Y(new_n11501_));
  AOI21X1  g09065(.A0(new_n11501_), .A1(new_n10708_), .B0(new_n11500_), .Y(new_n11502_));
  OAI21X1  g09066(.A0(new_n10483_), .A1(new_n5033_), .B0(new_n8747_), .Y(new_n11503_));
  OAI22X1  g09067(.A0(new_n10601_), .A1(pi0168), .B0(new_n10483_), .B1(new_n5033_), .Y(new_n11504_));
  NAND2X1  g09068(.A(new_n11504_), .B(pi0151), .Y(new_n11505_));
  NOR3X1   g09069(.A(new_n11394_), .B(new_n10922_), .C(pi0151), .Y(new_n11506_));
  NOR2X1   g09070(.A(new_n11506_), .B(new_n8747_), .Y(new_n11507_));
  AOI21X1  g09071(.A0(new_n11507_), .A1(new_n11505_), .B0(new_n2953_), .Y(new_n11508_));
  OAI21X1  g09072(.A0(new_n11503_), .A1(new_n11502_), .B0(new_n11508_), .Y(new_n11509_));
  AOI22X1  g09073(.A0(new_n10484_), .A1(new_n5057_), .B0(new_n9989_), .B1(pi0051), .Y(new_n11510_));
  OAI21X1  g09074(.A0(new_n10708_), .A1(pi0182), .B0(new_n11510_), .Y(new_n11511_));
  AND2X1   g09075(.A(new_n10922_), .B(pi0182), .Y(new_n11512_));
  OR4X1    g09076(.A(new_n11468_), .B(new_n10483_), .C(pi0299), .D(pi0190), .Y(new_n11513_));
  OAI21X1  g09077(.A0(new_n11513_), .A1(new_n11512_), .B0(pi0232), .Y(new_n11514_));
  AOI21X1  g09078(.A0(new_n11511_), .A1(new_n11451_), .B0(new_n11514_), .Y(new_n11515_));
  OAI21X1  g09079(.A0(new_n10484_), .A1(pi0232), .B0(new_n2959_), .Y(new_n11516_));
  AOI21X1  g09080(.A0(new_n11515_), .A1(new_n11509_), .B0(new_n11516_), .Y(new_n11517_));
  NOR2X1   g09081(.A(new_n11517_), .B(new_n5792_), .Y(new_n11518_));
  NAND3X1  g09082(.A(new_n11472_), .B(new_n11208_), .C(new_n5821_), .Y(new_n11519_));
  AOI21X1  g09083(.A0(new_n11518_), .A1(new_n11498_), .B0(new_n11519_), .Y(new_n11520_));
  AOI22X1  g09084(.A0(new_n11396_), .A1(new_n11395_), .B0(new_n6850_), .B1(pi0087), .Y(new_n11521_));
  OAI21X1  g09085(.A0(new_n11474_), .A1(new_n10646_), .B0(new_n11521_), .Y(new_n11522_));
  OAI21X1  g09086(.A0(new_n11522_), .A1(new_n11520_), .B0(new_n6520_), .Y(new_n11523_));
  OAI21X1  g09087(.A0(new_n11523_), .A1(new_n11477_), .B0(new_n11401_), .Y(po0289));
  AOI21X1  g09088(.A0(new_n10503_), .A1(new_n5057_), .B0(new_n10521_), .Y(new_n11525_));
  AND2X1   g09089(.A(pi0176), .B(new_n2959_), .Y(new_n11526_));
  OAI21X1  g09090(.A0(new_n10503_), .A1(new_n7189_), .B0(new_n11526_), .Y(new_n11527_));
  AOI21X1  g09091(.A0(new_n11525_), .A1(new_n7189_), .B0(new_n11527_), .Y(new_n11528_));
  NOR3X1   g09092(.A(new_n2953_), .B(new_n5237_), .C(new_n3158_), .Y(new_n11529_));
  NOR2X1   g09093(.A(pi0176), .B(pi0039), .Y(new_n11530_));
  OAI21X1  g09094(.A0(new_n11529_), .A1(new_n10503_), .B0(new_n11530_), .Y(new_n11531_));
  AOI21X1  g09095(.A0(new_n11529_), .A1(new_n11525_), .B0(new_n11531_), .Y(new_n11532_));
  INVX1    g09096(.A(new_n10850_), .Y(new_n11533_));
  NAND2X1  g09097(.A(new_n10690_), .B(new_n6278_), .Y(new_n11534_));
  OAI22X1  g09098(.A0(new_n10602_), .A1(new_n7347_), .B0(new_n2437_), .B1(pi0216), .Y(new_n11535_));
  AOI21X1  g09099(.A0(new_n6278_), .A1(new_n5224_), .B0(pi0299), .Y(new_n11536_));
  AOI22X1  g09100(.A0(new_n11536_), .A1(new_n11534_), .B0(new_n11535_), .B1(new_n5352_), .Y(new_n11537_));
  OAI21X1  g09101(.A0(new_n11537_), .A1(new_n3074_), .B0(pi0232), .Y(new_n11538_));
  AOI21X1  g09102(.A0(new_n11538_), .A1(new_n11533_), .B0(new_n2959_), .Y(new_n11539_));
  OR4X1    g09103(.A(new_n11539_), .B(new_n11532_), .C(new_n11528_), .D(new_n8508_), .Y(new_n11540_));
  AOI21X1  g09104(.A0(new_n10432_), .A1(new_n10766_), .B0(pi0133), .Y(new_n11541_));
  AND2X1   g09105(.A(new_n11541_), .B(new_n3156_), .Y(new_n11542_));
  NOR2X1   g09106(.A(new_n10995_), .B(pi0299), .Y(new_n11543_));
  OAI21X1  g09107(.A0(new_n10625_), .A1(new_n5224_), .B0(new_n11543_), .Y(new_n11544_));
  NAND2X1  g09108(.A(new_n10582_), .B(new_n6893_), .Y(new_n11545_));
  AOI21X1  g09109(.A0(new_n10594_), .A1(pi0197), .B0(new_n11545_), .Y(new_n11546_));
  OAI21X1  g09110(.A0(new_n11546_), .A1(new_n10459_), .B0(pi0299), .Y(new_n11547_));
  AND2X1   g09111(.A(new_n11547_), .B(new_n11544_), .Y(new_n11548_));
  OAI21X1  g09112(.A0(new_n11548_), .A1(new_n5237_), .B0(new_n11020_), .Y(new_n11549_));
  AND2X1   g09113(.A(new_n10440_), .B(new_n2959_), .Y(new_n11550_));
  OAI21X1  g09114(.A0(new_n10539_), .A1(new_n7192_), .B0(new_n11550_), .Y(new_n11551_));
  NAND3X1  g09115(.A(new_n11551_), .B(new_n11549_), .C(new_n2996_), .Y(new_n11552_));
  AOI21X1  g09116(.A0(new_n11552_), .A1(new_n10460_), .B0(new_n10643_), .Y(new_n11553_));
  AOI21X1  g09117(.A0(new_n10645_), .A1(new_n10459_), .B0(new_n11553_), .Y(new_n11554_));
  MX2X1    g09118(.A(pi0183), .B(pi0149), .S0(pi0299), .Y(new_n11555_));
  AND2X1   g09119(.A(new_n11555_), .B(new_n5930_), .Y(new_n11556_));
  OAI22X1  g09120(.A0(new_n11556_), .A1(new_n3156_), .B0(new_n11554_), .B1(new_n11541_), .Y(new_n11557_));
  AOI21X1  g09121(.A0(new_n11542_), .A1(new_n11540_), .B0(new_n11557_), .Y(new_n11558_));
  NOR3X1   g09122(.A(new_n11541_), .B(new_n10459_), .C(pi0087), .Y(new_n11559_));
  NAND4X1  g09123(.A(new_n5033_), .B(pi0232), .C(pi0149), .D(pi0087), .Y(new_n11560_));
  OAI21X1  g09124(.A0(new_n5118_), .A1(pi0057), .B0(new_n11560_), .Y(new_n11561_));
  OAI22X1  g09125(.A0(new_n11561_), .A1(new_n11559_), .B0(new_n11558_), .B1(po1038), .Y(po0290));
  INVX1    g09126(.A(pi0134), .Y(new_n11563_));
  INVX1    g09127(.A(pi0135), .Y(new_n11564_));
  NOR4X1   g09128(.A(new_n11337_), .B(pi0136), .C(pi0132), .D(pi0130), .Y(new_n11565_));
  AOI21X1  g09129(.A0(new_n11565_), .A1(new_n11564_), .B0(new_n11563_), .Y(new_n11566_));
  NAND3X1  g09130(.A(po1038), .B(new_n3156_), .C(new_n2516_), .Y(new_n11567_));
  NOR4X1   g09131(.A(new_n10437_), .B(pi0468), .C(pi0332), .D(new_n3774_), .Y(new_n11568_));
  AOI21X1  g09132(.A0(new_n11568_), .A1(pi0232), .B0(new_n11567_), .Y(new_n11569_));
  OAI21X1  g09133(.A0(new_n11566_), .A1(new_n10438_), .B0(new_n11569_), .Y(new_n11570_));
  AND2X1   g09134(.A(new_n11298_), .B(new_n5237_), .Y(new_n11571_));
  AND2X1   g09135(.A(pi0186), .B(pi0039), .Y(new_n11572_));
  AND2X1   g09136(.A(new_n2953_), .B(pi0192), .Y(new_n11573_));
  NAND3X1  g09137(.A(new_n11008_), .B(new_n10602_), .C(new_n2516_), .Y(new_n11574_));
  NOR2X1   g09138(.A(pi0299), .B(pi0192), .Y(new_n11575_));
  INVX1    g09139(.A(new_n11575_), .Y(new_n11576_));
  AOI21X1  g09140(.A0(new_n11319_), .A1(new_n11318_), .B0(new_n11576_), .Y(new_n11577_));
  AOI21X1  g09141(.A0(new_n11574_), .A1(new_n11573_), .B0(new_n11577_), .Y(new_n11578_));
  AND2X1   g09142(.A(new_n5033_), .B(pi0171), .Y(new_n11579_));
  OAI21X1  g09143(.A0(new_n11579_), .A1(new_n11314_), .B0(pi0299), .Y(new_n11580_));
  INVX1    g09144(.A(new_n11580_), .Y(new_n11581_));
  NOR3X1   g09145(.A(new_n5057_), .B(new_n3630_), .C(new_n3774_), .Y(new_n11582_));
  OAI21X1  g09146(.A0(new_n11579_), .A1(new_n10603_), .B0(new_n6893_), .Y(new_n11583_));
  OAI21X1  g09147(.A0(new_n11583_), .A1(new_n11582_), .B0(new_n11581_), .Y(new_n11584_));
  AOI21X1  g09148(.A0(new_n11584_), .A1(new_n11578_), .B0(new_n5237_), .Y(new_n11585_));
  OAI21X1  g09149(.A0(new_n11585_), .A1(new_n11571_), .B0(new_n11572_), .Y(new_n11586_));
  AND2X1   g09150(.A(new_n6861_), .B(pi0039), .Y(new_n11587_));
  INVX1    g09151(.A(new_n11319_), .Y(new_n11588_));
  INVX1    g09152(.A(new_n11573_), .Y(new_n11589_));
  AOI21X1  g09153(.A0(new_n11008_), .A1(new_n2516_), .B0(new_n11589_), .Y(new_n11590_));
  AOI21X1  g09154(.A0(new_n11575_), .A1(new_n11588_), .B0(new_n11590_), .Y(new_n11591_));
  AOI21X1  g09155(.A0(new_n11591_), .A1(new_n11584_), .B0(new_n5237_), .Y(new_n11592_));
  OAI21X1  g09156(.A0(new_n11592_), .A1(new_n11571_), .B0(new_n11587_), .Y(new_n11593_));
  INVX1    g09157(.A(pi0192), .Y(new_n11594_));
  MX2X1    g09158(.A(new_n11594_), .B(new_n3774_), .S0(pi0299), .Y(new_n11595_));
  INVX1    g09159(.A(new_n11595_), .Y(new_n11596_));
  AOI21X1  g09160(.A0(new_n11596_), .A1(new_n5930_), .B0(new_n11156_), .Y(new_n11597_));
  OR2X1    g09161(.A(new_n11597_), .B(pi0039), .Y(new_n11598_));
  NAND4X1  g09162(.A(new_n11598_), .B(new_n11593_), .C(new_n11586_), .D(new_n7223_), .Y(new_n11599_));
  NOR2X1   g09163(.A(new_n11304_), .B(new_n3774_), .Y(new_n11600_));
  OAI21X1  g09164(.A0(new_n11002_), .A1(pi0171), .B0(new_n6893_), .Y(new_n11601_));
  OAI21X1  g09165(.A0(new_n11601_), .A1(new_n11600_), .B0(new_n11581_), .Y(new_n11602_));
  AOI21X1  g09166(.A0(new_n11602_), .A1(new_n11578_), .B0(new_n5237_), .Y(new_n11603_));
  OAI21X1  g09167(.A0(new_n11603_), .A1(new_n11571_), .B0(new_n11572_), .Y(new_n11604_));
  AOI21X1  g09168(.A0(new_n11602_), .A1(new_n11591_), .B0(new_n5237_), .Y(new_n11605_));
  OAI21X1  g09169(.A0(new_n11605_), .A1(new_n11571_), .B0(new_n11587_), .Y(new_n11606_));
  NAND4X1  g09170(.A(new_n11606_), .B(new_n11604_), .C(new_n11598_), .D(pi0164), .Y(new_n11607_));
  NAND3X1  g09171(.A(new_n11607_), .B(new_n11599_), .C(new_n3277_), .Y(new_n11608_));
  NOR3X1   g09172(.A(new_n11597_), .B(new_n11104_), .C(new_n3277_), .Y(new_n11609_));
  NOR3X1   g09173(.A(new_n11609_), .B(new_n11207_), .C(new_n10641_), .Y(new_n11610_));
  AND2X1   g09174(.A(new_n11597_), .B(new_n10645_), .Y(new_n11611_));
  OR2X1    g09175(.A(new_n11611_), .B(new_n11566_), .Y(new_n11612_));
  AOI21X1  g09176(.A0(new_n11610_), .A1(new_n11608_), .B0(new_n11612_), .Y(new_n11613_));
  OR2X1    g09177(.A(new_n11609_), .B(new_n10641_), .Y(new_n11614_));
  NOR2X1   g09178(.A(new_n11568_), .B(pi0051), .Y(new_n11615_));
  AOI21X1  g09179(.A0(pi0216), .A1(new_n7223_), .B0(new_n5242_), .Y(new_n11616_));
  OR4X1    g09180(.A(new_n10583_), .B(pi0468), .C(pi0332), .D(new_n3774_), .Y(new_n11617_));
  OAI21X1  g09181(.A0(new_n11579_), .A1(new_n10589_), .B0(new_n11617_), .Y(new_n11618_));
  OR2X1    g09182(.A(new_n10860_), .B(pi0051), .Y(new_n11619_));
  OR2X1    g09183(.A(new_n11619_), .B(pi0171), .Y(new_n11620_));
  NAND2X1  g09184(.A(pi0216), .B(pi0164), .Y(new_n11621_));
  AOI21X1  g09185(.A0(new_n11341_), .A1(pi0171), .B0(new_n11621_), .Y(new_n11622_));
  AOI22X1  g09186(.A0(new_n11622_), .A1(new_n11620_), .B0(new_n11618_), .B1(new_n2438_), .Y(new_n11623_));
  OAI22X1  g09187(.A0(new_n11623_), .A1(new_n5242_), .B0(new_n11616_), .B1(new_n11615_), .Y(new_n11624_));
  AOI21X1  g09188(.A0(new_n11575_), .A1(new_n11363_), .B0(new_n11572_), .Y(new_n11625_));
  OAI21X1  g09189(.A0(new_n11589_), .A1(new_n11345_), .B0(new_n11625_), .Y(new_n11626_));
  INVX1    g09190(.A(new_n11360_), .Y(new_n11627_));
  AOI21X1  g09191(.A0(new_n11575_), .A1(new_n11627_), .B0(new_n6861_), .Y(new_n11628_));
  OAI21X1  g09192(.A0(new_n11589_), .A1(new_n11344_), .B0(new_n11628_), .Y(new_n11629_));
  AOI22X1  g09193(.A0(new_n11629_), .A1(new_n11626_), .B0(new_n11624_), .B1(pi0299), .Y(new_n11630_));
  OAI21X1  g09194(.A0(new_n11630_), .A1(new_n5237_), .B0(new_n11369_), .Y(new_n11631_));
  NAND3X1  g09195(.A(new_n11596_), .B(new_n11372_), .C(pi0232), .Y(new_n11632_));
  OAI22X1  g09196(.A0(new_n11595_), .A1(new_n5237_), .B0(new_n10516_), .B1(new_n10491_), .Y(new_n11633_));
  AND2X1   g09197(.A(new_n11633_), .B(new_n2959_), .Y(new_n11634_));
  AOI21X1  g09198(.A0(new_n11634_), .A1(new_n11632_), .B0(new_n5792_), .Y(new_n11635_));
  AOI21X1  g09199(.A0(new_n11635_), .A1(new_n11631_), .B0(new_n11614_), .Y(new_n11636_));
  OAI21X1  g09200(.A0(new_n11597_), .A1(new_n11104_), .B0(new_n10645_), .Y(new_n11637_));
  NAND2X1  g09201(.A(new_n11637_), .B(new_n11566_), .Y(new_n11638_));
  OAI21X1  g09202(.A0(new_n11638_), .A1(new_n11636_), .B0(new_n6520_), .Y(new_n11639_));
  OAI21X1  g09203(.A0(new_n11639_), .A1(new_n11613_), .B0(new_n11570_), .Y(po0291));
  INVX1    g09204(.A(pi0194), .Y(new_n11641_));
  AND2X1   g09205(.A(pi0299), .B(pi0232), .Y(new_n11642_));
  AND2X1   g09206(.A(new_n5033_), .B(pi0170), .Y(new_n11643_));
  AND2X1   g09207(.A(new_n11643_), .B(new_n11642_), .Y(new_n11644_));
  NOR2X1   g09208(.A(new_n11644_), .B(new_n11156_), .Y(new_n11645_));
  OAI21X1  g09209(.A0(new_n6862_), .A1(new_n11641_), .B0(new_n11645_), .Y(new_n11646_));
  AND2X1   g09210(.A(new_n11646_), .B(new_n11105_), .Y(new_n11647_));
  AOI21X1  g09211(.A0(new_n11647_), .A1(pi0100), .B0(new_n10641_), .Y(new_n11648_));
  AOI21X1  g09212(.A0(new_n11349_), .A1(pi0170), .B0(new_n6284_), .Y(new_n11649_));
  OAI21X1  g09213(.A0(new_n11643_), .A1(new_n10589_), .B0(new_n11649_), .Y(new_n11650_));
  NAND2X1  g09214(.A(new_n11650_), .B(new_n6905_), .Y(new_n11651_));
  NOR3X1   g09215(.A(new_n10860_), .B(pi0170), .C(pi0051), .Y(new_n11652_));
  NAND3X1  g09216(.A(new_n10889_), .B(new_n10992_), .C(pi0170), .Y(new_n11653_));
  NAND2X1  g09217(.A(new_n11653_), .B(pi0216), .Y(new_n11654_));
  OAI21X1  g09218(.A0(new_n11654_), .A1(new_n11652_), .B0(new_n11651_), .Y(new_n11655_));
  NAND2X1  g09219(.A(pi0299), .B(pi0150), .Y(new_n11656_));
  AOI21X1  g09220(.A0(new_n11643_), .A1(new_n10438_), .B0(pi0051), .Y(new_n11657_));
  AOI21X1  g09221(.A0(new_n11657_), .A1(new_n5242_), .B0(new_n11656_), .Y(new_n11658_));
  OR2X1    g09222(.A(new_n2953_), .B(pi0150), .Y(new_n11659_));
  AOI21X1  g09223(.A0(new_n11657_), .A1(new_n6284_), .B0(new_n11659_), .Y(new_n11660_));
  AOI22X1  g09224(.A0(new_n11660_), .A1(new_n11650_), .B0(new_n11658_), .B1(new_n11655_), .Y(new_n11661_));
  AOI21X1  g09225(.A0(new_n11362_), .A1(new_n9996_), .B0(pi0299), .Y(new_n11662_));
  OAI21X1  g09226(.A0(new_n11627_), .A1(new_n9996_), .B0(new_n11662_), .Y(new_n11663_));
  AOI21X1  g09227(.A0(new_n11663_), .A1(new_n11661_), .B0(new_n5237_), .Y(new_n11664_));
  NOR2X1   g09228(.A(new_n10795_), .B(pi0299), .Y(new_n11665_));
  NOR2X1   g09229(.A(new_n11372_), .B(new_n3917_), .Y(new_n11666_));
  OAI21X1  g09230(.A0(new_n11370_), .A1(pi0170), .B0(new_n11642_), .Y(new_n11667_));
  OAI21X1  g09231(.A0(new_n11667_), .A1(new_n11666_), .B0(new_n11371_), .Y(new_n11668_));
  OAI22X1  g09232(.A0(new_n11668_), .A1(new_n11665_), .B0(new_n11664_), .B1(new_n11368_), .Y(new_n11669_));
  OAI21X1  g09233(.A0(new_n11645_), .A1(new_n11104_), .B0(pi0038), .Y(new_n11670_));
  NAND2X1  g09234(.A(new_n11670_), .B(new_n11641_), .Y(new_n11671_));
  AOI21X1  g09235(.A0(new_n11669_), .A1(new_n2996_), .B0(new_n11671_), .Y(new_n11672_));
  AND2X1   g09236(.A(new_n11344_), .B(pi0185), .Y(new_n11673_));
  OAI21X1  g09237(.A0(new_n11346_), .A1(pi0185), .B0(new_n2953_), .Y(new_n11674_));
  OAI21X1  g09238(.A0(new_n11674_), .A1(new_n11673_), .B0(new_n11661_), .Y(new_n11675_));
  AND2X1   g09239(.A(new_n11675_), .B(pi0232), .Y(new_n11676_));
  AND2X1   g09240(.A(new_n11372_), .B(new_n7946_), .Y(new_n11677_));
  OAI22X1  g09241(.A0(new_n11677_), .A1(new_n11668_), .B0(new_n11676_), .B1(new_n11368_), .Y(new_n11678_));
  OAI21X1  g09242(.A0(new_n2953_), .A1(pi0170), .B0(new_n5930_), .Y(new_n11679_));
  AOI21X1  g09243(.A0(new_n11679_), .A1(new_n11155_), .B0(new_n11104_), .Y(new_n11680_));
  OAI21X1  g09244(.A0(new_n11680_), .A1(new_n2996_), .B0(pi0194), .Y(new_n11681_));
  AOI21X1  g09245(.A0(new_n11678_), .A1(new_n2996_), .B0(new_n11681_), .Y(new_n11682_));
  OAI21X1  g09246(.A0(new_n11682_), .A1(new_n11672_), .B0(new_n3026_), .Y(new_n11683_));
  NOR2X1   g09247(.A(new_n11565_), .B(new_n11564_), .Y(new_n11684_));
  INVX1    g09248(.A(new_n11338_), .Y(new_n11685_));
  NOR4X1   g09249(.A(new_n11685_), .B(pi0136), .C(pi0135), .D(new_n11563_), .Y(new_n11686_));
  OAI22X1  g09250(.A0(new_n11686_), .A1(new_n11684_), .B0(new_n11647_), .B1(new_n10720_), .Y(new_n11687_));
  AOI21X1  g09251(.A0(new_n11683_), .A1(new_n11648_), .B0(new_n11687_), .Y(new_n11688_));
  NOR3X1   g09252(.A(new_n11644_), .B(new_n11156_), .C(new_n8244_), .Y(new_n11689_));
  OR2X1    g09253(.A(new_n11689_), .B(pi0194), .Y(new_n11690_));
  NAND3X1  g09254(.A(new_n11679_), .B(new_n11155_), .C(new_n9590_), .Y(new_n11691_));
  AND2X1   g09255(.A(new_n11691_), .B(pi0194), .Y(new_n11692_));
  INVX1    g09256(.A(new_n11692_), .Y(new_n11693_));
  AND2X1   g09257(.A(new_n11693_), .B(new_n11690_), .Y(new_n11694_));
  AOI21X1  g09258(.A0(new_n11003_), .A1(pi0185), .B0(new_n11588_), .Y(new_n11695_));
  AND2X1   g09259(.A(new_n11301_), .B(new_n9996_), .Y(new_n11696_));
  NAND2X1  g09260(.A(new_n11692_), .B(new_n11574_), .Y(new_n11697_));
  OAI22X1  g09261(.A0(new_n11697_), .A1(new_n11696_), .B0(new_n11690_), .B1(new_n11695_), .Y(new_n11698_));
  NOR2X1   g09262(.A(new_n11304_), .B(new_n3917_), .Y(new_n11699_));
  OAI21X1  g09263(.A0(new_n11002_), .A1(pi0170), .B0(new_n6893_), .Y(new_n11700_));
  NOR2X1   g09264(.A(new_n11700_), .B(new_n11699_), .Y(new_n11701_));
  AND2X1   g09265(.A(new_n3074_), .B(pi0170), .Y(new_n11702_));
  OAI21X1  g09266(.A0(new_n11643_), .A1(new_n10603_), .B0(new_n6893_), .Y(new_n11703_));
  AOI21X1  g09267(.A0(new_n5033_), .A1(new_n11702_), .B0(new_n11703_), .Y(new_n11704_));
  OAI22X1  g09268(.A0(new_n11704_), .A1(new_n11659_), .B0(new_n11701_), .B1(new_n11656_), .Y(new_n11705_));
  INVX1    g09269(.A(new_n11643_), .Y(new_n11706_));
  AOI22X1  g09270(.A0(new_n11693_), .A1(new_n11690_), .B0(new_n11706_), .B1(new_n11313_), .Y(new_n11707_));
  AOI22X1  g09271(.A0(new_n11707_), .A1(new_n11705_), .B0(new_n11698_), .B1(new_n2953_), .Y(new_n11708_));
  OAI22X1  g09272(.A0(new_n11708_), .A1(new_n5237_), .B0(new_n11694_), .B1(new_n11299_), .Y(new_n11709_));
  OAI21X1  g09273(.A0(new_n10459_), .A1(new_n3026_), .B0(new_n11648_), .Y(new_n11710_));
  AOI21X1  g09274(.A0(new_n11709_), .A1(new_n3026_), .B0(new_n11710_), .Y(new_n11711_));
  NOR2X1   g09275(.A(new_n11686_), .B(new_n11684_), .Y(new_n11712_));
  OAI21X1  g09276(.A0(new_n11646_), .A1(new_n10720_), .B0(new_n11712_), .Y(new_n11713_));
  OAI21X1  g09277(.A0(new_n11713_), .A1(new_n11711_), .B0(new_n6520_), .Y(new_n11714_));
  NAND2X1  g09278(.A(new_n11712_), .B(new_n10437_), .Y(new_n11715_));
  NOR4X1   g09279(.A(pi0468), .B(pi0332), .C(new_n5237_), .D(new_n3917_), .Y(new_n11716_));
  AOI21X1  g09280(.A0(new_n11716_), .A1(new_n10438_), .B0(new_n11567_), .Y(new_n11717_));
  NAND2X1  g09281(.A(new_n11717_), .B(new_n11715_), .Y(new_n11718_));
  OAI21X1  g09282(.A0(new_n11714_), .A1(new_n11688_), .B0(new_n11718_), .Y(po0292));
  NOR3X1   g09283(.A(pi0136), .B(pi0135), .C(pi0134), .Y(new_n11720_));
  XOR2X1   g09284(.A(new_n11685_), .B(pi0136), .Y(new_n11721_));
  NOR2X1   g09285(.A(new_n11721_), .B(new_n11720_), .Y(new_n11722_));
  NAND3X1  g09286(.A(new_n5033_), .B(pi0232), .C(pi0148), .Y(new_n11723_));
  AOI22X1  g09287(.A0(new_n11723_), .A1(new_n10438_), .B0(new_n11722_), .B1(new_n11156_), .Y(new_n11724_));
  INVX1    g09288(.A(new_n11371_), .Y(new_n11725_));
  OR2X1    g09289(.A(new_n11372_), .B(new_n7383_), .Y(new_n11726_));
  AOI21X1  g09290(.A0(new_n10795_), .A1(new_n7383_), .B0(new_n5237_), .Y(new_n11727_));
  AND2X1   g09291(.A(new_n11727_), .B(new_n11726_), .Y(new_n11728_));
  AND2X1   g09292(.A(new_n2953_), .B(pi0141), .Y(new_n11729_));
  OAI21X1  g09293(.A0(new_n11346_), .A1(pi0184), .B0(new_n11729_), .Y(new_n11730_));
  AOI21X1  g09294(.A0(new_n11344_), .A1(pi0184), .B0(new_n11730_), .Y(new_n11731_));
  AND2X1   g09295(.A(new_n11360_), .B(pi0184), .Y(new_n11732_));
  NOR2X1   g09296(.A(pi0299), .B(pi0141), .Y(new_n11733_));
  OAI21X1  g09297(.A0(new_n11363_), .A1(pi0184), .B0(new_n11733_), .Y(new_n11734_));
  NAND4X1  g09298(.A(new_n10889_), .B(new_n10992_), .C(new_n5241_), .D(pi0163), .Y(new_n11735_));
  OR2X1    g09299(.A(new_n11104_), .B(new_n6283_), .Y(new_n11736_));
  AOI22X1  g09300(.A0(new_n11736_), .A1(new_n8705_), .B0(new_n11104_), .B1(new_n5242_), .Y(new_n11737_));
  AOI21X1  g09301(.A0(new_n11737_), .A1(new_n11735_), .B0(new_n4036_), .Y(new_n11738_));
  OAI21X1  g09302(.A0(new_n11342_), .A1(new_n6284_), .B0(new_n11738_), .Y(new_n11739_));
  NOR4X1   g09303(.A(pi0468), .B(pi0332), .C(pi0287), .D(new_n8705_), .Y(new_n11740_));
  OAI21X1  g09304(.A0(new_n11740_), .A1(new_n2438_), .B0(new_n5241_), .Y(new_n11741_));
  OR4X1    g09305(.A(new_n11741_), .B(new_n3256_), .C(new_n2555_), .D(pi0096), .Y(new_n11742_));
  NAND3X1  g09306(.A(new_n11742_), .B(new_n4036_), .C(new_n2516_), .Y(new_n11743_));
  NAND3X1  g09307(.A(new_n11743_), .B(new_n11739_), .C(pi0299), .Y(new_n11744_));
  OAI21X1  g09308(.A0(new_n11734_), .A1(new_n11732_), .B0(new_n11744_), .Y(new_n11745_));
  OAI21X1  g09309(.A0(new_n11745_), .A1(new_n11731_), .B0(pi0232), .Y(new_n11746_));
  AOI21X1  g09310(.A0(new_n11746_), .A1(new_n11369_), .B0(new_n5792_), .Y(new_n11747_));
  OAI21X1  g09311(.A0(new_n11728_), .A1(new_n11725_), .B0(new_n11747_), .Y(new_n11748_));
  OAI21X1  g09312(.A0(new_n10437_), .A1(new_n7385_), .B0(new_n2516_), .Y(new_n11749_));
  AOI21X1  g09313(.A0(new_n11749_), .A1(new_n5792_), .B0(new_n10641_), .Y(new_n11750_));
  OAI21X1  g09314(.A0(new_n11749_), .A1(new_n10720_), .B0(new_n11722_), .Y(new_n11751_));
  AOI21X1  g09315(.A0(new_n11750_), .A1(new_n11748_), .B0(new_n11751_), .Y(new_n11752_));
  NOR4X1   g09316(.A(new_n10437_), .B(new_n8339_), .C(new_n7384_), .D(pi0051), .Y(new_n11753_));
  INVX1    g09317(.A(new_n11729_), .Y(new_n11754_));
  NAND2X1  g09318(.A(new_n10594_), .B(pi0184), .Y(new_n11755_));
  AOI21X1  g09319(.A0(new_n11755_), .A1(new_n11301_), .B0(new_n11754_), .Y(new_n11756_));
  INVX1    g09320(.A(new_n11733_), .Y(new_n11757_));
  OR4X1    g09321(.A(new_n10590_), .B(new_n5242_), .C(new_n2438_), .D(pi0051), .Y(new_n11758_));
  AOI21X1  g09322(.A0(new_n11313_), .A1(new_n5057_), .B0(new_n4036_), .Y(new_n11759_));
  INVX1    g09323(.A(new_n11740_), .Y(new_n11760_));
  OAI21X1  g09324(.A0(new_n11545_), .A1(pi0051), .B0(new_n4036_), .Y(new_n11761_));
  AOI22X1  g09325(.A0(new_n11761_), .A1(new_n11760_), .B0(new_n11155_), .B1(new_n4036_), .Y(new_n11762_));
  AOI21X1  g09326(.A0(new_n11759_), .A1(new_n11758_), .B0(new_n11762_), .Y(new_n11763_));
  AOI21X1  g09327(.A0(new_n11003_), .A1(pi0184), .B0(new_n11588_), .Y(new_n11764_));
  OAI22X1  g09328(.A0(new_n11764_), .A1(new_n11757_), .B0(new_n11763_), .B1(new_n2953_), .Y(new_n11765_));
  OAI21X1  g09329(.A0(new_n11765_), .A1(new_n11756_), .B0(pi0232), .Y(new_n11766_));
  AND2X1   g09330(.A(new_n11299_), .B(new_n3026_), .Y(new_n11767_));
  AOI21X1  g09331(.A0(new_n11767_), .A1(new_n11766_), .B0(new_n11753_), .Y(new_n11768_));
  NOR4X1   g09332(.A(new_n10720_), .B(new_n10437_), .C(new_n7384_), .D(pi0051), .Y(new_n11769_));
  NOR2X1   g09333(.A(new_n11769_), .B(new_n11722_), .Y(new_n11770_));
  OAI21X1  g09334(.A0(new_n11768_), .A1(new_n10641_), .B0(new_n11770_), .Y(new_n11771_));
  NAND2X1  g09335(.A(new_n11771_), .B(new_n6520_), .Y(new_n11772_));
  OAI22X1  g09336(.A0(new_n11772_), .A1(new_n11752_), .B0(new_n11724_), .B1(new_n11567_), .Y(po0293));
  OR4X1    g09337(.A(new_n10761_), .B(new_n3003_), .C(new_n2555_), .D(new_n7862_), .Y(new_n11774_));
  NAND4X1  g09338(.A(new_n7783_), .B(new_n4515_), .C(pi0299), .D(new_n2766_), .Y(new_n11775_));
  AND2X1   g09339(.A(new_n6520_), .B(new_n2953_), .Y(new_n11776_));
  INVX1    g09340(.A(new_n11776_), .Y(new_n11777_));
  NAND3X1  g09341(.A(new_n5033_), .B(new_n2980_), .C(new_n2973_), .Y(new_n11778_));
  OAI21X1  g09342(.A0(new_n11778_), .A1(new_n11777_), .B0(new_n11775_), .Y(new_n11779_));
  NOR3X1   g09343(.A(new_n8682_), .B(new_n6520_), .C(pi0210), .Y(new_n11780_));
  AOI21X1  g09344(.A0(new_n11779_), .A1(new_n11774_), .B0(new_n11780_), .Y(new_n11781_));
  OAI22X1  g09345(.A0(new_n11781_), .A1(new_n7892_), .B0(new_n2453_), .B1(pi0039), .Y(po0294));
  NOR3X1   g09346(.A(new_n7230_), .B(new_n7502_), .C(new_n6832_), .Y(new_n11783_));
  OAI21X1  g09347(.A0(new_n11783_), .A1(new_n3100_), .B0(new_n3135_), .Y(new_n11784_));
  INVX1    g09348(.A(new_n11784_), .Y(new_n11785_));
  AOI21X1  g09349(.A0(new_n7181_), .A1(pi0087), .B0(pi0075), .Y(new_n11786_));
  INVX1    g09350(.A(new_n11786_), .Y(new_n11787_));
  NOR3X1   g09351(.A(new_n7110_), .B(new_n6990_), .C(new_n6935_), .Y(new_n11788_));
  NOR2X1   g09352(.A(new_n11788_), .B(new_n2953_), .Y(new_n11789_));
  NOR2X1   g09353(.A(new_n7419_), .B(pi0299), .Y(new_n11790_));
  NOR3X1   g09354(.A(new_n11790_), .B(new_n11789_), .C(pi0232), .Y(new_n11791_));
  NOR2X1   g09355(.A(new_n11791_), .B(pi0039), .Y(new_n11792_));
  MX2X1    g09356(.A(new_n7419_), .B(new_n6978_), .S0(new_n5033_), .Y(new_n11793_));
  NOR3X1   g09357(.A(new_n11793_), .B(pi0299), .C(new_n7382_), .Y(new_n11794_));
  NOR2X1   g09358(.A(new_n7114_), .B(new_n5057_), .Y(new_n11795_));
  AOI21X1  g09359(.A0(new_n5033_), .A1(pi0148), .B0(new_n11788_), .Y(new_n11796_));
  AOI21X1  g09360(.A0(new_n11795_), .A1(pi0148), .B0(new_n11796_), .Y(new_n11797_));
  AOI21X1  g09361(.A0(new_n11790_), .A1(new_n7382_), .B0(new_n5237_), .Y(new_n11798_));
  OAI21X1  g09362(.A0(new_n11797_), .A1(new_n2953_), .B0(new_n11798_), .Y(new_n11799_));
  OAI21X1  g09363(.A0(new_n11799_), .A1(new_n11794_), .B0(new_n11792_), .Y(new_n11800_));
  NAND3X1  g09364(.A(new_n6915_), .B(new_n6886_), .C(new_n6869_), .Y(new_n11801_));
  NOR2X1   g09365(.A(new_n8915_), .B(new_n6902_), .Y(new_n11802_));
  NOR2X1   g09366(.A(new_n11802_), .B(new_n11801_), .Y(new_n11803_));
  NOR2X1   g09367(.A(new_n11803_), .B(new_n10022_), .Y(new_n11804_));
  NOR2X1   g09368(.A(new_n6902_), .B(new_n5070_), .Y(new_n11805_));
  NOR3X1   g09369(.A(new_n11805_), .B(new_n11802_), .C(new_n6905_), .Y(new_n11806_));
  NOR2X1   g09370(.A(new_n11806_), .B(new_n6922_), .Y(new_n11807_));
  OAI21X1  g09371(.A0(new_n11807_), .A1(new_n11804_), .B0(new_n5237_), .Y(new_n11808_));
  AOI21X1  g09372(.A0(new_n6898_), .A1(new_n5071_), .B0(new_n11802_), .Y(new_n11809_));
  INVX1    g09373(.A(new_n11809_), .Y(new_n11810_));
  AOI21X1  g09374(.A0(new_n11810_), .A1(new_n6894_), .B0(new_n4036_), .Y(new_n11811_));
  AOI21X1  g09375(.A0(pi0299), .A1(pi0148), .B0(new_n11807_), .Y(new_n11812_));
  NOR2X1   g09376(.A(new_n11812_), .B(new_n11811_), .Y(new_n11813_));
  NOR3X1   g09377(.A(new_n11802_), .B(new_n6923_), .C(new_n11801_), .Y(new_n11814_));
  NOR2X1   g09378(.A(new_n11814_), .B(new_n10022_), .Y(new_n11815_));
  MX2X1    g09379(.A(new_n11815_), .B(new_n11804_), .S0(new_n7382_), .Y(new_n11816_));
  OAI21X1  g09380(.A0(new_n11816_), .A1(new_n11813_), .B0(pi0232), .Y(new_n11817_));
  AOI21X1  g09381(.A0(new_n11817_), .A1(new_n11808_), .B0(new_n2959_), .Y(new_n11818_));
  NOR2X1   g09382(.A(new_n11818_), .B(new_n5792_), .Y(new_n11819_));
  AOI21X1  g09383(.A0(new_n11819_), .A1(new_n11800_), .B0(pi0087), .Y(new_n11820_));
  OAI21X1  g09384(.A0(new_n11820_), .A1(new_n11787_), .B0(new_n3100_), .Y(new_n11821_));
  AOI21X1  g09385(.A0(new_n11821_), .A1(new_n11785_), .B0(pi0055), .Y(new_n11822_));
  OAI21X1  g09386(.A0(new_n10045_), .A1(new_n7368_), .B0(pi0055), .Y(new_n11823_));
  INVX1    g09387(.A(new_n11823_), .Y(new_n11824_));
  OAI21X1  g09388(.A0(new_n11824_), .A1(new_n11822_), .B0(new_n3148_), .Y(new_n11825_));
  NAND3X1  g09389(.A(new_n11825_), .B(new_n7369_), .C(pi0138), .Y(new_n11826_));
  AND2X1   g09390(.A(new_n8575_), .B(new_n5237_), .Y(new_n11827_));
  INVX1    g09391(.A(new_n11827_), .Y(new_n11828_));
  NAND2X1  g09392(.A(pi0299), .B(pi0148), .Y(new_n11829_));
  AND2X1   g09393(.A(new_n5261_), .B(new_n6269_), .Y(new_n11830_));
  AND2X1   g09394(.A(new_n11830_), .B(new_n6886_), .Y(new_n11831_));
  OAI22X1  g09395(.A0(new_n11831_), .A1(new_n11754_), .B0(new_n11829_), .B1(new_n6269_), .Y(new_n11832_));
  AOI21X1  g09396(.A0(new_n8575_), .A1(new_n11754_), .B0(new_n11832_), .Y(new_n11833_));
  OR2X1    g09397(.A(new_n11833_), .B(new_n5237_), .Y(new_n11834_));
  AOI21X1  g09398(.A0(new_n11834_), .A1(new_n11828_), .B0(new_n2959_), .Y(new_n11835_));
  AOI21X1  g09399(.A0(new_n10091_), .A1(new_n7385_), .B0(pi0039), .Y(new_n11836_));
  OR4X1    g09400(.A(new_n11836_), .B(new_n11835_), .C(new_n7690_), .D(pi0138), .Y(new_n11837_));
  NAND2X1  g09401(.A(new_n10057_), .B(new_n6817_), .Y(new_n11838_));
  NOR2X1   g09402(.A(new_n11838_), .B(pi0139), .Y(new_n11839_));
  INVX1    g09403(.A(new_n11839_), .Y(new_n11840_));
  AND2X1   g09404(.A(new_n11840_), .B(new_n11837_), .Y(new_n11841_));
  INVX1    g09405(.A(pi0195), .Y(new_n11842_));
  INVX1    g09406(.A(pi0196), .Y(new_n11843_));
  AOI21X1  g09407(.A0(new_n11843_), .A1(new_n11842_), .B0(pi0138), .Y(new_n11844_));
  NAND3X1  g09408(.A(new_n11844_), .B(new_n11825_), .C(new_n7369_), .Y(new_n11845_));
  OR4X1    g09409(.A(new_n11844_), .B(new_n11836_), .C(new_n11835_), .D(new_n7690_), .Y(new_n11846_));
  AND2X1   g09410(.A(new_n11846_), .B(new_n11839_), .Y(new_n11847_));
  AOI22X1  g09411(.A0(new_n11847_), .A1(new_n11845_), .B0(new_n11841_), .B1(new_n11826_), .Y(po0295));
  NOR3X1   g09412(.A(new_n11793_), .B(pi0299), .C(new_n6844_), .Y(new_n11849_));
  INVX1    g09413(.A(new_n11788_), .Y(new_n11850_));
  AOI22X1  g09414(.A0(new_n11310_), .A1(new_n11850_), .B0(new_n11795_), .B1(pi0169), .Y(new_n11851_));
  AOI21X1  g09415(.A0(new_n11790_), .A1(new_n6844_), .B0(new_n5237_), .Y(new_n11852_));
  OAI21X1  g09416(.A0(new_n11851_), .A1(new_n2953_), .B0(new_n11852_), .Y(new_n11853_));
  OAI21X1  g09417(.A0(new_n11853_), .A1(new_n11849_), .B0(new_n11792_), .Y(new_n11854_));
  OAI21X1  g09418(.A0(new_n7474_), .A1(pi0169), .B0(new_n11810_), .Y(new_n11855_));
  AOI21X1  g09419(.A0(new_n11855_), .A1(new_n6893_), .B0(new_n6922_), .Y(new_n11856_));
  MX2X1    g09420(.A(new_n11815_), .B(new_n11804_), .S0(new_n6844_), .Y(new_n11857_));
  OAI21X1  g09421(.A0(new_n11857_), .A1(new_n11856_), .B0(pi0232), .Y(new_n11858_));
  AOI21X1  g09422(.A0(new_n11858_), .A1(new_n11808_), .B0(new_n2959_), .Y(new_n11859_));
  NOR2X1   g09423(.A(new_n11859_), .B(new_n5792_), .Y(new_n11860_));
  AOI21X1  g09424(.A0(new_n11860_), .A1(new_n11854_), .B0(pi0087), .Y(new_n11861_));
  OAI21X1  g09425(.A0(new_n11861_), .A1(new_n11787_), .B0(new_n3100_), .Y(new_n11862_));
  AOI21X1  g09426(.A0(new_n11862_), .A1(new_n11785_), .B0(pi0055), .Y(new_n11863_));
  OAI21X1  g09427(.A0(new_n11863_), .A1(new_n11824_), .B0(new_n3148_), .Y(new_n11864_));
  NAND3X1  g09428(.A(new_n11864_), .B(new_n7369_), .C(pi0139), .Y(new_n11865_));
  INVX1    g09429(.A(pi0139), .Y(new_n11866_));
  NOR3X1   g09430(.A(new_n6269_), .B(new_n2953_), .C(new_n4210_), .Y(new_n11867_));
  NOR3X1   g09431(.A(new_n8571_), .B(pi0299), .C(pi0191), .Y(new_n11868_));
  NOR3X1   g09432(.A(new_n11831_), .B(pi0299), .C(new_n6844_), .Y(new_n11869_));
  OR4X1    g09433(.A(new_n11869_), .B(new_n11868_), .C(new_n11867_), .D(new_n8573_), .Y(new_n11870_));
  MX2X1    g09434(.A(new_n11870_), .B(new_n8575_), .S0(new_n5237_), .Y(new_n11871_));
  AOI21X1  g09435(.A0(new_n11324_), .A1(new_n10091_), .B0(pi0039), .Y(new_n11872_));
  OR2X1    g09436(.A(new_n11872_), .B(new_n7690_), .Y(new_n11873_));
  AOI21X1  g09437(.A0(new_n11871_), .A1(pi0039), .B0(new_n11873_), .Y(new_n11874_));
  AOI22X1  g09438(.A0(new_n11874_), .A1(new_n11866_), .B0(new_n10057_), .B1(new_n6817_), .Y(new_n11875_));
  NOR3X1   g09439(.A(pi0196), .B(pi0195), .C(pi0138), .Y(new_n11876_));
  NOR2X1   g09440(.A(new_n11876_), .B(pi0139), .Y(new_n11877_));
  NAND3X1  g09441(.A(new_n11877_), .B(new_n11864_), .C(new_n7369_), .Y(new_n11878_));
  INVX1    g09442(.A(new_n11877_), .Y(new_n11879_));
  AOI21X1  g09443(.A0(new_n11879_), .A1(new_n11874_), .B0(new_n11838_), .Y(new_n11880_));
  AOI22X1  g09444(.A0(new_n11880_), .A1(new_n11878_), .B0(new_n11875_), .B1(new_n11865_), .Y(po0296));
  INVX1    g09445(.A(pi1160), .Y(new_n11882_));
  INVX1    g09446(.A(pi0787), .Y(new_n11883_));
  INVX1    g09447(.A(pi0792), .Y(new_n11884_));
  INVX1    g09448(.A(pi0788), .Y(new_n11885_));
  INVX1    g09449(.A(pi0789), .Y(new_n11886_));
  INVX1    g09450(.A(pi0781), .Y(new_n11887_));
  INVX1    g09451(.A(pi0785), .Y(new_n11888_));
  INVX1    g09452(.A(pi0778), .Y(new_n11889_));
  INVX1    g09453(.A(pi0761), .Y(new_n11890_));
  AND2X1   g09454(.A(new_n8453_), .B(new_n2578_), .Y(new_n11891_));
  NOR3X1   g09455(.A(new_n11891_), .B(new_n2603_), .C(pi0098), .Y(new_n11892_));
  NOR3X1   g09456(.A(new_n8252_), .B(new_n2476_), .C(pi0088), .Y(new_n11893_));
  AND2X1   g09457(.A(new_n6972_), .B(new_n6769_), .Y(new_n11894_));
  NAND3X1  g09458(.A(new_n11894_), .B(new_n11893_), .C(new_n11892_), .Y(new_n11895_));
  AOI21X1  g09459(.A0(new_n11895_), .A1(new_n2549_), .B0(new_n7750_), .Y(new_n11896_));
  OR2X1    g09460(.A(new_n11896_), .B(pi0252), .Y(new_n11897_));
  NOR3X1   g09461(.A(new_n2570_), .B(new_n2744_), .C(pi0091), .Y(new_n11898_));
  INVX1    g09462(.A(new_n11893_), .Y(new_n11899_));
  OR4X1    g09463(.A(new_n11899_), .B(new_n11891_), .C(new_n2603_), .D(pi0098), .Y(new_n11900_));
  OAI21X1  g09464(.A0(new_n11900_), .A1(new_n10474_), .B0(new_n2567_), .Y(new_n11901_));
  NOR3X1   g09465(.A(new_n7731_), .B(new_n2583_), .C(new_n7734_), .Y(new_n11902_));
  OAI21X1  g09466(.A0(new_n11902_), .A1(new_n11901_), .B0(new_n11898_), .Y(new_n11903_));
  NAND2X1  g09467(.A(new_n7744_), .B(new_n2549_), .Y(new_n11904_));
  AOI21X1  g09468(.A0(new_n11903_), .A1(new_n2518_), .B0(new_n11904_), .Y(new_n11905_));
  NAND2X1  g09469(.A(new_n7639_), .B(pi0252), .Y(new_n11906_));
  OAI21X1  g09470(.A0(new_n11906_), .A1(new_n11905_), .B0(new_n11897_), .Y(new_n11907_));
  OR4X1    g09471(.A(new_n11907_), .B(new_n9046_), .C(new_n7272_), .D(new_n2755_), .Y(new_n11908_));
  INVX1    g09472(.A(new_n2569_), .Y(new_n11909_));
  OAI21X1  g09473(.A0(new_n11892_), .A1(pi0088), .B0(new_n8260_), .Y(new_n11910_));
  NOR2X1   g09474(.A(new_n11910_), .B(new_n11909_), .Y(new_n11911_));
  OR2X1    g09475(.A(new_n11902_), .B(pi0047), .Y(new_n11912_));
  OAI21X1  g09476(.A0(new_n11912_), .A1(new_n11911_), .B0(new_n11898_), .Y(new_n11913_));
  NAND2X1  g09477(.A(new_n7744_), .B(pi0252), .Y(new_n11914_));
  AOI21X1  g09478(.A0(new_n11913_), .A1(new_n2518_), .B0(new_n11914_), .Y(new_n11915_));
  NOR2X1   g09479(.A(new_n7057_), .B(pi0252), .Y(new_n11916_));
  INVX1    g09480(.A(new_n11916_), .Y(new_n11917_));
  OAI21X1  g09481(.A0(new_n11917_), .A1(new_n11910_), .B0(new_n2549_), .Y(new_n11918_));
  NOR2X1   g09482(.A(new_n7750_), .B(new_n5939_), .Y(new_n11919_));
  OAI21X1  g09483(.A0(new_n11918_), .A1(new_n11915_), .B0(new_n11919_), .Y(new_n11920_));
  AOI21X1  g09484(.A0(new_n11920_), .A1(new_n11908_), .B0(new_n2756_), .Y(new_n11921_));
  OR2X1    g09485(.A(new_n11907_), .B(new_n7272_), .Y(new_n11922_));
  INVX1    g09486(.A(new_n2781_), .Y(new_n11923_));
  NOR4X1   g09487(.A(new_n11923_), .B(new_n2755_), .C(new_n2780_), .D(pi0833), .Y(po1106));
  INVX1    g09488(.A(po1106), .Y(new_n11925_));
  OAI21X1  g09489(.A0(new_n11925_), .A1(new_n11922_), .B0(new_n2724_), .Y(new_n11926_));
  OAI21X1  g09490(.A0(new_n11921_), .A1(new_n2829_), .B0(new_n11926_), .Y(new_n11927_));
  NAND2X1  g09491(.A(new_n11921_), .B(new_n2722_), .Y(new_n11928_));
  NAND3X1  g09492(.A(new_n11928_), .B(new_n11927_), .C(new_n2766_), .Y(new_n11929_));
  NOR4X1   g09493(.A(new_n11907_), .B(new_n9046_), .C(new_n7272_), .D(new_n2755_), .Y(new_n11930_));
  OAI22X1  g09494(.A0(new_n11918_), .A1(new_n11915_), .B0(new_n2545_), .B1(new_n2549_), .Y(new_n11931_));
  NOR3X1   g09495(.A(new_n5194_), .B(new_n2768_), .C(new_n5193_), .Y(new_n11932_));
  AND2X1   g09496(.A(new_n2783_), .B(new_n2540_), .Y(new_n11933_));
  OAI21X1  g09497(.A0(new_n11932_), .A1(new_n2456_), .B0(new_n11933_), .Y(new_n11934_));
  AOI21X1  g09498(.A0(new_n11931_), .A1(new_n2456_), .B0(new_n11934_), .Y(new_n11935_));
  AOI21X1  g09499(.A0(new_n11935_), .A1(pi0824), .B0(new_n11930_), .Y(new_n11936_));
  OR2X1    g09500(.A(new_n11936_), .B(new_n5983_), .Y(new_n11937_));
  AOI21X1  g09501(.A0(new_n11907_), .A1(new_n2456_), .B0(new_n11934_), .Y(new_n11938_));
  NAND3X1  g09502(.A(new_n11938_), .B(pi0829), .C(new_n5251_), .Y(new_n11939_));
  AOI21X1  g09503(.A0(new_n11939_), .A1(new_n11936_), .B0(new_n2756_), .Y(new_n11940_));
  OAI21X1  g09504(.A0(new_n11940_), .A1(new_n2829_), .B0(new_n11926_), .Y(new_n11941_));
  NAND3X1  g09505(.A(new_n11941_), .B(new_n11937_), .C(pi0210), .Y(new_n11942_));
  AND2X1   g09506(.A(new_n11942_), .B(new_n11929_), .Y(new_n11943_));
  NAND3X1  g09507(.A(new_n11928_), .B(new_n11927_), .C(new_n2973_), .Y(new_n11944_));
  NAND3X1  g09508(.A(new_n11941_), .B(new_n11937_), .C(pi0198), .Y(new_n11945_));
  AND2X1   g09509(.A(new_n11945_), .B(new_n11944_), .Y(new_n11946_));
  MX2X1    g09510(.A(new_n11946_), .B(new_n11943_), .S0(pi0299), .Y(new_n11947_));
  INVX1    g09511(.A(new_n11947_), .Y(new_n11948_));
  INVX1    g09512(.A(pi0681), .Y(new_n11949_));
  INVX1    g09513(.A(pi0616), .Y(new_n11950_));
  OR4X1    g09514(.A(new_n7691_), .B(new_n3003_), .C(new_n2555_), .D(pi0287), .Y(new_n11951_));
  MX2X1    g09515(.A(new_n11951_), .B(new_n3074_), .S0(pi0120), .Y(new_n11952_));
  OR2X1    g09516(.A(new_n11952_), .B(new_n2740_), .Y(new_n11953_));
  OAI21X1  g09517(.A0(new_n11951_), .A1(new_n2740_), .B0(new_n10174_), .Y(new_n11954_));
  NOR2X1   g09518(.A(new_n10339_), .B(new_n5040_), .Y(new_n11955_));
  OR4X1    g09519(.A(new_n11955_), .B(new_n3003_), .C(new_n2740_), .D(new_n2555_), .Y(new_n11956_));
  AOI21X1  g09520(.A0(new_n11956_), .A1(pi0120), .B0(new_n2722_), .Y(new_n11957_));
  AND2X1   g09521(.A(new_n11957_), .B(new_n11954_), .Y(new_n11958_));
  NOR4X1   g09522(.A(new_n7691_), .B(new_n3003_), .C(new_n2555_), .D(pi0287), .Y(new_n11959_));
  AOI21X1  g09523(.A0(new_n11959_), .A1(new_n2739_), .B0(pi0120), .Y(new_n11960_));
  NOR3X1   g09524(.A(new_n3003_), .B(new_n2740_), .C(new_n2555_), .Y(new_n11961_));
  OAI21X1  g09525(.A0(new_n11961_), .A1(new_n10174_), .B0(new_n2722_), .Y(new_n11962_));
  NOR3X1   g09526(.A(new_n5040_), .B(new_n5251_), .C(new_n10174_), .Y(new_n11963_));
  NOR3X1   g09527(.A(new_n11963_), .B(new_n11962_), .C(new_n11960_), .Y(new_n11964_));
  NOR2X1   g09528(.A(new_n11964_), .B(new_n11958_), .Y(new_n11965_));
  MX2X1    g09529(.A(new_n11965_), .B(new_n11953_), .S0(new_n5057_), .Y(new_n11966_));
  OAI22X1  g09530(.A0(new_n11952_), .A1(new_n2740_), .B0(pi0642), .B1(new_n5027_), .Y(new_n11967_));
  INVX1    g09531(.A(pi0642), .Y(new_n11968_));
  AND2X1   g09532(.A(new_n11968_), .B(pi0603), .Y(new_n11969_));
  NOR3X1   g09533(.A(new_n11964_), .B(new_n11958_), .C(new_n5033_), .Y(new_n11970_));
  AND2X1   g09534(.A(new_n11953_), .B(new_n5033_), .Y(new_n11971_));
  OAI21X1  g09535(.A0(new_n11971_), .A1(new_n11970_), .B0(new_n11969_), .Y(new_n11972_));
  AOI21X1  g09536(.A0(new_n11972_), .A1(new_n11967_), .B0(pi0614), .Y(new_n11973_));
  AOI21X1  g09537(.A0(new_n11973_), .A1(new_n11950_), .B0(new_n11966_), .Y(new_n11974_));
  NOR2X1   g09538(.A(new_n11974_), .B(new_n11949_), .Y(new_n11975_));
  INVX1    g09539(.A(pi0661), .Y(new_n11976_));
  INVX1    g09540(.A(pi0662), .Y(new_n11977_));
  AND2X1   g09541(.A(pi0680), .B(new_n11977_), .Y(new_n11978_));
  OAI21X1  g09542(.A0(new_n11952_), .A1(new_n2740_), .B0(pi0616), .Y(new_n11979_));
  AND2X1   g09543(.A(new_n11953_), .B(pi0614), .Y(new_n11980_));
  OAI21X1  g09544(.A0(new_n11980_), .A1(new_n11973_), .B0(new_n11950_), .Y(new_n11981_));
  AOI21X1  g09545(.A0(new_n11981_), .A1(new_n11979_), .B0(new_n11978_), .Y(new_n11982_));
  INVX1    g09546(.A(new_n11978_), .Y(new_n11983_));
  NOR3X1   g09547(.A(new_n11964_), .B(new_n11958_), .C(new_n11983_), .Y(new_n11984_));
  OR2X1    g09548(.A(new_n11984_), .B(new_n5033_), .Y(new_n11985_));
  OAI22X1  g09549(.A0(new_n11985_), .A1(new_n11982_), .B0(new_n11965_), .B1(new_n5057_), .Y(new_n11986_));
  AND2X1   g09550(.A(new_n11973_), .B(new_n11950_), .Y(new_n11987_));
  OR2X1    g09551(.A(new_n11987_), .B(new_n11966_), .Y(new_n11988_));
  OAI21X1  g09552(.A0(new_n11988_), .A1(new_n11976_), .B0(new_n11949_), .Y(new_n11989_));
  AOI21X1  g09553(.A0(new_n11986_), .A1(new_n11976_), .B0(new_n11989_), .Y(new_n11990_));
  OR2X1    g09554(.A(new_n11990_), .B(new_n11975_), .Y(new_n11991_));
  AOI21X1  g09555(.A0(new_n11981_), .A1(new_n11979_), .B0(new_n11949_), .Y(new_n11992_));
  NOR3X1   g09556(.A(pi0681), .B(pi0662), .C(pi0661), .Y(new_n11993_));
  NOR2X1   g09557(.A(new_n11993_), .B(pi0616), .Y(new_n11994_));
  INVX1    g09558(.A(new_n11994_), .Y(new_n11995_));
  NOR3X1   g09559(.A(new_n11995_), .B(new_n11980_), .C(new_n11973_), .Y(new_n11996_));
  OR2X1    g09560(.A(new_n11980_), .B(new_n11973_), .Y(new_n11997_));
  AND2X1   g09561(.A(new_n11997_), .B(new_n11950_), .Y(new_n11998_));
  OAI21X1  g09562(.A0(new_n11971_), .A1(new_n11970_), .B0(pi0680), .Y(new_n11999_));
  NOR4X1   g09563(.A(pi0681), .B(pi0662), .C(pi0661), .D(pi0616), .Y(new_n12000_));
  NAND2X1  g09564(.A(new_n12000_), .B(new_n11999_), .Y(new_n12001_));
  AOI21X1  g09565(.A0(new_n11998_), .A1(new_n5029_), .B0(new_n12001_), .Y(new_n12002_));
  INVX1    g09566(.A(new_n11999_), .Y(new_n12003_));
  OAI21X1  g09567(.A0(new_n11952_), .A1(new_n2740_), .B0(new_n5029_), .Y(new_n12004_));
  NAND3X1  g09568(.A(new_n12004_), .B(new_n11993_), .C(pi0616), .Y(new_n12005_));
  OR4X1    g09569(.A(new_n11952_), .B(new_n2756_), .C(new_n2755_), .D(new_n11950_), .Y(new_n12006_));
  OAI22X1  g09570(.A0(new_n12006_), .A1(new_n11993_), .B0(new_n12005_), .B1(new_n12003_), .Y(new_n12007_));
  NOR4X1   g09571(.A(new_n12007_), .B(new_n12002_), .C(new_n11996_), .D(pi0681), .Y(new_n12008_));
  OR2X1    g09572(.A(new_n12008_), .B(new_n11992_), .Y(new_n12009_));
  MX2X1    g09573(.A(new_n12009_), .B(new_n11991_), .S0(new_n5051_), .Y(new_n12010_));
  AND2X1   g09574(.A(new_n12010_), .B(pi0223), .Y(new_n12011_));
  INVX1    g09575(.A(new_n11953_), .Y(new_n12012_));
  NOR2X1   g09576(.A(new_n11961_), .B(new_n10174_), .Y(new_n12013_));
  OR2X1    g09577(.A(new_n11959_), .B(pi0824), .Y(new_n12014_));
  INVX1    g09578(.A(new_n8278_), .Y(new_n12015_));
  OR4X1    g09579(.A(new_n7694_), .B(new_n3003_), .C(new_n2555_), .D(pi0287), .Y(new_n12016_));
  OAI21X1  g09580(.A0(new_n12016_), .A1(new_n2755_), .B0(new_n12015_), .Y(new_n12017_));
  NAND3X1  g09581(.A(new_n12017_), .B(new_n12014_), .C(pi1093), .Y(new_n12018_));
  AND2X1   g09582(.A(new_n12018_), .B(new_n10174_), .Y(new_n12019_));
  OR2X1    g09583(.A(new_n12019_), .B(new_n11962_), .Y(new_n12020_));
  NAND3X1  g09584(.A(new_n11959_), .B(new_n2739_), .C(new_n2829_), .Y(new_n12021_));
  AOI21X1  g09585(.A0(new_n12017_), .A1(new_n12014_), .B0(pi0829), .Y(new_n12022_));
  NOR4X1   g09586(.A(new_n7694_), .B(new_n3003_), .C(new_n2555_), .D(pi0287), .Y(new_n12023_));
  AOI21X1  g09587(.A0(new_n12023_), .A1(pi1092), .B0(new_n5258_), .Y(new_n12024_));
  OR2X1    g09588(.A(new_n12024_), .B(new_n10308_), .Y(new_n12025_));
  OAI21X1  g09589(.A0(new_n12025_), .A1(new_n12022_), .B0(new_n12021_), .Y(new_n12026_));
  AOI21X1  g09590(.A0(new_n12026_), .A1(pi1091), .B0(pi0120), .Y(new_n12027_));
  OAI21X1  g09591(.A0(new_n12027_), .A1(new_n12013_), .B0(new_n12020_), .Y(new_n12028_));
  MX2X1    g09592(.A(new_n12028_), .B(new_n12012_), .S0(new_n5033_), .Y(new_n12029_));
  MX2X1    g09593(.A(new_n12029_), .B(new_n12012_), .S0(new_n5027_), .Y(new_n12030_));
  OAI21X1  g09594(.A0(new_n12030_), .A1(pi0642), .B0(new_n11967_), .Y(new_n12031_));
  MX2X1    g09595(.A(new_n12031_), .B(new_n11953_), .S0(pi0614), .Y(new_n12032_));
  MX2X1    g09596(.A(new_n12032_), .B(new_n11953_), .S0(pi0616), .Y(new_n12033_));
  NOR2X1   g09597(.A(new_n5030_), .B(pi0614), .Y(new_n12034_));
  NAND2X1  g09598(.A(new_n12034_), .B(new_n11979_), .Y(new_n12035_));
  AOI21X1  g09599(.A0(new_n12031_), .A1(new_n11950_), .B0(new_n12035_), .Y(new_n12036_));
  INVX1    g09600(.A(new_n12013_), .Y(new_n12037_));
  AOI21X1  g09601(.A0(new_n12018_), .A1(new_n10174_), .B0(new_n11962_), .Y(new_n12038_));
  NOR3X1   g09602(.A(new_n11951_), .B(new_n2740_), .C(new_n8273_), .Y(new_n12039_));
  AND2X1   g09603(.A(new_n11951_), .B(new_n5251_), .Y(new_n12040_));
  AOI21X1  g09604(.A0(new_n12023_), .A1(pi1092), .B0(new_n8278_), .Y(new_n12041_));
  OAI21X1  g09605(.A0(new_n12041_), .A1(new_n12040_), .B0(new_n5258_), .Y(new_n12042_));
  NOR2X1   g09606(.A(new_n12024_), .B(new_n10308_), .Y(new_n12043_));
  AOI21X1  g09607(.A0(new_n12043_), .A1(new_n12042_), .B0(new_n12039_), .Y(new_n12044_));
  OAI21X1  g09608(.A0(new_n12044_), .A1(new_n2722_), .B0(new_n10174_), .Y(new_n12045_));
  AOI21X1  g09609(.A0(new_n12045_), .A1(new_n12037_), .B0(new_n12038_), .Y(new_n12046_));
  MX2X1    g09610(.A(new_n12046_), .B(new_n11953_), .S0(new_n5033_), .Y(new_n12047_));
  NOR3X1   g09611(.A(new_n12047_), .B(new_n5282_), .C(pi0614), .Y(new_n12048_));
  NAND3X1  g09612(.A(new_n12004_), .B(new_n11993_), .C(pi0614), .Y(new_n12049_));
  AOI21X1  g09613(.A0(new_n12047_), .A1(pi0680), .B0(new_n12049_), .Y(new_n12050_));
  INVX1    g09614(.A(pi0614), .Y(new_n12051_));
  NOR4X1   g09615(.A(new_n11993_), .B(new_n11952_), .C(new_n2740_), .D(new_n12051_), .Y(new_n12052_));
  OR2X1    g09616(.A(new_n12052_), .B(new_n12050_), .Y(new_n12053_));
  NOR4X1   g09617(.A(new_n12053_), .B(new_n12048_), .C(new_n12036_), .D(pi0681), .Y(new_n12054_));
  AOI21X1  g09618(.A0(new_n12033_), .A1(pi0681), .B0(new_n12054_), .Y(new_n12055_));
  MX2X1    g09619(.A(new_n12028_), .B(new_n12012_), .S0(new_n5057_), .Y(new_n12056_));
  MX2X1    g09620(.A(new_n12056_), .B(new_n12028_), .S0(new_n5028_), .Y(new_n12057_));
  NOR2X1   g09621(.A(new_n12057_), .B(new_n11949_), .Y(new_n12058_));
  NOR3X1   g09622(.A(new_n5029_), .B(pi0662), .C(pi0661), .Y(new_n12059_));
  INVX1    g09623(.A(new_n12059_), .Y(new_n12060_));
  OAI21X1  g09624(.A0(new_n12046_), .A1(new_n12060_), .B0(new_n11949_), .Y(new_n12061_));
  AOI21X1  g09625(.A0(new_n12057_), .A1(new_n12060_), .B0(new_n12061_), .Y(new_n12062_));
  NOR2X1   g09626(.A(new_n12062_), .B(new_n12058_), .Y(new_n12063_));
  MX2X1    g09627(.A(new_n12063_), .B(new_n12055_), .S0(new_n5050_), .Y(new_n12064_));
  NOR3X1   g09628(.A(new_n11952_), .B(new_n2971_), .C(new_n2740_), .Y(new_n12065_));
  OR2X1    g09629(.A(new_n12065_), .B(pi0223), .Y(new_n12066_));
  AOI21X1  g09630(.A0(new_n12064_), .A1(new_n2971_), .B0(new_n12066_), .Y(new_n12067_));
  OAI21X1  g09631(.A0(new_n12067_), .A1(new_n12011_), .B0(new_n2953_), .Y(new_n12068_));
  INVX1    g09632(.A(new_n5069_), .Y(new_n12069_));
  AOI21X1  g09633(.A0(new_n12031_), .A1(new_n12051_), .B0(new_n11980_), .Y(new_n12070_));
  MX2X1    g09634(.A(new_n12070_), .B(new_n12012_), .S0(pi0616), .Y(new_n12071_));
  OR4X1    g09635(.A(new_n12053_), .B(new_n12048_), .C(new_n12036_), .D(pi0681), .Y(new_n12072_));
  OAI21X1  g09636(.A0(new_n12071_), .A1(new_n11949_), .B0(new_n12072_), .Y(new_n12073_));
  OAI21X1  g09637(.A0(new_n12063_), .A1(new_n12069_), .B0(new_n5064_), .Y(new_n12074_));
  AOI21X1  g09638(.A0(new_n12073_), .A1(new_n12069_), .B0(new_n12074_), .Y(new_n12075_));
  NOR4X1   g09639(.A(new_n12062_), .B(new_n12058_), .C(new_n5064_), .D(new_n10136_), .Y(new_n12076_));
  NOR3X1   g09640(.A(new_n11952_), .B(new_n10137_), .C(new_n2740_), .Y(new_n12077_));
  OR2X1    g09641(.A(new_n12077_), .B(pi0215), .Y(new_n12078_));
  OR2X1    g09642(.A(new_n12078_), .B(new_n12076_), .Y(new_n12079_));
  AOI21X1  g09643(.A0(new_n12075_), .A1(new_n10137_), .B0(new_n12079_), .Y(new_n12080_));
  OR2X1    g09644(.A(new_n11991_), .B(new_n5064_), .Y(new_n12081_));
  NOR2X1   g09645(.A(new_n11990_), .B(new_n11975_), .Y(new_n12082_));
  NOR2X1   g09646(.A(new_n12082_), .B(new_n12069_), .Y(new_n12083_));
  NOR2X1   g09647(.A(new_n12008_), .B(new_n11992_), .Y(new_n12084_));
  OAI21X1  g09648(.A0(new_n12084_), .A1(new_n5069_), .B0(new_n5064_), .Y(new_n12085_));
  OAI21X1  g09649(.A0(new_n12085_), .A1(new_n12083_), .B0(new_n12081_), .Y(new_n12086_));
  NOR2X1   g09650(.A(new_n12086_), .B(new_n2954_), .Y(new_n12087_));
  OAI21X1  g09651(.A0(new_n12087_), .A1(new_n12080_), .B0(pi0299), .Y(new_n12088_));
  NAND2X1  g09652(.A(new_n12088_), .B(new_n12068_), .Y(new_n12089_));
  MX2X1    g09653(.A(new_n12089_), .B(new_n11948_), .S0(new_n2959_), .Y(new_n12090_));
  NAND2X1  g09654(.A(new_n11942_), .B(new_n11929_), .Y(new_n12091_));
  INVX1    g09655(.A(pi0621), .Y(new_n12092_));
  NOR2X1   g09656(.A(new_n11927_), .B(new_n12092_), .Y(new_n12093_));
  INVX1    g09657(.A(new_n12093_), .Y(new_n12094_));
  OR2X1    g09658(.A(new_n11941_), .B(new_n12092_), .Y(new_n12095_));
  MX2X1    g09659(.A(new_n12095_), .B(new_n12094_), .S0(new_n2766_), .Y(new_n12096_));
  AOI21X1  g09660(.A0(new_n12096_), .A1(pi0603), .B0(new_n12091_), .Y(new_n12097_));
  MX2X1    g09661(.A(new_n12095_), .B(new_n12094_), .S0(new_n2973_), .Y(new_n12098_));
  OAI21X1  g09662(.A0(new_n11927_), .A1(pi0621), .B0(new_n11928_), .Y(new_n12099_));
  AND2X1   g09663(.A(new_n12099_), .B(new_n2973_), .Y(new_n12100_));
  OAI21X1  g09664(.A0(new_n11941_), .A1(pi0621), .B0(new_n11937_), .Y(new_n12101_));
  AOI21X1  g09665(.A0(new_n12101_), .A1(pi0198), .B0(new_n12100_), .Y(new_n12102_));
  OAI21X1  g09666(.A0(new_n12102_), .A1(pi0603), .B0(new_n12098_), .Y(new_n12103_));
  MX2X1    g09667(.A(new_n12103_), .B(new_n12097_), .S0(pi0299), .Y(new_n12104_));
  NOR2X1   g09668(.A(new_n12104_), .B(pi0039), .Y(new_n12105_));
  MX2X1    g09669(.A(new_n12057_), .B(new_n12028_), .S0(new_n5030_), .Y(new_n12106_));
  MX2X1    g09670(.A(new_n12046_), .B(new_n11953_), .S0(new_n5057_), .Y(new_n12107_));
  AND2X1   g09671(.A(pi1091), .B(pi0621), .Y(new_n12108_));
  INVX1    g09672(.A(new_n12108_), .Y(new_n12109_));
  NOR4X1   g09673(.A(new_n12109_), .B(new_n12027_), .C(new_n12013_), .D(new_n5057_), .Y(new_n12110_));
  NOR4X1   g09674(.A(new_n12109_), .B(new_n11952_), .C(new_n5033_), .D(new_n2740_), .Y(new_n12111_));
  OR2X1    g09675(.A(new_n12111_), .B(new_n5027_), .Y(new_n12112_));
  NOR2X1   g09676(.A(new_n12112_), .B(new_n12110_), .Y(new_n12113_));
  AOI21X1  g09677(.A0(new_n12107_), .A1(new_n5027_), .B0(new_n12113_), .Y(new_n12114_));
  NAND3X1  g09678(.A(new_n12108_), .B(new_n12045_), .C(new_n12037_), .Y(new_n12115_));
  OAI21X1  g09679(.A0(new_n12038_), .A1(new_n12092_), .B0(new_n12028_), .Y(new_n12116_));
  OAI21X1  g09680(.A0(new_n12116_), .A1(pi0603), .B0(new_n12115_), .Y(new_n12117_));
  OR2X1    g09681(.A(new_n12117_), .B(new_n12114_), .Y(new_n12118_));
  AOI21X1  g09682(.A0(new_n12118_), .A1(new_n12106_), .B0(new_n5070_), .Y(new_n12119_));
  NOR2X1   g09683(.A(new_n12108_), .B(new_n5027_), .Y(new_n12120_));
  OR4X1    g09684(.A(new_n12120_), .B(new_n11952_), .C(new_n2756_), .D(new_n2755_), .Y(new_n12121_));
  OR4X1    g09685(.A(new_n12109_), .B(new_n11952_), .C(new_n2756_), .D(new_n2755_), .Y(new_n12122_));
  MX2X1    g09686(.A(new_n12122_), .B(new_n12115_), .S0(new_n5057_), .Y(new_n12123_));
  AOI21X1  g09687(.A0(new_n12123_), .A1(pi0603), .B0(new_n12047_), .Y(new_n12124_));
  NOR3X1   g09688(.A(pi0642), .B(pi0616), .C(pi0614), .Y(new_n12125_));
  NOR4X1   g09689(.A(new_n12120_), .B(new_n12125_), .C(new_n11952_), .D(new_n2740_), .Y(new_n12126_));
  INVX1    g09690(.A(new_n12125_), .Y(new_n12127_));
  AOI21X1  g09691(.A0(new_n11953_), .A1(new_n5027_), .B0(new_n12127_), .Y(new_n12128_));
  INVX1    g09692(.A(new_n12128_), .Y(new_n12129_));
  AOI21X1  g09693(.A0(new_n12123_), .A1(pi0603), .B0(new_n12129_), .Y(new_n12130_));
  OR2X1    g09694(.A(new_n12130_), .B(new_n12126_), .Y(new_n12131_));
  MX2X1    g09695(.A(new_n12131_), .B(new_n12124_), .S0(new_n5030_), .Y(new_n12132_));
  OAI21X1  g09696(.A0(new_n12132_), .A1(new_n5071_), .B0(new_n10137_), .Y(new_n12133_));
  OAI22X1  g09697(.A0(new_n12133_), .A1(new_n12119_), .B0(new_n12121_), .B1(new_n10137_), .Y(new_n12134_));
  NOR2X1   g09698(.A(new_n11971_), .B(new_n11970_), .Y(new_n12135_));
  AND2X1   g09699(.A(new_n12122_), .B(new_n5033_), .Y(new_n12136_));
  NAND3X1  g09700(.A(new_n11957_), .B(new_n11954_), .C(pi0621), .Y(new_n12137_));
  AOI21X1  g09701(.A0(new_n12137_), .A1(new_n5057_), .B0(new_n12136_), .Y(new_n12138_));
  OR2X1    g09702(.A(new_n12138_), .B(new_n5027_), .Y(new_n12139_));
  NAND3X1  g09703(.A(new_n12139_), .B(new_n12135_), .C(new_n5030_), .Y(new_n12140_));
  AOI21X1  g09704(.A0(new_n12139_), .A1(new_n12128_), .B0(new_n12126_), .Y(new_n12141_));
  OAI21X1  g09705(.A0(new_n12141_), .A1(new_n5030_), .B0(new_n12140_), .Y(new_n12142_));
  OR2X1    g09706(.A(new_n12142_), .B(new_n5071_), .Y(new_n12143_));
  OR2X1    g09707(.A(new_n11964_), .B(new_n11958_), .Y(new_n12144_));
  MX2X1    g09708(.A(new_n12144_), .B(new_n12012_), .S0(new_n5057_), .Y(new_n12145_));
  NOR2X1   g09709(.A(new_n12120_), .B(new_n2740_), .Y(new_n12146_));
  AND2X1   g09710(.A(new_n12146_), .B(new_n12145_), .Y(new_n12147_));
  OAI21X1  g09711(.A0(new_n11958_), .A1(new_n5367_), .B0(new_n12147_), .Y(new_n12148_));
  OAI21X1  g09712(.A0(new_n11964_), .A1(new_n11958_), .B0(new_n12146_), .Y(new_n12149_));
  AND2X1   g09713(.A(new_n12149_), .B(new_n5030_), .Y(new_n12150_));
  AOI21X1  g09714(.A0(new_n12148_), .A1(new_n5282_), .B0(new_n12150_), .Y(new_n12151_));
  INVX1    g09715(.A(new_n12151_), .Y(new_n12152_));
  AOI21X1  g09716(.A0(new_n12152_), .A1(new_n5071_), .B0(new_n2954_), .Y(new_n12153_));
  AOI22X1  g09717(.A0(new_n12153_), .A1(new_n12143_), .B0(new_n12134_), .B1(new_n2954_), .Y(new_n12154_));
  AOI21X1  g09718(.A0(new_n12118_), .A1(new_n12106_), .B0(new_n5050_), .Y(new_n12155_));
  OAI21X1  g09719(.A0(new_n12132_), .A1(new_n5051_), .B0(new_n2971_), .Y(new_n12156_));
  OAI22X1  g09720(.A0(new_n12156_), .A1(new_n12155_), .B0(new_n12121_), .B1(new_n2971_), .Y(new_n12157_));
  OR2X1    g09721(.A(new_n12142_), .B(new_n5051_), .Y(new_n12158_));
  AOI21X1  g09722(.A0(new_n12152_), .A1(new_n5051_), .B0(new_n2964_), .Y(new_n12159_));
  AOI22X1  g09723(.A0(new_n12159_), .A1(new_n12158_), .B0(new_n12157_), .B1(new_n2964_), .Y(new_n12160_));
  MX2X1    g09724(.A(new_n12160_), .B(new_n12154_), .S0(pi0299), .Y(new_n12161_));
  AOI21X1  g09725(.A0(new_n12161_), .A1(pi0039), .B0(new_n12105_), .Y(new_n12162_));
  AOI21X1  g09726(.A0(new_n12162_), .A1(new_n11890_), .B0(pi0140), .Y(new_n12163_));
  OAI21X1  g09727(.A0(new_n12090_), .A1(new_n11890_), .B0(new_n12163_), .Y(new_n12164_));
  NOR2X1   g09728(.A(new_n12102_), .B(new_n5027_), .Y(new_n12165_));
  MX2X1    g09729(.A(new_n12101_), .B(new_n12099_), .S0(new_n2766_), .Y(new_n12166_));
  AND2X1   g09730(.A(new_n12166_), .B(pi0603), .Y(new_n12167_));
  MX2X1    g09731(.A(new_n12167_), .B(new_n12165_), .S0(new_n2953_), .Y(new_n12168_));
  NOR2X1   g09732(.A(new_n12168_), .B(pi0039), .Y(new_n12169_));
  AND2X1   g09733(.A(new_n12120_), .B(new_n12029_), .Y(new_n12170_));
  INVX1    g09734(.A(new_n12120_), .Y(new_n12171_));
  NOR3X1   g09735(.A(new_n12171_), .B(new_n11952_), .C(new_n2740_), .Y(new_n12172_));
  MX2X1    g09736(.A(new_n12172_), .B(new_n12170_), .S0(new_n12125_), .Y(new_n12173_));
  MX2X1    g09737(.A(new_n12173_), .B(new_n12170_), .S0(new_n5030_), .Y(new_n12174_));
  NAND2X1  g09738(.A(new_n12120_), .B(new_n12106_), .Y(new_n12175_));
  AOI21X1  g09739(.A0(new_n12175_), .A1(new_n5071_), .B0(new_n10136_), .Y(new_n12176_));
  OAI21X1  g09740(.A0(new_n12174_), .A1(new_n5071_), .B0(new_n12176_), .Y(new_n12177_));
  NOR4X1   g09741(.A(new_n12108_), .B(new_n2756_), .C(new_n2755_), .D(new_n5027_), .Y(new_n12178_));
  NOR2X1   g09742(.A(new_n11952_), .B(new_n10137_), .Y(new_n12179_));
  AOI21X1  g09743(.A0(new_n12179_), .A1(new_n12178_), .B0(pi0215), .Y(new_n12180_));
  INVX1    g09744(.A(new_n12172_), .Y(new_n12181_));
  NOR2X1   g09745(.A(new_n12181_), .B(new_n11970_), .Y(new_n12182_));
  INVX1    g09746(.A(new_n12182_), .Y(new_n12183_));
  OR4X1    g09747(.A(new_n12127_), .B(new_n11964_), .C(new_n11958_), .D(new_n5033_), .Y(new_n12184_));
  NAND4X1  g09748(.A(new_n12184_), .B(new_n12172_), .C(new_n12145_), .D(new_n5282_), .Y(new_n12185_));
  AND2X1   g09749(.A(new_n11966_), .B(new_n5071_), .Y(new_n12186_));
  AOI21X1  g09750(.A0(new_n12185_), .A1(new_n12183_), .B0(new_n12186_), .Y(new_n12187_));
  OAI21X1  g09751(.A0(new_n12187_), .A1(new_n2954_), .B0(pi0299), .Y(new_n12188_));
  AOI21X1  g09752(.A0(new_n12180_), .A1(new_n12177_), .B0(new_n12188_), .Y(new_n12189_));
  NOR4X1   g09753(.A(new_n12171_), .B(new_n11952_), .C(new_n2971_), .D(new_n2740_), .Y(new_n12190_));
  NOR2X1   g09754(.A(new_n12190_), .B(pi0223), .Y(new_n12191_));
  AOI21X1  g09755(.A0(new_n12175_), .A1(new_n5051_), .B0(new_n2970_), .Y(new_n12192_));
  OAI21X1  g09756(.A0(new_n12174_), .A1(new_n5051_), .B0(new_n12192_), .Y(new_n12193_));
  AND2X1   g09757(.A(new_n11966_), .B(new_n5051_), .Y(new_n12194_));
  AOI21X1  g09758(.A0(new_n12185_), .A1(new_n12183_), .B0(new_n12194_), .Y(new_n12195_));
  OAI21X1  g09759(.A0(new_n12195_), .A1(new_n2964_), .B0(new_n2953_), .Y(new_n12196_));
  AOI21X1  g09760(.A0(new_n12193_), .A1(new_n12191_), .B0(new_n12196_), .Y(new_n12197_));
  NOR2X1   g09761(.A(new_n12197_), .B(new_n12189_), .Y(new_n12198_));
  AOI21X1  g09762(.A0(new_n12198_), .A1(pi0039), .B0(new_n12169_), .Y(new_n12199_));
  NAND3X1  g09763(.A(new_n12199_), .B(new_n11890_), .C(pi0140), .Y(new_n12200_));
  AND2X1   g09764(.A(new_n12200_), .B(new_n12164_), .Y(new_n12201_));
  NOR4X1   g09765(.A(new_n3003_), .B(new_n2740_), .C(new_n2555_), .D(pi0039), .Y(new_n12202_));
  NOR2X1   g09766(.A(new_n12202_), .B(pi0140), .Y(new_n12203_));
  INVX1    g09767(.A(new_n12178_), .Y(new_n12204_));
  NOR4X1   g09768(.A(new_n12204_), .B(new_n3003_), .C(new_n2555_), .D(pi0039), .Y(new_n12205_));
  AOI21X1  g09769(.A0(new_n12205_), .A1(new_n11890_), .B0(new_n12203_), .Y(new_n12206_));
  OR2X1    g09770(.A(new_n12206_), .B(new_n2996_), .Y(new_n12207_));
  OAI21X1  g09771(.A0(new_n12201_), .A1(pi0038), .B0(new_n12207_), .Y(new_n12208_));
  NOR2X1   g09772(.A(new_n11993_), .B(new_n5029_), .Y(new_n12209_));
  AND2X1   g09773(.A(pi1091), .B(pi0665), .Y(new_n12210_));
  NOR2X1   g09774(.A(new_n12210_), .B(new_n12120_), .Y(new_n12211_));
  OR4X1    g09775(.A(new_n12211_), .B(new_n11952_), .C(new_n2756_), .D(new_n2755_), .Y(new_n12212_));
  AND2X1   g09776(.A(new_n12212_), .B(pi0616), .Y(new_n12213_));
  AND2X1   g09777(.A(new_n12212_), .B(pi0614), .Y(new_n12214_));
  INVX1    g09778(.A(new_n12214_), .Y(new_n12215_));
  AND2X1   g09779(.A(new_n12212_), .B(pi0642), .Y(new_n12216_));
  AND2X1   g09780(.A(new_n11958_), .B(pi0665), .Y(new_n12217_));
  AOI21X1  g09781(.A0(new_n12172_), .A1(new_n12144_), .B0(new_n12217_), .Y(new_n12218_));
  INVX1    g09782(.A(new_n12210_), .Y(new_n12219_));
  NOR4X1   g09783(.A(new_n12219_), .B(new_n11952_), .C(new_n5033_), .D(new_n2740_), .Y(new_n12220_));
  INVX1    g09784(.A(new_n12220_), .Y(new_n12221_));
  OAI21X1  g09785(.A0(new_n12221_), .A1(pi0603), .B0(new_n12218_), .Y(new_n12222_));
  NOR3X1   g09786(.A(new_n12219_), .B(new_n11952_), .C(new_n2740_), .Y(new_n12223_));
  MX2X1    g09787(.A(new_n12223_), .B(new_n12217_), .S0(new_n5057_), .Y(new_n12224_));
  NOR4X1   g09788(.A(new_n12224_), .B(new_n12222_), .C(new_n12182_), .D(pi0642), .Y(new_n12225_));
  OAI21X1  g09789(.A0(new_n12225_), .A1(new_n12216_), .B0(new_n12051_), .Y(new_n12226_));
  AOI21X1  g09790(.A0(new_n12226_), .A1(new_n12215_), .B0(pi0616), .Y(new_n12227_));
  OAI21X1  g09791(.A0(new_n12227_), .A1(new_n12213_), .B0(new_n12209_), .Y(new_n12228_));
  AND2X1   g09792(.A(new_n11981_), .B(new_n11979_), .Y(new_n12229_));
  INVX1    g09793(.A(new_n12229_), .Y(new_n12230_));
  NOR3X1   g09794(.A(new_n12224_), .B(new_n12182_), .C(new_n5282_), .Y(new_n12231_));
  AOI21X1  g09795(.A0(new_n12230_), .A1(new_n5029_), .B0(new_n12231_), .Y(new_n12232_));
  AOI21X1  g09796(.A0(new_n12232_), .A1(new_n12228_), .B0(new_n5051_), .Y(new_n12233_));
  NOR2X1   g09797(.A(new_n11974_), .B(pi0680), .Y(new_n12234_));
  INVX1    g09798(.A(new_n12209_), .Y(new_n12235_));
  NAND2X1  g09799(.A(new_n12218_), .B(new_n5030_), .Y(new_n12236_));
  AOI21X1  g09800(.A0(new_n11958_), .A1(pi0665), .B0(new_n12220_), .Y(new_n12237_));
  OAI21X1  g09801(.A0(new_n12181_), .A1(new_n11966_), .B0(new_n12237_), .Y(new_n12238_));
  MX2X1    g09802(.A(new_n12238_), .B(new_n12222_), .S0(new_n12125_), .Y(new_n12239_));
  OAI21X1  g09803(.A0(new_n12239_), .A1(new_n12235_), .B0(new_n12236_), .Y(new_n12240_));
  NOR2X1   g09804(.A(new_n12240_), .B(new_n12234_), .Y(new_n12241_));
  OAI21X1  g09805(.A0(new_n12241_), .A1(new_n5050_), .B0(pi0223), .Y(new_n12242_));
  OR2X1    g09806(.A(new_n12242_), .B(new_n12233_), .Y(new_n12243_));
  INVX1    g09807(.A(new_n12213_), .Y(new_n12244_));
  INVX1    g09808(.A(new_n12216_), .Y(new_n12245_));
  MX2X1    g09809(.A(new_n12047_), .B(new_n11953_), .S0(new_n5027_), .Y(new_n12246_));
  OAI21X1  g09810(.A0(new_n12211_), .A1(new_n12246_), .B0(new_n11968_), .Y(new_n12247_));
  AOI21X1  g09811(.A0(new_n12247_), .A1(new_n12245_), .B0(pi0614), .Y(new_n12248_));
  OAI21X1  g09812(.A0(new_n12248_), .A1(new_n12214_), .B0(new_n11950_), .Y(new_n12249_));
  AOI21X1  g09813(.A0(new_n12249_), .A1(new_n12244_), .B0(new_n12235_), .Y(new_n12250_));
  AND2X1   g09814(.A(new_n12033_), .B(new_n5029_), .Y(new_n12251_));
  NOR3X1   g09815(.A(new_n12219_), .B(new_n12027_), .C(new_n12013_), .Y(new_n12252_));
  MX2X1    g09816(.A(new_n12252_), .B(new_n12223_), .S0(new_n5033_), .Y(new_n12253_));
  OR2X1    g09817(.A(new_n12253_), .B(pi0603), .Y(new_n12254_));
  INVX1    g09818(.A(pi0665), .Y(new_n12255_));
  AND2X1   g09819(.A(new_n12255_), .B(pi0603), .Y(new_n12256_));
  AOI22X1  g09820(.A0(new_n12256_), .A1(new_n12108_), .B0(new_n12047_), .B1(pi0603), .Y(new_n12257_));
  AOI21X1  g09821(.A0(new_n12257_), .A1(new_n12254_), .B0(new_n5282_), .Y(new_n12258_));
  NOR4X1   g09822(.A(new_n12258_), .B(new_n12251_), .C(new_n12250_), .D(new_n5051_), .Y(new_n12259_));
  MX2X1    g09823(.A(new_n12107_), .B(new_n12046_), .S0(new_n5028_), .Y(new_n12260_));
  OAI21X1  g09824(.A0(new_n12211_), .A1(new_n12260_), .B0(new_n12209_), .Y(new_n12261_));
  OR2X1    g09825(.A(new_n12116_), .B(new_n5027_), .Y(new_n12262_));
  AND2X1   g09826(.A(new_n12092_), .B(pi0603), .Y(new_n12263_));
  OR4X1    g09827(.A(new_n12263_), .B(new_n12219_), .C(new_n12027_), .D(new_n12013_), .Y(new_n12264_));
  AND2X1   g09828(.A(new_n12264_), .B(new_n5030_), .Y(new_n12265_));
  AOI22X1  g09829(.A0(new_n12265_), .A1(new_n12262_), .B0(new_n12260_), .B1(new_n5029_), .Y(new_n12266_));
  NAND3X1  g09830(.A(new_n12266_), .B(new_n12261_), .C(new_n5051_), .Y(new_n12267_));
  NAND2X1  g09831(.A(new_n12267_), .B(new_n2971_), .Y(new_n12268_));
  NOR3X1   g09832(.A(new_n12210_), .B(new_n12120_), .C(new_n5029_), .Y(new_n12269_));
  NOR3X1   g09833(.A(new_n12269_), .B(new_n11952_), .C(new_n2740_), .Y(new_n12270_));
  INVX1    g09834(.A(new_n12270_), .Y(new_n12271_));
  AOI21X1  g09835(.A0(new_n12271_), .A1(new_n2970_), .B0(pi0223), .Y(new_n12272_));
  OAI21X1  g09836(.A0(new_n12268_), .A1(new_n12259_), .B0(new_n12272_), .Y(new_n12273_));
  AND2X1   g09837(.A(new_n12273_), .B(new_n12243_), .Y(new_n12274_));
  AOI21X1  g09838(.A0(new_n12266_), .A1(new_n12261_), .B0(new_n5070_), .Y(new_n12275_));
  INVX1    g09839(.A(new_n12211_), .Y(new_n12276_));
  AOI21X1  g09840(.A0(new_n12276_), .A1(new_n12030_), .B0(pi0642), .Y(new_n12277_));
  OAI21X1  g09841(.A0(new_n12277_), .A1(new_n12216_), .B0(new_n12051_), .Y(new_n12278_));
  AOI21X1  g09842(.A0(new_n12278_), .A1(new_n12215_), .B0(pi0616), .Y(new_n12279_));
  OAI21X1  g09843(.A0(new_n12279_), .A1(new_n12213_), .B0(new_n12209_), .Y(new_n12280_));
  AOI21X1  g09844(.A0(new_n12033_), .A1(new_n5029_), .B0(new_n12258_), .Y(new_n12281_));
  AOI21X1  g09845(.A0(new_n12281_), .A1(new_n12280_), .B0(new_n5071_), .Y(new_n12282_));
  OAI21X1  g09846(.A0(new_n12282_), .A1(new_n12275_), .B0(new_n10137_), .Y(new_n12283_));
  AOI21X1  g09847(.A0(new_n12271_), .A1(new_n10136_), .B0(pi0215), .Y(new_n12284_));
  AOI21X1  g09848(.A0(new_n12232_), .A1(new_n12228_), .B0(new_n5071_), .Y(new_n12285_));
  OAI21X1  g09849(.A0(new_n12241_), .A1(new_n5070_), .B0(pi0215), .Y(new_n12286_));
  NOR2X1   g09850(.A(new_n12286_), .B(new_n12285_), .Y(new_n12287_));
  AOI21X1  g09851(.A0(new_n12284_), .A1(new_n12283_), .B0(new_n12287_), .Y(new_n12288_));
  MX2X1    g09852(.A(new_n12288_), .B(new_n12274_), .S0(new_n2953_), .Y(new_n12289_));
  INVX1    g09853(.A(new_n11993_), .Y(new_n12290_));
  OAI22X1  g09854(.A0(new_n12112_), .A1(new_n12110_), .B0(new_n12056_), .B1(pi0603), .Y(new_n12291_));
  NOR3X1   g09855(.A(new_n12210_), .B(new_n11952_), .C(new_n2740_), .Y(new_n12292_));
  OR2X1    g09856(.A(new_n12038_), .B(new_n12255_), .Y(new_n12293_));
  AOI21X1  g09857(.A0(new_n12293_), .A1(new_n12028_), .B0(new_n12292_), .Y(new_n12294_));
  OAI21X1  g09858(.A0(new_n12294_), .A1(new_n12291_), .B0(pi0616), .Y(new_n12295_));
  OR2X1    g09859(.A(new_n12294_), .B(new_n12291_), .Y(new_n12296_));
  NOR4X1   g09860(.A(new_n12109_), .B(new_n12027_), .C(new_n12013_), .D(pi0665), .Y(new_n12297_));
  OR2X1    g09861(.A(new_n12297_), .B(new_n5027_), .Y(new_n12298_));
  OAI21X1  g09862(.A0(new_n12294_), .A1(new_n12107_), .B0(new_n5027_), .Y(new_n12299_));
  AOI21X1  g09863(.A0(new_n12299_), .A1(new_n12298_), .B0(new_n12127_), .Y(new_n12300_));
  NOR2X1   g09864(.A(new_n12300_), .B(new_n12296_), .Y(new_n12301_));
  NOR2X1   g09865(.A(pi0642), .B(pi0614), .Y(new_n12302_));
  NAND3X1  g09866(.A(new_n12299_), .B(new_n12298_), .C(new_n12302_), .Y(new_n12303_));
  NAND2X1  g09867(.A(new_n12303_), .B(new_n11950_), .Y(new_n12304_));
  OAI21X1  g09868(.A0(new_n12304_), .A1(new_n12301_), .B0(new_n12295_), .Y(new_n12305_));
  NAND4X1  g09869(.A(new_n12298_), .B(new_n12293_), .C(new_n12028_), .D(new_n5030_), .Y(new_n12306_));
  AOI22X1  g09870(.A0(new_n12306_), .A1(new_n12235_), .B0(new_n12305_), .B1(new_n12290_), .Y(new_n12307_));
  NOR4X1   g09871(.A(new_n12210_), .B(new_n12120_), .C(new_n11952_), .D(new_n2740_), .Y(new_n12308_));
  OR2X1    g09872(.A(new_n12308_), .B(new_n11950_), .Y(new_n12309_));
  AND2X1   g09873(.A(new_n12309_), .B(new_n12209_), .Y(new_n12310_));
  INVX1    g09874(.A(new_n12302_), .Y(new_n12311_));
  AOI21X1  g09875(.A0(new_n12115_), .A1(new_n5057_), .B0(new_n12136_), .Y(new_n12312_));
  MX2X1    g09876(.A(new_n12292_), .B(new_n12255_), .S0(pi0603), .Y(new_n12313_));
  OAI21X1  g09877(.A0(new_n12312_), .A1(new_n5027_), .B0(new_n12313_), .Y(new_n12314_));
  AOI21X1  g09878(.A0(new_n12308_), .A1(new_n12311_), .B0(pi0616), .Y(new_n12315_));
  OAI21X1  g09879(.A0(new_n12314_), .A1(new_n12311_), .B0(new_n12315_), .Y(new_n12316_));
  AOI22X1  g09880(.A0(new_n12316_), .A1(new_n12310_), .B0(new_n12258_), .B1(new_n12029_), .Y(new_n12317_));
  AOI21X1  g09881(.A0(new_n12317_), .A1(new_n5070_), .B0(new_n10136_), .Y(new_n12318_));
  OAI21X1  g09882(.A0(new_n12307_), .A1(new_n5070_), .B0(new_n12318_), .Y(new_n12319_));
  AOI21X1  g09883(.A0(new_n12269_), .A1(new_n12077_), .B0(pi0215), .Y(new_n12320_));
  NAND3X1  g09884(.A(new_n12313_), .B(new_n12146_), .C(new_n12145_), .Y(new_n12321_));
  AND2X1   g09885(.A(new_n12321_), .B(pi0616), .Y(new_n12322_));
  NOR2X1   g09886(.A(pi0616), .B(pi0614), .Y(new_n12323_));
  INVX1    g09887(.A(new_n12323_), .Y(new_n12324_));
  AND2X1   g09888(.A(new_n12313_), .B(new_n12147_), .Y(new_n12325_));
  OR2X1    g09889(.A(pi0616), .B(new_n12051_), .Y(new_n12326_));
  OAI21X1  g09890(.A0(new_n12138_), .A1(new_n5027_), .B0(new_n12313_), .Y(new_n12327_));
  AOI21X1  g09891(.A0(new_n12327_), .A1(new_n11968_), .B0(new_n12321_), .Y(new_n12328_));
  OAI22X1  g09892(.A0(new_n12328_), .A1(new_n12324_), .B0(new_n12326_), .B1(new_n12325_), .Y(new_n12329_));
  OR2X1    g09893(.A(new_n12329_), .B(new_n12322_), .Y(new_n12330_));
  AOI21X1  g09894(.A0(new_n12269_), .A1(new_n12144_), .B0(new_n12209_), .Y(new_n12331_));
  AOI21X1  g09895(.A0(new_n12330_), .A1(new_n12290_), .B0(new_n12331_), .Y(new_n12332_));
  INVX1    g09896(.A(new_n12140_), .Y(new_n12333_));
  OAI21X1  g09897(.A0(new_n12210_), .A1(new_n12141_), .B0(new_n11950_), .Y(new_n12334_));
  AOI22X1  g09898(.A0(new_n12334_), .A1(new_n12310_), .B0(new_n12313_), .B1(new_n12333_), .Y(new_n12335_));
  OAI21X1  g09899(.A0(new_n12335_), .A1(new_n5071_), .B0(pi0215), .Y(new_n12336_));
  AOI21X1  g09900(.A0(new_n12332_), .A1(new_n5071_), .B0(new_n12336_), .Y(new_n12337_));
  AOI21X1  g09901(.A0(new_n12320_), .A1(new_n12319_), .B0(new_n12337_), .Y(new_n12338_));
  OAI21X1  g09902(.A0(new_n12317_), .A1(new_n5051_), .B0(new_n2971_), .Y(new_n12339_));
  AOI21X1  g09903(.A0(new_n12307_), .A1(new_n5051_), .B0(new_n12339_), .Y(new_n12340_));
  NOR2X1   g09904(.A(new_n12210_), .B(new_n5029_), .Y(new_n12341_));
  OAI21X1  g09905(.A0(new_n12341_), .A1(new_n12120_), .B0(new_n2739_), .Y(new_n12342_));
  NOR3X1   g09906(.A(new_n12342_), .B(new_n11952_), .C(new_n2740_), .Y(new_n12343_));
  NOR2X1   g09907(.A(new_n12343_), .B(new_n2971_), .Y(new_n12344_));
  NOR4X1   g09908(.A(new_n12344_), .B(new_n12340_), .C(new_n12190_), .D(pi0223), .Y(new_n12345_));
  AOI21X1  g09909(.A0(new_n12335_), .A1(new_n5050_), .B0(new_n2964_), .Y(new_n12346_));
  OAI21X1  g09910(.A0(new_n12332_), .A1(new_n5050_), .B0(new_n12346_), .Y(new_n12347_));
  NAND2X1  g09911(.A(new_n12347_), .B(new_n2953_), .Y(new_n12348_));
  OAI22X1  g09912(.A0(new_n12348_), .A1(new_n12345_), .B0(new_n12338_), .B1(new_n2953_), .Y(new_n12349_));
  OAI21X1  g09913(.A0(new_n12349_), .A1(new_n7398_), .B0(pi0761), .Y(new_n12350_));
  AOI21X1  g09914(.A0(new_n12289_), .A1(new_n7398_), .B0(new_n12350_), .Y(new_n12351_));
  NOR2X1   g09915(.A(new_n12116_), .B(new_n5027_), .Y(new_n12352_));
  AOI21X1  g09916(.A0(new_n12299_), .A1(new_n12298_), .B0(new_n12352_), .Y(new_n12353_));
  AOI21X1  g09917(.A0(new_n12294_), .A1(new_n12171_), .B0(new_n12107_), .Y(new_n12354_));
  AOI21X1  g09918(.A0(new_n12354_), .A1(new_n12127_), .B0(new_n12235_), .Y(new_n12355_));
  OAI21X1  g09919(.A0(new_n12353_), .A1(new_n12127_), .B0(new_n12355_), .Y(new_n12356_));
  NAND3X1  g09920(.A(new_n12293_), .B(new_n12028_), .C(new_n5030_), .Y(new_n12357_));
  NAND3X1  g09921(.A(new_n12357_), .B(new_n12235_), .C(new_n12175_), .Y(new_n12358_));
  NAND3X1  g09922(.A(new_n12358_), .B(new_n12356_), .C(new_n5051_), .Y(new_n12359_));
  NOR2X1   g09923(.A(new_n12263_), .B(new_n12219_), .Y(new_n12360_));
  NOR3X1   g09924(.A(new_n12360_), .B(new_n11952_), .C(new_n2740_), .Y(new_n12361_));
  AOI21X1  g09925(.A0(new_n12361_), .A1(new_n12127_), .B0(new_n12235_), .Y(new_n12362_));
  INVX1    g09926(.A(new_n12362_), .Y(new_n12363_));
  NAND2X1  g09927(.A(new_n12120_), .B(new_n12029_), .Y(new_n12364_));
  AOI21X1  g09928(.A0(new_n12314_), .A1(new_n12364_), .B0(new_n12127_), .Y(new_n12365_));
  OR2X1    g09929(.A(new_n12365_), .B(new_n12363_), .Y(new_n12366_));
  MX2X1    g09930(.A(new_n12181_), .B(new_n12364_), .S0(new_n12125_), .Y(new_n12367_));
  NOR2X1   g09931(.A(new_n12294_), .B(new_n12047_), .Y(new_n12368_));
  NOR3X1   g09932(.A(new_n12368_), .B(new_n12170_), .C(new_n5282_), .Y(new_n12369_));
  AOI21X1  g09933(.A0(new_n12367_), .A1(new_n5029_), .B0(new_n12369_), .Y(new_n12370_));
  NAND3X1  g09934(.A(new_n12370_), .B(new_n12366_), .C(new_n5050_), .Y(new_n12371_));
  AND2X1   g09935(.A(new_n12371_), .B(new_n2971_), .Y(new_n12372_));
  NAND2X1  g09936(.A(new_n12372_), .B(new_n12359_), .Y(new_n12373_));
  NOR2X1   g09937(.A(new_n12344_), .B(pi0223), .Y(new_n12374_));
  NAND2X1  g09938(.A(new_n12185_), .B(new_n12183_), .Y(new_n12375_));
  INVX1    g09939(.A(new_n12292_), .Y(new_n12376_));
  AOI21X1  g09940(.A0(new_n11970_), .A1(new_n5028_), .B0(new_n12376_), .Y(new_n12377_));
  INVX1    g09941(.A(new_n12377_), .Y(new_n12378_));
  AOI21X1  g09942(.A0(new_n12378_), .A1(new_n12183_), .B0(new_n12127_), .Y(new_n12379_));
  OAI21X1  g09943(.A0(new_n12376_), .A1(new_n11970_), .B0(new_n11993_), .Y(new_n12380_));
  AND2X1   g09944(.A(new_n12380_), .B(pi0680), .Y(new_n12381_));
  OAI22X1  g09945(.A0(new_n12381_), .A1(new_n12375_), .B0(new_n12379_), .B1(new_n12363_), .Y(new_n12382_));
  NAND2X1  g09946(.A(new_n12382_), .B(new_n5050_), .Y(new_n12383_));
  OAI21X1  g09947(.A0(new_n12181_), .A1(new_n11965_), .B0(new_n12185_), .Y(new_n12384_));
  OR2X1    g09948(.A(new_n12376_), .B(new_n11966_), .Y(new_n12385_));
  NAND3X1  g09949(.A(new_n12380_), .B(new_n12377_), .C(pi0680), .Y(new_n12386_));
  NOR2X1   g09950(.A(new_n12386_), .B(new_n12385_), .Y(new_n12387_));
  NOR2X1   g09951(.A(new_n12387_), .B(new_n12384_), .Y(new_n12388_));
  AOI21X1  g09952(.A0(new_n12388_), .A1(new_n5051_), .B0(new_n2964_), .Y(new_n12389_));
  AOI21X1  g09953(.A0(new_n12389_), .A1(new_n12383_), .B0(pi0299), .Y(new_n12390_));
  INVX1    g09954(.A(new_n12390_), .Y(new_n12391_));
  AOI21X1  g09955(.A0(new_n12374_), .A1(new_n12373_), .B0(new_n12391_), .Y(new_n12392_));
  NAND3X1  g09956(.A(new_n12358_), .B(new_n12356_), .C(new_n5071_), .Y(new_n12393_));
  NAND3X1  g09957(.A(new_n12370_), .B(new_n12366_), .C(new_n5070_), .Y(new_n12394_));
  AOI21X1  g09958(.A0(new_n12394_), .A1(new_n12393_), .B0(new_n10136_), .Y(new_n12395_));
  AOI21X1  g09959(.A0(new_n12343_), .A1(new_n10136_), .B0(pi0215), .Y(new_n12396_));
  INVX1    g09960(.A(new_n12396_), .Y(new_n12397_));
  NOR2X1   g09961(.A(new_n12382_), .B(new_n5071_), .Y(new_n12398_));
  OAI21X1  g09962(.A0(new_n12388_), .A1(new_n5070_), .B0(pi0215), .Y(new_n12399_));
  OAI22X1  g09963(.A0(new_n12399_), .A1(new_n12398_), .B0(new_n12397_), .B1(new_n12395_), .Y(new_n12400_));
  AOI21X1  g09964(.A0(new_n12400_), .A1(pi0299), .B0(new_n12392_), .Y(new_n12401_));
  AOI21X1  g09965(.A0(new_n12171_), .A1(new_n12057_), .B0(pi0680), .Y(new_n12402_));
  NAND3X1  g09966(.A(new_n12210_), .B(new_n12045_), .C(new_n12037_), .Y(new_n12403_));
  OAI22X1  g09967(.A0(new_n12403_), .A1(new_n5371_), .B0(new_n12221_), .B1(new_n5028_), .Y(new_n12404_));
  AOI21X1  g09968(.A0(new_n12404_), .A1(new_n12360_), .B0(new_n12235_), .Y(new_n12405_));
  OR4X1    g09969(.A(new_n12405_), .B(new_n12402_), .C(new_n12265_), .D(new_n5050_), .Y(new_n12406_));
  NOR3X1   g09970(.A(new_n12130_), .B(new_n12126_), .C(pi0680), .Y(new_n12407_));
  NOR4X1   g09971(.A(new_n12263_), .B(new_n12219_), .C(new_n11952_), .D(new_n2740_), .Y(new_n12408_));
  INVX1    g09972(.A(new_n12408_), .Y(new_n12409_));
  OAI21X1  g09973(.A0(new_n12409_), .A1(new_n12125_), .B0(new_n12209_), .Y(new_n12410_));
  AOI21X1  g09974(.A0(new_n12210_), .A1(new_n12130_), .B0(new_n12410_), .Y(new_n12411_));
  AOI21X1  g09975(.A0(new_n12360_), .A1(new_n12253_), .B0(new_n5282_), .Y(new_n12412_));
  OR4X1    g09976(.A(new_n12412_), .B(new_n12411_), .C(new_n12407_), .D(new_n5051_), .Y(new_n12413_));
  AOI21X1  g09977(.A0(new_n12413_), .A1(new_n12406_), .B0(new_n2970_), .Y(new_n12414_));
  AND2X1   g09978(.A(new_n11951_), .B(new_n10174_), .Y(new_n12415_));
  INVX1    g09979(.A(new_n11961_), .Y(new_n12416_));
  NOR4X1   g09980(.A(new_n12341_), .B(new_n12120_), .C(new_n12416_), .D(new_n12415_), .Y(new_n12417_));
  AOI21X1  g09981(.A0(new_n12417_), .A1(new_n2970_), .B0(pi0223), .Y(new_n12418_));
  INVX1    g09982(.A(new_n12418_), .Y(new_n12419_));
  NOR3X1   g09983(.A(new_n12341_), .B(new_n12141_), .C(new_n5030_), .Y(new_n12420_));
  NOR2X1   g09984(.A(new_n12263_), .B(new_n5282_), .Y(new_n12421_));
  AOI21X1  g09985(.A0(new_n12421_), .A1(new_n12224_), .B0(new_n12420_), .Y(new_n12422_));
  NOR2X1   g09986(.A(new_n12422_), .B(new_n5051_), .Y(new_n12423_));
  OAI21X1  g09987(.A0(new_n12237_), .A1(new_n12141_), .B0(new_n12209_), .Y(new_n12424_));
  AOI21X1  g09988(.A0(new_n11958_), .A1(pi0665), .B0(new_n5029_), .Y(new_n12425_));
  OR2X1    g09989(.A(new_n12425_), .B(new_n12263_), .Y(new_n12426_));
  AOI22X1  g09990(.A0(new_n12426_), .A1(new_n5030_), .B0(new_n12148_), .B1(new_n5029_), .Y(new_n12427_));
  NAND2X1  g09991(.A(new_n12427_), .B(new_n12424_), .Y(new_n12428_));
  OAI21X1  g09992(.A0(new_n12428_), .A1(new_n5050_), .B0(pi0223), .Y(new_n12429_));
  OAI22X1  g09993(.A0(new_n12429_), .A1(new_n12423_), .B0(new_n12419_), .B1(new_n12414_), .Y(new_n12430_));
  AND2X1   g09994(.A(new_n12430_), .B(new_n2953_), .Y(new_n12431_));
  OR4X1    g09995(.A(new_n12405_), .B(new_n12402_), .C(new_n12265_), .D(new_n5070_), .Y(new_n12432_));
  OR4X1    g09996(.A(new_n12412_), .B(new_n12411_), .C(new_n12407_), .D(new_n5071_), .Y(new_n12433_));
  AOI21X1  g09997(.A0(new_n12433_), .A1(new_n12432_), .B0(new_n10136_), .Y(new_n12434_));
  AOI21X1  g09998(.A0(new_n12417_), .A1(new_n10136_), .B0(pi0215), .Y(new_n12435_));
  INVX1    g09999(.A(new_n12435_), .Y(new_n12436_));
  NOR2X1   g10000(.A(new_n12422_), .B(new_n5071_), .Y(new_n12437_));
  OAI21X1  g10001(.A0(new_n12428_), .A1(new_n5070_), .B0(pi0215), .Y(new_n12438_));
  OAI22X1  g10002(.A0(new_n12438_), .A1(new_n12437_), .B0(new_n12436_), .B1(new_n12434_), .Y(new_n12439_));
  AOI21X1  g10003(.A0(new_n12439_), .A1(pi0299), .B0(new_n12431_), .Y(new_n12440_));
  OAI21X1  g10004(.A0(new_n12440_), .A1(pi0140), .B0(new_n11890_), .Y(new_n12441_));
  AOI21X1  g10005(.A0(new_n12401_), .A1(pi0140), .B0(new_n12441_), .Y(new_n12442_));
  OAI21X1  g10006(.A0(new_n12442_), .A1(new_n12351_), .B0(pi0039), .Y(new_n12443_));
  NAND2X1  g10007(.A(new_n11928_), .B(new_n11927_), .Y(new_n12444_));
  OAI21X1  g10008(.A0(new_n12444_), .A1(pi0198), .B0(new_n11945_), .Y(new_n12445_));
  OR2X1    g10009(.A(new_n11941_), .B(new_n12255_), .Y(new_n12446_));
  NOR2X1   g10010(.A(new_n11927_), .B(new_n12255_), .Y(new_n12447_));
  INVX1    g10011(.A(new_n12447_), .Y(new_n12448_));
  MX2X1    g10012(.A(new_n12448_), .B(new_n12446_), .S0(pi0198), .Y(new_n12449_));
  AOI21X1  g10013(.A0(new_n12449_), .A1(pi0680), .B0(new_n12445_), .Y(new_n12450_));
  MX2X1    g10014(.A(new_n12448_), .B(new_n12446_), .S0(pi0210), .Y(new_n12451_));
  AOI21X1  g10015(.A0(new_n12451_), .A1(pi0680), .B0(new_n12091_), .Y(new_n12452_));
  MX2X1    g10016(.A(new_n12452_), .B(new_n12450_), .S0(new_n2953_), .Y(new_n12453_));
  AOI21X1  g10017(.A0(new_n12168_), .A1(pi0680), .B0(new_n12453_), .Y(new_n12454_));
  OAI21X1  g10018(.A0(new_n11927_), .A1(pi0665), .B0(new_n11928_), .Y(new_n12455_));
  OR2X1    g10019(.A(new_n12455_), .B(pi0198), .Y(new_n12456_));
  OAI21X1  g10020(.A0(new_n11941_), .A1(pi0665), .B0(new_n11937_), .Y(new_n12457_));
  OAI21X1  g10021(.A0(new_n12457_), .A1(new_n2973_), .B0(new_n12456_), .Y(new_n12458_));
  NAND2X1  g10022(.A(new_n12458_), .B(new_n5027_), .Y(new_n12459_));
  AND2X1   g10023(.A(pi0665), .B(pi0603), .Y(new_n12460_));
  AOI21X1  g10024(.A0(new_n12098_), .A1(pi0603), .B0(new_n12460_), .Y(new_n12461_));
  NAND3X1  g10025(.A(new_n12461_), .B(new_n12459_), .C(pi0680), .Y(new_n12462_));
  MX2X1    g10026(.A(new_n12457_), .B(new_n12455_), .S0(new_n2766_), .Y(new_n12463_));
  OR2X1    g10027(.A(new_n12463_), .B(pi0603), .Y(new_n12464_));
  AOI21X1  g10028(.A0(new_n12096_), .A1(pi0603), .B0(new_n12460_), .Y(new_n12465_));
  NAND3X1  g10029(.A(new_n12465_), .B(new_n12464_), .C(pi0680), .Y(new_n12466_));
  MX2X1    g10030(.A(new_n12466_), .B(new_n12462_), .S0(new_n2953_), .Y(new_n12467_));
  AOI21X1  g10031(.A0(new_n12467_), .A1(pi0140), .B0(new_n11890_), .Y(new_n12468_));
  OAI21X1  g10032(.A0(new_n12454_), .A1(pi0140), .B0(new_n12468_), .Y(new_n12469_));
  NAND3X1  g10033(.A(new_n12453_), .B(new_n12104_), .C(new_n7398_), .Y(new_n12470_));
  NOR2X1   g10034(.A(new_n12458_), .B(new_n5029_), .Y(new_n12471_));
  AND2X1   g10035(.A(new_n12463_), .B(pi0680), .Y(new_n12472_));
  MX2X1    g10036(.A(new_n12472_), .B(new_n12471_), .S0(new_n2953_), .Y(new_n12473_));
  NOR2X1   g10037(.A(new_n12473_), .B(new_n12168_), .Y(new_n12474_));
  AOI21X1  g10038(.A0(new_n12474_), .A1(pi0140), .B0(pi0761), .Y(new_n12475_));
  AOI21X1  g10039(.A0(new_n12475_), .A1(new_n12470_), .B0(pi0039), .Y(new_n12476_));
  AOI21X1  g10040(.A0(new_n12476_), .A1(new_n12469_), .B0(pi0038), .Y(new_n12477_));
  NOR4X1   g10041(.A(new_n12341_), .B(new_n12120_), .C(new_n3074_), .D(new_n2740_), .Y(new_n12478_));
  OR4X1    g10042(.A(new_n12342_), .B(new_n3003_), .C(new_n2555_), .D(new_n7398_), .Y(new_n12479_));
  AND2X1   g10043(.A(new_n12479_), .B(new_n11890_), .Y(new_n12480_));
  OAI21X1  g10044(.A0(new_n12478_), .A1(pi0140), .B0(new_n12480_), .Y(new_n12481_));
  INVX1    g10045(.A(new_n12269_), .Y(new_n12482_));
  NOR4X1   g10046(.A(new_n12482_), .B(new_n3003_), .C(new_n2740_), .D(new_n2555_), .Y(new_n12483_));
  NOR2X1   g10047(.A(new_n12483_), .B(new_n11890_), .Y(new_n12484_));
  OAI21X1  g10048(.A0(new_n11961_), .A1(pi0140), .B0(new_n12484_), .Y(new_n12485_));
  AOI21X1  g10049(.A0(new_n12485_), .A1(new_n12481_), .B0(pi0039), .Y(new_n12486_));
  AND2X1   g10050(.A(pi0140), .B(pi0039), .Y(new_n12487_));
  NOR3X1   g10051(.A(new_n12487_), .B(new_n12486_), .C(new_n2996_), .Y(new_n12488_));
  AOI21X1  g10052(.A0(new_n12477_), .A1(new_n12443_), .B0(new_n12488_), .Y(new_n12489_));
  OAI21X1  g10053(.A0(new_n12489_), .A1(pi0738), .B0(new_n3129_), .Y(new_n12490_));
  AOI21X1  g10054(.A0(new_n12208_), .A1(pi0738), .B0(new_n12490_), .Y(new_n12491_));
  AOI21X1  g10055(.A0(new_n3810_), .A1(pi0140), .B0(new_n12491_), .Y(new_n12492_));
  INVX1    g10056(.A(pi0625), .Y(new_n12493_));
  INVX1    g10057(.A(pi1153), .Y(new_n12494_));
  MX2X1    g10058(.A(new_n12206_), .B(new_n12201_), .S0(new_n2996_), .Y(new_n12495_));
  MX2X1    g10059(.A(new_n12495_), .B(pi0140), .S0(new_n3810_), .Y(new_n12496_));
  OAI21X1  g10060(.A0(new_n12496_), .A1(new_n12493_), .B0(new_n12494_), .Y(new_n12497_));
  AOI21X1  g10061(.A0(new_n12492_), .A1(new_n12493_), .B0(new_n12497_), .Y(new_n12498_));
  INVX1    g10062(.A(new_n12341_), .Y(new_n12499_));
  OR4X1    g10063(.A(new_n12499_), .B(new_n11952_), .C(new_n2971_), .D(new_n2740_), .Y(new_n12500_));
  OR2X1    g10064(.A(new_n12294_), .B(new_n12047_), .Y(new_n12501_));
  MX2X1    g10065(.A(new_n12501_), .B(new_n12376_), .S0(new_n5367_), .Y(new_n12502_));
  OAI21X1  g10066(.A0(new_n12368_), .A1(new_n12290_), .B0(pi0680), .Y(new_n12503_));
  AOI21X1  g10067(.A0(new_n12502_), .A1(new_n12290_), .B0(new_n12503_), .Y(new_n12504_));
  NOR2X1   g10068(.A(new_n12504_), .B(new_n5051_), .Y(new_n12505_));
  OR2X1    g10069(.A(new_n12499_), .B(new_n12260_), .Y(new_n12506_));
  OAI21X1  g10070(.A0(new_n12506_), .A1(new_n11993_), .B0(new_n12357_), .Y(new_n12507_));
  OAI21X1  g10071(.A0(new_n12507_), .A1(new_n5050_), .B0(new_n2971_), .Y(new_n12508_));
  OAI21X1  g10072(.A0(new_n12508_), .A1(new_n12505_), .B0(new_n12500_), .Y(new_n12509_));
  NOR3X1   g10073(.A(new_n12378_), .B(new_n12194_), .C(new_n5029_), .Y(new_n12510_));
  AND2X1   g10074(.A(new_n12380_), .B(pi0223), .Y(new_n12511_));
  AND2X1   g10075(.A(new_n12511_), .B(new_n12510_), .Y(new_n12512_));
  AOI21X1  g10076(.A0(new_n12509_), .A1(new_n2964_), .B0(new_n12512_), .Y(new_n12513_));
  NOR2X1   g10077(.A(new_n12507_), .B(new_n5070_), .Y(new_n12514_));
  OAI21X1  g10078(.A0(new_n12504_), .A1(new_n5071_), .B0(new_n10137_), .Y(new_n12515_));
  OR4X1    g10079(.A(new_n12499_), .B(new_n11952_), .C(new_n10137_), .D(new_n2740_), .Y(new_n12516_));
  OAI21X1  g10080(.A0(new_n12515_), .A1(new_n12514_), .B0(new_n12516_), .Y(new_n12517_));
  NOR3X1   g10081(.A(new_n12378_), .B(new_n12186_), .C(new_n5029_), .Y(new_n12518_));
  AND2X1   g10082(.A(new_n12380_), .B(pi0215), .Y(new_n12519_));
  AND2X1   g10083(.A(new_n12519_), .B(new_n12518_), .Y(new_n12520_));
  AOI21X1  g10084(.A0(new_n12517_), .A1(new_n2954_), .B0(new_n12520_), .Y(new_n12521_));
  MX2X1    g10085(.A(new_n12521_), .B(new_n12513_), .S0(new_n2953_), .Y(new_n12522_));
  OR2X1    g10086(.A(new_n12522_), .B(new_n7398_), .Y(new_n12523_));
  NAND2X1  g10087(.A(new_n12033_), .B(new_n5029_), .Y(new_n12524_));
  AOI21X1  g10088(.A0(new_n12223_), .A1(new_n5367_), .B0(new_n5029_), .Y(new_n12525_));
  INVX1    g10089(.A(new_n12525_), .Y(new_n12526_));
  AOI21X1  g10090(.A0(new_n12253_), .A1(new_n5028_), .B0(new_n12526_), .Y(new_n12527_));
  AOI21X1  g10091(.A0(new_n12033_), .A1(new_n5029_), .B0(new_n12527_), .Y(new_n12528_));
  OR2X1    g10092(.A(new_n12253_), .B(new_n5029_), .Y(new_n12529_));
  AND2X1   g10093(.A(new_n12529_), .B(new_n11993_), .Y(new_n12530_));
  AOI22X1  g10094(.A0(new_n12530_), .A1(new_n12524_), .B0(new_n12528_), .B1(new_n12290_), .Y(new_n12531_));
  OAI21X1  g10095(.A0(new_n12403_), .A1(new_n12290_), .B0(pi0680), .Y(new_n12532_));
  AOI21X1  g10096(.A0(new_n12404_), .A1(new_n12290_), .B0(new_n12532_), .Y(new_n12533_));
  AOI21X1  g10097(.A0(new_n12260_), .A1(new_n5029_), .B0(new_n12533_), .Y(new_n12534_));
  INVX1    g10098(.A(new_n12534_), .Y(new_n12535_));
  AOI21X1  g10099(.A0(new_n12535_), .A1(new_n5051_), .B0(new_n2970_), .Y(new_n12536_));
  INVX1    g10100(.A(new_n12536_), .Y(new_n12537_));
  AOI21X1  g10101(.A0(new_n12531_), .A1(new_n5050_), .B0(new_n12537_), .Y(new_n12538_));
  AOI21X1  g10102(.A0(new_n12499_), .A1(new_n12065_), .B0(pi0223), .Y(new_n12539_));
  INVX1    g10103(.A(new_n12539_), .Y(new_n12540_));
  AOI21X1  g10104(.A0(new_n12526_), .A1(new_n5282_), .B0(new_n12224_), .Y(new_n12541_));
  AOI21X1  g10105(.A0(new_n12230_), .A1(new_n5029_), .B0(new_n12541_), .Y(new_n12542_));
  AND2X1   g10106(.A(new_n12542_), .B(new_n5050_), .Y(new_n12543_));
  OAI21X1  g10107(.A0(new_n12221_), .A1(new_n5028_), .B0(new_n12425_), .Y(new_n12544_));
  OAI21X1  g10108(.A0(new_n11974_), .A1(pi0680), .B0(new_n12544_), .Y(new_n12545_));
  NOR2X1   g10109(.A(new_n12545_), .B(new_n12541_), .Y(new_n12546_));
  AOI21X1  g10110(.A0(new_n12546_), .A1(new_n5051_), .B0(new_n2964_), .Y(new_n12547_));
  INVX1    g10111(.A(new_n12547_), .Y(new_n12548_));
  OAI22X1  g10112(.A0(new_n12548_), .A1(new_n12543_), .B0(new_n12540_), .B1(new_n12538_), .Y(new_n12549_));
  AOI21X1  g10113(.A0(new_n12535_), .A1(new_n5071_), .B0(new_n10136_), .Y(new_n12550_));
  INVX1    g10114(.A(new_n12550_), .Y(new_n12551_));
  AOI21X1  g10115(.A0(new_n12531_), .A1(new_n5070_), .B0(new_n12551_), .Y(new_n12552_));
  OR4X1    g10116(.A(new_n12341_), .B(new_n11952_), .C(new_n10137_), .D(new_n2740_), .Y(new_n12553_));
  AND2X1   g10117(.A(new_n12553_), .B(new_n2954_), .Y(new_n12554_));
  INVX1    g10118(.A(new_n12554_), .Y(new_n12555_));
  AND2X1   g10119(.A(new_n12542_), .B(new_n5070_), .Y(new_n12556_));
  AOI21X1  g10120(.A0(new_n12546_), .A1(new_n5071_), .B0(new_n2954_), .Y(new_n12557_));
  INVX1    g10121(.A(new_n12557_), .Y(new_n12558_));
  OAI22X1  g10122(.A0(new_n12558_), .A1(new_n12556_), .B0(new_n12555_), .B1(new_n12552_), .Y(new_n12559_));
  MX2X1    g10123(.A(new_n12559_), .B(new_n12549_), .S0(new_n2953_), .Y(new_n12560_));
  AOI21X1  g10124(.A0(new_n12560_), .A1(new_n7398_), .B0(new_n2959_), .Y(new_n12561_));
  OAI21X1  g10125(.A0(new_n12453_), .A1(pi0140), .B0(new_n2959_), .Y(new_n12562_));
  AOI21X1  g10126(.A0(new_n12473_), .A1(pi0140), .B0(new_n12562_), .Y(new_n12563_));
  AOI21X1  g10127(.A0(new_n12561_), .A1(new_n12523_), .B0(new_n12563_), .Y(new_n12564_));
  INVX1    g10128(.A(pi0738), .Y(new_n12565_));
  NOR4X1   g10129(.A(new_n12210_), .B(new_n2756_), .C(new_n2755_), .D(new_n5029_), .Y(new_n12566_));
  AOI21X1  g10130(.A0(new_n12566_), .A1(new_n6857_), .B0(new_n2996_), .Y(new_n12567_));
  INVX1    g10131(.A(new_n12567_), .Y(new_n12568_));
  OAI21X1  g10132(.A0(new_n12568_), .A1(new_n12203_), .B0(new_n12565_), .Y(new_n12569_));
  INVX1    g10133(.A(new_n12569_), .Y(new_n12570_));
  OAI21X1  g10134(.A0(new_n12564_), .A1(pi0038), .B0(new_n12570_), .Y(new_n12571_));
  AND2X1   g10135(.A(new_n4995_), .B(new_n2739_), .Y(new_n12572_));
  INVX1    g10136(.A(new_n12572_), .Y(new_n12573_));
  MX2X1    g10137(.A(new_n12573_), .B(new_n12090_), .S0(new_n2996_), .Y(new_n12574_));
  AND2X1   g10138(.A(pi0738), .B(new_n7398_), .Y(new_n12575_));
  AOI21X1  g10139(.A0(new_n12575_), .A1(new_n12574_), .B0(new_n3810_), .Y(new_n12576_));
  AOI22X1  g10140(.A0(new_n12576_), .A1(new_n12571_), .B0(new_n3810_), .B1(pi0140), .Y(new_n12577_));
  OAI21X1  g10141(.A0(new_n12574_), .A1(new_n3810_), .B0(new_n7398_), .Y(new_n12578_));
  OAI21X1  g10142(.A0(new_n12578_), .A1(pi0625), .B0(pi1153), .Y(new_n12579_));
  AOI21X1  g10143(.A0(new_n12577_), .A1(pi0625), .B0(new_n12579_), .Y(new_n12580_));
  OR2X1    g10144(.A(new_n12580_), .B(pi0608), .Y(new_n12581_));
  OAI21X1  g10145(.A0(new_n12496_), .A1(pi0625), .B0(pi1153), .Y(new_n12582_));
  AOI21X1  g10146(.A0(new_n12492_), .A1(pi0625), .B0(new_n12582_), .Y(new_n12583_));
  INVX1    g10147(.A(pi0608), .Y(new_n12584_));
  OAI21X1  g10148(.A0(new_n12578_), .A1(new_n12493_), .B0(new_n12494_), .Y(new_n12585_));
  AOI21X1  g10149(.A0(new_n12577_), .A1(new_n12493_), .B0(new_n12585_), .Y(new_n12586_));
  OR2X1    g10150(.A(new_n12586_), .B(new_n12584_), .Y(new_n12587_));
  OAI22X1  g10151(.A0(new_n12587_), .A1(new_n12583_), .B0(new_n12581_), .B1(new_n12498_), .Y(new_n12588_));
  MX2X1    g10152(.A(new_n12588_), .B(new_n12492_), .S0(new_n11889_), .Y(new_n12589_));
  INVX1    g10153(.A(pi0609), .Y(new_n12590_));
  INVX1    g10154(.A(pi1155), .Y(new_n12591_));
  OAI21X1  g10155(.A0(new_n12586_), .A1(new_n12580_), .B0(pi0778), .Y(new_n12592_));
  OAI21X1  g10156(.A0(new_n12577_), .A1(pi0778), .B0(new_n12592_), .Y(new_n12593_));
  OAI21X1  g10157(.A0(new_n12593_), .A1(new_n12590_), .B0(new_n12591_), .Y(new_n12594_));
  AOI21X1  g10158(.A0(new_n12589_), .A1(new_n12590_), .B0(new_n12594_), .Y(new_n12595_));
  INVX1    g10159(.A(pi0660), .Y(new_n12596_));
  INVX1    g10160(.A(new_n12578_), .Y(new_n12597_));
  XOR2X1   g10161(.A(pi1153), .B(pi0608), .Y(new_n12598_));
  AOI21X1  g10162(.A0(new_n12598_), .A1(pi0778), .B0(new_n12590_), .Y(new_n12599_));
  MX2X1    g10163(.A(new_n12208_), .B(new_n7398_), .S0(new_n3810_), .Y(new_n12600_));
  AND2X1   g10164(.A(new_n12598_), .B(pi0778), .Y(new_n12601_));
  OR2X1    g10165(.A(new_n12601_), .B(new_n12600_), .Y(new_n12602_));
  OAI22X1  g10166(.A0(new_n12602_), .A1(new_n12590_), .B0(new_n12599_), .B1(new_n12597_), .Y(new_n12603_));
  NAND2X1  g10167(.A(new_n12603_), .B(pi1155), .Y(new_n12604_));
  NAND2X1  g10168(.A(new_n12604_), .B(new_n12596_), .Y(new_n12605_));
  OAI21X1  g10169(.A0(new_n12593_), .A1(pi0609), .B0(pi1155), .Y(new_n12606_));
  AOI21X1  g10170(.A0(new_n12589_), .A1(pi0609), .B0(new_n12606_), .Y(new_n12607_));
  AOI21X1  g10171(.A0(new_n12598_), .A1(pi0778), .B0(pi0609), .Y(new_n12608_));
  OAI22X1  g10172(.A0(new_n12608_), .A1(new_n12597_), .B0(new_n12602_), .B1(pi0609), .Y(new_n12609_));
  NAND2X1  g10173(.A(new_n12609_), .B(new_n12591_), .Y(new_n12610_));
  NAND2X1  g10174(.A(new_n12610_), .B(pi0660), .Y(new_n12611_));
  OAI22X1  g10175(.A0(new_n12611_), .A1(new_n12607_), .B0(new_n12605_), .B1(new_n12595_), .Y(new_n12612_));
  MX2X1    g10176(.A(new_n12612_), .B(new_n12589_), .S0(new_n11888_), .Y(new_n12613_));
  INVX1    g10177(.A(pi0618), .Y(new_n12614_));
  INVX1    g10178(.A(pi1154), .Y(new_n12615_));
  AND2X1   g10179(.A(pi1155), .B(pi0660), .Y(new_n12616_));
  NOR2X1   g10180(.A(pi1155), .B(pi0660), .Y(new_n12617_));
  NOR3X1   g10181(.A(new_n12617_), .B(new_n12616_), .C(new_n11888_), .Y(new_n12618_));
  MX2X1    g10182(.A(new_n12593_), .B(new_n12578_), .S0(new_n12618_), .Y(new_n12619_));
  OAI21X1  g10183(.A0(new_n12619_), .A1(new_n12614_), .B0(new_n12615_), .Y(new_n12620_));
  AOI21X1  g10184(.A0(new_n12613_), .A1(new_n12614_), .B0(new_n12620_), .Y(new_n12621_));
  INVX1    g10185(.A(pi0627), .Y(new_n12622_));
  INVX1    g10186(.A(new_n12601_), .Y(new_n12623_));
  MX2X1    g10187(.A(new_n12578_), .B(new_n12496_), .S0(new_n12623_), .Y(new_n12624_));
  MX2X1    g10188(.A(new_n12609_), .B(new_n12603_), .S0(pi1155), .Y(new_n12625_));
  MX2X1    g10189(.A(new_n12625_), .B(new_n12624_), .S0(new_n11888_), .Y(new_n12626_));
  AOI21X1  g10190(.A0(new_n12597_), .A1(new_n12614_), .B0(new_n12615_), .Y(new_n12627_));
  OAI21X1  g10191(.A0(new_n12626_), .A1(new_n12614_), .B0(new_n12627_), .Y(new_n12628_));
  NAND2X1  g10192(.A(new_n12628_), .B(new_n12622_), .Y(new_n12629_));
  OAI21X1  g10193(.A0(new_n12619_), .A1(pi0618), .B0(pi1154), .Y(new_n12630_));
  AOI21X1  g10194(.A0(new_n12613_), .A1(pi0618), .B0(new_n12630_), .Y(new_n12631_));
  AOI21X1  g10195(.A0(new_n12597_), .A1(pi0618), .B0(pi1154), .Y(new_n12632_));
  OAI21X1  g10196(.A0(new_n12626_), .A1(pi0618), .B0(new_n12632_), .Y(new_n12633_));
  NAND2X1  g10197(.A(new_n12633_), .B(pi0627), .Y(new_n12634_));
  OAI22X1  g10198(.A0(new_n12634_), .A1(new_n12631_), .B0(new_n12629_), .B1(new_n12621_), .Y(new_n12635_));
  MX2X1    g10199(.A(new_n12635_), .B(new_n12613_), .S0(new_n11887_), .Y(new_n12636_));
  INVX1    g10200(.A(pi0619), .Y(new_n12637_));
  INVX1    g10201(.A(pi1159), .Y(new_n12638_));
  AND2X1   g10202(.A(pi1154), .B(pi0627), .Y(new_n12639_));
  OAI21X1  g10203(.A0(pi1154), .A1(pi0627), .B0(pi0781), .Y(new_n12640_));
  NOR2X1   g10204(.A(new_n12640_), .B(new_n12639_), .Y(new_n12641_));
  MX2X1    g10205(.A(new_n12619_), .B(new_n12578_), .S0(new_n12641_), .Y(new_n12642_));
  OAI21X1  g10206(.A0(new_n12642_), .A1(new_n12637_), .B0(new_n12638_), .Y(new_n12643_));
  AOI21X1  g10207(.A0(new_n12636_), .A1(new_n12637_), .B0(new_n12643_), .Y(new_n12644_));
  INVX1    g10208(.A(pi0648), .Y(new_n12645_));
  NAND2X1  g10209(.A(new_n12633_), .B(new_n12628_), .Y(new_n12646_));
  MX2X1    g10210(.A(new_n12646_), .B(new_n12626_), .S0(new_n11887_), .Y(new_n12647_));
  AOI21X1  g10211(.A0(new_n12597_), .A1(new_n12637_), .B0(new_n12638_), .Y(new_n12648_));
  OAI21X1  g10212(.A0(new_n12647_), .A1(new_n12637_), .B0(new_n12648_), .Y(new_n12649_));
  NAND2X1  g10213(.A(new_n12649_), .B(new_n12645_), .Y(new_n12650_));
  OAI21X1  g10214(.A0(new_n12642_), .A1(pi0619), .B0(pi1159), .Y(new_n12651_));
  AOI21X1  g10215(.A0(new_n12636_), .A1(pi0619), .B0(new_n12651_), .Y(new_n12652_));
  AOI21X1  g10216(.A0(new_n12597_), .A1(pi0619), .B0(pi1159), .Y(new_n12653_));
  OAI21X1  g10217(.A0(new_n12647_), .A1(pi0619), .B0(new_n12653_), .Y(new_n12654_));
  NAND2X1  g10218(.A(new_n12654_), .B(pi0648), .Y(new_n12655_));
  OAI22X1  g10219(.A0(new_n12655_), .A1(new_n12652_), .B0(new_n12650_), .B1(new_n12644_), .Y(new_n12656_));
  MX2X1    g10220(.A(new_n12656_), .B(new_n12636_), .S0(new_n11886_), .Y(new_n12657_));
  XOR2X1   g10221(.A(pi1159), .B(new_n12645_), .Y(new_n12658_));
  NOR2X1   g10222(.A(new_n12658_), .B(new_n11886_), .Y(new_n12659_));
  MX2X1    g10223(.A(new_n12642_), .B(new_n12578_), .S0(new_n12659_), .Y(new_n12660_));
  AOI21X1  g10224(.A0(new_n12660_), .A1(pi0626), .B0(pi0641), .Y(new_n12661_));
  OAI21X1  g10225(.A0(new_n12657_), .A1(pi0626), .B0(new_n12661_), .Y(new_n12662_));
  NOR2X1   g10226(.A(pi1158), .B(pi0641), .Y(new_n12663_));
  INVX1    g10227(.A(pi0626), .Y(new_n12664_));
  AND2X1   g10228(.A(new_n12647_), .B(new_n11886_), .Y(new_n12665_));
  AOI21X1  g10229(.A0(new_n12654_), .A1(new_n12649_), .B0(new_n11886_), .Y(new_n12666_));
  NOR2X1   g10230(.A(new_n12666_), .B(new_n12665_), .Y(new_n12667_));
  AOI21X1  g10231(.A0(new_n12597_), .A1(pi0626), .B0(pi1158), .Y(new_n12668_));
  INVX1    g10232(.A(new_n12668_), .Y(new_n12669_));
  AOI21X1  g10233(.A0(new_n12667_), .A1(new_n12664_), .B0(new_n12669_), .Y(new_n12670_));
  OR2X1    g10234(.A(new_n12670_), .B(new_n12663_), .Y(new_n12671_));
  INVX1    g10235(.A(pi0641), .Y(new_n12672_));
  AOI21X1  g10236(.A0(new_n12660_), .A1(new_n12664_), .B0(new_n12672_), .Y(new_n12673_));
  OAI21X1  g10237(.A0(new_n12657_), .A1(new_n12664_), .B0(new_n12673_), .Y(new_n12674_));
  AND2X1   g10238(.A(pi1158), .B(pi0641), .Y(new_n12675_));
  INVX1    g10239(.A(pi1158), .Y(new_n12676_));
  AOI21X1  g10240(.A0(new_n12597_), .A1(new_n12664_), .B0(new_n12676_), .Y(new_n12677_));
  INVX1    g10241(.A(new_n12677_), .Y(new_n12678_));
  AOI21X1  g10242(.A0(new_n12667_), .A1(pi0626), .B0(new_n12678_), .Y(new_n12679_));
  OR2X1    g10243(.A(new_n12679_), .B(new_n12675_), .Y(new_n12680_));
  AOI22X1  g10244(.A0(new_n12680_), .A1(new_n12674_), .B0(new_n12671_), .B1(new_n12662_), .Y(new_n12681_));
  MX2X1    g10245(.A(new_n12681_), .B(new_n12657_), .S0(new_n11885_), .Y(new_n12682_));
  INVX1    g10246(.A(pi0628), .Y(new_n12683_));
  INVX1    g10247(.A(pi1156), .Y(new_n12684_));
  OAI21X1  g10248(.A0(new_n12679_), .A1(new_n12670_), .B0(pi0788), .Y(new_n12685_));
  OAI21X1  g10249(.A0(new_n12667_), .A1(pi0788), .B0(new_n12685_), .Y(new_n12686_));
  OAI21X1  g10250(.A0(new_n12686_), .A1(new_n12683_), .B0(new_n12684_), .Y(new_n12687_));
  AOI21X1  g10251(.A0(new_n12682_), .A1(new_n12683_), .B0(new_n12687_), .Y(new_n12688_));
  INVX1    g10252(.A(pi0629), .Y(new_n12689_));
  XOR2X1   g10253(.A(pi1158), .B(new_n12672_), .Y(new_n12690_));
  NOR2X1   g10254(.A(new_n12690_), .B(new_n11885_), .Y(new_n12691_));
  MX2X1    g10255(.A(new_n12660_), .B(new_n12578_), .S0(new_n12691_), .Y(new_n12692_));
  AOI21X1  g10256(.A0(new_n12597_), .A1(new_n12683_), .B0(new_n12684_), .Y(new_n12693_));
  OAI21X1  g10257(.A0(new_n12692_), .A1(new_n12683_), .B0(new_n12693_), .Y(new_n12694_));
  AND2X1   g10258(.A(new_n12694_), .B(new_n12689_), .Y(new_n12695_));
  INVX1    g10259(.A(new_n12695_), .Y(new_n12696_));
  OAI21X1  g10260(.A0(new_n12686_), .A1(pi0628), .B0(pi1156), .Y(new_n12697_));
  AOI21X1  g10261(.A0(new_n12682_), .A1(pi0628), .B0(new_n12697_), .Y(new_n12698_));
  AOI21X1  g10262(.A0(new_n12597_), .A1(pi0628), .B0(pi1156), .Y(new_n12699_));
  OAI21X1  g10263(.A0(new_n12692_), .A1(pi0628), .B0(new_n12699_), .Y(new_n12700_));
  AND2X1   g10264(.A(new_n12700_), .B(pi0629), .Y(new_n12701_));
  INVX1    g10265(.A(new_n12701_), .Y(new_n12702_));
  OAI22X1  g10266(.A0(new_n12702_), .A1(new_n12698_), .B0(new_n12696_), .B1(new_n12688_), .Y(new_n12703_));
  MX2X1    g10267(.A(new_n12703_), .B(new_n12682_), .S0(new_n11884_), .Y(new_n12704_));
  INVX1    g10268(.A(pi0647), .Y(new_n12705_));
  INVX1    g10269(.A(pi1157), .Y(new_n12706_));
  AND2X1   g10270(.A(pi1156), .B(new_n12689_), .Y(new_n12707_));
  INVX1    g10271(.A(new_n12707_), .Y(new_n12708_));
  AND2X1   g10272(.A(new_n12684_), .B(pi0629), .Y(new_n12709_));
  INVX1    g10273(.A(new_n12709_), .Y(new_n12710_));
  AOI21X1  g10274(.A0(new_n12710_), .A1(new_n12708_), .B0(new_n11884_), .Y(new_n12711_));
  MX2X1    g10275(.A(new_n12686_), .B(new_n12578_), .S0(new_n12711_), .Y(new_n12712_));
  OAI21X1  g10276(.A0(new_n12712_), .A1(new_n12705_), .B0(new_n12706_), .Y(new_n12713_));
  AOI21X1  g10277(.A0(new_n12704_), .A1(new_n12705_), .B0(new_n12713_), .Y(new_n12714_));
  AOI21X1  g10278(.A0(new_n12700_), .A1(new_n12694_), .B0(new_n11884_), .Y(new_n12715_));
  AOI21X1  g10279(.A0(new_n12692_), .A1(new_n11884_), .B0(new_n12715_), .Y(new_n12716_));
  OAI21X1  g10280(.A0(new_n12578_), .A1(pi0647), .B0(pi1157), .Y(new_n12717_));
  AOI21X1  g10281(.A0(new_n12716_), .A1(pi0647), .B0(new_n12717_), .Y(new_n12718_));
  NOR2X1   g10282(.A(new_n12718_), .B(pi0630), .Y(new_n12719_));
  INVX1    g10283(.A(new_n12719_), .Y(new_n12720_));
  OAI21X1  g10284(.A0(new_n12712_), .A1(pi0647), .B0(pi1157), .Y(new_n12721_));
  AOI21X1  g10285(.A0(new_n12704_), .A1(pi0647), .B0(new_n12721_), .Y(new_n12722_));
  INVX1    g10286(.A(pi0630), .Y(new_n12723_));
  OAI21X1  g10287(.A0(new_n12578_), .A1(new_n12705_), .B0(new_n12706_), .Y(new_n12724_));
  AOI21X1  g10288(.A0(new_n12716_), .A1(new_n12705_), .B0(new_n12724_), .Y(new_n12725_));
  NOR2X1   g10289(.A(new_n12725_), .B(new_n12723_), .Y(new_n12726_));
  INVX1    g10290(.A(new_n12726_), .Y(new_n12727_));
  OAI22X1  g10291(.A0(new_n12727_), .A1(new_n12722_), .B0(new_n12720_), .B1(new_n12714_), .Y(new_n12728_));
  MX2X1    g10292(.A(new_n12728_), .B(new_n12704_), .S0(new_n11883_), .Y(new_n12729_));
  OAI21X1  g10293(.A0(new_n12725_), .A1(new_n12718_), .B0(pi0787), .Y(new_n12730_));
  OAI21X1  g10294(.A0(new_n12716_), .A1(pi0787), .B0(new_n12730_), .Y(new_n12731_));
  OAI21X1  g10295(.A0(new_n12731_), .A1(pi0644), .B0(pi0715), .Y(new_n12732_));
  AOI21X1  g10296(.A0(new_n12729_), .A1(pi0644), .B0(new_n12732_), .Y(new_n12733_));
  XOR2X1   g10297(.A(pi1157), .B(new_n12723_), .Y(new_n12734_));
  NOR2X1   g10298(.A(new_n12734_), .B(new_n11883_), .Y(new_n12735_));
  INVX1    g10299(.A(new_n12735_), .Y(new_n12736_));
  AND2X1   g10300(.A(new_n12735_), .B(new_n12578_), .Y(new_n12737_));
  AOI21X1  g10301(.A0(new_n12736_), .A1(new_n12712_), .B0(new_n12737_), .Y(new_n12738_));
  INVX1    g10302(.A(pi0715), .Y(new_n12739_));
  OAI21X1  g10303(.A0(new_n12578_), .A1(pi0644), .B0(new_n12739_), .Y(new_n12740_));
  AOI21X1  g10304(.A0(new_n12738_), .A1(pi0644), .B0(new_n12740_), .Y(new_n12741_));
  NOR3X1   g10305(.A(new_n12741_), .B(new_n12733_), .C(new_n11882_), .Y(new_n12742_));
  INVX1    g10306(.A(pi0644), .Y(new_n12743_));
  OAI21X1  g10307(.A0(new_n12731_), .A1(new_n12743_), .B0(new_n12739_), .Y(new_n12744_));
  AOI21X1  g10308(.A0(new_n12729_), .A1(new_n12743_), .B0(new_n12744_), .Y(new_n12745_));
  OAI21X1  g10309(.A0(new_n12578_), .A1(new_n12743_), .B0(pi0715), .Y(new_n12746_));
  AOI21X1  g10310(.A0(new_n12738_), .A1(new_n12743_), .B0(new_n12746_), .Y(new_n12747_));
  OR2X1    g10311(.A(new_n12747_), .B(pi1160), .Y(new_n12748_));
  OAI21X1  g10312(.A0(new_n12748_), .A1(new_n12745_), .B0(pi0790), .Y(new_n12749_));
  OR2X1    g10313(.A(new_n12729_), .B(pi0790), .Y(new_n12750_));
  AND2X1   g10314(.A(new_n12750_), .B(new_n6520_), .Y(new_n12751_));
  OAI21X1  g10315(.A0(new_n12749_), .A1(new_n12742_), .B0(new_n12751_), .Y(new_n12752_));
  AOI21X1  g10316(.A0(po1038), .A1(new_n7398_), .B0(pi0832), .Y(new_n12753_));
  AOI21X1  g10317(.A0(pi1093), .A1(pi1092), .B0(pi0140), .Y(new_n12754_));
  AOI21X1  g10318(.A0(new_n12566_), .A1(new_n12565_), .B0(new_n12754_), .Y(new_n12755_));
  AND2X1   g10319(.A(new_n12566_), .B(new_n12565_), .Y(new_n12756_));
  AND2X1   g10320(.A(new_n12756_), .B(new_n12493_), .Y(new_n12757_));
  MX2X1    g10321(.A(new_n12754_), .B(pi0625), .S0(new_n12756_), .Y(new_n12758_));
  OR2X1    g10322(.A(new_n12754_), .B(pi1153), .Y(new_n12759_));
  OAI22X1  g10323(.A0(new_n12759_), .A1(new_n12757_), .B0(new_n12758_), .B1(new_n12494_), .Y(new_n12760_));
  MX2X1    g10324(.A(new_n12760_), .B(new_n12755_), .S0(new_n11889_), .Y(new_n12761_));
  AND2X1   g10325(.A(new_n12618_), .B(new_n2739_), .Y(new_n12762_));
  OR2X1    g10326(.A(new_n12762_), .B(new_n12761_), .Y(new_n12763_));
  NOR4X1   g10327(.A(new_n12640_), .B(new_n12639_), .C(new_n2756_), .D(new_n2755_), .Y(new_n12764_));
  NOR3X1   g10328(.A(new_n12658_), .B(new_n2740_), .C(new_n11886_), .Y(new_n12765_));
  XOR2X1   g10329(.A(pi1158), .B(pi0626), .Y(new_n12766_));
  XOR2X1   g10330(.A(pi0641), .B(new_n12664_), .Y(new_n12767_));
  INVX1    g10331(.A(new_n12767_), .Y(new_n12768_));
  AND2X1   g10332(.A(new_n12768_), .B(new_n12766_), .Y(new_n12769_));
  INVX1    g10333(.A(new_n12769_), .Y(new_n12770_));
  NOR4X1   g10334(.A(new_n12770_), .B(new_n12765_), .C(new_n12764_), .D(new_n12763_), .Y(new_n12771_));
  AOI21X1  g10335(.A0(new_n12178_), .A1(new_n11890_), .B0(new_n12754_), .Y(new_n12772_));
  AOI21X1  g10336(.A0(new_n12601_), .A1(new_n2739_), .B0(new_n12772_), .Y(new_n12773_));
  INVX1    g10337(.A(new_n12772_), .Y(new_n12774_));
  NOR2X1   g10338(.A(new_n12599_), .B(new_n2740_), .Y(new_n12775_));
  INVX1    g10339(.A(new_n12775_), .Y(new_n12776_));
  AOI21X1  g10340(.A0(new_n12776_), .A1(new_n12774_), .B0(new_n12591_), .Y(new_n12777_));
  AND2X1   g10341(.A(new_n2739_), .B(pi0609), .Y(new_n12778_));
  INVX1    g10342(.A(new_n12778_), .Y(new_n12779_));
  AOI21X1  g10343(.A0(new_n12779_), .A1(new_n12773_), .B0(pi1155), .Y(new_n12780_));
  OAI21X1  g10344(.A0(new_n12780_), .A1(new_n12777_), .B0(pi0785), .Y(new_n12781_));
  OAI21X1  g10345(.A0(new_n12773_), .A1(pi0785), .B0(new_n12781_), .Y(new_n12782_));
  INVX1    g10346(.A(new_n12782_), .Y(new_n12783_));
  AND2X1   g10347(.A(new_n2739_), .B(new_n12614_), .Y(new_n12784_));
  INVX1    g10348(.A(new_n12784_), .Y(new_n12785_));
  AOI21X1  g10349(.A0(new_n12785_), .A1(new_n12783_), .B0(new_n12615_), .Y(new_n12786_));
  AND2X1   g10350(.A(new_n2739_), .B(pi0618), .Y(new_n12787_));
  INVX1    g10351(.A(new_n12787_), .Y(new_n12788_));
  AOI21X1  g10352(.A0(new_n12788_), .A1(new_n12783_), .B0(pi1154), .Y(new_n12789_));
  OR2X1    g10353(.A(new_n12789_), .B(new_n12786_), .Y(new_n12790_));
  MX2X1    g10354(.A(new_n12790_), .B(new_n12782_), .S0(new_n11887_), .Y(new_n12791_));
  AOI21X1  g10355(.A0(new_n12754_), .A1(new_n12637_), .B0(new_n12638_), .Y(new_n12792_));
  OAI21X1  g10356(.A0(new_n12791_), .A1(new_n12637_), .B0(new_n12792_), .Y(new_n12793_));
  AOI21X1  g10357(.A0(new_n12754_), .A1(pi0619), .B0(pi1159), .Y(new_n12794_));
  OAI21X1  g10358(.A0(new_n12791_), .A1(pi0619), .B0(new_n12794_), .Y(new_n12795_));
  AOI21X1  g10359(.A0(new_n12795_), .A1(new_n12793_), .B0(new_n11886_), .Y(new_n12796_));
  AOI21X1  g10360(.A0(new_n12791_), .A1(new_n11886_), .B0(new_n12796_), .Y(new_n12797_));
  INVX1    g10361(.A(new_n12754_), .Y(new_n12798_));
  OAI21X1  g10362(.A0(new_n12798_), .A1(pi0626), .B0(pi1158), .Y(new_n12799_));
  AOI21X1  g10363(.A0(new_n12797_), .A1(pi0626), .B0(new_n12799_), .Y(new_n12800_));
  OAI21X1  g10364(.A0(new_n12798_), .A1(new_n12664_), .B0(new_n12676_), .Y(new_n12801_));
  AOI21X1  g10365(.A0(new_n12797_), .A1(new_n12664_), .B0(new_n12801_), .Y(new_n12802_));
  NOR3X1   g10366(.A(new_n12802_), .B(new_n12800_), .C(new_n12690_), .Y(new_n12803_));
  OAI21X1  g10367(.A0(new_n12803_), .A1(new_n12771_), .B0(pi0788), .Y(new_n12804_));
  OAI21X1  g10368(.A0(new_n12755_), .A1(new_n12120_), .B0(new_n12772_), .Y(new_n12805_));
  NOR2X1   g10369(.A(new_n12755_), .B(new_n12120_), .Y(new_n12806_));
  MX2X1    g10370(.A(new_n12774_), .B(new_n12493_), .S0(new_n12806_), .Y(new_n12807_));
  NOR2X1   g10371(.A(new_n12807_), .B(new_n12759_), .Y(new_n12808_));
  OAI21X1  g10372(.A0(new_n12758_), .A1(new_n12494_), .B0(new_n12584_), .Y(new_n12809_));
  NOR3X1   g10373(.A(new_n12755_), .B(new_n12120_), .C(new_n12493_), .Y(new_n12810_));
  NOR3X1   g10374(.A(new_n12810_), .B(new_n12774_), .C(new_n12494_), .Y(new_n12811_));
  OAI21X1  g10375(.A0(new_n12759_), .A1(new_n12757_), .B0(pi0608), .Y(new_n12812_));
  OAI22X1  g10376(.A0(new_n12812_), .A1(new_n12811_), .B0(new_n12809_), .B1(new_n12808_), .Y(new_n12813_));
  MX2X1    g10377(.A(new_n12813_), .B(new_n12805_), .S0(new_n11889_), .Y(new_n12814_));
  OAI21X1  g10378(.A0(new_n12761_), .A1(new_n12590_), .B0(new_n12591_), .Y(new_n12815_));
  AOI21X1  g10379(.A0(new_n12814_), .A1(new_n12590_), .B0(new_n12815_), .Y(new_n12816_));
  OR2X1    g10380(.A(new_n12777_), .B(pi0660), .Y(new_n12817_));
  OAI21X1  g10381(.A0(new_n12761_), .A1(pi0609), .B0(pi1155), .Y(new_n12818_));
  AOI21X1  g10382(.A0(new_n12814_), .A1(pi0609), .B0(new_n12818_), .Y(new_n12819_));
  OR2X1    g10383(.A(new_n12780_), .B(new_n12596_), .Y(new_n12820_));
  OAI22X1  g10384(.A0(new_n12820_), .A1(new_n12819_), .B0(new_n12817_), .B1(new_n12816_), .Y(new_n12821_));
  MX2X1    g10385(.A(new_n12821_), .B(new_n12814_), .S0(new_n11888_), .Y(new_n12822_));
  OAI21X1  g10386(.A0(new_n12763_), .A1(new_n12614_), .B0(new_n12615_), .Y(new_n12823_));
  AOI21X1  g10387(.A0(new_n12822_), .A1(new_n12614_), .B0(new_n12823_), .Y(new_n12824_));
  OR2X1    g10388(.A(new_n12786_), .B(pi0627), .Y(new_n12825_));
  OAI21X1  g10389(.A0(new_n12763_), .A1(pi0618), .B0(pi1154), .Y(new_n12826_));
  AOI21X1  g10390(.A0(new_n12822_), .A1(pi0618), .B0(new_n12826_), .Y(new_n12827_));
  OR2X1    g10391(.A(new_n12789_), .B(new_n12622_), .Y(new_n12828_));
  OAI22X1  g10392(.A0(new_n12828_), .A1(new_n12827_), .B0(new_n12825_), .B1(new_n12824_), .Y(new_n12829_));
  MX2X1    g10393(.A(new_n12829_), .B(new_n12822_), .S0(new_n11887_), .Y(new_n12830_));
  NAND2X1  g10394(.A(new_n12830_), .B(new_n12637_), .Y(new_n12831_));
  NOR3X1   g10395(.A(new_n12764_), .B(new_n12762_), .C(new_n12761_), .Y(new_n12832_));
  AOI21X1  g10396(.A0(new_n12832_), .A1(pi0619), .B0(pi1159), .Y(new_n12833_));
  NAND2X1  g10397(.A(new_n12793_), .B(new_n12645_), .Y(new_n12834_));
  AOI21X1  g10398(.A0(new_n12833_), .A1(new_n12831_), .B0(new_n12834_), .Y(new_n12835_));
  NAND2X1  g10399(.A(new_n12830_), .B(pi0619), .Y(new_n12836_));
  AOI21X1  g10400(.A0(new_n12832_), .A1(new_n12637_), .B0(new_n12638_), .Y(new_n12837_));
  NAND2X1  g10401(.A(new_n12795_), .B(pi0648), .Y(new_n12838_));
  AOI21X1  g10402(.A0(new_n12837_), .A1(new_n12836_), .B0(new_n12838_), .Y(new_n12839_));
  NOR3X1   g10403(.A(new_n12839_), .B(new_n12835_), .C(new_n11886_), .Y(new_n12840_));
  AND2X1   g10404(.A(new_n12766_), .B(pi0788), .Y(new_n12841_));
  NOR2X1   g10405(.A(new_n12841_), .B(new_n12691_), .Y(new_n12842_));
  OAI21X1  g10406(.A0(new_n12830_), .A1(pi0789), .B0(new_n12842_), .Y(new_n12843_));
  OAI21X1  g10407(.A0(new_n12843_), .A1(new_n12840_), .B0(new_n12804_), .Y(new_n12844_));
  NOR2X1   g10408(.A(new_n12802_), .B(new_n12800_), .Y(new_n12845_));
  MX2X1    g10409(.A(new_n12845_), .B(new_n12797_), .S0(new_n11885_), .Y(new_n12846_));
  INVX1    g10410(.A(new_n12846_), .Y(new_n12847_));
  OAI21X1  g10411(.A0(new_n12847_), .A1(new_n12683_), .B0(new_n12684_), .Y(new_n12848_));
  AOI21X1  g10412(.A0(new_n12844_), .A1(new_n12683_), .B0(new_n12848_), .Y(new_n12849_));
  INVX1    g10413(.A(new_n12765_), .Y(new_n12850_));
  NOR3X1   g10414(.A(new_n12690_), .B(new_n2740_), .C(new_n11885_), .Y(new_n12851_));
  INVX1    g10415(.A(new_n12851_), .Y(new_n12852_));
  NAND3X1  g10416(.A(new_n12852_), .B(new_n12850_), .C(new_n12832_), .Y(new_n12853_));
  AOI21X1  g10417(.A0(new_n2739_), .A1(new_n12683_), .B0(new_n12853_), .Y(new_n12854_));
  OAI21X1  g10418(.A0(new_n12854_), .A1(new_n12684_), .B0(new_n12689_), .Y(new_n12855_));
  OAI21X1  g10419(.A0(new_n12847_), .A1(pi0628), .B0(pi1156), .Y(new_n12856_));
  AOI21X1  g10420(.A0(new_n12844_), .A1(pi0628), .B0(new_n12856_), .Y(new_n12857_));
  AOI21X1  g10421(.A0(new_n2739_), .A1(pi0628), .B0(new_n12853_), .Y(new_n12858_));
  OAI21X1  g10422(.A0(new_n12858_), .A1(pi1156), .B0(pi0629), .Y(new_n12859_));
  OAI22X1  g10423(.A0(new_n12859_), .A1(new_n12857_), .B0(new_n12855_), .B1(new_n12849_), .Y(new_n12860_));
  MX2X1    g10424(.A(new_n12860_), .B(new_n12844_), .S0(new_n11884_), .Y(new_n12861_));
  MX2X1    g10425(.A(new_n12847_), .B(new_n12798_), .S0(new_n12711_), .Y(new_n12862_));
  OAI21X1  g10426(.A0(new_n12862_), .A1(new_n12705_), .B0(new_n12706_), .Y(new_n12863_));
  AOI21X1  g10427(.A0(new_n12861_), .A1(new_n12705_), .B0(new_n12863_), .Y(new_n12864_));
  AND2X1   g10428(.A(pi1156), .B(new_n12683_), .Y(new_n12865_));
  INVX1    g10429(.A(new_n12865_), .Y(new_n12866_));
  AND2X1   g10430(.A(new_n12684_), .B(pi0628), .Y(new_n12867_));
  INVX1    g10431(.A(new_n12867_), .Y(new_n12868_));
  AOI21X1  g10432(.A0(new_n12868_), .A1(new_n12866_), .B0(new_n11884_), .Y(new_n12869_));
  AND2X1   g10433(.A(new_n12869_), .B(new_n2739_), .Y(new_n12870_));
  NOR2X1   g10434(.A(new_n12870_), .B(new_n12853_), .Y(new_n12871_));
  OAI21X1  g10435(.A0(new_n12798_), .A1(pi0647), .B0(pi1157), .Y(new_n12872_));
  AOI21X1  g10436(.A0(new_n12871_), .A1(pi0647), .B0(new_n12872_), .Y(new_n12873_));
  OR2X1    g10437(.A(new_n12873_), .B(pi0630), .Y(new_n12874_));
  OAI21X1  g10438(.A0(new_n12862_), .A1(pi0647), .B0(pi1157), .Y(new_n12875_));
  AOI21X1  g10439(.A0(new_n12861_), .A1(pi0647), .B0(new_n12875_), .Y(new_n12876_));
  OAI21X1  g10440(.A0(new_n12798_), .A1(new_n12705_), .B0(new_n12706_), .Y(new_n12877_));
  AOI21X1  g10441(.A0(new_n12871_), .A1(new_n12705_), .B0(new_n12877_), .Y(new_n12878_));
  OR2X1    g10442(.A(new_n12878_), .B(new_n12723_), .Y(new_n12879_));
  OAI22X1  g10443(.A0(new_n12879_), .A1(new_n12876_), .B0(new_n12874_), .B1(new_n12864_), .Y(new_n12880_));
  MX2X1    g10444(.A(new_n12880_), .B(new_n12861_), .S0(new_n11883_), .Y(new_n12881_));
  OAI21X1  g10445(.A0(new_n12878_), .A1(new_n12873_), .B0(pi0787), .Y(new_n12882_));
  OAI21X1  g10446(.A0(new_n12871_), .A1(pi0787), .B0(new_n12882_), .Y(new_n12883_));
  OAI21X1  g10447(.A0(new_n12883_), .A1(pi0644), .B0(pi0715), .Y(new_n12884_));
  AOI21X1  g10448(.A0(new_n12881_), .A1(pi0644), .B0(new_n12884_), .Y(new_n12885_));
  NOR3X1   g10449(.A(new_n12754_), .B(new_n12734_), .C(new_n11883_), .Y(new_n12886_));
  AOI21X1  g10450(.A0(new_n12862_), .A1(new_n12736_), .B0(new_n12886_), .Y(new_n12887_));
  OAI21X1  g10451(.A0(new_n12798_), .A1(pi0644), .B0(new_n12739_), .Y(new_n12888_));
  AOI21X1  g10452(.A0(new_n12887_), .A1(pi0644), .B0(new_n12888_), .Y(new_n12889_));
  NOR3X1   g10453(.A(new_n12889_), .B(new_n12885_), .C(new_n11882_), .Y(new_n12890_));
  OAI21X1  g10454(.A0(new_n12883_), .A1(new_n12743_), .B0(new_n12739_), .Y(new_n12891_));
  AOI21X1  g10455(.A0(new_n12881_), .A1(new_n12743_), .B0(new_n12891_), .Y(new_n12892_));
  OAI21X1  g10456(.A0(new_n12798_), .A1(new_n12743_), .B0(pi0715), .Y(new_n12893_));
  AOI21X1  g10457(.A0(new_n12887_), .A1(new_n12743_), .B0(new_n12893_), .Y(new_n12894_));
  NOR3X1   g10458(.A(new_n12894_), .B(new_n12892_), .C(pi1160), .Y(new_n12895_));
  OAI21X1  g10459(.A0(new_n12895_), .A1(new_n12890_), .B0(pi0790), .Y(new_n12896_));
  INVX1    g10460(.A(pi0790), .Y(new_n12897_));
  INVX1    g10461(.A(pi0832), .Y(new_n12898_));
  AOI21X1  g10462(.A0(new_n12881_), .A1(new_n12897_), .B0(new_n12898_), .Y(new_n12899_));
  AOI22X1  g10463(.A0(new_n12899_), .A1(new_n12896_), .B0(new_n12753_), .B1(new_n12752_), .Y(po0297));
  INVX1    g10464(.A(new_n12202_), .Y(new_n12901_));
  AOI22X1  g10465(.A0(new_n12205_), .A1(pi0749), .B0(new_n12901_), .B1(new_n7382_), .Y(new_n12902_));
  NOR2X1   g10466(.A(new_n12902_), .B(new_n2996_), .Y(new_n12903_));
  INVX1    g10467(.A(new_n12198_), .Y(new_n12904_));
  OAI22X1  g10468(.A0(new_n12904_), .A1(new_n7382_), .B0(new_n12089_), .B1(pi0749), .Y(new_n12905_));
  NAND2X1  g10469(.A(new_n12905_), .B(pi0039), .Y(new_n12906_));
  NOR2X1   g10470(.A(new_n12097_), .B(new_n2953_), .Y(new_n12907_));
  NOR2X1   g10471(.A(new_n12103_), .B(pi0299), .Y(new_n12908_));
  OR2X1    g10472(.A(new_n12908_), .B(new_n12907_), .Y(new_n12909_));
  MX2X1    g10473(.A(new_n12161_), .B(new_n12909_), .S0(new_n2959_), .Y(new_n12910_));
  INVX1    g10474(.A(pi0749), .Y(new_n12911_));
  AOI21X1  g10475(.A0(new_n12169_), .A1(pi0141), .B0(new_n12911_), .Y(new_n12912_));
  OAI21X1  g10476(.A0(new_n12910_), .A1(pi0141), .B0(new_n12912_), .Y(new_n12913_));
  NAND2X1  g10477(.A(new_n11947_), .B(new_n2959_), .Y(new_n12914_));
  NAND3X1  g10478(.A(new_n12914_), .B(new_n12911_), .C(new_n7382_), .Y(new_n12915_));
  AOI21X1  g10479(.A0(new_n12915_), .A1(new_n12913_), .B0(pi0038), .Y(new_n12916_));
  AOI21X1  g10480(.A0(new_n12916_), .A1(new_n12906_), .B0(new_n12903_), .Y(new_n12917_));
  OR2X1    g10481(.A(new_n12917_), .B(pi0706), .Y(new_n12918_));
  OAI21X1  g10482(.A0(new_n12349_), .A1(new_n7382_), .B0(new_n12911_), .Y(new_n12919_));
  AOI21X1  g10483(.A0(new_n12289_), .A1(new_n7382_), .B0(new_n12919_), .Y(new_n12920_));
  OAI21X1  g10484(.A0(new_n12440_), .A1(pi0141), .B0(pi0749), .Y(new_n12921_));
  AOI21X1  g10485(.A0(new_n12401_), .A1(pi0141), .B0(new_n12921_), .Y(new_n12922_));
  OR2X1    g10486(.A(new_n12922_), .B(new_n2959_), .Y(new_n12923_));
  AND2X1   g10487(.A(new_n12454_), .B(new_n7382_), .Y(new_n12924_));
  OAI21X1  g10488(.A0(new_n12467_), .A1(new_n7382_), .B0(new_n12911_), .Y(new_n12925_));
  OR2X1    g10489(.A(new_n12925_), .B(new_n12924_), .Y(new_n12926_));
  NAND2X1  g10490(.A(new_n12453_), .B(new_n12104_), .Y(new_n12927_));
  NAND2X1  g10491(.A(new_n12927_), .B(new_n7382_), .Y(new_n12928_));
  OR2X1    g10492(.A(new_n12473_), .B(new_n12168_), .Y(new_n12929_));
  AOI21X1  g10493(.A0(new_n12929_), .A1(pi0141), .B0(new_n12911_), .Y(new_n12930_));
  AOI21X1  g10494(.A0(new_n12930_), .A1(new_n12928_), .B0(pi0039), .Y(new_n12931_));
  AOI21X1  g10495(.A0(new_n12931_), .A1(new_n12926_), .B0(pi0038), .Y(new_n12932_));
  OAI21X1  g10496(.A0(new_n12923_), .A1(new_n12920_), .B0(new_n12932_), .Y(new_n12933_));
  INVX1    g10497(.A(pi0706), .Y(new_n12934_));
  AOI21X1  g10498(.A0(new_n12483_), .A1(new_n2959_), .B0(new_n2996_), .Y(new_n12935_));
  AOI21X1  g10499(.A0(new_n12935_), .A1(new_n12902_), .B0(new_n12934_), .Y(new_n12936_));
  AOI21X1  g10500(.A0(new_n12936_), .A1(new_n12933_), .B0(new_n3810_), .Y(new_n12937_));
  AOI22X1  g10501(.A0(new_n12937_), .A1(new_n12918_), .B0(new_n3810_), .B1(pi0141), .Y(new_n12938_));
  MX2X1    g10502(.A(new_n12917_), .B(pi0141), .S0(new_n3810_), .Y(new_n12939_));
  OAI21X1  g10503(.A0(new_n12939_), .A1(new_n12493_), .B0(new_n12494_), .Y(new_n12940_));
  AOI21X1  g10504(.A0(new_n12938_), .A1(new_n12493_), .B0(new_n12940_), .Y(new_n12941_));
  INVX1    g10505(.A(new_n12527_), .Y(new_n12942_));
  OAI21X1  g10506(.A0(new_n12071_), .A1(pi0680), .B0(new_n12942_), .Y(new_n12943_));
  OAI21X1  g10507(.A0(new_n12071_), .A1(pi0680), .B0(new_n12530_), .Y(new_n12944_));
  OAI21X1  g10508(.A0(new_n12943_), .A1(new_n11993_), .B0(new_n12944_), .Y(new_n12945_));
  OAI21X1  g10509(.A0(new_n12945_), .A1(new_n5051_), .B0(new_n12536_), .Y(new_n12946_));
  NOR2X1   g10510(.A(new_n12548_), .B(new_n12543_), .Y(new_n12947_));
  AOI21X1  g10511(.A0(new_n12539_), .A1(new_n12946_), .B0(new_n12947_), .Y(new_n12948_));
  OAI21X1  g10512(.A0(new_n12945_), .A1(new_n5071_), .B0(new_n12550_), .Y(new_n12949_));
  NOR2X1   g10513(.A(new_n12558_), .B(new_n12556_), .Y(new_n12950_));
  AOI21X1  g10514(.A0(new_n12554_), .A1(new_n12949_), .B0(new_n12950_), .Y(new_n12951_));
  MX2X1    g10515(.A(new_n12951_), .B(new_n12948_), .S0(new_n2953_), .Y(new_n12952_));
  MX2X1    g10516(.A(new_n12952_), .B(new_n12453_), .S0(new_n2959_), .Y(new_n12953_));
  NAND2X1  g10517(.A(new_n12473_), .B(new_n2959_), .Y(new_n12954_));
  OAI21X1  g10518(.A0(new_n12522_), .A1(new_n2959_), .B0(new_n12954_), .Y(new_n12955_));
  AOI21X1  g10519(.A0(new_n12955_), .A1(pi0141), .B0(pi0038), .Y(new_n12956_));
  OAI21X1  g10520(.A0(new_n12953_), .A1(pi0141), .B0(new_n12956_), .Y(new_n12957_));
  OR2X1    g10521(.A(new_n12202_), .B(pi0141), .Y(new_n12958_));
  AOI21X1  g10522(.A0(new_n12958_), .A1(new_n12567_), .B0(new_n12934_), .Y(new_n12959_));
  NAND2X1  g10523(.A(new_n12959_), .B(new_n12957_), .Y(new_n12960_));
  NOR2X1   g10524(.A(pi0706), .B(pi0141), .Y(new_n12961_));
  AOI21X1  g10525(.A0(new_n12961_), .A1(new_n12574_), .B0(new_n3810_), .Y(new_n12962_));
  AOI22X1  g10526(.A0(new_n12962_), .A1(new_n12960_), .B0(new_n3810_), .B1(pi0141), .Y(new_n12963_));
  OAI21X1  g10527(.A0(new_n12574_), .A1(new_n3810_), .B0(new_n7382_), .Y(new_n12964_));
  OAI21X1  g10528(.A0(new_n12964_), .A1(pi0625), .B0(pi1153), .Y(new_n12965_));
  AOI21X1  g10529(.A0(new_n12963_), .A1(pi0625), .B0(new_n12965_), .Y(new_n12966_));
  OR2X1    g10530(.A(new_n12966_), .B(pi0608), .Y(new_n12967_));
  OAI21X1  g10531(.A0(new_n12939_), .A1(pi0625), .B0(pi1153), .Y(new_n12968_));
  AOI21X1  g10532(.A0(new_n12938_), .A1(pi0625), .B0(new_n12968_), .Y(new_n12969_));
  OAI21X1  g10533(.A0(new_n12964_), .A1(new_n12493_), .B0(new_n12494_), .Y(new_n12970_));
  AOI21X1  g10534(.A0(new_n12963_), .A1(new_n12493_), .B0(new_n12970_), .Y(new_n12971_));
  OR2X1    g10535(.A(new_n12971_), .B(new_n12584_), .Y(new_n12972_));
  OAI22X1  g10536(.A0(new_n12972_), .A1(new_n12969_), .B0(new_n12967_), .B1(new_n12941_), .Y(new_n12973_));
  MX2X1    g10537(.A(new_n12973_), .B(new_n12938_), .S0(new_n11889_), .Y(new_n12974_));
  OAI21X1  g10538(.A0(new_n12971_), .A1(new_n12966_), .B0(pi0778), .Y(new_n12975_));
  OAI21X1  g10539(.A0(new_n12963_), .A1(pi0778), .B0(new_n12975_), .Y(new_n12976_));
  OAI21X1  g10540(.A0(new_n12976_), .A1(new_n12590_), .B0(new_n12591_), .Y(new_n12977_));
  AOI21X1  g10541(.A0(new_n12974_), .A1(new_n12590_), .B0(new_n12977_), .Y(new_n12978_));
  INVX1    g10542(.A(new_n12964_), .Y(new_n12979_));
  NAND2X1  g10543(.A(new_n12939_), .B(new_n12623_), .Y(new_n12980_));
  OAI22X1  g10544(.A0(new_n12980_), .A1(new_n12590_), .B0(new_n12979_), .B1(new_n12599_), .Y(new_n12981_));
  NAND2X1  g10545(.A(new_n12981_), .B(pi1155), .Y(new_n12982_));
  NAND2X1  g10546(.A(new_n12982_), .B(new_n12596_), .Y(new_n12983_));
  OAI21X1  g10547(.A0(new_n12976_), .A1(pi0609), .B0(pi1155), .Y(new_n12984_));
  AOI21X1  g10548(.A0(new_n12974_), .A1(pi0609), .B0(new_n12984_), .Y(new_n12985_));
  OAI22X1  g10549(.A0(new_n12980_), .A1(pi0609), .B0(new_n12979_), .B1(new_n12608_), .Y(new_n12986_));
  NAND2X1  g10550(.A(new_n12986_), .B(new_n12591_), .Y(new_n12987_));
  NAND2X1  g10551(.A(new_n12987_), .B(pi0660), .Y(new_n12988_));
  OAI22X1  g10552(.A0(new_n12988_), .A1(new_n12985_), .B0(new_n12983_), .B1(new_n12978_), .Y(new_n12989_));
  MX2X1    g10553(.A(new_n12989_), .B(new_n12974_), .S0(new_n11888_), .Y(new_n12990_));
  MX2X1    g10554(.A(new_n12976_), .B(new_n12964_), .S0(new_n12618_), .Y(new_n12991_));
  OAI21X1  g10555(.A0(new_n12991_), .A1(new_n12614_), .B0(new_n12615_), .Y(new_n12992_));
  AOI21X1  g10556(.A0(new_n12990_), .A1(new_n12614_), .B0(new_n12992_), .Y(new_n12993_));
  MX2X1    g10557(.A(new_n12964_), .B(new_n12939_), .S0(new_n12623_), .Y(new_n12994_));
  AOI21X1  g10558(.A0(new_n12987_), .A1(new_n12982_), .B0(new_n11888_), .Y(new_n12995_));
  AOI21X1  g10559(.A0(new_n12994_), .A1(new_n11888_), .B0(new_n12995_), .Y(new_n12996_));
  AOI21X1  g10560(.A0(new_n12979_), .A1(new_n12614_), .B0(new_n12615_), .Y(new_n12997_));
  INVX1    g10561(.A(new_n12997_), .Y(new_n12998_));
  AOI21X1  g10562(.A0(new_n12996_), .A1(pi0618), .B0(new_n12998_), .Y(new_n12999_));
  OR2X1    g10563(.A(new_n12999_), .B(pi0627), .Y(new_n13000_));
  OAI21X1  g10564(.A0(new_n12991_), .A1(pi0618), .B0(pi1154), .Y(new_n13001_));
  AOI21X1  g10565(.A0(new_n12990_), .A1(pi0618), .B0(new_n13001_), .Y(new_n13002_));
  AOI21X1  g10566(.A0(new_n12979_), .A1(pi0618), .B0(pi1154), .Y(new_n13003_));
  INVX1    g10567(.A(new_n13003_), .Y(new_n13004_));
  AOI21X1  g10568(.A0(new_n12996_), .A1(new_n12614_), .B0(new_n13004_), .Y(new_n13005_));
  OR2X1    g10569(.A(new_n13005_), .B(new_n12622_), .Y(new_n13006_));
  OAI22X1  g10570(.A0(new_n13006_), .A1(new_n13002_), .B0(new_n13000_), .B1(new_n12993_), .Y(new_n13007_));
  MX2X1    g10571(.A(new_n13007_), .B(new_n12990_), .S0(new_n11887_), .Y(new_n13008_));
  MX2X1    g10572(.A(new_n12991_), .B(new_n12964_), .S0(new_n12641_), .Y(new_n13009_));
  OAI21X1  g10573(.A0(new_n13009_), .A1(new_n12637_), .B0(new_n12638_), .Y(new_n13010_));
  AOI21X1  g10574(.A0(new_n13008_), .A1(new_n12637_), .B0(new_n13010_), .Y(new_n13011_));
  OAI21X1  g10575(.A0(new_n13005_), .A1(new_n12999_), .B0(pi0781), .Y(new_n13012_));
  OAI21X1  g10576(.A0(new_n12996_), .A1(pi0781), .B0(new_n13012_), .Y(new_n13013_));
  AOI21X1  g10577(.A0(new_n12979_), .A1(new_n12637_), .B0(new_n12638_), .Y(new_n13014_));
  OAI21X1  g10578(.A0(new_n13013_), .A1(new_n12637_), .B0(new_n13014_), .Y(new_n13015_));
  NAND2X1  g10579(.A(new_n13015_), .B(new_n12645_), .Y(new_n13016_));
  OAI21X1  g10580(.A0(new_n13009_), .A1(pi0619), .B0(pi1159), .Y(new_n13017_));
  AOI21X1  g10581(.A0(new_n13008_), .A1(pi0619), .B0(new_n13017_), .Y(new_n13018_));
  AOI21X1  g10582(.A0(new_n12979_), .A1(pi0619), .B0(pi1159), .Y(new_n13019_));
  OAI21X1  g10583(.A0(new_n13013_), .A1(pi0619), .B0(new_n13019_), .Y(new_n13020_));
  NAND2X1  g10584(.A(new_n13020_), .B(pi0648), .Y(new_n13021_));
  OAI22X1  g10585(.A0(new_n13021_), .A1(new_n13018_), .B0(new_n13016_), .B1(new_n13011_), .Y(new_n13022_));
  MX2X1    g10586(.A(new_n13022_), .B(new_n13008_), .S0(new_n11886_), .Y(new_n13023_));
  MX2X1    g10587(.A(new_n13009_), .B(new_n12964_), .S0(new_n12659_), .Y(new_n13024_));
  AOI21X1  g10588(.A0(new_n13024_), .A1(pi0626), .B0(pi0641), .Y(new_n13025_));
  OAI21X1  g10589(.A0(new_n13023_), .A1(pi0626), .B0(new_n13025_), .Y(new_n13026_));
  INVX1    g10590(.A(new_n12663_), .Y(new_n13027_));
  NAND2X1  g10591(.A(new_n13020_), .B(new_n13015_), .Y(new_n13028_));
  MX2X1    g10592(.A(new_n13028_), .B(new_n13013_), .S0(new_n11886_), .Y(new_n13029_));
  AOI21X1  g10593(.A0(new_n12979_), .A1(pi0626), .B0(pi1158), .Y(new_n13030_));
  OAI21X1  g10594(.A0(new_n13029_), .A1(pi0626), .B0(new_n13030_), .Y(new_n13031_));
  NAND2X1  g10595(.A(new_n13031_), .B(new_n13027_), .Y(new_n13032_));
  AOI21X1  g10596(.A0(new_n13024_), .A1(new_n12664_), .B0(new_n12672_), .Y(new_n13033_));
  OAI21X1  g10597(.A0(new_n13023_), .A1(new_n12664_), .B0(new_n13033_), .Y(new_n13034_));
  INVX1    g10598(.A(new_n12675_), .Y(new_n13035_));
  AOI21X1  g10599(.A0(new_n12979_), .A1(new_n12664_), .B0(new_n12676_), .Y(new_n13036_));
  OAI21X1  g10600(.A0(new_n13029_), .A1(new_n12664_), .B0(new_n13036_), .Y(new_n13037_));
  NAND2X1  g10601(.A(new_n13037_), .B(new_n13035_), .Y(new_n13038_));
  AOI22X1  g10602(.A0(new_n13038_), .A1(new_n13034_), .B0(new_n13032_), .B1(new_n13026_), .Y(new_n13039_));
  MX2X1    g10603(.A(new_n13039_), .B(new_n13023_), .S0(new_n11885_), .Y(new_n13040_));
  NAND2X1  g10604(.A(new_n13040_), .B(new_n12683_), .Y(new_n13041_));
  NAND2X1  g10605(.A(new_n13037_), .B(new_n13031_), .Y(new_n13042_));
  MX2X1    g10606(.A(new_n13042_), .B(new_n13029_), .S0(new_n11885_), .Y(new_n13043_));
  INVX1    g10607(.A(new_n13043_), .Y(new_n13044_));
  AOI21X1  g10608(.A0(new_n13044_), .A1(pi0628), .B0(pi1156), .Y(new_n13045_));
  MX2X1    g10609(.A(new_n13024_), .B(new_n12964_), .S0(new_n12691_), .Y(new_n13046_));
  AOI21X1  g10610(.A0(new_n12979_), .A1(new_n12683_), .B0(new_n12684_), .Y(new_n13047_));
  OAI21X1  g10611(.A0(new_n13046_), .A1(new_n12683_), .B0(new_n13047_), .Y(new_n13048_));
  NAND2X1  g10612(.A(new_n13048_), .B(new_n12689_), .Y(new_n13049_));
  AOI21X1  g10613(.A0(new_n13045_), .A1(new_n13041_), .B0(new_n13049_), .Y(new_n13050_));
  NAND2X1  g10614(.A(new_n13040_), .B(pi0628), .Y(new_n13051_));
  AOI21X1  g10615(.A0(new_n13044_), .A1(new_n12683_), .B0(new_n12684_), .Y(new_n13052_));
  AOI21X1  g10616(.A0(new_n12979_), .A1(pi0628), .B0(pi1156), .Y(new_n13053_));
  OAI21X1  g10617(.A0(new_n13046_), .A1(pi0628), .B0(new_n13053_), .Y(new_n13054_));
  NAND2X1  g10618(.A(new_n13054_), .B(pi0629), .Y(new_n13055_));
  AOI21X1  g10619(.A0(new_n13052_), .A1(new_n13051_), .B0(new_n13055_), .Y(new_n13056_));
  OAI21X1  g10620(.A0(new_n13056_), .A1(new_n13050_), .B0(pi0792), .Y(new_n13057_));
  NAND2X1  g10621(.A(new_n13040_), .B(new_n11884_), .Y(new_n13058_));
  AND2X1   g10622(.A(new_n13058_), .B(new_n13057_), .Y(new_n13059_));
  AOI21X1  g10623(.A0(new_n13058_), .A1(new_n13057_), .B0(pi0647), .Y(new_n13060_));
  MX2X1    g10624(.A(new_n13043_), .B(new_n12964_), .S0(new_n12711_), .Y(new_n13061_));
  OAI21X1  g10625(.A0(new_n13061_), .A1(new_n12705_), .B0(new_n12706_), .Y(new_n13062_));
  INVX1    g10626(.A(new_n13046_), .Y(new_n13063_));
  AND2X1   g10627(.A(new_n13054_), .B(new_n13048_), .Y(new_n13064_));
  MX2X1    g10628(.A(new_n13064_), .B(new_n13063_), .S0(new_n11884_), .Y(new_n13065_));
  INVX1    g10629(.A(new_n13065_), .Y(new_n13066_));
  AOI21X1  g10630(.A0(new_n12979_), .A1(new_n12705_), .B0(new_n12706_), .Y(new_n13067_));
  OAI21X1  g10631(.A0(new_n13066_), .A1(new_n12705_), .B0(new_n13067_), .Y(new_n13068_));
  AND2X1   g10632(.A(new_n13068_), .B(new_n12723_), .Y(new_n13069_));
  OAI21X1  g10633(.A0(new_n13062_), .A1(new_n13060_), .B0(new_n13069_), .Y(new_n13070_));
  AOI21X1  g10634(.A0(new_n13058_), .A1(new_n13057_), .B0(new_n12705_), .Y(new_n13071_));
  OAI21X1  g10635(.A0(new_n13061_), .A1(pi0647), .B0(pi1157), .Y(new_n13072_));
  AOI21X1  g10636(.A0(new_n12979_), .A1(pi0647), .B0(pi1157), .Y(new_n13073_));
  OAI21X1  g10637(.A0(new_n13066_), .A1(pi0647), .B0(new_n13073_), .Y(new_n13074_));
  AND2X1   g10638(.A(new_n13074_), .B(pi0630), .Y(new_n13075_));
  OAI21X1  g10639(.A0(new_n13072_), .A1(new_n13071_), .B0(new_n13075_), .Y(new_n13076_));
  AND2X1   g10640(.A(new_n13076_), .B(new_n13070_), .Y(new_n13077_));
  MX2X1    g10641(.A(new_n13077_), .B(new_n13059_), .S0(new_n11883_), .Y(new_n13078_));
  AND2X1   g10642(.A(new_n13074_), .B(new_n13068_), .Y(new_n13079_));
  MX2X1    g10643(.A(new_n13079_), .B(new_n13065_), .S0(new_n11883_), .Y(new_n13080_));
  AOI21X1  g10644(.A0(new_n13080_), .A1(new_n12743_), .B0(new_n12739_), .Y(new_n13081_));
  OAI21X1  g10645(.A0(new_n13078_), .A1(new_n12743_), .B0(new_n13081_), .Y(new_n13082_));
  AND2X1   g10646(.A(new_n12964_), .B(new_n12735_), .Y(new_n13083_));
  AOI21X1  g10647(.A0(new_n13061_), .A1(new_n12736_), .B0(new_n13083_), .Y(new_n13084_));
  OAI21X1  g10648(.A0(new_n12964_), .A1(pi0644), .B0(new_n12739_), .Y(new_n13085_));
  AOI21X1  g10649(.A0(new_n13084_), .A1(pi0644), .B0(new_n13085_), .Y(new_n13086_));
  NOR2X1   g10650(.A(new_n13086_), .B(new_n11882_), .Y(new_n13087_));
  AND2X1   g10651(.A(new_n13087_), .B(new_n13082_), .Y(new_n13088_));
  OR2X1    g10652(.A(new_n13059_), .B(pi0787), .Y(new_n13089_));
  OAI21X1  g10653(.A0(new_n13077_), .A1(new_n11883_), .B0(new_n13089_), .Y(new_n13090_));
  AND2X1   g10654(.A(new_n13080_), .B(pi0644), .Y(new_n13091_));
  OR2X1    g10655(.A(new_n13091_), .B(pi0715), .Y(new_n13092_));
  AOI21X1  g10656(.A0(new_n13090_), .A1(new_n12743_), .B0(new_n13092_), .Y(new_n13093_));
  OAI21X1  g10657(.A0(new_n12964_), .A1(new_n12743_), .B0(pi0715), .Y(new_n13094_));
  AOI21X1  g10658(.A0(new_n13084_), .A1(new_n12743_), .B0(new_n13094_), .Y(new_n13095_));
  OR2X1    g10659(.A(new_n13095_), .B(pi1160), .Y(new_n13096_));
  OAI21X1  g10660(.A0(new_n13096_), .A1(new_n13093_), .B0(pi0790), .Y(new_n13097_));
  AOI21X1  g10661(.A0(new_n13078_), .A1(new_n12897_), .B0(po1038), .Y(new_n13098_));
  OAI21X1  g10662(.A0(new_n13097_), .A1(new_n13088_), .B0(new_n13098_), .Y(new_n13099_));
  AOI21X1  g10663(.A0(po1038), .A1(new_n7382_), .B0(pi0832), .Y(new_n13100_));
  AOI21X1  g10664(.A0(pi1093), .A1(pi1092), .B0(pi0141), .Y(new_n13101_));
  AOI21X1  g10665(.A0(new_n12566_), .A1(pi0706), .B0(new_n13101_), .Y(new_n13102_));
  AND2X1   g10666(.A(new_n12566_), .B(pi0706), .Y(new_n13103_));
  AND2X1   g10667(.A(new_n13103_), .B(new_n12493_), .Y(new_n13104_));
  MX2X1    g10668(.A(new_n13101_), .B(pi0625), .S0(new_n13103_), .Y(new_n13105_));
  OR2X1    g10669(.A(new_n13101_), .B(pi1153), .Y(new_n13106_));
  OAI22X1  g10670(.A0(new_n13106_), .A1(new_n13104_), .B0(new_n13105_), .B1(new_n12494_), .Y(new_n13107_));
  MX2X1    g10671(.A(new_n13107_), .B(new_n13102_), .S0(new_n11889_), .Y(new_n13108_));
  OR2X1    g10672(.A(new_n13108_), .B(new_n12762_), .Y(new_n13109_));
  NOR4X1   g10673(.A(new_n13109_), .B(new_n12770_), .C(new_n12765_), .D(new_n12764_), .Y(new_n13110_));
  AOI21X1  g10674(.A0(new_n12178_), .A1(pi0749), .B0(new_n13101_), .Y(new_n13111_));
  AOI21X1  g10675(.A0(new_n12601_), .A1(new_n2739_), .B0(new_n13111_), .Y(new_n13112_));
  INVX1    g10676(.A(new_n13111_), .Y(new_n13113_));
  AOI21X1  g10677(.A0(new_n13113_), .A1(new_n12776_), .B0(new_n12591_), .Y(new_n13114_));
  AOI21X1  g10678(.A0(new_n13112_), .A1(new_n12779_), .B0(pi1155), .Y(new_n13115_));
  OAI21X1  g10679(.A0(new_n13115_), .A1(new_n13114_), .B0(pi0785), .Y(new_n13116_));
  OAI21X1  g10680(.A0(new_n13112_), .A1(pi0785), .B0(new_n13116_), .Y(new_n13117_));
  INVX1    g10681(.A(new_n13117_), .Y(new_n13118_));
  AOI21X1  g10682(.A0(new_n13118_), .A1(new_n12785_), .B0(new_n12615_), .Y(new_n13119_));
  AOI21X1  g10683(.A0(new_n13118_), .A1(new_n12788_), .B0(pi1154), .Y(new_n13120_));
  OR2X1    g10684(.A(new_n13120_), .B(new_n13119_), .Y(new_n13121_));
  MX2X1    g10685(.A(new_n13121_), .B(new_n13117_), .S0(new_n11887_), .Y(new_n13122_));
  AOI21X1  g10686(.A0(new_n13101_), .A1(new_n12637_), .B0(new_n12638_), .Y(new_n13123_));
  OAI21X1  g10687(.A0(new_n13122_), .A1(new_n12637_), .B0(new_n13123_), .Y(new_n13124_));
  AOI21X1  g10688(.A0(new_n13101_), .A1(pi0619), .B0(pi1159), .Y(new_n13125_));
  OAI21X1  g10689(.A0(new_n13122_), .A1(pi0619), .B0(new_n13125_), .Y(new_n13126_));
  AOI21X1  g10690(.A0(new_n13126_), .A1(new_n13124_), .B0(new_n11886_), .Y(new_n13127_));
  AOI21X1  g10691(.A0(new_n13122_), .A1(new_n11886_), .B0(new_n13127_), .Y(new_n13128_));
  INVX1    g10692(.A(new_n13101_), .Y(new_n13129_));
  OAI21X1  g10693(.A0(new_n13129_), .A1(pi0626), .B0(pi1158), .Y(new_n13130_));
  AOI21X1  g10694(.A0(new_n13128_), .A1(pi0626), .B0(new_n13130_), .Y(new_n13131_));
  OAI21X1  g10695(.A0(new_n13129_), .A1(new_n12664_), .B0(new_n12676_), .Y(new_n13132_));
  AOI21X1  g10696(.A0(new_n13128_), .A1(new_n12664_), .B0(new_n13132_), .Y(new_n13133_));
  NOR3X1   g10697(.A(new_n13133_), .B(new_n13131_), .C(new_n12690_), .Y(new_n13134_));
  OAI21X1  g10698(.A0(new_n13134_), .A1(new_n13110_), .B0(pi0788), .Y(new_n13135_));
  OAI21X1  g10699(.A0(new_n13102_), .A1(new_n12120_), .B0(new_n13111_), .Y(new_n13136_));
  NOR2X1   g10700(.A(new_n13102_), .B(new_n12120_), .Y(new_n13137_));
  MX2X1    g10701(.A(new_n13113_), .B(new_n12493_), .S0(new_n13137_), .Y(new_n13138_));
  NOR2X1   g10702(.A(new_n13138_), .B(new_n13106_), .Y(new_n13139_));
  OAI21X1  g10703(.A0(new_n13105_), .A1(new_n12494_), .B0(new_n12584_), .Y(new_n13140_));
  NOR3X1   g10704(.A(new_n13102_), .B(new_n12120_), .C(new_n12493_), .Y(new_n13141_));
  NOR3X1   g10705(.A(new_n13141_), .B(new_n13113_), .C(new_n12494_), .Y(new_n13142_));
  OAI21X1  g10706(.A0(new_n13106_), .A1(new_n13104_), .B0(pi0608), .Y(new_n13143_));
  OAI22X1  g10707(.A0(new_n13143_), .A1(new_n13142_), .B0(new_n13140_), .B1(new_n13139_), .Y(new_n13144_));
  MX2X1    g10708(.A(new_n13144_), .B(new_n13136_), .S0(new_n11889_), .Y(new_n13145_));
  OAI21X1  g10709(.A0(new_n13108_), .A1(new_n12590_), .B0(new_n12591_), .Y(new_n13146_));
  AOI21X1  g10710(.A0(new_n13145_), .A1(new_n12590_), .B0(new_n13146_), .Y(new_n13147_));
  OR2X1    g10711(.A(new_n13114_), .B(pi0660), .Y(new_n13148_));
  OAI21X1  g10712(.A0(new_n13108_), .A1(pi0609), .B0(pi1155), .Y(new_n13149_));
  AOI21X1  g10713(.A0(new_n13145_), .A1(pi0609), .B0(new_n13149_), .Y(new_n13150_));
  OR2X1    g10714(.A(new_n13115_), .B(new_n12596_), .Y(new_n13151_));
  OAI22X1  g10715(.A0(new_n13151_), .A1(new_n13150_), .B0(new_n13148_), .B1(new_n13147_), .Y(new_n13152_));
  MX2X1    g10716(.A(new_n13152_), .B(new_n13145_), .S0(new_n11888_), .Y(new_n13153_));
  OAI21X1  g10717(.A0(new_n13109_), .A1(new_n12614_), .B0(new_n12615_), .Y(new_n13154_));
  AOI21X1  g10718(.A0(new_n13153_), .A1(new_n12614_), .B0(new_n13154_), .Y(new_n13155_));
  OR2X1    g10719(.A(new_n13119_), .B(pi0627), .Y(new_n13156_));
  OAI21X1  g10720(.A0(new_n13109_), .A1(pi0618), .B0(pi1154), .Y(new_n13157_));
  AOI21X1  g10721(.A0(new_n13153_), .A1(pi0618), .B0(new_n13157_), .Y(new_n13158_));
  OR2X1    g10722(.A(new_n13120_), .B(new_n12622_), .Y(new_n13159_));
  OAI22X1  g10723(.A0(new_n13159_), .A1(new_n13158_), .B0(new_n13156_), .B1(new_n13155_), .Y(new_n13160_));
  MX2X1    g10724(.A(new_n13160_), .B(new_n13153_), .S0(new_n11887_), .Y(new_n13161_));
  NAND2X1  g10725(.A(new_n13161_), .B(new_n12637_), .Y(new_n13162_));
  NOR3X1   g10726(.A(new_n13108_), .B(new_n12764_), .C(new_n12762_), .Y(new_n13163_));
  AOI21X1  g10727(.A0(new_n13163_), .A1(pi0619), .B0(pi1159), .Y(new_n13164_));
  NAND2X1  g10728(.A(new_n13124_), .B(new_n12645_), .Y(new_n13165_));
  AOI21X1  g10729(.A0(new_n13164_), .A1(new_n13162_), .B0(new_n13165_), .Y(new_n13166_));
  NAND2X1  g10730(.A(new_n13161_), .B(pi0619), .Y(new_n13167_));
  AOI21X1  g10731(.A0(new_n13163_), .A1(new_n12637_), .B0(new_n12638_), .Y(new_n13168_));
  NAND2X1  g10732(.A(new_n13126_), .B(pi0648), .Y(new_n13169_));
  AOI21X1  g10733(.A0(new_n13168_), .A1(new_n13167_), .B0(new_n13169_), .Y(new_n13170_));
  NOR3X1   g10734(.A(new_n13170_), .B(new_n13166_), .C(new_n11886_), .Y(new_n13171_));
  OAI21X1  g10735(.A0(new_n13161_), .A1(pi0789), .B0(new_n12842_), .Y(new_n13172_));
  OAI21X1  g10736(.A0(new_n13172_), .A1(new_n13171_), .B0(new_n13135_), .Y(new_n13173_));
  NOR2X1   g10737(.A(new_n13133_), .B(new_n13131_), .Y(new_n13174_));
  MX2X1    g10738(.A(new_n13174_), .B(new_n13128_), .S0(new_n11885_), .Y(new_n13175_));
  INVX1    g10739(.A(new_n13175_), .Y(new_n13176_));
  OAI21X1  g10740(.A0(new_n13176_), .A1(new_n12683_), .B0(new_n12684_), .Y(new_n13177_));
  AOI21X1  g10741(.A0(new_n13173_), .A1(new_n12683_), .B0(new_n13177_), .Y(new_n13178_));
  NAND3X1  g10742(.A(new_n13163_), .B(new_n12852_), .C(new_n12850_), .Y(new_n13179_));
  AOI21X1  g10743(.A0(new_n2739_), .A1(new_n12683_), .B0(new_n13179_), .Y(new_n13180_));
  OAI21X1  g10744(.A0(new_n13180_), .A1(new_n12684_), .B0(new_n12689_), .Y(new_n13181_));
  OAI21X1  g10745(.A0(new_n13176_), .A1(pi0628), .B0(pi1156), .Y(new_n13182_));
  AOI21X1  g10746(.A0(new_n13173_), .A1(pi0628), .B0(new_n13182_), .Y(new_n13183_));
  AOI21X1  g10747(.A0(new_n2739_), .A1(pi0628), .B0(new_n13179_), .Y(new_n13184_));
  OAI21X1  g10748(.A0(new_n13184_), .A1(pi1156), .B0(pi0629), .Y(new_n13185_));
  OAI22X1  g10749(.A0(new_n13185_), .A1(new_n13183_), .B0(new_n13181_), .B1(new_n13178_), .Y(new_n13186_));
  MX2X1    g10750(.A(new_n13186_), .B(new_n13173_), .S0(new_n11884_), .Y(new_n13187_));
  MX2X1    g10751(.A(new_n13176_), .B(new_n13129_), .S0(new_n12711_), .Y(new_n13188_));
  OAI21X1  g10752(.A0(new_n13188_), .A1(new_n12705_), .B0(new_n12706_), .Y(new_n13189_));
  AOI21X1  g10753(.A0(new_n13187_), .A1(new_n12705_), .B0(new_n13189_), .Y(new_n13190_));
  NOR2X1   g10754(.A(new_n13179_), .B(new_n12870_), .Y(new_n13191_));
  OAI21X1  g10755(.A0(new_n13129_), .A1(pi0647), .B0(pi1157), .Y(new_n13192_));
  AOI21X1  g10756(.A0(new_n13191_), .A1(pi0647), .B0(new_n13192_), .Y(new_n13193_));
  OR2X1    g10757(.A(new_n13193_), .B(pi0630), .Y(new_n13194_));
  OAI21X1  g10758(.A0(new_n13188_), .A1(pi0647), .B0(pi1157), .Y(new_n13195_));
  AOI21X1  g10759(.A0(new_n13187_), .A1(pi0647), .B0(new_n13195_), .Y(new_n13196_));
  OAI21X1  g10760(.A0(new_n13129_), .A1(new_n12705_), .B0(new_n12706_), .Y(new_n13197_));
  AOI21X1  g10761(.A0(new_n13191_), .A1(new_n12705_), .B0(new_n13197_), .Y(new_n13198_));
  OR2X1    g10762(.A(new_n13198_), .B(new_n12723_), .Y(new_n13199_));
  OAI22X1  g10763(.A0(new_n13199_), .A1(new_n13196_), .B0(new_n13194_), .B1(new_n13190_), .Y(new_n13200_));
  MX2X1    g10764(.A(new_n13200_), .B(new_n13187_), .S0(new_n11883_), .Y(new_n13201_));
  OAI21X1  g10765(.A0(new_n13198_), .A1(new_n13193_), .B0(pi0787), .Y(new_n13202_));
  OAI21X1  g10766(.A0(new_n13191_), .A1(pi0787), .B0(new_n13202_), .Y(new_n13203_));
  OAI21X1  g10767(.A0(new_n13203_), .A1(pi0644), .B0(pi0715), .Y(new_n13204_));
  AOI21X1  g10768(.A0(new_n13201_), .A1(pi0644), .B0(new_n13204_), .Y(new_n13205_));
  NOR3X1   g10769(.A(new_n13101_), .B(new_n12734_), .C(new_n11883_), .Y(new_n13206_));
  AOI21X1  g10770(.A0(new_n13188_), .A1(new_n12736_), .B0(new_n13206_), .Y(new_n13207_));
  OAI21X1  g10771(.A0(new_n13129_), .A1(pi0644), .B0(new_n12739_), .Y(new_n13208_));
  AOI21X1  g10772(.A0(new_n13207_), .A1(pi0644), .B0(new_n13208_), .Y(new_n13209_));
  NOR3X1   g10773(.A(new_n13209_), .B(new_n13205_), .C(new_n11882_), .Y(new_n13210_));
  OAI21X1  g10774(.A0(new_n13203_), .A1(new_n12743_), .B0(new_n12739_), .Y(new_n13211_));
  AOI21X1  g10775(.A0(new_n13201_), .A1(new_n12743_), .B0(new_n13211_), .Y(new_n13212_));
  OAI21X1  g10776(.A0(new_n13129_), .A1(new_n12743_), .B0(pi0715), .Y(new_n13213_));
  AOI21X1  g10777(.A0(new_n13207_), .A1(new_n12743_), .B0(new_n13213_), .Y(new_n13214_));
  NOR3X1   g10778(.A(new_n13214_), .B(new_n13212_), .C(pi1160), .Y(new_n13215_));
  OAI21X1  g10779(.A0(new_n13215_), .A1(new_n13210_), .B0(pi0790), .Y(new_n13216_));
  AOI21X1  g10780(.A0(new_n13201_), .A1(new_n12897_), .B0(new_n12898_), .Y(new_n13217_));
  AOI22X1  g10781(.A0(new_n13217_), .A1(new_n13216_), .B0(new_n13100_), .B1(new_n13099_), .Y(po0298));
  NOR2X1   g10782(.A(new_n3129_), .B(new_n2972_), .Y(new_n13219_));
  INVX1    g10783(.A(pi0743), .Y(new_n13220_));
  NAND3X1  g10784(.A(new_n12450_), .B(new_n12103_), .C(pi0142), .Y(new_n13221_));
  OR2X1    g10785(.A(new_n12102_), .B(new_n5027_), .Y(new_n13222_));
  AND2X1   g10786(.A(new_n13222_), .B(new_n2972_), .Y(new_n13223_));
  OAI21X1  g10787(.A0(new_n12458_), .A1(new_n5029_), .B0(new_n13223_), .Y(new_n13224_));
  AOI21X1  g10788(.A0(new_n13224_), .A1(new_n13221_), .B0(new_n13220_), .Y(new_n13225_));
  NAND4X1  g10789(.A(new_n12461_), .B(new_n12459_), .C(pi0680), .D(new_n2972_), .Y(new_n13226_));
  NOR2X1   g10790(.A(new_n11941_), .B(new_n12255_), .Y(new_n13227_));
  MX2X1    g10791(.A(new_n12447_), .B(new_n13227_), .S0(pi0198), .Y(new_n13228_));
  OAI21X1  g10792(.A0(new_n13228_), .A1(new_n5029_), .B0(new_n11946_), .Y(new_n13229_));
  NAND3X1  g10793(.A(new_n13229_), .B(new_n13222_), .C(pi0142), .Y(new_n13230_));
  NAND3X1  g10794(.A(new_n13230_), .B(new_n13226_), .C(new_n13220_), .Y(new_n13231_));
  NAND2X1  g10795(.A(new_n13231_), .B(new_n2953_), .Y(new_n13232_));
  NAND2X1  g10796(.A(new_n12451_), .B(pi0680), .Y(new_n13233_));
  NOR3X1   g10797(.A(new_n12472_), .B(new_n12167_), .C(pi0142), .Y(new_n13234_));
  AND2X1   g10798(.A(new_n12097_), .B(pi0142), .Y(new_n13235_));
  AOI21X1  g10799(.A0(new_n13235_), .A1(new_n13233_), .B0(new_n13234_), .Y(new_n13236_));
  NOR2X1   g10800(.A(new_n13236_), .B(new_n13220_), .Y(new_n13237_));
  NAND4X1  g10801(.A(new_n12465_), .B(new_n12464_), .C(pi0680), .D(new_n2972_), .Y(new_n13238_));
  NAND2X1  g10802(.A(new_n12166_), .B(pi0603), .Y(new_n13239_));
  MX2X1    g10803(.A(new_n12447_), .B(new_n13227_), .S0(pi0210), .Y(new_n13240_));
  OAI21X1  g10804(.A0(new_n13240_), .A1(new_n5029_), .B0(new_n11943_), .Y(new_n13241_));
  NAND3X1  g10805(.A(new_n13241_), .B(new_n13239_), .C(pi0142), .Y(new_n13242_));
  NAND3X1  g10806(.A(new_n13242_), .B(new_n13238_), .C(new_n13220_), .Y(new_n13243_));
  NAND2X1  g10807(.A(new_n13243_), .B(pi0299), .Y(new_n13244_));
  OAI22X1  g10808(.A0(new_n13244_), .A1(new_n13237_), .B0(new_n13232_), .B1(new_n13225_), .Y(new_n13245_));
  AND2X1   g10809(.A(new_n12103_), .B(pi0142), .Y(new_n13246_));
  NOR3X1   g10810(.A(new_n13223_), .B(new_n13246_), .C(new_n13220_), .Y(new_n13247_));
  OR2X1    g10811(.A(pi0743), .B(new_n2972_), .Y(new_n13248_));
  OAI21X1  g10812(.A0(new_n13248_), .A1(new_n11946_), .B0(new_n2953_), .Y(new_n13249_));
  AOI21X1  g10813(.A0(new_n12166_), .A1(pi0603), .B0(pi0142), .Y(new_n13250_));
  AOI21X1  g10814(.A0(new_n12091_), .A1(pi0142), .B0(pi0743), .Y(new_n13251_));
  NOR3X1   g10815(.A(new_n13251_), .B(new_n13235_), .C(new_n13250_), .Y(new_n13252_));
  OAI22X1  g10816(.A0(new_n13252_), .A1(new_n2953_), .B0(new_n13249_), .B1(new_n13247_), .Y(new_n13253_));
  OAI21X1  g10817(.A0(new_n13253_), .A1(pi0735), .B0(new_n2959_), .Y(new_n13254_));
  AOI21X1  g10818(.A0(new_n13245_), .A1(pi0735), .B0(new_n13254_), .Y(new_n13255_));
  NAND3X1  g10819(.A(new_n12427_), .B(new_n12424_), .C(pi0142), .Y(new_n13256_));
  AOI21X1  g10820(.A0(new_n12388_), .A1(new_n2972_), .B0(new_n13220_), .Y(new_n13257_));
  AND2X1   g10821(.A(new_n13257_), .B(new_n13256_), .Y(new_n13258_));
  NOR2X1   g10822(.A(new_n12332_), .B(pi0142), .Y(new_n13259_));
  NOR3X1   g10823(.A(new_n12240_), .B(new_n12234_), .C(new_n2972_), .Y(new_n13260_));
  NOR3X1   g10824(.A(new_n13260_), .B(new_n13259_), .C(pi0743), .Y(new_n13261_));
  OR2X1    g10825(.A(new_n13261_), .B(new_n13258_), .Y(new_n13262_));
  OAI21X1  g10826(.A0(new_n11990_), .A1(new_n11975_), .B0(pi0142), .Y(new_n13263_));
  NOR2X1   g10827(.A(new_n12384_), .B(new_n13220_), .Y(new_n13264_));
  OAI21X1  g10828(.A0(new_n12151_), .A1(new_n2972_), .B0(new_n13264_), .Y(new_n13265_));
  INVX1    g10829(.A(new_n13265_), .Y(new_n13266_));
  AOI21X1  g10830(.A0(new_n13263_), .A1(new_n13220_), .B0(new_n13266_), .Y(new_n13267_));
  MX2X1    g10831(.A(new_n13267_), .B(new_n13262_), .S0(pi0735), .Y(new_n13268_));
  OAI21X1  g10832(.A0(new_n12422_), .A1(new_n2972_), .B0(pi0743), .Y(new_n13269_));
  AOI21X1  g10833(.A0(new_n12382_), .A1(new_n2972_), .B0(new_n13269_), .Y(new_n13270_));
  NAND3X1  g10834(.A(new_n12232_), .B(new_n12228_), .C(pi0142), .Y(new_n13271_));
  AOI21X1  g10835(.A0(new_n12335_), .A1(new_n2972_), .B0(pi0743), .Y(new_n13272_));
  AOI21X1  g10836(.A0(new_n13272_), .A1(new_n13271_), .B0(new_n13270_), .Y(new_n13273_));
  AOI21X1  g10837(.A0(new_n12009_), .A1(pi0142), .B0(pi0743), .Y(new_n13274_));
  NOR2X1   g10838(.A(new_n12142_), .B(new_n2972_), .Y(new_n13275_));
  NOR3X1   g10839(.A(new_n13275_), .B(new_n12375_), .C(new_n13220_), .Y(new_n13276_));
  OR2X1    g10840(.A(new_n13276_), .B(new_n13274_), .Y(new_n13277_));
  MX2X1    g10841(.A(new_n13277_), .B(new_n13273_), .S0(pi0735), .Y(new_n13278_));
  AOI21X1  g10842(.A0(new_n13278_), .A1(new_n5050_), .B0(new_n2964_), .Y(new_n13279_));
  OAI21X1  g10843(.A0(new_n13268_), .A1(new_n5050_), .B0(new_n13279_), .Y(new_n13280_));
  NOR4X1   g10844(.A(new_n12412_), .B(new_n12411_), .C(new_n12407_), .D(new_n2972_), .Y(new_n13281_));
  AOI21X1  g10845(.A0(new_n12370_), .A1(new_n12366_), .B0(pi0142), .Y(new_n13282_));
  OR2X1    g10846(.A(new_n13282_), .B(new_n13220_), .Y(new_n13283_));
  NOR4X1   g10847(.A(new_n12258_), .B(new_n12251_), .C(new_n12250_), .D(new_n2972_), .Y(new_n13284_));
  AND2X1   g10848(.A(new_n12317_), .B(new_n2972_), .Y(new_n13285_));
  OR2X1    g10849(.A(new_n13285_), .B(pi0743), .Y(new_n13286_));
  OAI22X1  g10850(.A0(new_n13286_), .A1(new_n13284_), .B0(new_n13283_), .B1(new_n13281_), .Y(new_n13287_));
  NOR2X1   g10851(.A(new_n12174_), .B(pi0142), .Y(new_n13288_));
  AOI21X1  g10852(.A0(new_n12132_), .A1(pi0142), .B0(new_n13288_), .Y(new_n13289_));
  NOR2X1   g10853(.A(new_n12055_), .B(new_n2972_), .Y(new_n13290_));
  MX2X1    g10854(.A(new_n13290_), .B(new_n13289_), .S0(pi0743), .Y(new_n13291_));
  MX2X1    g10855(.A(new_n13291_), .B(new_n13287_), .S0(pi0735), .Y(new_n13292_));
  AND2X1   g10856(.A(new_n13292_), .B(new_n5050_), .Y(new_n13293_));
  INVX1    g10857(.A(pi0735), .Y(new_n13294_));
  AOI21X1  g10858(.A0(new_n12358_), .A1(new_n12356_), .B0(pi0142), .Y(new_n13295_));
  NOR4X1   g10859(.A(new_n12405_), .B(new_n12402_), .C(new_n12265_), .D(new_n2972_), .Y(new_n13296_));
  OR2X1    g10860(.A(new_n13296_), .B(new_n13220_), .Y(new_n13297_));
  OR2X1    g10861(.A(new_n13297_), .B(new_n13295_), .Y(new_n13298_));
  NAND3X1  g10862(.A(new_n12266_), .B(new_n12261_), .C(pi0142), .Y(new_n13299_));
  AND2X1   g10863(.A(new_n13299_), .B(new_n13220_), .Y(new_n13300_));
  OAI21X1  g10864(.A0(new_n12307_), .A1(pi0142), .B0(new_n13300_), .Y(new_n13301_));
  AOI21X1  g10865(.A0(new_n13301_), .A1(new_n13298_), .B0(new_n13294_), .Y(new_n13302_));
  NOR2X1   g10866(.A(new_n12063_), .B(new_n2972_), .Y(new_n13303_));
  AOI21X1  g10867(.A0(new_n12118_), .A1(new_n12106_), .B0(new_n2972_), .Y(new_n13304_));
  NAND2X1  g10868(.A(new_n12175_), .B(pi0743), .Y(new_n13305_));
  OAI22X1  g10869(.A0(new_n13305_), .A1(new_n13304_), .B0(new_n13303_), .B1(pi0743), .Y(new_n13306_));
  INVX1    g10870(.A(new_n13306_), .Y(new_n13307_));
  AOI21X1  g10871(.A0(new_n13307_), .A1(new_n13294_), .B0(new_n13302_), .Y(new_n13308_));
  OAI21X1  g10872(.A0(new_n13308_), .A1(new_n5050_), .B0(new_n2971_), .Y(new_n13309_));
  AND2X1   g10873(.A(new_n11953_), .B(pi0142), .Y(new_n13310_));
  AOI22X1  g10874(.A0(new_n12172_), .A1(pi0743), .B0(new_n11953_), .B1(pi0142), .Y(new_n13311_));
  NAND2X1  g10875(.A(new_n13311_), .B(new_n13294_), .Y(new_n13312_));
  NAND2X1  g10876(.A(new_n12178_), .B(pi0743), .Y(new_n13313_));
  OAI22X1  g10877(.A0(new_n13313_), .A1(new_n3074_), .B0(new_n11961_), .B1(new_n2972_), .Y(new_n13314_));
  OAI22X1  g10878(.A0(new_n13314_), .A1(new_n12483_), .B0(new_n11959_), .B1(pi0120), .Y(new_n13315_));
  NAND2X1  g10879(.A(new_n13315_), .B(pi0735), .Y(new_n13316_));
  OAI21X1  g10880(.A0(new_n13316_), .A1(new_n13310_), .B0(new_n13312_), .Y(new_n13317_));
  AOI21X1  g10881(.A0(new_n13317_), .A1(new_n2970_), .B0(pi0223), .Y(new_n13318_));
  OAI21X1  g10882(.A0(new_n13309_), .A1(new_n13293_), .B0(new_n13318_), .Y(new_n13319_));
  AOI21X1  g10883(.A0(new_n13319_), .A1(new_n13280_), .B0(pi0299), .Y(new_n13320_));
  AOI21X1  g10884(.A0(new_n13278_), .A1(new_n5070_), .B0(new_n2954_), .Y(new_n13321_));
  OAI21X1  g10885(.A0(new_n13268_), .A1(new_n5070_), .B0(new_n13321_), .Y(new_n13322_));
  AND2X1   g10886(.A(new_n13292_), .B(new_n5070_), .Y(new_n13323_));
  OAI21X1  g10887(.A0(new_n13308_), .A1(new_n5070_), .B0(new_n10137_), .Y(new_n13324_));
  AOI21X1  g10888(.A0(new_n13317_), .A1(new_n10136_), .B0(pi0215), .Y(new_n13325_));
  OAI21X1  g10889(.A0(new_n13324_), .A1(new_n13323_), .B0(new_n13325_), .Y(new_n13326_));
  AOI21X1  g10890(.A0(new_n13326_), .A1(new_n13322_), .B0(new_n2953_), .Y(new_n13327_));
  NOR3X1   g10891(.A(new_n13327_), .B(new_n13320_), .C(new_n2959_), .Y(new_n13328_));
  OAI21X1  g10892(.A0(new_n13328_), .A1(new_n13255_), .B0(new_n2996_), .Y(new_n13329_));
  AOI21X1  g10893(.A0(pi0142), .A1(pi0039), .B0(new_n2996_), .Y(new_n13330_));
  AND2X1   g10894(.A(new_n12483_), .B(pi0735), .Y(new_n13331_));
  OAI21X1  g10895(.A0(new_n13331_), .A1(new_n13314_), .B0(new_n2959_), .Y(new_n13332_));
  AOI21X1  g10896(.A0(new_n13332_), .A1(new_n13330_), .B0(new_n3810_), .Y(new_n13333_));
  AOI21X1  g10897(.A0(new_n13333_), .A1(new_n13329_), .B0(new_n13219_), .Y(new_n13334_));
  MX2X1    g10898(.A(new_n13307_), .B(new_n13291_), .S0(new_n5070_), .Y(new_n13335_));
  OAI21X1  g10899(.A0(new_n13311_), .A1(new_n10137_), .B0(new_n2954_), .Y(new_n13336_));
  AOI21X1  g10900(.A0(new_n13335_), .A1(new_n10137_), .B0(new_n13336_), .Y(new_n13337_));
  OAI21X1  g10901(.A0(new_n13277_), .A1(new_n5071_), .B0(pi0215), .Y(new_n13338_));
  AOI21X1  g10902(.A0(new_n13267_), .A1(new_n5071_), .B0(new_n13338_), .Y(new_n13339_));
  OAI21X1  g10903(.A0(new_n13339_), .A1(new_n13337_), .B0(pi0299), .Y(new_n13340_));
  AND2X1   g10904(.A(new_n13291_), .B(new_n5050_), .Y(new_n13341_));
  OAI21X1  g10905(.A0(new_n13306_), .A1(new_n5050_), .B0(new_n2971_), .Y(new_n13342_));
  AOI21X1  g10906(.A0(new_n13311_), .A1(new_n2970_), .B0(pi0223), .Y(new_n13343_));
  OAI21X1  g10907(.A0(new_n13342_), .A1(new_n13341_), .B0(new_n13343_), .Y(new_n13344_));
  OR2X1    g10908(.A(new_n13267_), .B(new_n5050_), .Y(new_n13345_));
  OAI21X1  g10909(.A0(new_n13276_), .A1(new_n13274_), .B0(new_n5050_), .Y(new_n13346_));
  NAND3X1  g10910(.A(new_n13346_), .B(new_n13345_), .C(pi0223), .Y(new_n13347_));
  AND2X1   g10911(.A(new_n13347_), .B(new_n2953_), .Y(new_n13348_));
  AOI21X1  g10912(.A0(new_n13348_), .A1(new_n13344_), .B0(new_n2959_), .Y(new_n13349_));
  OAI21X1  g10913(.A0(new_n13253_), .A1(pi0039), .B0(new_n2996_), .Y(new_n13350_));
  AOI21X1  g10914(.A0(new_n13349_), .A1(new_n13340_), .B0(new_n13350_), .Y(new_n13351_));
  INVX1    g10915(.A(new_n13330_), .Y(new_n13352_));
  AOI21X1  g10916(.A0(new_n13314_), .A1(new_n2959_), .B0(new_n13352_), .Y(new_n13353_));
  OR2X1    g10917(.A(new_n13353_), .B(new_n3810_), .Y(new_n13354_));
  OAI22X1  g10918(.A0(new_n13354_), .A1(new_n13351_), .B0(new_n3129_), .B1(new_n2972_), .Y(new_n13355_));
  OAI21X1  g10919(.A0(new_n13355_), .A1(pi0625), .B0(pi1153), .Y(new_n13356_));
  AOI21X1  g10920(.A0(new_n13334_), .A1(pi0625), .B0(new_n13356_), .Y(new_n13357_));
  MX2X1    g10921(.A(new_n12531_), .B(new_n12504_), .S0(new_n2972_), .Y(new_n13358_));
  OAI21X1  g10922(.A0(new_n12055_), .A1(new_n2972_), .B0(new_n13294_), .Y(new_n13359_));
  OAI21X1  g10923(.A0(new_n13358_), .A1(new_n13294_), .B0(new_n13359_), .Y(new_n13360_));
  MX2X1    g10924(.A(new_n12535_), .B(new_n12507_), .S0(new_n2972_), .Y(new_n13361_));
  MX2X1    g10925(.A(new_n13361_), .B(new_n13303_), .S0(new_n13294_), .Y(new_n13362_));
  AOI21X1  g10926(.A0(new_n13362_), .A1(new_n5071_), .B0(new_n10136_), .Y(new_n13363_));
  OAI21X1  g10927(.A0(new_n13360_), .A1(new_n5071_), .B0(new_n13363_), .Y(new_n13364_));
  INVX1    g10928(.A(new_n11952_), .Y(new_n13365_));
  AND2X1   g10929(.A(new_n12566_), .B(pi0735), .Y(new_n13366_));
  AOI22X1  g10930(.A0(new_n13366_), .A1(new_n13365_), .B0(new_n11953_), .B1(pi0142), .Y(new_n13367_));
  AOI21X1  g10931(.A0(new_n13367_), .A1(new_n10136_), .B0(pi0215), .Y(new_n13368_));
  NOR2X1   g10932(.A(new_n12546_), .B(new_n2972_), .Y(new_n13369_));
  NAND4X1  g10933(.A(new_n12380_), .B(new_n12377_), .C(pi0680), .D(new_n2972_), .Y(new_n13370_));
  OAI21X1  g10934(.A0(new_n13370_), .A1(new_n12385_), .B0(pi0735), .Y(new_n13371_));
  NOR2X1   g10935(.A(new_n13371_), .B(new_n13369_), .Y(new_n13372_));
  AOI21X1  g10936(.A0(new_n13263_), .A1(new_n13294_), .B0(new_n13372_), .Y(new_n13373_));
  OAI21X1  g10937(.A0(new_n12084_), .A1(new_n2972_), .B0(new_n13294_), .Y(new_n13374_));
  AND2X1   g10938(.A(new_n13370_), .B(pi0735), .Y(new_n13375_));
  OAI21X1  g10939(.A0(new_n12542_), .A1(new_n2972_), .B0(new_n13375_), .Y(new_n13376_));
  NAND2X1  g10940(.A(new_n13376_), .B(new_n13374_), .Y(new_n13377_));
  AOI21X1  g10941(.A0(new_n13377_), .A1(new_n5070_), .B0(new_n2954_), .Y(new_n13378_));
  OAI21X1  g10942(.A0(new_n13373_), .A1(new_n5070_), .B0(new_n13378_), .Y(new_n13379_));
  NAND2X1  g10943(.A(new_n13379_), .B(pi0299), .Y(new_n13380_));
  AOI21X1  g10944(.A0(new_n13368_), .A1(new_n13364_), .B0(new_n13380_), .Y(new_n13381_));
  AOI21X1  g10945(.A0(new_n13362_), .A1(new_n5051_), .B0(new_n2970_), .Y(new_n13382_));
  OAI21X1  g10946(.A0(new_n13360_), .A1(new_n5051_), .B0(new_n13382_), .Y(new_n13383_));
  AOI21X1  g10947(.A0(new_n13367_), .A1(new_n2970_), .B0(pi0223), .Y(new_n13384_));
  AOI21X1  g10948(.A0(new_n13377_), .A1(new_n5050_), .B0(new_n2964_), .Y(new_n13385_));
  OAI21X1  g10949(.A0(new_n13373_), .A1(new_n5050_), .B0(new_n13385_), .Y(new_n13386_));
  NAND2X1  g10950(.A(new_n13386_), .B(new_n2953_), .Y(new_n13387_));
  AOI21X1  g10951(.A0(new_n13384_), .A1(new_n13383_), .B0(new_n13387_), .Y(new_n13388_));
  NOR3X1   g10952(.A(new_n13388_), .B(new_n13381_), .C(new_n2959_), .Y(new_n13389_));
  NOR2X1   g10953(.A(new_n12473_), .B(pi0142), .Y(new_n13390_));
  MX2X1    g10954(.A(new_n13241_), .B(new_n13229_), .S0(new_n2953_), .Y(new_n13391_));
  OAI21X1  g10955(.A0(new_n13391_), .A1(new_n2972_), .B0(pi0735), .Y(new_n13392_));
  NAND3X1  g10956(.A(new_n11948_), .B(new_n13294_), .C(pi0142), .Y(new_n13393_));
  OAI21X1  g10957(.A0(new_n13392_), .A1(new_n13390_), .B0(new_n13393_), .Y(new_n13394_));
  AND2X1   g10958(.A(new_n13394_), .B(new_n2959_), .Y(new_n13395_));
  NOR3X1   g10959(.A(new_n13395_), .B(new_n13389_), .C(pi0038), .Y(new_n13396_));
  AOI22X1  g10960(.A0(new_n13366_), .A1(new_n3630_), .B0(new_n12416_), .B1(pi0142), .Y(new_n13397_));
  OAI21X1  g10961(.A0(new_n13397_), .A1(pi0039), .B0(new_n13330_), .Y(new_n13398_));
  NAND2X1  g10962(.A(new_n13398_), .B(new_n3129_), .Y(new_n13399_));
  OAI22X1  g10963(.A0(new_n13399_), .A1(new_n13396_), .B0(new_n3129_), .B1(new_n2972_), .Y(new_n13400_));
  NOR2X1   g10964(.A(new_n13400_), .B(pi0625), .Y(new_n13401_));
  AOI21X1  g10965(.A0(new_n4995_), .A1(new_n2739_), .B0(new_n2996_), .Y(new_n13402_));
  NOR2X1   g10966(.A(new_n13402_), .B(new_n3810_), .Y(new_n13403_));
  NAND2X1  g10967(.A(new_n12068_), .B(pi0039), .Y(new_n13404_));
  AOI21X1  g10968(.A0(new_n11947_), .A1(new_n2959_), .B0(new_n2972_), .Y(new_n13405_));
  NAND2X1  g10969(.A(new_n13263_), .B(new_n5071_), .Y(new_n13406_));
  OAI21X1  g10970(.A0(new_n12084_), .A1(new_n2972_), .B0(new_n5070_), .Y(new_n13407_));
  NAND3X1  g10971(.A(new_n13407_), .B(new_n13406_), .C(pi0215), .Y(new_n13408_));
  MX2X1    g10972(.A(new_n13303_), .B(new_n13290_), .S0(new_n5070_), .Y(new_n13409_));
  OAI21X1  g10973(.A0(new_n13310_), .A1(new_n10137_), .B0(new_n2954_), .Y(new_n13410_));
  INVX1    g10974(.A(new_n13410_), .Y(new_n13411_));
  OAI21X1  g10975(.A0(new_n13409_), .A1(new_n10136_), .B0(new_n13411_), .Y(new_n13412_));
  NAND2X1  g10976(.A(pi0299), .B(pi0039), .Y(new_n13413_));
  AOI21X1  g10977(.A0(new_n13412_), .A1(new_n13408_), .B0(new_n13413_), .Y(new_n13414_));
  AOI21X1  g10978(.A0(new_n13405_), .A1(new_n13404_), .B0(new_n13414_), .Y(new_n13415_));
  OAI22X1  g10979(.A0(new_n13415_), .A1(new_n10761_), .B0(new_n13403_), .B1(new_n2972_), .Y(new_n13416_));
  OAI21X1  g10980(.A0(new_n13416_), .A1(new_n12493_), .B0(new_n12494_), .Y(new_n13417_));
  OAI21X1  g10981(.A0(new_n13417_), .A1(new_n13401_), .B0(pi0608), .Y(new_n13418_));
  OAI21X1  g10982(.A0(new_n13355_), .A1(new_n12493_), .B0(new_n12494_), .Y(new_n13419_));
  AOI21X1  g10983(.A0(new_n13334_), .A1(new_n12493_), .B0(new_n13419_), .Y(new_n13420_));
  NOR2X1   g10984(.A(new_n13400_), .B(new_n12493_), .Y(new_n13421_));
  OAI21X1  g10985(.A0(new_n13416_), .A1(pi0625), .B0(pi1153), .Y(new_n13422_));
  OAI21X1  g10986(.A0(new_n13422_), .A1(new_n13421_), .B0(new_n12584_), .Y(new_n13423_));
  OAI22X1  g10987(.A0(new_n13423_), .A1(new_n13420_), .B0(new_n13418_), .B1(new_n13357_), .Y(new_n13424_));
  MX2X1    g10988(.A(new_n13424_), .B(new_n13334_), .S0(new_n11889_), .Y(new_n13425_));
  OAI22X1  g10989(.A0(new_n13422_), .A1(new_n13421_), .B0(new_n13417_), .B1(new_n13401_), .Y(new_n13426_));
  MX2X1    g10990(.A(new_n13426_), .B(new_n13400_), .S0(new_n11889_), .Y(new_n13427_));
  OAI21X1  g10991(.A0(new_n13427_), .A1(new_n12590_), .B0(new_n12591_), .Y(new_n13428_));
  AOI21X1  g10992(.A0(new_n13425_), .A1(new_n12590_), .B0(new_n13428_), .Y(new_n13429_));
  INVX1    g10993(.A(new_n12599_), .Y(new_n13430_));
  AND2X1   g10994(.A(new_n13355_), .B(new_n12623_), .Y(new_n13431_));
  AOI22X1  g10995(.A0(new_n13431_), .A1(pi0609), .B0(new_n13416_), .B1(new_n13430_), .Y(new_n13432_));
  OAI21X1  g10996(.A0(new_n13432_), .A1(new_n12591_), .B0(new_n12596_), .Y(new_n13433_));
  OAI21X1  g10997(.A0(new_n13427_), .A1(pi0609), .B0(pi1155), .Y(new_n13434_));
  AOI21X1  g10998(.A0(new_n13425_), .A1(pi0609), .B0(new_n13434_), .Y(new_n13435_));
  INVX1    g10999(.A(new_n12608_), .Y(new_n13436_));
  AOI22X1  g11000(.A0(new_n13431_), .A1(new_n12590_), .B0(new_n13416_), .B1(new_n13436_), .Y(new_n13437_));
  OAI21X1  g11001(.A0(new_n13437_), .A1(pi1155), .B0(pi0660), .Y(new_n13438_));
  OAI22X1  g11002(.A0(new_n13438_), .A1(new_n13435_), .B0(new_n13433_), .B1(new_n13429_), .Y(new_n13439_));
  MX2X1    g11003(.A(new_n13439_), .B(new_n13425_), .S0(new_n11888_), .Y(new_n13440_));
  MX2X1    g11004(.A(new_n13427_), .B(new_n13416_), .S0(new_n12618_), .Y(new_n13441_));
  OAI21X1  g11005(.A0(new_n13441_), .A1(new_n12614_), .B0(new_n12615_), .Y(new_n13442_));
  AOI21X1  g11006(.A0(new_n13440_), .A1(new_n12614_), .B0(new_n13442_), .Y(new_n13443_));
  AOI21X1  g11007(.A0(new_n13416_), .A1(new_n12601_), .B0(new_n13431_), .Y(new_n13444_));
  MX2X1    g11008(.A(new_n13437_), .B(new_n13432_), .S0(pi1155), .Y(new_n13445_));
  MX2X1    g11009(.A(new_n13445_), .B(new_n13444_), .S0(new_n11888_), .Y(new_n13446_));
  OAI21X1  g11010(.A0(new_n13416_), .A1(pi0618), .B0(pi1154), .Y(new_n13447_));
  AOI21X1  g11011(.A0(new_n13446_), .A1(pi0618), .B0(new_n13447_), .Y(new_n13448_));
  OR2X1    g11012(.A(new_n13448_), .B(pi0627), .Y(new_n13449_));
  OAI21X1  g11013(.A0(new_n13441_), .A1(pi0618), .B0(pi1154), .Y(new_n13450_));
  AOI21X1  g11014(.A0(new_n13440_), .A1(pi0618), .B0(new_n13450_), .Y(new_n13451_));
  OAI21X1  g11015(.A0(new_n13416_), .A1(new_n12614_), .B0(new_n12615_), .Y(new_n13452_));
  AOI21X1  g11016(.A0(new_n13446_), .A1(new_n12614_), .B0(new_n13452_), .Y(new_n13453_));
  OR2X1    g11017(.A(new_n13453_), .B(new_n12622_), .Y(new_n13454_));
  OAI22X1  g11018(.A0(new_n13454_), .A1(new_n13451_), .B0(new_n13449_), .B1(new_n13443_), .Y(new_n13455_));
  MX2X1    g11019(.A(new_n13455_), .B(new_n13440_), .S0(new_n11887_), .Y(new_n13456_));
  MX2X1    g11020(.A(new_n13441_), .B(new_n13416_), .S0(new_n12641_), .Y(new_n13457_));
  OAI21X1  g11021(.A0(new_n13457_), .A1(new_n12637_), .B0(new_n12638_), .Y(new_n13458_));
  AOI21X1  g11022(.A0(new_n13456_), .A1(new_n12637_), .B0(new_n13458_), .Y(new_n13459_));
  NOR2X1   g11023(.A(new_n13453_), .B(new_n13448_), .Y(new_n13460_));
  MX2X1    g11024(.A(new_n13460_), .B(new_n13446_), .S0(new_n11887_), .Y(new_n13461_));
  OAI21X1  g11025(.A0(new_n13416_), .A1(pi0619), .B0(pi1159), .Y(new_n13462_));
  AOI21X1  g11026(.A0(new_n13461_), .A1(pi0619), .B0(new_n13462_), .Y(new_n13463_));
  OR2X1    g11027(.A(new_n13463_), .B(pi0648), .Y(new_n13464_));
  OAI21X1  g11028(.A0(new_n13457_), .A1(pi0619), .B0(pi1159), .Y(new_n13465_));
  AOI21X1  g11029(.A0(new_n13456_), .A1(pi0619), .B0(new_n13465_), .Y(new_n13466_));
  OAI21X1  g11030(.A0(new_n13416_), .A1(new_n12637_), .B0(new_n12638_), .Y(new_n13467_));
  AOI21X1  g11031(.A0(new_n13461_), .A1(new_n12637_), .B0(new_n13467_), .Y(new_n13468_));
  OR2X1    g11032(.A(new_n13468_), .B(new_n12645_), .Y(new_n13469_));
  OAI22X1  g11033(.A0(new_n13469_), .A1(new_n13466_), .B0(new_n13464_), .B1(new_n13459_), .Y(new_n13470_));
  MX2X1    g11034(.A(new_n13470_), .B(new_n13456_), .S0(new_n11886_), .Y(new_n13471_));
  MX2X1    g11035(.A(new_n13457_), .B(new_n13416_), .S0(new_n12659_), .Y(new_n13472_));
  AOI21X1  g11036(.A0(new_n13472_), .A1(pi0626), .B0(pi0641), .Y(new_n13473_));
  OAI21X1  g11037(.A0(new_n13471_), .A1(pi0626), .B0(new_n13473_), .Y(new_n13474_));
  NOR2X1   g11038(.A(new_n13468_), .B(new_n13463_), .Y(new_n13475_));
  MX2X1    g11039(.A(new_n13475_), .B(new_n13461_), .S0(new_n11886_), .Y(new_n13476_));
  OAI21X1  g11040(.A0(new_n13416_), .A1(new_n12664_), .B0(new_n12676_), .Y(new_n13477_));
  AOI21X1  g11041(.A0(new_n13476_), .A1(new_n12664_), .B0(new_n13477_), .Y(new_n13478_));
  OR2X1    g11042(.A(new_n13478_), .B(new_n12663_), .Y(new_n13479_));
  AOI21X1  g11043(.A0(new_n13472_), .A1(new_n12664_), .B0(new_n12672_), .Y(new_n13480_));
  OAI21X1  g11044(.A0(new_n13471_), .A1(new_n12664_), .B0(new_n13480_), .Y(new_n13481_));
  OAI21X1  g11045(.A0(new_n13416_), .A1(pi0626), .B0(pi1158), .Y(new_n13482_));
  AOI21X1  g11046(.A0(new_n13476_), .A1(pi0626), .B0(new_n13482_), .Y(new_n13483_));
  OR2X1    g11047(.A(new_n13483_), .B(new_n12675_), .Y(new_n13484_));
  AOI22X1  g11048(.A0(new_n13484_), .A1(new_n13481_), .B0(new_n13479_), .B1(new_n13474_), .Y(new_n13485_));
  MX2X1    g11049(.A(new_n13485_), .B(new_n13471_), .S0(new_n11885_), .Y(new_n13486_));
  OAI21X1  g11050(.A0(new_n13483_), .A1(new_n13478_), .B0(pi0788), .Y(new_n13487_));
  OAI21X1  g11051(.A0(new_n13476_), .A1(pi0788), .B0(new_n13487_), .Y(new_n13488_));
  OAI21X1  g11052(.A0(new_n13488_), .A1(new_n12683_), .B0(new_n12684_), .Y(new_n13489_));
  AOI21X1  g11053(.A0(new_n13486_), .A1(new_n12683_), .B0(new_n13489_), .Y(new_n13490_));
  MX2X1    g11054(.A(new_n13472_), .B(new_n13416_), .S0(new_n12691_), .Y(new_n13491_));
  INVX1    g11055(.A(new_n13416_), .Y(new_n13492_));
  AOI21X1  g11056(.A0(new_n13492_), .A1(new_n12683_), .B0(new_n12684_), .Y(new_n13493_));
  OAI21X1  g11057(.A0(new_n13491_), .A1(new_n12683_), .B0(new_n13493_), .Y(new_n13494_));
  NAND2X1  g11058(.A(new_n13494_), .B(new_n12689_), .Y(new_n13495_));
  OAI21X1  g11059(.A0(new_n13488_), .A1(pi0628), .B0(pi1156), .Y(new_n13496_));
  AOI21X1  g11060(.A0(new_n13486_), .A1(pi0628), .B0(new_n13496_), .Y(new_n13497_));
  AOI21X1  g11061(.A0(new_n13492_), .A1(pi0628), .B0(pi1156), .Y(new_n13498_));
  OAI21X1  g11062(.A0(new_n13491_), .A1(pi0628), .B0(new_n13498_), .Y(new_n13499_));
  NAND2X1  g11063(.A(new_n13499_), .B(pi0629), .Y(new_n13500_));
  OAI22X1  g11064(.A0(new_n13500_), .A1(new_n13497_), .B0(new_n13495_), .B1(new_n13490_), .Y(new_n13501_));
  MX2X1    g11065(.A(new_n13501_), .B(new_n13486_), .S0(new_n11884_), .Y(new_n13502_));
  MX2X1    g11066(.A(new_n13488_), .B(new_n13416_), .S0(new_n12711_), .Y(new_n13503_));
  OAI21X1  g11067(.A0(new_n13503_), .A1(new_n12705_), .B0(new_n12706_), .Y(new_n13504_));
  AOI21X1  g11068(.A0(new_n13502_), .A1(new_n12705_), .B0(new_n13504_), .Y(new_n13505_));
  AOI21X1  g11069(.A0(new_n13499_), .A1(new_n13494_), .B0(new_n11884_), .Y(new_n13506_));
  AOI21X1  g11070(.A0(new_n13491_), .A1(new_n11884_), .B0(new_n13506_), .Y(new_n13507_));
  OAI21X1  g11071(.A0(new_n13416_), .A1(pi0647), .B0(pi1157), .Y(new_n13508_));
  AOI21X1  g11072(.A0(new_n13507_), .A1(pi0647), .B0(new_n13508_), .Y(new_n13509_));
  OR2X1    g11073(.A(new_n13509_), .B(pi0630), .Y(new_n13510_));
  OAI21X1  g11074(.A0(new_n13503_), .A1(pi0647), .B0(pi1157), .Y(new_n13511_));
  AOI21X1  g11075(.A0(new_n13502_), .A1(pi0647), .B0(new_n13511_), .Y(new_n13512_));
  OAI21X1  g11076(.A0(new_n13416_), .A1(new_n12705_), .B0(new_n12706_), .Y(new_n13513_));
  AOI21X1  g11077(.A0(new_n13507_), .A1(new_n12705_), .B0(new_n13513_), .Y(new_n13514_));
  OR2X1    g11078(.A(new_n13514_), .B(new_n12723_), .Y(new_n13515_));
  OAI22X1  g11079(.A0(new_n13515_), .A1(new_n13512_), .B0(new_n13510_), .B1(new_n13505_), .Y(new_n13516_));
  MX2X1    g11080(.A(new_n13516_), .B(new_n13502_), .S0(new_n11883_), .Y(new_n13517_));
  OAI21X1  g11081(.A0(new_n13514_), .A1(new_n13509_), .B0(pi0787), .Y(new_n13518_));
  OAI21X1  g11082(.A0(new_n13507_), .A1(pi0787), .B0(new_n13518_), .Y(new_n13519_));
  OAI21X1  g11083(.A0(new_n13519_), .A1(pi0644), .B0(pi0715), .Y(new_n13520_));
  AOI21X1  g11084(.A0(new_n13517_), .A1(pi0644), .B0(new_n13520_), .Y(new_n13521_));
  AND2X1   g11085(.A(new_n13416_), .B(new_n12735_), .Y(new_n13522_));
  AOI21X1  g11086(.A0(new_n13503_), .A1(new_n12736_), .B0(new_n13522_), .Y(new_n13523_));
  OAI21X1  g11087(.A0(new_n13416_), .A1(pi0644), .B0(new_n12739_), .Y(new_n13524_));
  AOI21X1  g11088(.A0(new_n13523_), .A1(pi0644), .B0(new_n13524_), .Y(new_n13525_));
  NOR3X1   g11089(.A(new_n13525_), .B(new_n13521_), .C(new_n11882_), .Y(new_n13526_));
  OAI21X1  g11090(.A0(new_n13519_), .A1(new_n12743_), .B0(new_n12739_), .Y(new_n13527_));
  AOI21X1  g11091(.A0(new_n13517_), .A1(new_n12743_), .B0(new_n13527_), .Y(new_n13528_));
  OAI21X1  g11092(.A0(new_n13416_), .A1(new_n12743_), .B0(pi0715), .Y(new_n13529_));
  AOI21X1  g11093(.A0(new_n13523_), .A1(new_n12743_), .B0(new_n13529_), .Y(new_n13530_));
  NOR3X1   g11094(.A(new_n13530_), .B(new_n13528_), .C(pi1160), .Y(new_n13531_));
  NOR3X1   g11095(.A(new_n13531_), .B(new_n13526_), .C(new_n12897_), .Y(new_n13532_));
  OAI21X1  g11096(.A0(new_n13517_), .A1(pi0790), .B0(new_n5117_), .Y(new_n13533_));
  AOI21X1  g11097(.A0(new_n5118_), .A1(new_n2972_), .B0(pi0057), .Y(new_n13534_));
  OAI21X1  g11098(.A0(new_n13533_), .A1(new_n13532_), .B0(new_n13534_), .Y(new_n13535_));
  AOI21X1  g11099(.A0(pi0142), .A1(pi0057), .B0(pi0832), .Y(new_n13536_));
  INVX1    g11100(.A(new_n12690_), .Y(new_n13537_));
  NOR3X1   g11101(.A(new_n13313_), .B(new_n12601_), .C(new_n12590_), .Y(new_n13538_));
  NOR2X1   g11102(.A(new_n2739_), .B(new_n2972_), .Y(new_n13539_));
  NOR3X1   g11103(.A(new_n13539_), .B(new_n13538_), .C(new_n12591_), .Y(new_n13540_));
  NOR3X1   g11104(.A(new_n13313_), .B(new_n12601_), .C(pi0609), .Y(new_n13541_));
  NOR3X1   g11105(.A(new_n13541_), .B(new_n13539_), .C(pi1155), .Y(new_n13542_));
  OAI21X1  g11106(.A0(new_n13542_), .A1(new_n13540_), .B0(pi0785), .Y(new_n13543_));
  NOR2X1   g11107(.A(new_n13539_), .B(pi0785), .Y(new_n13544_));
  OAI21X1  g11108(.A0(new_n13313_), .A1(new_n12601_), .B0(new_n13544_), .Y(new_n13545_));
  AOI21X1  g11109(.A0(new_n13545_), .A1(new_n13543_), .B0(pi0781), .Y(new_n13546_));
  AND2X1   g11110(.A(new_n13545_), .B(new_n13543_), .Y(new_n13547_));
  INVX1    g11111(.A(new_n13547_), .Y(new_n13548_));
  AOI21X1  g11112(.A0(new_n13539_), .A1(new_n12614_), .B0(new_n12615_), .Y(new_n13549_));
  OAI21X1  g11113(.A0(new_n13548_), .A1(new_n12614_), .B0(new_n13549_), .Y(new_n13550_));
  AOI21X1  g11114(.A0(new_n13539_), .A1(pi0618), .B0(pi1154), .Y(new_n13551_));
  OAI21X1  g11115(.A0(new_n13548_), .A1(pi0618), .B0(new_n13551_), .Y(new_n13552_));
  AOI21X1  g11116(.A0(new_n13552_), .A1(new_n13550_), .B0(new_n11887_), .Y(new_n13553_));
  NOR2X1   g11117(.A(new_n13553_), .B(new_n13546_), .Y(new_n13554_));
  INVX1    g11118(.A(new_n13554_), .Y(new_n13555_));
  AOI21X1  g11119(.A0(new_n13539_), .A1(new_n12637_), .B0(new_n12638_), .Y(new_n13556_));
  OAI21X1  g11120(.A0(new_n13555_), .A1(new_n12637_), .B0(new_n13556_), .Y(new_n13557_));
  AOI21X1  g11121(.A0(new_n13539_), .A1(pi0619), .B0(pi1159), .Y(new_n13558_));
  OAI21X1  g11122(.A0(new_n13555_), .A1(pi0619), .B0(new_n13558_), .Y(new_n13559_));
  AND2X1   g11123(.A(new_n13559_), .B(new_n13557_), .Y(new_n13560_));
  MX2X1    g11124(.A(new_n13560_), .B(new_n13554_), .S0(new_n11886_), .Y(new_n13561_));
  INVX1    g11125(.A(new_n13539_), .Y(new_n13562_));
  OAI21X1  g11126(.A0(new_n13562_), .A1(pi0626), .B0(pi1158), .Y(new_n13563_));
  AOI21X1  g11127(.A0(new_n13561_), .A1(pi0626), .B0(new_n13563_), .Y(new_n13564_));
  OAI21X1  g11128(.A0(new_n13562_), .A1(new_n12664_), .B0(new_n12676_), .Y(new_n13565_));
  AOI21X1  g11129(.A0(new_n13561_), .A1(new_n12664_), .B0(new_n13565_), .Y(new_n13566_));
  NOR2X1   g11130(.A(new_n13566_), .B(new_n13564_), .Y(new_n13567_));
  XOR2X1   g11131(.A(pi1153), .B(pi0625), .Y(new_n13568_));
  AND2X1   g11132(.A(new_n13568_), .B(pi0778), .Y(new_n13569_));
  INVX1    g11133(.A(new_n13569_), .Y(new_n13570_));
  AOI21X1  g11134(.A0(new_n13570_), .A1(new_n13366_), .B0(new_n13539_), .Y(new_n13571_));
  NOR3X1   g11135(.A(new_n13571_), .B(new_n12641_), .C(new_n12618_), .Y(new_n13572_));
  OR2X1    g11136(.A(new_n13572_), .B(new_n13539_), .Y(new_n13573_));
  AOI21X1  g11137(.A0(new_n13562_), .A1(new_n12659_), .B0(new_n12770_), .Y(new_n13574_));
  AOI22X1  g11138(.A0(new_n13574_), .A1(new_n13573_), .B0(new_n13567_), .B1(new_n13537_), .Y(new_n13575_));
  NOR4X1   g11139(.A(new_n12210_), .B(new_n12120_), .C(new_n2740_), .D(new_n5029_), .Y(new_n13576_));
  NAND2X1  g11140(.A(new_n13576_), .B(pi0735), .Y(new_n13577_));
  NAND3X1  g11141(.A(new_n13577_), .B(new_n13562_), .C(new_n13313_), .Y(new_n13578_));
  NAND3X1  g11142(.A(new_n13576_), .B(pi0735), .C(pi0625), .Y(new_n13579_));
  AOI21X1  g11143(.A0(new_n13578_), .A1(new_n13579_), .B0(pi1153), .Y(new_n13580_));
  OAI21X1  g11144(.A0(new_n2739_), .A1(new_n2972_), .B0(pi1153), .Y(new_n13581_));
  AOI21X1  g11145(.A0(new_n13366_), .A1(pi0625), .B0(new_n13581_), .Y(new_n13582_));
  OR2X1    g11146(.A(new_n13582_), .B(pi0608), .Y(new_n13583_));
  AOI21X1  g11147(.A0(new_n13579_), .A1(new_n13313_), .B0(new_n12494_), .Y(new_n13584_));
  INVX1    g11148(.A(new_n12566_), .Y(new_n13585_));
  NOR4X1   g11149(.A(new_n13585_), .B(pi1153), .C(new_n13294_), .D(pi0625), .Y(new_n13586_));
  NOR3X1   g11150(.A(new_n13586_), .B(new_n13584_), .C(new_n13539_), .Y(new_n13587_));
  OAI22X1  g11151(.A0(new_n13587_), .A1(new_n12584_), .B0(new_n13583_), .B1(new_n13580_), .Y(new_n13588_));
  MX2X1    g11152(.A(new_n13588_), .B(new_n13578_), .S0(new_n11889_), .Y(new_n13589_));
  OAI21X1  g11153(.A0(new_n13571_), .A1(new_n12590_), .B0(new_n12591_), .Y(new_n13590_));
  AOI21X1  g11154(.A0(new_n13589_), .A1(new_n12590_), .B0(new_n13590_), .Y(new_n13591_));
  OR2X1    g11155(.A(new_n13540_), .B(pi0660), .Y(new_n13592_));
  OAI21X1  g11156(.A0(new_n13571_), .A1(pi0609), .B0(pi1155), .Y(new_n13593_));
  AOI21X1  g11157(.A0(new_n13589_), .A1(pi0609), .B0(new_n13593_), .Y(new_n13594_));
  OR2X1    g11158(.A(new_n13542_), .B(new_n12596_), .Y(new_n13595_));
  OAI22X1  g11159(.A0(new_n13595_), .A1(new_n13594_), .B0(new_n13592_), .B1(new_n13591_), .Y(new_n13596_));
  MX2X1    g11160(.A(new_n13596_), .B(new_n13589_), .S0(new_n11888_), .Y(new_n13597_));
  INVX1    g11161(.A(new_n12618_), .Y(new_n13598_));
  AND2X1   g11162(.A(new_n13570_), .B(new_n13366_), .Y(new_n13599_));
  AOI21X1  g11163(.A0(new_n13599_), .A1(new_n13598_), .B0(new_n13539_), .Y(new_n13600_));
  OAI21X1  g11164(.A0(new_n13600_), .A1(new_n12614_), .B0(new_n12615_), .Y(new_n13601_));
  AOI21X1  g11165(.A0(new_n13597_), .A1(new_n12614_), .B0(new_n13601_), .Y(new_n13602_));
  NAND2X1  g11166(.A(new_n13550_), .B(new_n12622_), .Y(new_n13603_));
  OAI21X1  g11167(.A0(new_n13600_), .A1(pi0618), .B0(pi1154), .Y(new_n13604_));
  AOI21X1  g11168(.A0(new_n13597_), .A1(pi0618), .B0(new_n13604_), .Y(new_n13605_));
  NAND2X1  g11169(.A(new_n13552_), .B(pi0627), .Y(new_n13606_));
  OAI22X1  g11170(.A0(new_n13606_), .A1(new_n13605_), .B0(new_n13603_), .B1(new_n13602_), .Y(new_n13607_));
  MX2X1    g11171(.A(new_n13607_), .B(new_n13597_), .S0(new_n11887_), .Y(new_n13608_));
  NAND2X1  g11172(.A(new_n13608_), .B(new_n12637_), .Y(new_n13609_));
  AOI21X1  g11173(.A0(new_n13573_), .A1(pi0619), .B0(pi1159), .Y(new_n13610_));
  NAND2X1  g11174(.A(new_n13557_), .B(new_n12645_), .Y(new_n13611_));
  AOI21X1  g11175(.A0(new_n13610_), .A1(new_n13609_), .B0(new_n13611_), .Y(new_n13612_));
  NAND2X1  g11176(.A(new_n13608_), .B(pi0619), .Y(new_n13613_));
  AOI21X1  g11177(.A0(new_n13573_), .A1(new_n12637_), .B0(new_n12638_), .Y(new_n13614_));
  NAND2X1  g11178(.A(new_n13559_), .B(pi0648), .Y(new_n13615_));
  AOI21X1  g11179(.A0(new_n13614_), .A1(new_n13613_), .B0(new_n13615_), .Y(new_n13616_));
  NOR3X1   g11180(.A(new_n13616_), .B(new_n13612_), .C(new_n11886_), .Y(new_n13617_));
  OAI21X1  g11181(.A0(new_n13608_), .A1(pi0789), .B0(new_n12842_), .Y(new_n13618_));
  OAI22X1  g11182(.A0(new_n13618_), .A1(new_n13617_), .B0(new_n13575_), .B1(new_n11885_), .Y(new_n13619_));
  MX2X1    g11183(.A(new_n13567_), .B(new_n13561_), .S0(new_n11885_), .Y(new_n13620_));
  INVX1    g11184(.A(new_n13620_), .Y(new_n13621_));
  AOI21X1  g11185(.A0(new_n13621_), .A1(pi0628), .B0(pi1156), .Y(new_n13622_));
  OAI21X1  g11186(.A0(new_n13619_), .A1(pi0628), .B0(new_n13622_), .Y(new_n13623_));
  OR4X1    g11187(.A(new_n12691_), .B(new_n12659_), .C(new_n12641_), .D(new_n12618_), .Y(new_n13624_));
  OR2X1    g11188(.A(new_n13624_), .B(new_n13571_), .Y(new_n13625_));
  OAI21X1  g11189(.A0(new_n13625_), .A1(new_n12683_), .B0(new_n13562_), .Y(new_n13626_));
  AOI21X1  g11190(.A0(new_n13626_), .A1(pi1156), .B0(pi0629), .Y(new_n13627_));
  AOI21X1  g11191(.A0(new_n13621_), .A1(new_n12683_), .B0(new_n12684_), .Y(new_n13628_));
  OAI21X1  g11192(.A0(new_n13619_), .A1(new_n12683_), .B0(new_n13628_), .Y(new_n13629_));
  OAI21X1  g11193(.A0(new_n13625_), .A1(pi0628), .B0(new_n13562_), .Y(new_n13630_));
  AOI21X1  g11194(.A0(new_n13630_), .A1(new_n12684_), .B0(new_n12689_), .Y(new_n13631_));
  AOI22X1  g11195(.A0(new_n13631_), .A1(new_n13629_), .B0(new_n13627_), .B1(new_n13623_), .Y(new_n13632_));
  MX2X1    g11196(.A(new_n13632_), .B(new_n13619_), .S0(new_n11884_), .Y(new_n13633_));
  MX2X1    g11197(.A(new_n13621_), .B(new_n13562_), .S0(new_n12711_), .Y(new_n13634_));
  OAI21X1  g11198(.A0(new_n13634_), .A1(new_n12705_), .B0(new_n12706_), .Y(new_n13635_));
  AOI21X1  g11199(.A0(new_n13633_), .A1(new_n12705_), .B0(new_n13635_), .Y(new_n13636_));
  AND2X1   g11200(.A(pi1156), .B(pi0628), .Y(new_n13637_));
  OAI21X1  g11201(.A0(pi1156), .A1(pi0628), .B0(pi0792), .Y(new_n13638_));
  NOR2X1   g11202(.A(new_n13638_), .B(new_n13637_), .Y(new_n13639_));
  NOR4X1   g11203(.A(new_n13639_), .B(new_n13624_), .C(new_n13571_), .D(new_n12705_), .Y(new_n13640_));
  OAI21X1  g11204(.A0(new_n2739_), .A1(new_n2972_), .B0(pi1157), .Y(new_n13641_));
  OAI21X1  g11205(.A0(new_n13641_), .A1(new_n13640_), .B0(new_n12723_), .Y(new_n13642_));
  OAI21X1  g11206(.A0(new_n13634_), .A1(pi0647), .B0(pi1157), .Y(new_n13643_));
  AOI21X1  g11207(.A0(new_n13633_), .A1(pi0647), .B0(new_n13643_), .Y(new_n13644_));
  NOR4X1   g11208(.A(new_n13639_), .B(new_n13624_), .C(new_n13571_), .D(pi0647), .Y(new_n13645_));
  OAI21X1  g11209(.A0(new_n2739_), .A1(new_n2972_), .B0(new_n12706_), .Y(new_n13646_));
  OAI21X1  g11210(.A0(new_n13646_), .A1(new_n13645_), .B0(pi0630), .Y(new_n13647_));
  OAI22X1  g11211(.A0(new_n13647_), .A1(new_n13644_), .B0(new_n13642_), .B1(new_n13636_), .Y(new_n13648_));
  MX2X1    g11212(.A(new_n13648_), .B(new_n13633_), .S0(new_n11883_), .Y(new_n13649_));
  XOR2X1   g11213(.A(pi1157), .B(new_n12705_), .Y(new_n13650_));
  NOR2X1   g11214(.A(new_n13650_), .B(new_n11883_), .Y(new_n13651_));
  OR4X1    g11215(.A(new_n13651_), .B(new_n13639_), .C(new_n13624_), .D(new_n13571_), .Y(new_n13652_));
  AND2X1   g11216(.A(new_n13652_), .B(new_n13562_), .Y(new_n13653_));
  OAI21X1  g11217(.A0(new_n13653_), .A1(pi0644), .B0(pi0715), .Y(new_n13654_));
  AOI21X1  g11218(.A0(new_n13649_), .A1(pi0644), .B0(new_n13654_), .Y(new_n13655_));
  NOR3X1   g11219(.A(new_n13539_), .B(new_n12734_), .C(new_n11883_), .Y(new_n13656_));
  AOI21X1  g11220(.A0(new_n13634_), .A1(new_n12736_), .B0(new_n13656_), .Y(new_n13657_));
  OAI21X1  g11221(.A0(new_n13562_), .A1(pi0644), .B0(new_n12739_), .Y(new_n13658_));
  AOI21X1  g11222(.A0(new_n13657_), .A1(pi0644), .B0(new_n13658_), .Y(new_n13659_));
  NOR3X1   g11223(.A(new_n13659_), .B(new_n13655_), .C(new_n11882_), .Y(new_n13660_));
  OAI21X1  g11224(.A0(new_n13653_), .A1(new_n12743_), .B0(new_n12739_), .Y(new_n13661_));
  AOI21X1  g11225(.A0(new_n13649_), .A1(new_n12743_), .B0(new_n13661_), .Y(new_n13662_));
  OAI21X1  g11226(.A0(new_n13562_), .A1(new_n12743_), .B0(pi0715), .Y(new_n13663_));
  AOI21X1  g11227(.A0(new_n13657_), .A1(new_n12743_), .B0(new_n13663_), .Y(new_n13664_));
  NOR3X1   g11228(.A(new_n13664_), .B(new_n13662_), .C(pi1160), .Y(new_n13665_));
  OAI21X1  g11229(.A0(new_n13665_), .A1(new_n13660_), .B0(pi0790), .Y(new_n13666_));
  AOI21X1  g11230(.A0(new_n13649_), .A1(new_n12897_), .B0(new_n12898_), .Y(new_n13667_));
  AOI22X1  g11231(.A0(new_n13667_), .A1(new_n13666_), .B0(new_n13536_), .B1(new_n13535_), .Y(po0299));
  AND2X1   g11232(.A(new_n12482_), .B(new_n12202_), .Y(new_n13669_));
  INVX1    g11233(.A(new_n13669_), .Y(new_n13670_));
  MX2X1    g11234(.A(new_n12454_), .B(new_n12289_), .S0(pi0039), .Y(new_n13671_));
  MX2X1    g11235(.A(new_n13671_), .B(new_n13670_), .S0(pi0038), .Y(new_n13672_));
  MX2X1    g11236(.A(new_n12467_), .B(new_n12349_), .S0(pi0039), .Y(new_n13673_));
  OR2X1    g11237(.A(new_n13673_), .B(pi0038), .Y(new_n13674_));
  INVX1    g11238(.A(pi0774), .Y(new_n13675_));
  NOR4X1   g11239(.A(new_n12482_), .B(new_n12416_), .C(pi0039), .D(new_n2996_), .Y(new_n13676_));
  NOR2X1   g11240(.A(new_n13676_), .B(new_n13675_), .Y(new_n13677_));
  OAI21X1  g11241(.A0(new_n13674_), .A1(new_n9960_), .B0(new_n13677_), .Y(new_n13678_));
  AOI21X1  g11242(.A0(new_n13672_), .A1(new_n9960_), .B0(new_n13678_), .Y(new_n13679_));
  INVX1    g11243(.A(pi0687), .Y(new_n13680_));
  OR4X1    g11244(.A(new_n12342_), .B(new_n3003_), .C(new_n2555_), .D(pi0039), .Y(new_n13681_));
  AND2X1   g11245(.A(new_n13681_), .B(pi0038), .Y(new_n13682_));
  MX2X1    g11246(.A(new_n13239_), .B(new_n13222_), .S0(new_n2953_), .Y(new_n13683_));
  OAI21X1  g11247(.A0(new_n12458_), .A1(new_n5029_), .B0(new_n2953_), .Y(new_n13684_));
  OAI21X1  g11248(.A0(new_n12472_), .A1(new_n2953_), .B0(new_n13684_), .Y(new_n13685_));
  NAND3X1  g11249(.A(new_n13685_), .B(new_n13683_), .C(new_n2959_), .Y(new_n13686_));
  OAI21X1  g11250(.A0(new_n12401_), .A1(new_n2959_), .B0(new_n13686_), .Y(new_n13687_));
  AOI21X1  g11251(.A0(new_n13687_), .A1(new_n2996_), .B0(new_n13682_), .Y(new_n13688_));
  MX2X1    g11252(.A(new_n12439_), .B(new_n12430_), .S0(new_n2953_), .Y(new_n13689_));
  AND2X1   g11253(.A(new_n13689_), .B(pi0039), .Y(new_n13690_));
  AOI21X1  g11254(.A0(new_n12453_), .A1(new_n12104_), .B0(pi0039), .Y(new_n13691_));
  NAND4X1  g11255(.A(new_n12499_), .B(new_n12171_), .C(new_n11961_), .D(new_n2959_), .Y(new_n13692_));
  MX2X1    g11256(.A(new_n13692_), .B(new_n13691_), .S0(new_n2996_), .Y(new_n13693_));
  NOR2X1   g11257(.A(new_n13693_), .B(new_n13690_), .Y(new_n13694_));
  OAI21X1  g11258(.A0(new_n13694_), .A1(pi0143), .B0(new_n13675_), .Y(new_n13695_));
  AOI21X1  g11259(.A0(new_n13688_), .A1(pi0143), .B0(new_n13695_), .Y(new_n13696_));
  OR2X1    g11260(.A(new_n13696_), .B(new_n13680_), .Y(new_n13697_));
  OR2X1    g11261(.A(new_n13697_), .B(new_n13679_), .Y(new_n13698_));
  AOI21X1  g11262(.A0(new_n12090_), .A1(new_n2996_), .B0(new_n13402_), .Y(new_n13699_));
  OAI21X1  g11263(.A0(new_n13699_), .A1(pi0143), .B0(pi0774), .Y(new_n13700_));
  NOR4X1   g11264(.A(new_n12204_), .B(new_n3015_), .C(pi0039), .D(new_n2996_), .Y(new_n13701_));
  AOI21X1  g11265(.A0(new_n12199_), .A1(new_n2996_), .B0(new_n9960_), .Y(new_n13702_));
  AOI21X1  g11266(.A0(new_n12146_), .A1(new_n6857_), .B0(new_n2996_), .Y(new_n13703_));
  AOI21X1  g11267(.A0(new_n12910_), .A1(new_n2996_), .B0(new_n13703_), .Y(new_n13704_));
  NOR2X1   g11268(.A(pi0774), .B(pi0143), .Y(new_n13705_));
  AOI21X1  g11269(.A0(new_n13705_), .A1(new_n13704_), .B0(new_n13702_), .Y(new_n13706_));
  OR2X1    g11270(.A(new_n13706_), .B(new_n13701_), .Y(new_n13707_));
  AND2X1   g11271(.A(new_n13707_), .B(new_n13700_), .Y(new_n13708_));
  AOI21X1  g11272(.A0(new_n13708_), .A1(new_n13680_), .B0(new_n3810_), .Y(new_n13709_));
  AOI22X1  g11273(.A0(new_n13709_), .A1(new_n13698_), .B0(new_n3810_), .B1(pi0143), .Y(new_n13710_));
  NAND2X1  g11274(.A(new_n13707_), .B(new_n13700_), .Y(new_n13711_));
  MX2X1    g11275(.A(new_n13711_), .B(pi0143), .S0(new_n3810_), .Y(new_n13712_));
  OAI21X1  g11276(.A0(new_n13712_), .A1(new_n12493_), .B0(new_n12494_), .Y(new_n13713_));
  AOI21X1  g11277(.A0(new_n13710_), .A1(new_n12493_), .B0(new_n13713_), .Y(new_n13714_));
  NAND3X1  g11278(.A(new_n12574_), .B(new_n13680_), .C(new_n9960_), .Y(new_n13715_));
  AOI21X1  g11279(.A0(new_n12955_), .A1(pi0143), .B0(pi0038), .Y(new_n13716_));
  OAI21X1  g11280(.A0(new_n12953_), .A1(pi0143), .B0(new_n13716_), .Y(new_n13717_));
  OR2X1    g11281(.A(new_n12202_), .B(pi0143), .Y(new_n13718_));
  AOI21X1  g11282(.A0(new_n13718_), .A1(new_n12567_), .B0(new_n13680_), .Y(new_n13719_));
  AOI21X1  g11283(.A0(new_n13719_), .A1(new_n13717_), .B0(new_n3810_), .Y(new_n13720_));
  AOI22X1  g11284(.A0(new_n13720_), .A1(new_n13715_), .B0(new_n3810_), .B1(pi0143), .Y(new_n13721_));
  OAI21X1  g11285(.A0(new_n12574_), .A1(new_n3810_), .B0(new_n9960_), .Y(new_n13722_));
  OAI21X1  g11286(.A0(new_n13722_), .A1(pi0625), .B0(pi1153), .Y(new_n13723_));
  AOI21X1  g11287(.A0(new_n13721_), .A1(pi0625), .B0(new_n13723_), .Y(new_n13724_));
  OR2X1    g11288(.A(new_n13724_), .B(pi0608), .Y(new_n13725_));
  OAI21X1  g11289(.A0(new_n13712_), .A1(pi0625), .B0(pi1153), .Y(new_n13726_));
  AOI21X1  g11290(.A0(new_n13710_), .A1(pi0625), .B0(new_n13726_), .Y(new_n13727_));
  OAI21X1  g11291(.A0(new_n13722_), .A1(new_n12493_), .B0(new_n12494_), .Y(new_n13728_));
  AOI21X1  g11292(.A0(new_n13721_), .A1(new_n12493_), .B0(new_n13728_), .Y(new_n13729_));
  OR2X1    g11293(.A(new_n13729_), .B(new_n12584_), .Y(new_n13730_));
  OAI22X1  g11294(.A0(new_n13730_), .A1(new_n13727_), .B0(new_n13725_), .B1(new_n13714_), .Y(new_n13731_));
  MX2X1    g11295(.A(new_n13731_), .B(new_n13710_), .S0(new_n11889_), .Y(new_n13732_));
  OAI21X1  g11296(.A0(new_n13729_), .A1(new_n13724_), .B0(pi0778), .Y(new_n13733_));
  OAI21X1  g11297(.A0(new_n13721_), .A1(pi0778), .B0(new_n13733_), .Y(new_n13734_));
  OAI21X1  g11298(.A0(new_n13734_), .A1(new_n12590_), .B0(new_n12591_), .Y(new_n13735_));
  AOI21X1  g11299(.A0(new_n13732_), .A1(new_n12590_), .B0(new_n13735_), .Y(new_n13736_));
  INVX1    g11300(.A(new_n13722_), .Y(new_n13737_));
  NAND2X1  g11301(.A(new_n13712_), .B(new_n12623_), .Y(new_n13738_));
  OAI22X1  g11302(.A0(new_n13738_), .A1(new_n12590_), .B0(new_n13737_), .B1(new_n12599_), .Y(new_n13739_));
  NAND2X1  g11303(.A(new_n13739_), .B(pi1155), .Y(new_n13740_));
  NAND2X1  g11304(.A(new_n13740_), .B(new_n12596_), .Y(new_n13741_));
  OAI21X1  g11305(.A0(new_n13734_), .A1(pi0609), .B0(pi1155), .Y(new_n13742_));
  AOI21X1  g11306(.A0(new_n13732_), .A1(pi0609), .B0(new_n13742_), .Y(new_n13743_));
  OAI22X1  g11307(.A0(new_n13738_), .A1(pi0609), .B0(new_n13737_), .B1(new_n12608_), .Y(new_n13744_));
  NAND2X1  g11308(.A(new_n13744_), .B(new_n12591_), .Y(new_n13745_));
  NAND2X1  g11309(.A(new_n13745_), .B(pi0660), .Y(new_n13746_));
  OAI22X1  g11310(.A0(new_n13746_), .A1(new_n13743_), .B0(new_n13741_), .B1(new_n13736_), .Y(new_n13747_));
  MX2X1    g11311(.A(new_n13747_), .B(new_n13732_), .S0(new_n11888_), .Y(new_n13748_));
  MX2X1    g11312(.A(new_n13734_), .B(new_n13722_), .S0(new_n12618_), .Y(new_n13749_));
  OAI21X1  g11313(.A0(new_n13749_), .A1(new_n12614_), .B0(new_n12615_), .Y(new_n13750_));
  AOI21X1  g11314(.A0(new_n13748_), .A1(new_n12614_), .B0(new_n13750_), .Y(new_n13751_));
  MX2X1    g11315(.A(new_n13722_), .B(new_n13712_), .S0(new_n12623_), .Y(new_n13752_));
  AOI21X1  g11316(.A0(new_n13745_), .A1(new_n13740_), .B0(new_n11888_), .Y(new_n13753_));
  AOI21X1  g11317(.A0(new_n13752_), .A1(new_n11888_), .B0(new_n13753_), .Y(new_n13754_));
  OAI21X1  g11318(.A0(new_n13722_), .A1(pi0618), .B0(pi1154), .Y(new_n13755_));
  AOI21X1  g11319(.A0(new_n13754_), .A1(pi0618), .B0(new_n13755_), .Y(new_n13756_));
  OR2X1    g11320(.A(new_n13756_), .B(pi0627), .Y(new_n13757_));
  OAI21X1  g11321(.A0(new_n13749_), .A1(pi0618), .B0(pi1154), .Y(new_n13758_));
  AOI21X1  g11322(.A0(new_n13748_), .A1(pi0618), .B0(new_n13758_), .Y(new_n13759_));
  OAI21X1  g11323(.A0(new_n13722_), .A1(new_n12614_), .B0(new_n12615_), .Y(new_n13760_));
  AOI21X1  g11324(.A0(new_n13754_), .A1(new_n12614_), .B0(new_n13760_), .Y(new_n13761_));
  OR2X1    g11325(.A(new_n13761_), .B(new_n12622_), .Y(new_n13762_));
  OAI22X1  g11326(.A0(new_n13762_), .A1(new_n13759_), .B0(new_n13757_), .B1(new_n13751_), .Y(new_n13763_));
  MX2X1    g11327(.A(new_n13763_), .B(new_n13748_), .S0(new_n11887_), .Y(new_n13764_));
  MX2X1    g11328(.A(new_n13749_), .B(new_n13722_), .S0(new_n12641_), .Y(new_n13765_));
  OAI21X1  g11329(.A0(new_n13765_), .A1(new_n12637_), .B0(new_n12638_), .Y(new_n13766_));
  AOI21X1  g11330(.A0(new_n13764_), .A1(new_n12637_), .B0(new_n13766_), .Y(new_n13767_));
  NOR2X1   g11331(.A(new_n13761_), .B(new_n13756_), .Y(new_n13768_));
  MX2X1    g11332(.A(new_n13768_), .B(new_n13754_), .S0(new_n11887_), .Y(new_n13769_));
  OAI21X1  g11333(.A0(new_n13722_), .A1(pi0619), .B0(pi1159), .Y(new_n13770_));
  AOI21X1  g11334(.A0(new_n13769_), .A1(pi0619), .B0(new_n13770_), .Y(new_n13771_));
  OR2X1    g11335(.A(new_n13771_), .B(pi0648), .Y(new_n13772_));
  OAI21X1  g11336(.A0(new_n13765_), .A1(pi0619), .B0(pi1159), .Y(new_n13773_));
  AOI21X1  g11337(.A0(new_n13764_), .A1(pi0619), .B0(new_n13773_), .Y(new_n13774_));
  OAI21X1  g11338(.A0(new_n13722_), .A1(new_n12637_), .B0(new_n12638_), .Y(new_n13775_));
  AOI21X1  g11339(.A0(new_n13769_), .A1(new_n12637_), .B0(new_n13775_), .Y(new_n13776_));
  OR2X1    g11340(.A(new_n13776_), .B(new_n12645_), .Y(new_n13777_));
  OAI22X1  g11341(.A0(new_n13777_), .A1(new_n13774_), .B0(new_n13772_), .B1(new_n13767_), .Y(new_n13778_));
  MX2X1    g11342(.A(new_n13778_), .B(new_n13764_), .S0(new_n11886_), .Y(new_n13779_));
  MX2X1    g11343(.A(new_n13765_), .B(new_n13722_), .S0(new_n12659_), .Y(new_n13780_));
  AOI21X1  g11344(.A0(new_n13780_), .A1(pi0626), .B0(pi0641), .Y(new_n13781_));
  OAI21X1  g11345(.A0(new_n13779_), .A1(pi0626), .B0(new_n13781_), .Y(new_n13782_));
  OR2X1    g11346(.A(new_n13769_), .B(pi0789), .Y(new_n13783_));
  OAI21X1  g11347(.A0(new_n13776_), .A1(new_n13771_), .B0(pi0789), .Y(new_n13784_));
  NAND3X1  g11348(.A(new_n13784_), .B(new_n13783_), .C(new_n12664_), .Y(new_n13785_));
  AOI21X1  g11349(.A0(new_n13737_), .A1(pi0626), .B0(pi1158), .Y(new_n13786_));
  AND2X1   g11350(.A(new_n13786_), .B(new_n13785_), .Y(new_n13787_));
  OR2X1    g11351(.A(new_n13787_), .B(new_n12663_), .Y(new_n13788_));
  AOI21X1  g11352(.A0(new_n13780_), .A1(new_n12664_), .B0(new_n12672_), .Y(new_n13789_));
  OAI21X1  g11353(.A0(new_n13779_), .A1(new_n12664_), .B0(new_n13789_), .Y(new_n13790_));
  NAND3X1  g11354(.A(new_n13784_), .B(new_n13783_), .C(pi0626), .Y(new_n13791_));
  AOI21X1  g11355(.A0(new_n13737_), .A1(new_n12664_), .B0(new_n12676_), .Y(new_n13792_));
  AND2X1   g11356(.A(new_n13792_), .B(new_n13791_), .Y(new_n13793_));
  OR2X1    g11357(.A(new_n13793_), .B(new_n12675_), .Y(new_n13794_));
  AOI22X1  g11358(.A0(new_n13794_), .A1(new_n13790_), .B0(new_n13788_), .B1(new_n13782_), .Y(new_n13795_));
  MX2X1    g11359(.A(new_n13795_), .B(new_n13779_), .S0(new_n11885_), .Y(new_n13796_));
  AND2X1   g11360(.A(new_n13784_), .B(new_n13783_), .Y(new_n13797_));
  OAI21X1  g11361(.A0(new_n13793_), .A1(new_n13787_), .B0(pi0788), .Y(new_n13798_));
  OAI21X1  g11362(.A0(new_n13797_), .A1(pi0788), .B0(new_n13798_), .Y(new_n13799_));
  OAI21X1  g11363(.A0(new_n13799_), .A1(new_n12683_), .B0(new_n12684_), .Y(new_n13800_));
  AOI21X1  g11364(.A0(new_n13796_), .A1(new_n12683_), .B0(new_n13800_), .Y(new_n13801_));
  MX2X1    g11365(.A(new_n13780_), .B(new_n13722_), .S0(new_n12691_), .Y(new_n13802_));
  AOI21X1  g11366(.A0(new_n13737_), .A1(new_n12683_), .B0(new_n12684_), .Y(new_n13803_));
  OAI21X1  g11367(.A0(new_n13802_), .A1(new_n12683_), .B0(new_n13803_), .Y(new_n13804_));
  AND2X1   g11368(.A(new_n13804_), .B(new_n12689_), .Y(new_n13805_));
  INVX1    g11369(.A(new_n13805_), .Y(new_n13806_));
  OAI21X1  g11370(.A0(new_n13799_), .A1(pi0628), .B0(pi1156), .Y(new_n13807_));
  AOI21X1  g11371(.A0(new_n13796_), .A1(pi0628), .B0(new_n13807_), .Y(new_n13808_));
  AOI21X1  g11372(.A0(new_n13737_), .A1(pi0628), .B0(pi1156), .Y(new_n13809_));
  OAI21X1  g11373(.A0(new_n13802_), .A1(pi0628), .B0(new_n13809_), .Y(new_n13810_));
  AND2X1   g11374(.A(new_n13810_), .B(pi0629), .Y(new_n13811_));
  INVX1    g11375(.A(new_n13811_), .Y(new_n13812_));
  OAI22X1  g11376(.A0(new_n13812_), .A1(new_n13808_), .B0(new_n13806_), .B1(new_n13801_), .Y(new_n13813_));
  MX2X1    g11377(.A(new_n13813_), .B(new_n13796_), .S0(new_n11884_), .Y(new_n13814_));
  MX2X1    g11378(.A(new_n13799_), .B(new_n13722_), .S0(new_n12711_), .Y(new_n13815_));
  OAI21X1  g11379(.A0(new_n13815_), .A1(new_n12705_), .B0(new_n12706_), .Y(new_n13816_));
  AOI21X1  g11380(.A0(new_n13814_), .A1(new_n12705_), .B0(new_n13816_), .Y(new_n13817_));
  AOI21X1  g11381(.A0(new_n13810_), .A1(new_n13804_), .B0(new_n11884_), .Y(new_n13818_));
  AOI21X1  g11382(.A0(new_n13802_), .A1(new_n11884_), .B0(new_n13818_), .Y(new_n13819_));
  OAI21X1  g11383(.A0(new_n13722_), .A1(pi0647), .B0(pi1157), .Y(new_n13820_));
  AOI21X1  g11384(.A0(new_n13819_), .A1(pi0647), .B0(new_n13820_), .Y(new_n13821_));
  NOR2X1   g11385(.A(new_n13821_), .B(pi0630), .Y(new_n13822_));
  INVX1    g11386(.A(new_n13822_), .Y(new_n13823_));
  OAI21X1  g11387(.A0(new_n13815_), .A1(pi0647), .B0(pi1157), .Y(new_n13824_));
  AOI21X1  g11388(.A0(new_n13814_), .A1(pi0647), .B0(new_n13824_), .Y(new_n13825_));
  OAI21X1  g11389(.A0(new_n13722_), .A1(new_n12705_), .B0(new_n12706_), .Y(new_n13826_));
  AOI21X1  g11390(.A0(new_n13819_), .A1(new_n12705_), .B0(new_n13826_), .Y(new_n13827_));
  NOR2X1   g11391(.A(new_n13827_), .B(new_n12723_), .Y(new_n13828_));
  INVX1    g11392(.A(new_n13828_), .Y(new_n13829_));
  OAI22X1  g11393(.A0(new_n13829_), .A1(new_n13825_), .B0(new_n13823_), .B1(new_n13817_), .Y(new_n13830_));
  MX2X1    g11394(.A(new_n13830_), .B(new_n13814_), .S0(new_n11883_), .Y(new_n13831_));
  OAI21X1  g11395(.A0(new_n13827_), .A1(new_n13821_), .B0(pi0787), .Y(new_n13832_));
  OAI21X1  g11396(.A0(new_n13819_), .A1(pi0787), .B0(new_n13832_), .Y(new_n13833_));
  OAI21X1  g11397(.A0(new_n13833_), .A1(pi0644), .B0(pi0715), .Y(new_n13834_));
  AOI21X1  g11398(.A0(new_n13831_), .A1(pi0644), .B0(new_n13834_), .Y(new_n13835_));
  AND2X1   g11399(.A(new_n13722_), .B(new_n12735_), .Y(new_n13836_));
  AOI21X1  g11400(.A0(new_n13815_), .A1(new_n12736_), .B0(new_n13836_), .Y(new_n13837_));
  OAI21X1  g11401(.A0(new_n13722_), .A1(pi0644), .B0(new_n12739_), .Y(new_n13838_));
  AOI21X1  g11402(.A0(new_n13837_), .A1(pi0644), .B0(new_n13838_), .Y(new_n13839_));
  NOR3X1   g11403(.A(new_n13839_), .B(new_n13835_), .C(new_n11882_), .Y(new_n13840_));
  OAI21X1  g11404(.A0(new_n13833_), .A1(new_n12743_), .B0(new_n12739_), .Y(new_n13841_));
  AOI21X1  g11405(.A0(new_n13831_), .A1(new_n12743_), .B0(new_n13841_), .Y(new_n13842_));
  OAI21X1  g11406(.A0(new_n13722_), .A1(new_n12743_), .B0(pi0715), .Y(new_n13843_));
  AOI21X1  g11407(.A0(new_n13837_), .A1(new_n12743_), .B0(new_n13843_), .Y(new_n13844_));
  OR2X1    g11408(.A(new_n13844_), .B(pi1160), .Y(new_n13845_));
  OAI21X1  g11409(.A0(new_n13845_), .A1(new_n13842_), .B0(pi0790), .Y(new_n13846_));
  OR2X1    g11410(.A(new_n13831_), .B(pi0790), .Y(new_n13847_));
  AND2X1   g11411(.A(new_n13847_), .B(new_n6520_), .Y(new_n13848_));
  OAI21X1  g11412(.A0(new_n13846_), .A1(new_n13840_), .B0(new_n13848_), .Y(new_n13849_));
  AOI21X1  g11413(.A0(po1038), .A1(new_n9960_), .B0(pi0832), .Y(new_n13850_));
  AOI21X1  g11414(.A0(pi1093), .A1(pi1092), .B0(pi0143), .Y(new_n13851_));
  AOI21X1  g11415(.A0(new_n12566_), .A1(pi0687), .B0(new_n13851_), .Y(new_n13852_));
  AND2X1   g11416(.A(new_n12566_), .B(pi0687), .Y(new_n13853_));
  AND2X1   g11417(.A(new_n13853_), .B(new_n12493_), .Y(new_n13854_));
  MX2X1    g11418(.A(new_n13851_), .B(pi0625), .S0(new_n13853_), .Y(new_n13855_));
  OR2X1    g11419(.A(new_n13851_), .B(pi1153), .Y(new_n13856_));
  OAI22X1  g11420(.A0(new_n13856_), .A1(new_n13854_), .B0(new_n13855_), .B1(new_n12494_), .Y(new_n13857_));
  MX2X1    g11421(.A(new_n13857_), .B(new_n13852_), .S0(new_n11889_), .Y(new_n13858_));
  OR2X1    g11422(.A(new_n13858_), .B(new_n12762_), .Y(new_n13859_));
  NOR4X1   g11423(.A(new_n13859_), .B(new_n12770_), .C(new_n12765_), .D(new_n12764_), .Y(new_n13860_));
  AOI21X1  g11424(.A0(new_n12178_), .A1(new_n13675_), .B0(new_n13851_), .Y(new_n13861_));
  AOI21X1  g11425(.A0(new_n12601_), .A1(new_n2739_), .B0(new_n13861_), .Y(new_n13862_));
  INVX1    g11426(.A(new_n13861_), .Y(new_n13863_));
  AOI21X1  g11427(.A0(new_n13863_), .A1(new_n12776_), .B0(new_n12591_), .Y(new_n13864_));
  AOI21X1  g11428(.A0(new_n13862_), .A1(new_n12779_), .B0(pi1155), .Y(new_n13865_));
  OAI21X1  g11429(.A0(new_n13865_), .A1(new_n13864_), .B0(pi0785), .Y(new_n13866_));
  OAI21X1  g11430(.A0(new_n13862_), .A1(pi0785), .B0(new_n13866_), .Y(new_n13867_));
  INVX1    g11431(.A(new_n13867_), .Y(new_n13868_));
  AOI21X1  g11432(.A0(new_n13868_), .A1(new_n12785_), .B0(new_n12615_), .Y(new_n13869_));
  AOI21X1  g11433(.A0(new_n13868_), .A1(new_n12788_), .B0(pi1154), .Y(new_n13870_));
  OR2X1    g11434(.A(new_n13870_), .B(new_n13869_), .Y(new_n13871_));
  MX2X1    g11435(.A(new_n13871_), .B(new_n13867_), .S0(new_n11887_), .Y(new_n13872_));
  AOI21X1  g11436(.A0(new_n13851_), .A1(new_n12637_), .B0(new_n12638_), .Y(new_n13873_));
  OAI21X1  g11437(.A0(new_n13872_), .A1(new_n12637_), .B0(new_n13873_), .Y(new_n13874_));
  AOI21X1  g11438(.A0(new_n13851_), .A1(pi0619), .B0(pi1159), .Y(new_n13875_));
  OAI21X1  g11439(.A0(new_n13872_), .A1(pi0619), .B0(new_n13875_), .Y(new_n13876_));
  AOI21X1  g11440(.A0(new_n13876_), .A1(new_n13874_), .B0(new_n11886_), .Y(new_n13877_));
  AOI21X1  g11441(.A0(new_n13872_), .A1(new_n11886_), .B0(new_n13877_), .Y(new_n13878_));
  INVX1    g11442(.A(new_n13851_), .Y(new_n13879_));
  OAI21X1  g11443(.A0(new_n13879_), .A1(pi0626), .B0(pi1158), .Y(new_n13880_));
  AOI21X1  g11444(.A0(new_n13878_), .A1(pi0626), .B0(new_n13880_), .Y(new_n13881_));
  OAI21X1  g11445(.A0(new_n13879_), .A1(new_n12664_), .B0(new_n12676_), .Y(new_n13882_));
  AOI21X1  g11446(.A0(new_n13878_), .A1(new_n12664_), .B0(new_n13882_), .Y(new_n13883_));
  NOR3X1   g11447(.A(new_n13883_), .B(new_n13881_), .C(new_n12690_), .Y(new_n13884_));
  OAI21X1  g11448(.A0(new_n13884_), .A1(new_n13860_), .B0(pi0788), .Y(new_n13885_));
  OAI21X1  g11449(.A0(new_n13852_), .A1(new_n12120_), .B0(new_n13861_), .Y(new_n13886_));
  NOR2X1   g11450(.A(new_n13852_), .B(new_n12120_), .Y(new_n13887_));
  MX2X1    g11451(.A(new_n13863_), .B(new_n12493_), .S0(new_n13887_), .Y(new_n13888_));
  NOR2X1   g11452(.A(new_n13888_), .B(new_n13856_), .Y(new_n13889_));
  OAI21X1  g11453(.A0(new_n13855_), .A1(new_n12494_), .B0(new_n12584_), .Y(new_n13890_));
  NOR3X1   g11454(.A(new_n13852_), .B(new_n12120_), .C(new_n12493_), .Y(new_n13891_));
  NOR3X1   g11455(.A(new_n13891_), .B(new_n13863_), .C(new_n12494_), .Y(new_n13892_));
  OAI21X1  g11456(.A0(new_n13856_), .A1(new_n13854_), .B0(pi0608), .Y(new_n13893_));
  OAI22X1  g11457(.A0(new_n13893_), .A1(new_n13892_), .B0(new_n13890_), .B1(new_n13889_), .Y(new_n13894_));
  MX2X1    g11458(.A(new_n13894_), .B(new_n13886_), .S0(new_n11889_), .Y(new_n13895_));
  OAI21X1  g11459(.A0(new_n13858_), .A1(new_n12590_), .B0(new_n12591_), .Y(new_n13896_));
  AOI21X1  g11460(.A0(new_n13895_), .A1(new_n12590_), .B0(new_n13896_), .Y(new_n13897_));
  OR2X1    g11461(.A(new_n13864_), .B(pi0660), .Y(new_n13898_));
  OAI21X1  g11462(.A0(new_n13858_), .A1(pi0609), .B0(pi1155), .Y(new_n13899_));
  AOI21X1  g11463(.A0(new_n13895_), .A1(pi0609), .B0(new_n13899_), .Y(new_n13900_));
  OR2X1    g11464(.A(new_n13865_), .B(new_n12596_), .Y(new_n13901_));
  OAI22X1  g11465(.A0(new_n13901_), .A1(new_n13900_), .B0(new_n13898_), .B1(new_n13897_), .Y(new_n13902_));
  MX2X1    g11466(.A(new_n13902_), .B(new_n13895_), .S0(new_n11888_), .Y(new_n13903_));
  OAI21X1  g11467(.A0(new_n13859_), .A1(new_n12614_), .B0(new_n12615_), .Y(new_n13904_));
  AOI21X1  g11468(.A0(new_n13903_), .A1(new_n12614_), .B0(new_n13904_), .Y(new_n13905_));
  OR2X1    g11469(.A(new_n13869_), .B(pi0627), .Y(new_n13906_));
  OAI21X1  g11470(.A0(new_n13859_), .A1(pi0618), .B0(pi1154), .Y(new_n13907_));
  AOI21X1  g11471(.A0(new_n13903_), .A1(pi0618), .B0(new_n13907_), .Y(new_n13908_));
  OR2X1    g11472(.A(new_n13870_), .B(new_n12622_), .Y(new_n13909_));
  OAI22X1  g11473(.A0(new_n13909_), .A1(new_n13908_), .B0(new_n13906_), .B1(new_n13905_), .Y(new_n13910_));
  MX2X1    g11474(.A(new_n13910_), .B(new_n13903_), .S0(new_n11887_), .Y(new_n13911_));
  NAND2X1  g11475(.A(new_n13911_), .B(new_n12637_), .Y(new_n13912_));
  NOR3X1   g11476(.A(new_n13858_), .B(new_n12764_), .C(new_n12762_), .Y(new_n13913_));
  AOI21X1  g11477(.A0(new_n13913_), .A1(pi0619), .B0(pi1159), .Y(new_n13914_));
  NAND2X1  g11478(.A(new_n13874_), .B(new_n12645_), .Y(new_n13915_));
  AOI21X1  g11479(.A0(new_n13914_), .A1(new_n13912_), .B0(new_n13915_), .Y(new_n13916_));
  NAND2X1  g11480(.A(new_n13911_), .B(pi0619), .Y(new_n13917_));
  AOI21X1  g11481(.A0(new_n13913_), .A1(new_n12637_), .B0(new_n12638_), .Y(new_n13918_));
  NAND2X1  g11482(.A(new_n13876_), .B(pi0648), .Y(new_n13919_));
  AOI21X1  g11483(.A0(new_n13918_), .A1(new_n13917_), .B0(new_n13919_), .Y(new_n13920_));
  NOR3X1   g11484(.A(new_n13920_), .B(new_n13916_), .C(new_n11886_), .Y(new_n13921_));
  OAI21X1  g11485(.A0(new_n13911_), .A1(pi0789), .B0(new_n12842_), .Y(new_n13922_));
  OAI21X1  g11486(.A0(new_n13922_), .A1(new_n13921_), .B0(new_n13885_), .Y(new_n13923_));
  NOR2X1   g11487(.A(new_n13883_), .B(new_n13881_), .Y(new_n13924_));
  MX2X1    g11488(.A(new_n13924_), .B(new_n13878_), .S0(new_n11885_), .Y(new_n13925_));
  INVX1    g11489(.A(new_n13925_), .Y(new_n13926_));
  OAI21X1  g11490(.A0(new_n13926_), .A1(new_n12683_), .B0(new_n12684_), .Y(new_n13927_));
  AOI21X1  g11491(.A0(new_n13923_), .A1(new_n12683_), .B0(new_n13927_), .Y(new_n13928_));
  NAND3X1  g11492(.A(new_n13913_), .B(new_n12852_), .C(new_n12850_), .Y(new_n13929_));
  AOI21X1  g11493(.A0(new_n2739_), .A1(new_n12683_), .B0(new_n13929_), .Y(new_n13930_));
  OAI21X1  g11494(.A0(new_n13930_), .A1(new_n12684_), .B0(new_n12689_), .Y(new_n13931_));
  OAI21X1  g11495(.A0(new_n13926_), .A1(pi0628), .B0(pi1156), .Y(new_n13932_));
  AOI21X1  g11496(.A0(new_n13923_), .A1(pi0628), .B0(new_n13932_), .Y(new_n13933_));
  AOI21X1  g11497(.A0(new_n2739_), .A1(pi0628), .B0(new_n13929_), .Y(new_n13934_));
  OAI21X1  g11498(.A0(new_n13934_), .A1(pi1156), .B0(pi0629), .Y(new_n13935_));
  OAI22X1  g11499(.A0(new_n13935_), .A1(new_n13933_), .B0(new_n13931_), .B1(new_n13928_), .Y(new_n13936_));
  MX2X1    g11500(.A(new_n13936_), .B(new_n13923_), .S0(new_n11884_), .Y(new_n13937_));
  MX2X1    g11501(.A(new_n13926_), .B(new_n13879_), .S0(new_n12711_), .Y(new_n13938_));
  OAI21X1  g11502(.A0(new_n13938_), .A1(new_n12705_), .B0(new_n12706_), .Y(new_n13939_));
  AOI21X1  g11503(.A0(new_n13937_), .A1(new_n12705_), .B0(new_n13939_), .Y(new_n13940_));
  NOR2X1   g11504(.A(new_n13929_), .B(new_n12870_), .Y(new_n13941_));
  OAI21X1  g11505(.A0(new_n13879_), .A1(pi0647), .B0(pi1157), .Y(new_n13942_));
  AOI21X1  g11506(.A0(new_n13941_), .A1(pi0647), .B0(new_n13942_), .Y(new_n13943_));
  OR2X1    g11507(.A(new_n13943_), .B(pi0630), .Y(new_n13944_));
  OAI21X1  g11508(.A0(new_n13938_), .A1(pi0647), .B0(pi1157), .Y(new_n13945_));
  AOI21X1  g11509(.A0(new_n13937_), .A1(pi0647), .B0(new_n13945_), .Y(new_n13946_));
  OAI21X1  g11510(.A0(new_n13879_), .A1(new_n12705_), .B0(new_n12706_), .Y(new_n13947_));
  AOI21X1  g11511(.A0(new_n13941_), .A1(new_n12705_), .B0(new_n13947_), .Y(new_n13948_));
  OR2X1    g11512(.A(new_n13948_), .B(new_n12723_), .Y(new_n13949_));
  OAI22X1  g11513(.A0(new_n13949_), .A1(new_n13946_), .B0(new_n13944_), .B1(new_n13940_), .Y(new_n13950_));
  MX2X1    g11514(.A(new_n13950_), .B(new_n13937_), .S0(new_n11883_), .Y(new_n13951_));
  OAI21X1  g11515(.A0(new_n13948_), .A1(new_n13943_), .B0(pi0787), .Y(new_n13952_));
  OAI21X1  g11516(.A0(new_n13941_), .A1(pi0787), .B0(new_n13952_), .Y(new_n13953_));
  OAI21X1  g11517(.A0(new_n13953_), .A1(pi0644), .B0(pi0715), .Y(new_n13954_));
  AOI21X1  g11518(.A0(new_n13951_), .A1(pi0644), .B0(new_n13954_), .Y(new_n13955_));
  NOR3X1   g11519(.A(new_n13851_), .B(new_n12734_), .C(new_n11883_), .Y(new_n13956_));
  AOI21X1  g11520(.A0(new_n13938_), .A1(new_n12736_), .B0(new_n13956_), .Y(new_n13957_));
  OAI21X1  g11521(.A0(new_n13879_), .A1(pi0644), .B0(new_n12739_), .Y(new_n13958_));
  AOI21X1  g11522(.A0(new_n13957_), .A1(pi0644), .B0(new_n13958_), .Y(new_n13959_));
  NOR3X1   g11523(.A(new_n13959_), .B(new_n13955_), .C(new_n11882_), .Y(new_n13960_));
  OAI21X1  g11524(.A0(new_n13953_), .A1(new_n12743_), .B0(new_n12739_), .Y(new_n13961_));
  AOI21X1  g11525(.A0(new_n13951_), .A1(new_n12743_), .B0(new_n13961_), .Y(new_n13962_));
  OAI21X1  g11526(.A0(new_n13879_), .A1(new_n12743_), .B0(pi0715), .Y(new_n13963_));
  AOI21X1  g11527(.A0(new_n13957_), .A1(new_n12743_), .B0(new_n13963_), .Y(new_n13964_));
  NOR3X1   g11528(.A(new_n13964_), .B(new_n13962_), .C(pi1160), .Y(new_n13965_));
  OAI21X1  g11529(.A0(new_n13965_), .A1(new_n13960_), .B0(pi0790), .Y(new_n13966_));
  AOI21X1  g11530(.A0(new_n13951_), .A1(new_n12897_), .B0(new_n12898_), .Y(new_n13967_));
  AOI22X1  g11531(.A0(new_n13967_), .A1(new_n13966_), .B0(new_n13850_), .B1(new_n13849_), .Y(po0300));
  INVX1    g11532(.A(pi0736), .Y(new_n13969_));
  AOI21X1  g11533(.A0(new_n12088_), .A1(new_n12068_), .B0(pi0758), .Y(new_n13970_));
  AND2X1   g11534(.A(new_n12161_), .B(pi0758), .Y(new_n13971_));
  OAI21X1  g11535(.A0(new_n13971_), .A1(new_n13970_), .B0(pi0039), .Y(new_n13972_));
  INVX1    g11536(.A(pi0758), .Y(new_n13973_));
  AOI21X1  g11537(.A0(new_n11947_), .A1(new_n13973_), .B0(pi0039), .Y(new_n13974_));
  OAI21X1  g11538(.A0(new_n12909_), .A1(new_n13973_), .B0(new_n13974_), .Y(new_n13975_));
  AOI21X1  g11539(.A0(new_n13975_), .A1(new_n13972_), .B0(new_n7548_), .Y(new_n13976_));
  MX2X1    g11540(.A(new_n12198_), .B(new_n13683_), .S0(new_n2959_), .Y(new_n13977_));
  NOR3X1   g11541(.A(new_n13977_), .B(new_n13973_), .C(pi0144), .Y(new_n13978_));
  OAI21X1  g11542(.A0(new_n13978_), .A1(new_n13976_), .B0(new_n2996_), .Y(new_n13979_));
  NOR2X1   g11543(.A(new_n12202_), .B(pi0144), .Y(new_n13980_));
  AOI21X1  g11544(.A0(new_n12120_), .A1(pi0758), .B0(new_n12901_), .Y(new_n13981_));
  NOR3X1   g11545(.A(new_n13981_), .B(new_n13980_), .C(new_n2996_), .Y(new_n13982_));
  INVX1    g11546(.A(new_n13982_), .Y(new_n13983_));
  NAND3X1  g11547(.A(new_n13983_), .B(new_n13979_), .C(new_n13969_), .Y(new_n13984_));
  OR2X1    g11548(.A(new_n12288_), .B(new_n2953_), .Y(new_n13985_));
  OAI21X1  g11549(.A0(new_n12274_), .A1(pi0299), .B0(new_n13985_), .Y(new_n13986_));
  OR2X1    g11550(.A(new_n12338_), .B(new_n2953_), .Y(new_n13987_));
  OR2X1    g11551(.A(new_n12348_), .B(new_n12345_), .Y(new_n13988_));
  AND2X1   g11552(.A(new_n13988_), .B(new_n13987_), .Y(new_n13989_));
  OAI21X1  g11553(.A0(new_n13989_), .A1(pi0144), .B0(new_n13973_), .Y(new_n13990_));
  AOI21X1  g11554(.A0(new_n13986_), .A1(pi0144), .B0(new_n13990_), .Y(new_n13991_));
  AOI21X1  g11555(.A0(new_n12440_), .A1(pi0144), .B0(new_n13973_), .Y(new_n13992_));
  OAI21X1  g11556(.A0(new_n12401_), .A1(pi0144), .B0(new_n13992_), .Y(new_n13993_));
  NAND2X1  g11557(.A(new_n13993_), .B(pi0039), .Y(new_n13994_));
  INVX1    g11558(.A(new_n12467_), .Y(new_n13995_));
  OAI21X1  g11559(.A0(new_n13683_), .A1(new_n5029_), .B0(new_n13391_), .Y(new_n13996_));
  AOI21X1  g11560(.A0(new_n13996_), .A1(pi0144), .B0(pi0758), .Y(new_n13997_));
  OAI21X1  g11561(.A0(new_n13995_), .A1(pi0144), .B0(new_n13997_), .Y(new_n13998_));
  NAND3X1  g11562(.A(new_n12453_), .B(new_n12104_), .C(pi0144), .Y(new_n13999_));
  AOI21X1  g11563(.A0(new_n12474_), .A1(new_n7548_), .B0(new_n13973_), .Y(new_n14000_));
  AOI21X1  g11564(.A0(new_n14000_), .A1(new_n13999_), .B0(pi0039), .Y(new_n14001_));
  AOI21X1  g11565(.A0(new_n14001_), .A1(new_n13998_), .B0(pi0038), .Y(new_n14002_));
  OAI21X1  g11566(.A0(new_n13994_), .A1(new_n13991_), .B0(new_n14002_), .Y(new_n14003_));
  NOR3X1   g11567(.A(new_n13982_), .B(new_n13676_), .C(new_n13969_), .Y(new_n14004_));
  AOI21X1  g11568(.A0(new_n14004_), .A1(new_n14003_), .B0(new_n3810_), .Y(new_n14005_));
  AOI22X1  g11569(.A0(new_n14005_), .A1(new_n13984_), .B0(new_n3810_), .B1(pi0144), .Y(new_n14006_));
  AND2X1   g11570(.A(new_n14006_), .B(new_n12493_), .Y(new_n14007_));
  NAND2X1  g11571(.A(new_n13983_), .B(new_n13979_), .Y(new_n14008_));
  MX2X1    g11572(.A(new_n14008_), .B(pi0144), .S0(new_n3810_), .Y(new_n14009_));
  OAI21X1  g11573(.A0(new_n14009_), .A1(new_n12493_), .B0(new_n12494_), .Y(new_n14010_));
  OAI21X1  g11574(.A0(new_n12574_), .A1(new_n3810_), .B0(pi0144), .Y(new_n14011_));
  NOR4X1   g11575(.A(new_n3125_), .B(new_n13969_), .C(pi0100), .D(pi0087), .Y(new_n14012_));
  INVX1    g11576(.A(new_n14012_), .Y(new_n14013_));
  OAI21X1  g11577(.A0(new_n12955_), .A1(pi0144), .B0(new_n2996_), .Y(new_n14014_));
  AOI21X1  g11578(.A0(new_n12953_), .A1(pi0144), .B0(new_n14014_), .Y(new_n14015_));
  AOI21X1  g11579(.A0(new_n12499_), .A1(new_n12202_), .B0(new_n2996_), .Y(new_n14016_));
  INVX1    g11580(.A(new_n14016_), .Y(new_n14017_));
  OAI21X1  g11581(.A0(new_n14017_), .A1(new_n13980_), .B0(new_n14012_), .Y(new_n14018_));
  NOR2X1   g11582(.A(new_n14018_), .B(new_n14015_), .Y(new_n14019_));
  AOI21X1  g11583(.A0(new_n14013_), .A1(new_n14011_), .B0(new_n14019_), .Y(new_n14020_));
  AOI21X1  g11584(.A0(new_n14011_), .A1(new_n12493_), .B0(new_n12494_), .Y(new_n14021_));
  OAI21X1  g11585(.A0(new_n14020_), .A1(new_n12493_), .B0(new_n14021_), .Y(new_n14022_));
  AND2X1   g11586(.A(new_n14022_), .B(new_n12584_), .Y(new_n14023_));
  OAI21X1  g11587(.A0(new_n14010_), .A1(new_n14007_), .B0(new_n14023_), .Y(new_n14024_));
  AND2X1   g11588(.A(new_n14006_), .B(pi0625), .Y(new_n14025_));
  OAI21X1  g11589(.A0(new_n14009_), .A1(pi0625), .B0(pi1153), .Y(new_n14026_));
  AOI21X1  g11590(.A0(new_n14011_), .A1(pi0625), .B0(pi1153), .Y(new_n14027_));
  OAI21X1  g11591(.A0(new_n14020_), .A1(pi0625), .B0(new_n14027_), .Y(new_n14028_));
  AND2X1   g11592(.A(new_n14028_), .B(pi0608), .Y(new_n14029_));
  OAI21X1  g11593(.A0(new_n14026_), .A1(new_n14025_), .B0(new_n14029_), .Y(new_n14030_));
  AOI21X1  g11594(.A0(new_n14030_), .A1(new_n14024_), .B0(new_n11889_), .Y(new_n14031_));
  AND2X1   g11595(.A(new_n14006_), .B(new_n11889_), .Y(new_n14032_));
  OAI21X1  g11596(.A0(new_n14032_), .A1(new_n14031_), .B0(new_n12590_), .Y(new_n14033_));
  AND2X1   g11597(.A(new_n14020_), .B(new_n11889_), .Y(new_n14034_));
  NAND2X1  g11598(.A(new_n14028_), .B(new_n14022_), .Y(new_n14035_));
  AOI21X1  g11599(.A0(new_n14035_), .A1(pi0778), .B0(new_n14034_), .Y(new_n14036_));
  AOI21X1  g11600(.A0(new_n14036_), .A1(pi0609), .B0(pi1155), .Y(new_n14037_));
  NAND2X1  g11601(.A(new_n14011_), .B(new_n12601_), .Y(new_n14038_));
  OAI21X1  g11602(.A0(new_n14009_), .A1(new_n12601_), .B0(new_n14038_), .Y(new_n14039_));
  INVX1    g11603(.A(new_n14011_), .Y(new_n14040_));
  OAI21X1  g11604(.A0(new_n14040_), .A1(pi0609), .B0(pi1155), .Y(new_n14041_));
  AOI21X1  g11605(.A0(new_n14039_), .A1(pi0609), .B0(new_n14041_), .Y(new_n14042_));
  OR2X1    g11606(.A(new_n14042_), .B(pi0660), .Y(new_n14043_));
  AOI21X1  g11607(.A0(new_n14037_), .A1(new_n14033_), .B0(new_n14043_), .Y(new_n14044_));
  OAI21X1  g11608(.A0(new_n14032_), .A1(new_n14031_), .B0(pi0609), .Y(new_n14045_));
  AOI21X1  g11609(.A0(new_n14036_), .A1(new_n12590_), .B0(new_n12591_), .Y(new_n14046_));
  OAI21X1  g11610(.A0(new_n14040_), .A1(new_n12590_), .B0(new_n12591_), .Y(new_n14047_));
  AOI21X1  g11611(.A0(new_n14039_), .A1(new_n12590_), .B0(new_n14047_), .Y(new_n14048_));
  OR2X1    g11612(.A(new_n14048_), .B(new_n12596_), .Y(new_n14049_));
  AOI21X1  g11613(.A0(new_n14046_), .A1(new_n14045_), .B0(new_n14049_), .Y(new_n14050_));
  OAI21X1  g11614(.A0(new_n14050_), .A1(new_n14044_), .B0(pi0785), .Y(new_n14051_));
  OAI21X1  g11615(.A0(new_n14032_), .A1(new_n14031_), .B0(new_n11888_), .Y(new_n14052_));
  AOI21X1  g11616(.A0(new_n14052_), .A1(new_n14051_), .B0(pi0618), .Y(new_n14053_));
  AND2X1   g11617(.A(new_n14011_), .B(new_n12618_), .Y(new_n14054_));
  AOI21X1  g11618(.A0(new_n14036_), .A1(new_n13598_), .B0(new_n14054_), .Y(new_n14055_));
  OAI21X1  g11619(.A0(new_n14055_), .A1(new_n12614_), .B0(new_n12615_), .Y(new_n14056_));
  OAI21X1  g11620(.A0(new_n14048_), .A1(new_n14042_), .B0(pi0785), .Y(new_n14057_));
  OAI21X1  g11621(.A0(new_n14039_), .A1(pi0785), .B0(new_n14057_), .Y(new_n14058_));
  AOI21X1  g11622(.A0(new_n14011_), .A1(new_n12614_), .B0(new_n12615_), .Y(new_n14059_));
  OAI21X1  g11623(.A0(new_n14058_), .A1(new_n12614_), .B0(new_n14059_), .Y(new_n14060_));
  AND2X1   g11624(.A(new_n14060_), .B(new_n12622_), .Y(new_n14061_));
  OAI21X1  g11625(.A0(new_n14056_), .A1(new_n14053_), .B0(new_n14061_), .Y(new_n14062_));
  AOI21X1  g11626(.A0(new_n14052_), .A1(new_n14051_), .B0(new_n12614_), .Y(new_n14063_));
  OAI21X1  g11627(.A0(new_n14055_), .A1(pi0618), .B0(pi1154), .Y(new_n14064_));
  AOI21X1  g11628(.A0(new_n14011_), .A1(pi0618), .B0(pi1154), .Y(new_n14065_));
  OAI21X1  g11629(.A0(new_n14058_), .A1(pi0618), .B0(new_n14065_), .Y(new_n14066_));
  AND2X1   g11630(.A(new_n14066_), .B(pi0627), .Y(new_n14067_));
  OAI21X1  g11631(.A0(new_n14064_), .A1(new_n14063_), .B0(new_n14067_), .Y(new_n14068_));
  AOI21X1  g11632(.A0(new_n14068_), .A1(new_n14062_), .B0(new_n11887_), .Y(new_n14069_));
  AOI21X1  g11633(.A0(new_n14052_), .A1(new_n14051_), .B0(pi0781), .Y(new_n14070_));
  OAI21X1  g11634(.A0(new_n14070_), .A1(new_n14069_), .B0(new_n12637_), .Y(new_n14071_));
  MX2X1    g11635(.A(new_n14055_), .B(new_n14040_), .S0(new_n12641_), .Y(new_n14072_));
  INVX1    g11636(.A(new_n14072_), .Y(new_n14073_));
  AOI21X1  g11637(.A0(new_n14073_), .A1(pi0619), .B0(pi1159), .Y(new_n14074_));
  AOI21X1  g11638(.A0(new_n14066_), .A1(new_n14060_), .B0(new_n11887_), .Y(new_n14075_));
  AOI21X1  g11639(.A0(new_n14058_), .A1(new_n11887_), .B0(new_n14075_), .Y(new_n14076_));
  OAI21X1  g11640(.A0(new_n14040_), .A1(pi0619), .B0(pi1159), .Y(new_n14077_));
  AOI21X1  g11641(.A0(new_n14076_), .A1(pi0619), .B0(new_n14077_), .Y(new_n14078_));
  OR2X1    g11642(.A(new_n14078_), .B(pi0648), .Y(new_n14079_));
  AOI21X1  g11643(.A0(new_n14074_), .A1(new_n14071_), .B0(new_n14079_), .Y(new_n14080_));
  OAI21X1  g11644(.A0(new_n14070_), .A1(new_n14069_), .B0(pi0619), .Y(new_n14081_));
  AOI21X1  g11645(.A0(new_n14073_), .A1(new_n12637_), .B0(new_n12638_), .Y(new_n14082_));
  OAI21X1  g11646(.A0(new_n14040_), .A1(new_n12637_), .B0(new_n12638_), .Y(new_n14083_));
  AOI21X1  g11647(.A0(new_n14076_), .A1(new_n12637_), .B0(new_n14083_), .Y(new_n14084_));
  OR2X1    g11648(.A(new_n14084_), .B(new_n12645_), .Y(new_n14085_));
  AOI21X1  g11649(.A0(new_n14082_), .A1(new_n14081_), .B0(new_n14085_), .Y(new_n14086_));
  OAI21X1  g11650(.A0(new_n14086_), .A1(new_n14080_), .B0(pi0789), .Y(new_n14087_));
  OAI21X1  g11651(.A0(new_n14070_), .A1(new_n14069_), .B0(new_n11886_), .Y(new_n14088_));
  NAND3X1  g11652(.A(new_n14088_), .B(new_n14087_), .C(new_n11885_), .Y(new_n14089_));
  NAND3X1  g11653(.A(new_n14088_), .B(new_n14087_), .C(new_n12664_), .Y(new_n14090_));
  MX2X1    g11654(.A(new_n14072_), .B(new_n14040_), .S0(new_n12659_), .Y(new_n14091_));
  AOI21X1  g11655(.A0(new_n14091_), .A1(pi0626), .B0(pi0641), .Y(new_n14092_));
  OAI21X1  g11656(.A0(new_n14084_), .A1(new_n14078_), .B0(pi0789), .Y(new_n14093_));
  OAI21X1  g11657(.A0(new_n14076_), .A1(pi0789), .B0(new_n14093_), .Y(new_n14094_));
  AOI21X1  g11658(.A0(new_n14011_), .A1(pi0626), .B0(pi1158), .Y(new_n14095_));
  OAI21X1  g11659(.A0(new_n14094_), .A1(pi0626), .B0(new_n14095_), .Y(new_n14096_));
  AOI22X1  g11660(.A0(new_n14096_), .A1(new_n13027_), .B0(new_n14092_), .B1(new_n14090_), .Y(new_n14097_));
  NAND3X1  g11661(.A(new_n14088_), .B(new_n14087_), .C(pi0626), .Y(new_n14098_));
  AOI21X1  g11662(.A0(new_n14091_), .A1(new_n12664_), .B0(new_n12672_), .Y(new_n14099_));
  AOI21X1  g11663(.A0(new_n14011_), .A1(new_n12664_), .B0(new_n12676_), .Y(new_n14100_));
  OAI21X1  g11664(.A0(new_n14094_), .A1(new_n12664_), .B0(new_n14100_), .Y(new_n14101_));
  AOI22X1  g11665(.A0(new_n14101_), .A1(new_n13035_), .B0(new_n14099_), .B1(new_n14098_), .Y(new_n14102_));
  OAI21X1  g11666(.A0(new_n14102_), .A1(new_n14097_), .B0(pi0788), .Y(new_n14103_));
  NAND3X1  g11667(.A(new_n14103_), .B(new_n14089_), .C(new_n12683_), .Y(new_n14104_));
  AOI21X1  g11668(.A0(new_n14101_), .A1(new_n14096_), .B0(new_n11885_), .Y(new_n14105_));
  AND2X1   g11669(.A(new_n14094_), .B(new_n11885_), .Y(new_n14106_));
  NOR2X1   g11670(.A(new_n14106_), .B(new_n14105_), .Y(new_n14107_));
  AOI21X1  g11671(.A0(new_n14107_), .A1(pi0628), .B0(pi1156), .Y(new_n14108_));
  MX2X1    g11672(.A(new_n14091_), .B(new_n14040_), .S0(new_n12691_), .Y(new_n14109_));
  AOI21X1  g11673(.A0(new_n14011_), .A1(new_n12683_), .B0(new_n12684_), .Y(new_n14110_));
  OAI21X1  g11674(.A0(new_n14109_), .A1(new_n12683_), .B0(new_n14110_), .Y(new_n14111_));
  NAND2X1  g11675(.A(new_n14111_), .B(new_n12689_), .Y(new_n14112_));
  AOI21X1  g11676(.A0(new_n14108_), .A1(new_n14104_), .B0(new_n14112_), .Y(new_n14113_));
  NAND3X1  g11677(.A(new_n14103_), .B(new_n14089_), .C(pi0628), .Y(new_n14114_));
  AOI21X1  g11678(.A0(new_n14107_), .A1(new_n12683_), .B0(new_n12684_), .Y(new_n14115_));
  AOI21X1  g11679(.A0(new_n14011_), .A1(pi0628), .B0(pi1156), .Y(new_n14116_));
  OAI21X1  g11680(.A0(new_n14109_), .A1(pi0628), .B0(new_n14116_), .Y(new_n14117_));
  NAND2X1  g11681(.A(new_n14117_), .B(pi0629), .Y(new_n14118_));
  AOI21X1  g11682(.A0(new_n14115_), .A1(new_n14114_), .B0(new_n14118_), .Y(new_n14119_));
  OAI21X1  g11683(.A0(new_n14119_), .A1(new_n14113_), .B0(pi0792), .Y(new_n14120_));
  NAND3X1  g11684(.A(new_n14103_), .B(new_n14089_), .C(new_n11884_), .Y(new_n14121_));
  AOI21X1  g11685(.A0(new_n14121_), .A1(new_n14120_), .B0(pi0647), .Y(new_n14122_));
  INVX1    g11686(.A(new_n12711_), .Y(new_n14123_));
  OR2X1    g11687(.A(new_n14011_), .B(new_n14123_), .Y(new_n14124_));
  OAI21X1  g11688(.A0(new_n14107_), .A1(new_n12711_), .B0(new_n14124_), .Y(new_n14125_));
  OAI21X1  g11689(.A0(new_n14125_), .A1(new_n12705_), .B0(new_n12706_), .Y(new_n14126_));
  AND2X1   g11690(.A(new_n14109_), .B(new_n11884_), .Y(new_n14127_));
  AOI21X1  g11691(.A0(new_n14117_), .A1(new_n14111_), .B0(new_n11884_), .Y(new_n14128_));
  NOR2X1   g11692(.A(new_n14128_), .B(new_n14127_), .Y(new_n14129_));
  INVX1    g11693(.A(new_n14129_), .Y(new_n14130_));
  AOI21X1  g11694(.A0(new_n14011_), .A1(new_n12705_), .B0(new_n12706_), .Y(new_n14131_));
  OAI21X1  g11695(.A0(new_n14130_), .A1(new_n12705_), .B0(new_n14131_), .Y(new_n14132_));
  AND2X1   g11696(.A(new_n14132_), .B(new_n12723_), .Y(new_n14133_));
  OAI21X1  g11697(.A0(new_n14126_), .A1(new_n14122_), .B0(new_n14133_), .Y(new_n14134_));
  AOI21X1  g11698(.A0(new_n14121_), .A1(new_n14120_), .B0(new_n12705_), .Y(new_n14135_));
  OAI21X1  g11699(.A0(new_n14125_), .A1(pi0647), .B0(pi1157), .Y(new_n14136_));
  AOI21X1  g11700(.A0(new_n14011_), .A1(pi0647), .B0(pi1157), .Y(new_n14137_));
  OAI21X1  g11701(.A0(new_n14130_), .A1(pi0647), .B0(new_n14137_), .Y(new_n14138_));
  AND2X1   g11702(.A(new_n14138_), .B(pi0630), .Y(new_n14139_));
  OAI21X1  g11703(.A0(new_n14136_), .A1(new_n14135_), .B0(new_n14139_), .Y(new_n14140_));
  AOI21X1  g11704(.A0(new_n14140_), .A1(new_n14134_), .B0(new_n11883_), .Y(new_n14141_));
  AOI21X1  g11705(.A0(new_n14121_), .A1(new_n14120_), .B0(pi0787), .Y(new_n14142_));
  OAI21X1  g11706(.A0(new_n14142_), .A1(new_n14141_), .B0(pi0644), .Y(new_n14143_));
  AND2X1   g11707(.A(new_n14138_), .B(new_n14132_), .Y(new_n14144_));
  MX2X1    g11708(.A(new_n14144_), .B(new_n14129_), .S0(new_n11883_), .Y(new_n14145_));
  AOI21X1  g11709(.A0(new_n14145_), .A1(new_n12743_), .B0(new_n12739_), .Y(new_n14146_));
  MX2X1    g11710(.A(new_n14125_), .B(new_n14040_), .S0(new_n12735_), .Y(new_n14147_));
  NOR2X1   g11711(.A(new_n14147_), .B(new_n12743_), .Y(new_n14148_));
  OAI21X1  g11712(.A0(new_n14040_), .A1(pi0644), .B0(new_n12739_), .Y(new_n14149_));
  OAI21X1  g11713(.A0(new_n14149_), .A1(new_n14148_), .B0(pi1160), .Y(new_n14150_));
  AOI21X1  g11714(.A0(new_n14146_), .A1(new_n14143_), .B0(new_n14150_), .Y(new_n14151_));
  OAI21X1  g11715(.A0(new_n14142_), .A1(new_n14141_), .B0(new_n12743_), .Y(new_n14152_));
  AOI21X1  g11716(.A0(new_n14145_), .A1(pi0644), .B0(pi0715), .Y(new_n14153_));
  NOR2X1   g11717(.A(new_n14147_), .B(pi0644), .Y(new_n14154_));
  OAI21X1  g11718(.A0(new_n14040_), .A1(new_n12743_), .B0(pi0715), .Y(new_n14155_));
  OAI21X1  g11719(.A0(new_n14155_), .A1(new_n14154_), .B0(new_n11882_), .Y(new_n14156_));
  AOI21X1  g11720(.A0(new_n14153_), .A1(new_n14152_), .B0(new_n14156_), .Y(new_n14157_));
  NOR3X1   g11721(.A(new_n14157_), .B(new_n14151_), .C(new_n12897_), .Y(new_n14158_));
  NOR3X1   g11722(.A(new_n14142_), .B(new_n14141_), .C(pi0790), .Y(new_n14159_));
  OR2X1    g11723(.A(new_n14159_), .B(new_n5118_), .Y(new_n14160_));
  AOI21X1  g11724(.A0(new_n5118_), .A1(new_n7548_), .B0(pi0057), .Y(new_n14161_));
  OAI21X1  g11725(.A0(new_n14160_), .A1(new_n14158_), .B0(new_n14161_), .Y(new_n14162_));
  AOI21X1  g11726(.A0(pi0144), .A1(pi0057), .B0(pi0832), .Y(new_n14163_));
  NOR2X1   g11727(.A(new_n2739_), .B(new_n7548_), .Y(new_n14164_));
  AOI21X1  g11728(.A0(new_n12566_), .A1(pi0736), .B0(new_n14164_), .Y(new_n14165_));
  INVX1    g11729(.A(new_n14165_), .Y(new_n14166_));
  NOR3X1   g11730(.A(new_n13585_), .B(new_n13969_), .C(new_n12493_), .Y(new_n14167_));
  OR2X1    g11731(.A(new_n14167_), .B(new_n14165_), .Y(new_n14168_));
  NOR3X1   g11732(.A(new_n14167_), .B(new_n14164_), .C(new_n12494_), .Y(new_n14169_));
  AOI21X1  g11733(.A0(new_n14168_), .A1(new_n12494_), .B0(new_n14169_), .Y(new_n14170_));
  MX2X1    g11734(.A(new_n14170_), .B(new_n14166_), .S0(new_n11889_), .Y(new_n14171_));
  INVX1    g11735(.A(new_n14171_), .Y(new_n14172_));
  NOR2X1   g11736(.A(new_n14172_), .B(new_n13624_), .Y(new_n14173_));
  AOI21X1  g11737(.A0(new_n14173_), .A1(new_n12683_), .B0(new_n12689_), .Y(new_n14174_));
  INVX1    g11738(.A(new_n12841_), .Y(new_n14175_));
  NOR2X1   g11739(.A(pi1155), .B(pi0609), .Y(new_n14176_));
  AND2X1   g11740(.A(pi1155), .B(pi0609), .Y(new_n14177_));
  NOR3X1   g11741(.A(new_n14177_), .B(new_n14176_), .C(new_n11888_), .Y(new_n14178_));
  XOR2X1   g11742(.A(pi1159), .B(pi0619), .Y(new_n14179_));
  AND2X1   g11743(.A(new_n14179_), .B(pi0789), .Y(new_n14180_));
  NOR2X1   g11744(.A(pi1154), .B(pi0618), .Y(new_n14181_));
  AND2X1   g11745(.A(pi1154), .B(pi0618), .Y(new_n14182_));
  NOR3X1   g11746(.A(new_n14182_), .B(new_n14181_), .C(new_n11887_), .Y(new_n14183_));
  OR2X1    g11747(.A(new_n14183_), .B(new_n12601_), .Y(new_n14184_));
  OR2X1    g11748(.A(new_n14184_), .B(new_n14180_), .Y(new_n14185_));
  NOR4X1   g11749(.A(new_n14185_), .B(new_n14178_), .C(new_n12204_), .D(new_n13973_), .Y(new_n14186_));
  AOI21X1  g11750(.A0(new_n14186_), .A1(new_n14175_), .B0(new_n12683_), .Y(new_n14187_));
  OAI21X1  g11751(.A0(new_n14187_), .A1(new_n14174_), .B0(new_n12684_), .Y(new_n14188_));
  INVX1    g11752(.A(new_n14173_), .Y(new_n14189_));
  AOI21X1  g11753(.A0(new_n14186_), .A1(new_n14175_), .B0(pi0628), .Y(new_n14190_));
  NOR2X1   g11754(.A(new_n14190_), .B(new_n12689_), .Y(new_n14191_));
  NOR2X1   g11755(.A(new_n14191_), .B(new_n12684_), .Y(new_n14192_));
  OAI21X1  g11756(.A0(new_n14189_), .A1(new_n12683_), .B0(new_n14192_), .Y(new_n14193_));
  AOI21X1  g11757(.A0(new_n14193_), .A1(new_n14188_), .B0(new_n14164_), .Y(new_n14194_));
  INVX1    g11758(.A(new_n14194_), .Y(new_n14195_));
  AND2X1   g11759(.A(pi1158), .B(new_n12664_), .Y(new_n14196_));
  INVX1    g11760(.A(new_n14164_), .Y(new_n14197_));
  INVX1    g11761(.A(new_n12641_), .Y(new_n14198_));
  NAND3X1  g11762(.A(new_n14171_), .B(new_n14198_), .C(new_n13598_), .Y(new_n14199_));
  OAI21X1  g11763(.A0(new_n14199_), .A1(new_n12659_), .B0(new_n14197_), .Y(new_n14200_));
  AOI21X1  g11764(.A0(new_n14186_), .A1(new_n12664_), .B0(new_n14164_), .Y(new_n14201_));
  OAI21X1  g11765(.A0(new_n14201_), .A1(pi1158), .B0(pi0641), .Y(new_n14202_));
  AOI21X1  g11766(.A0(new_n14200_), .A1(new_n14196_), .B0(new_n14202_), .Y(new_n14203_));
  AND2X1   g11767(.A(new_n12676_), .B(pi0626), .Y(new_n14204_));
  AOI21X1  g11768(.A0(new_n14186_), .A1(pi0626), .B0(new_n14164_), .Y(new_n14205_));
  OAI21X1  g11769(.A0(new_n14205_), .A1(new_n12676_), .B0(new_n12672_), .Y(new_n14206_));
  AOI21X1  g11770(.A0(new_n14200_), .A1(new_n14204_), .B0(new_n14206_), .Y(new_n14207_));
  NOR3X1   g11771(.A(new_n14207_), .B(new_n14203_), .C(new_n11885_), .Y(new_n14208_));
  INVX1    g11772(.A(new_n13576_), .Y(new_n14209_));
  AOI21X1  g11773(.A0(new_n12178_), .A1(pi0758), .B0(new_n14164_), .Y(new_n14210_));
  OAI21X1  g11774(.A0(new_n14209_), .A1(new_n13969_), .B0(new_n14210_), .Y(new_n14211_));
  NAND3X1  g11775(.A(new_n13576_), .B(pi0736), .C(pi0625), .Y(new_n14212_));
  AOI21X1  g11776(.A0(new_n14212_), .A1(new_n14211_), .B0(pi1153), .Y(new_n14213_));
  OR2X1    g11777(.A(new_n14169_), .B(pi0608), .Y(new_n14214_));
  OR2X1    g11778(.A(new_n14214_), .B(new_n14213_), .Y(new_n14215_));
  NAND3X1  g11779(.A(new_n14212_), .B(new_n14210_), .C(pi1153), .Y(new_n14216_));
  AOI21X1  g11780(.A0(new_n14168_), .A1(new_n12494_), .B0(new_n12584_), .Y(new_n14217_));
  NAND2X1  g11781(.A(new_n14217_), .B(new_n14216_), .Y(new_n14218_));
  AOI21X1  g11782(.A0(new_n14218_), .A1(new_n14215_), .B0(new_n11889_), .Y(new_n14219_));
  AOI21X1  g11783(.A0(new_n14211_), .A1(new_n11889_), .B0(new_n14219_), .Y(new_n14220_));
  AOI21X1  g11784(.A0(new_n14171_), .A1(pi0609), .B0(pi1155), .Y(new_n14221_));
  OAI21X1  g11785(.A0(new_n14220_), .A1(pi0609), .B0(new_n14221_), .Y(new_n14222_));
  NAND3X1  g11786(.A(new_n12599_), .B(new_n12178_), .C(pi0758), .Y(new_n14223_));
  NOR2X1   g11787(.A(new_n14164_), .B(new_n12591_), .Y(new_n14224_));
  AOI21X1  g11788(.A0(new_n14224_), .A1(new_n14223_), .B0(pi0660), .Y(new_n14225_));
  AOI21X1  g11789(.A0(new_n14171_), .A1(new_n12590_), .B0(new_n12591_), .Y(new_n14226_));
  OAI21X1  g11790(.A0(new_n14220_), .A1(new_n12590_), .B0(new_n14226_), .Y(new_n14227_));
  NAND3X1  g11791(.A(new_n12608_), .B(new_n12178_), .C(pi0758), .Y(new_n14228_));
  NOR2X1   g11792(.A(new_n14164_), .B(pi1155), .Y(new_n14229_));
  AOI21X1  g11793(.A0(new_n14229_), .A1(new_n14228_), .B0(new_n12596_), .Y(new_n14230_));
  AOI22X1  g11794(.A0(new_n14230_), .A1(new_n14227_), .B0(new_n14225_), .B1(new_n14222_), .Y(new_n14231_));
  MX2X1    g11795(.A(new_n14231_), .B(new_n14220_), .S0(new_n11888_), .Y(new_n14232_));
  AOI21X1  g11796(.A0(new_n14171_), .A1(new_n13598_), .B0(new_n14164_), .Y(new_n14233_));
  INVX1    g11797(.A(new_n14233_), .Y(new_n14234_));
  AOI21X1  g11798(.A0(new_n14234_), .A1(pi0618), .B0(pi1154), .Y(new_n14235_));
  OAI21X1  g11799(.A0(new_n14232_), .A1(pi0618), .B0(new_n14235_), .Y(new_n14236_));
  NOR3X1   g11800(.A(new_n14178_), .B(new_n12204_), .C(new_n13973_), .Y(new_n14237_));
  INVX1    g11801(.A(new_n14237_), .Y(new_n14238_));
  NOR3X1   g11802(.A(new_n14238_), .B(new_n12601_), .C(new_n12614_), .Y(new_n14239_));
  NOR3X1   g11803(.A(new_n14239_), .B(new_n14164_), .C(new_n12615_), .Y(new_n14240_));
  NOR2X1   g11804(.A(new_n14240_), .B(pi0627), .Y(new_n14241_));
  AOI21X1  g11805(.A0(new_n14234_), .A1(new_n12614_), .B0(new_n12615_), .Y(new_n14242_));
  OAI21X1  g11806(.A0(new_n14232_), .A1(new_n12614_), .B0(new_n14242_), .Y(new_n14243_));
  NOR3X1   g11807(.A(new_n14238_), .B(new_n12601_), .C(pi0618), .Y(new_n14244_));
  NOR3X1   g11808(.A(new_n14244_), .B(new_n14164_), .C(pi1154), .Y(new_n14245_));
  NOR2X1   g11809(.A(new_n14245_), .B(new_n12622_), .Y(new_n14246_));
  AOI22X1  g11810(.A0(new_n14246_), .A1(new_n14243_), .B0(new_n14241_), .B1(new_n14236_), .Y(new_n14247_));
  MX2X1    g11811(.A(new_n14247_), .B(new_n14232_), .S0(new_n11887_), .Y(new_n14248_));
  AND2X1   g11812(.A(new_n14199_), .B(new_n14197_), .Y(new_n14249_));
  INVX1    g11813(.A(new_n14249_), .Y(new_n14250_));
  AOI21X1  g11814(.A0(new_n14250_), .A1(pi0619), .B0(pi1159), .Y(new_n14251_));
  OAI21X1  g11815(.A0(new_n14248_), .A1(pi0619), .B0(new_n14251_), .Y(new_n14252_));
  NOR4X1   g11816(.A(new_n14183_), .B(new_n14238_), .C(new_n12601_), .D(new_n12637_), .Y(new_n14253_));
  NOR3X1   g11817(.A(new_n14253_), .B(new_n14164_), .C(new_n12638_), .Y(new_n14254_));
  NOR2X1   g11818(.A(new_n14254_), .B(pi0648), .Y(new_n14255_));
  AND2X1   g11819(.A(new_n14255_), .B(new_n14252_), .Y(new_n14256_));
  INVX1    g11820(.A(new_n14256_), .Y(new_n14257_));
  AOI21X1  g11821(.A0(new_n14250_), .A1(new_n12637_), .B0(new_n12638_), .Y(new_n14258_));
  OAI21X1  g11822(.A0(new_n14248_), .A1(new_n12637_), .B0(new_n14258_), .Y(new_n14259_));
  NOR4X1   g11823(.A(new_n14183_), .B(new_n14238_), .C(new_n12601_), .D(pi0619), .Y(new_n14260_));
  NOR3X1   g11824(.A(new_n14260_), .B(new_n14164_), .C(pi1159), .Y(new_n14261_));
  NOR2X1   g11825(.A(new_n14261_), .B(new_n12645_), .Y(new_n14262_));
  AOI21X1  g11826(.A0(new_n14262_), .A1(new_n14259_), .B0(new_n11886_), .Y(new_n14263_));
  INVX1    g11827(.A(new_n12842_), .Y(new_n14264_));
  AOI21X1  g11828(.A0(new_n14248_), .A1(new_n11886_), .B0(new_n14264_), .Y(new_n14265_));
  INVX1    g11829(.A(new_n14265_), .Y(new_n14266_));
  AOI21X1  g11830(.A0(new_n14263_), .A1(new_n14257_), .B0(new_n14266_), .Y(new_n14267_));
  OAI22X1  g11831(.A0(new_n14267_), .A1(new_n14208_), .B0(new_n14195_), .B1(new_n11884_), .Y(new_n14268_));
  AOI21X1  g11832(.A0(new_n13650_), .A1(new_n12734_), .B0(new_n11883_), .Y(new_n14269_));
  AND2X1   g11833(.A(new_n13637_), .B(pi0629), .Y(new_n14270_));
  NOR3X1   g11834(.A(pi1156), .B(pi0629), .C(pi0628), .Y(new_n14271_));
  OR2X1    g11835(.A(new_n14271_), .B(new_n11884_), .Y(new_n14272_));
  NOR2X1   g11836(.A(new_n14272_), .B(new_n14270_), .Y(new_n14273_));
  AOI21X1  g11837(.A0(new_n14273_), .A1(new_n14195_), .B0(new_n14269_), .Y(new_n14274_));
  NOR4X1   g11838(.A(new_n14185_), .B(new_n14238_), .C(new_n12841_), .D(new_n12711_), .Y(new_n14275_));
  AOI21X1  g11839(.A0(new_n14275_), .A1(new_n12723_), .B0(new_n12705_), .Y(new_n14276_));
  NOR3X1   g11840(.A(new_n14172_), .B(new_n13639_), .C(new_n13624_), .Y(new_n14277_));
  INVX1    g11841(.A(new_n14277_), .Y(new_n14278_));
  AOI21X1  g11842(.A0(new_n14278_), .A1(pi0630), .B0(new_n14276_), .Y(new_n14279_));
  AOI21X1  g11843(.A0(new_n14278_), .A1(new_n12723_), .B0(new_n12705_), .Y(new_n14280_));
  AOI21X1  g11844(.A0(new_n14275_), .A1(pi0630), .B0(new_n12706_), .Y(new_n14281_));
  INVX1    g11845(.A(new_n14281_), .Y(new_n14282_));
  OAI22X1  g11846(.A0(new_n14282_), .A1(new_n14280_), .B0(new_n14279_), .B1(pi1157), .Y(new_n14283_));
  NOR2X1   g11847(.A(new_n14164_), .B(new_n11883_), .Y(new_n14284_));
  AOI22X1  g11848(.A0(new_n14284_), .A1(new_n14283_), .B0(new_n14274_), .B1(new_n14268_), .Y(new_n14285_));
  INVX1    g11849(.A(new_n13651_), .Y(new_n14286_));
  AOI21X1  g11850(.A0(new_n14277_), .A1(new_n14286_), .B0(new_n14164_), .Y(new_n14287_));
  OAI21X1  g11851(.A0(new_n14287_), .A1(pi0644), .B0(pi0715), .Y(new_n14288_));
  AOI21X1  g11852(.A0(new_n14285_), .A1(pi0644), .B0(new_n14288_), .Y(new_n14289_));
  INVX1    g11853(.A(new_n14275_), .Y(new_n14290_));
  NOR3X1   g11854(.A(new_n14290_), .B(new_n12735_), .C(new_n12743_), .Y(new_n14291_));
  OAI21X1  g11855(.A0(new_n2739_), .A1(new_n7548_), .B0(new_n12739_), .Y(new_n14292_));
  OAI21X1  g11856(.A0(new_n14292_), .A1(new_n14291_), .B0(pi1160), .Y(new_n14293_));
  OAI21X1  g11857(.A0(new_n14287_), .A1(new_n12743_), .B0(new_n12739_), .Y(new_n14294_));
  AOI21X1  g11858(.A0(new_n14285_), .A1(new_n12743_), .B0(new_n14294_), .Y(new_n14295_));
  NOR3X1   g11859(.A(new_n14290_), .B(new_n12735_), .C(pi0644), .Y(new_n14296_));
  OAI21X1  g11860(.A0(new_n2739_), .A1(new_n7548_), .B0(pi0715), .Y(new_n14297_));
  OAI21X1  g11861(.A0(new_n14297_), .A1(new_n14296_), .B0(new_n11882_), .Y(new_n14298_));
  OAI22X1  g11862(.A0(new_n14298_), .A1(new_n14295_), .B0(new_n14293_), .B1(new_n14289_), .Y(new_n14299_));
  NAND2X1  g11863(.A(new_n14299_), .B(pi0790), .Y(new_n14300_));
  AOI21X1  g11864(.A0(new_n14285_), .A1(new_n12897_), .B0(new_n12898_), .Y(new_n14301_));
  AOI22X1  g11865(.A0(new_n14301_), .A1(new_n14300_), .B0(new_n14163_), .B1(new_n14162_), .Y(po0301));
  AOI21X1  g11866(.A0(new_n13699_), .A1(new_n3129_), .B0(pi0145), .Y(new_n14303_));
  INVX1    g11867(.A(new_n14303_), .Y(new_n14304_));
  OAI21X1  g11868(.A0(new_n3810_), .A1(pi0698), .B0(new_n14303_), .Y(new_n14305_));
  INVX1    g11869(.A(pi0698), .Y(new_n14306_));
  AOI21X1  g11870(.A0(new_n12955_), .A1(pi0145), .B0(pi0038), .Y(new_n14307_));
  OAI22X1  g11871(.A0(new_n14307_), .A1(new_n3810_), .B0(new_n12953_), .B1(pi0145), .Y(new_n14308_));
  OAI21X1  g11872(.A0(new_n12202_), .A1(pi0145), .B0(new_n12567_), .Y(new_n14309_));
  NAND3X1  g11873(.A(new_n14309_), .B(new_n14308_), .C(new_n14306_), .Y(new_n14310_));
  AND2X1   g11874(.A(new_n14310_), .B(new_n14305_), .Y(new_n14311_));
  AOI21X1  g11875(.A0(new_n14303_), .A1(new_n12493_), .B0(new_n12494_), .Y(new_n14312_));
  OAI21X1  g11876(.A0(new_n14311_), .A1(new_n12493_), .B0(new_n14312_), .Y(new_n14313_));
  AOI21X1  g11877(.A0(new_n14303_), .A1(pi0625), .B0(pi1153), .Y(new_n14314_));
  OAI21X1  g11878(.A0(new_n14311_), .A1(pi0625), .B0(new_n14314_), .Y(new_n14315_));
  AOI21X1  g11879(.A0(new_n14315_), .A1(new_n14313_), .B0(new_n11889_), .Y(new_n14316_));
  AOI21X1  g11880(.A0(new_n14311_), .A1(new_n11889_), .B0(new_n14316_), .Y(new_n14317_));
  MX2X1    g11881(.A(new_n14317_), .B(new_n14303_), .S0(new_n12618_), .Y(new_n14318_));
  MX2X1    g11882(.A(new_n14318_), .B(new_n14303_), .S0(new_n12641_), .Y(new_n14319_));
  MX2X1    g11883(.A(new_n14319_), .B(new_n14303_), .S0(new_n12659_), .Y(new_n14320_));
  INVX1    g11884(.A(new_n14320_), .Y(new_n14321_));
  MX2X1    g11885(.A(new_n14321_), .B(new_n14304_), .S0(new_n12691_), .Y(new_n14322_));
  AND2X1   g11886(.A(new_n14322_), .B(new_n11884_), .Y(new_n14323_));
  AOI21X1  g11887(.A0(new_n14303_), .A1(new_n12683_), .B0(new_n12684_), .Y(new_n14324_));
  OAI21X1  g11888(.A0(new_n14322_), .A1(new_n12683_), .B0(new_n14324_), .Y(new_n14325_));
  AOI21X1  g11889(.A0(new_n14303_), .A1(pi0628), .B0(pi1156), .Y(new_n14326_));
  OAI21X1  g11890(.A0(new_n14322_), .A1(pi0628), .B0(new_n14326_), .Y(new_n14327_));
  AOI21X1  g11891(.A0(new_n14327_), .A1(new_n14325_), .B0(new_n11884_), .Y(new_n14328_));
  NOR2X1   g11892(.A(new_n14328_), .B(new_n14323_), .Y(new_n14329_));
  MX2X1    g11893(.A(new_n14329_), .B(new_n14303_), .S0(pi0647), .Y(new_n14330_));
  MX2X1    g11894(.A(new_n14329_), .B(new_n14303_), .S0(new_n12705_), .Y(new_n14331_));
  MX2X1    g11895(.A(new_n14331_), .B(new_n14330_), .S0(new_n12706_), .Y(new_n14332_));
  NOR3X1   g11896(.A(new_n14328_), .B(new_n14323_), .C(pi0787), .Y(new_n14333_));
  AOI21X1  g11897(.A0(new_n14332_), .A1(pi0787), .B0(new_n14333_), .Y(new_n14334_));
  OAI21X1  g11898(.A0(new_n14334_), .A1(pi0644), .B0(pi0715), .Y(new_n14335_));
  INVX1    g11899(.A(pi0767), .Y(new_n14336_));
  AOI21X1  g11900(.A0(new_n12090_), .A1(new_n5224_), .B0(new_n14336_), .Y(new_n14337_));
  NOR2X1   g11901(.A(pi0767), .B(pi0145), .Y(new_n14338_));
  INVX1    g11902(.A(new_n14338_), .Y(new_n14339_));
  OAI22X1  g11903(.A0(new_n14339_), .A1(new_n12910_), .B0(new_n12199_), .B1(new_n5224_), .Y(new_n14340_));
  OAI21X1  g11904(.A0(new_n14340_), .A1(new_n14337_), .B0(new_n2996_), .Y(new_n14341_));
  INVX1    g11905(.A(new_n12205_), .Y(new_n14342_));
  AOI21X1  g11906(.A0(new_n12901_), .A1(new_n5224_), .B0(new_n2996_), .Y(new_n14343_));
  OAI21X1  g11907(.A0(new_n14342_), .A1(pi0767), .B0(new_n14343_), .Y(new_n14344_));
  AND2X1   g11908(.A(new_n14344_), .B(new_n14341_), .Y(new_n14345_));
  MX2X1    g11909(.A(new_n14345_), .B(new_n5224_), .S0(new_n3810_), .Y(new_n14346_));
  INVX1    g11910(.A(new_n14346_), .Y(new_n14347_));
  MX2X1    g11911(.A(new_n14347_), .B(new_n14304_), .S0(new_n12601_), .Y(new_n14348_));
  NOR2X1   g11912(.A(new_n14346_), .B(new_n12601_), .Y(new_n14349_));
  AOI22X1  g11913(.A0(new_n14349_), .A1(pi0609), .B0(new_n14304_), .B1(new_n13430_), .Y(new_n14350_));
  OR2X1    g11914(.A(new_n14350_), .B(new_n12591_), .Y(new_n14351_));
  AOI22X1  g11915(.A0(new_n14349_), .A1(new_n12590_), .B0(new_n14304_), .B1(new_n13436_), .Y(new_n14352_));
  OR2X1    g11916(.A(new_n14352_), .B(pi1155), .Y(new_n14353_));
  NAND2X1  g11917(.A(new_n14353_), .B(new_n14351_), .Y(new_n14354_));
  MX2X1    g11918(.A(new_n14354_), .B(new_n14348_), .S0(new_n11888_), .Y(new_n14355_));
  AOI21X1  g11919(.A0(new_n14303_), .A1(new_n12614_), .B0(new_n12615_), .Y(new_n14356_));
  OAI21X1  g11920(.A0(new_n14355_), .A1(new_n12614_), .B0(new_n14356_), .Y(new_n14357_));
  AOI21X1  g11921(.A0(new_n14303_), .A1(pi0618), .B0(pi1154), .Y(new_n14358_));
  OAI21X1  g11922(.A0(new_n14355_), .A1(pi0618), .B0(new_n14358_), .Y(new_n14359_));
  NAND2X1  g11923(.A(new_n14359_), .B(new_n14357_), .Y(new_n14360_));
  MX2X1    g11924(.A(new_n14360_), .B(new_n14355_), .S0(new_n11887_), .Y(new_n14361_));
  AND2X1   g11925(.A(new_n14361_), .B(new_n11886_), .Y(new_n14362_));
  AOI21X1  g11926(.A0(new_n14303_), .A1(new_n12637_), .B0(new_n12638_), .Y(new_n14363_));
  OAI21X1  g11927(.A0(new_n14361_), .A1(new_n12637_), .B0(new_n14363_), .Y(new_n14364_));
  AOI21X1  g11928(.A0(new_n14303_), .A1(pi0619), .B0(pi1159), .Y(new_n14365_));
  OAI21X1  g11929(.A0(new_n14361_), .A1(pi0619), .B0(new_n14365_), .Y(new_n14366_));
  AOI21X1  g11930(.A0(new_n14366_), .A1(new_n14364_), .B0(new_n11886_), .Y(new_n14367_));
  NOR2X1   g11931(.A(new_n14367_), .B(new_n14362_), .Y(new_n14368_));
  INVX1    g11932(.A(new_n14368_), .Y(new_n14369_));
  AOI21X1  g11933(.A0(new_n14303_), .A1(new_n12664_), .B0(new_n12676_), .Y(new_n14370_));
  OAI21X1  g11934(.A0(new_n14369_), .A1(new_n12664_), .B0(new_n14370_), .Y(new_n14371_));
  AOI21X1  g11935(.A0(new_n14303_), .A1(pi0626), .B0(pi1158), .Y(new_n14372_));
  OAI21X1  g11936(.A0(new_n14369_), .A1(pi0626), .B0(new_n14372_), .Y(new_n14373_));
  AND2X1   g11937(.A(new_n14373_), .B(new_n14371_), .Y(new_n14374_));
  MX2X1    g11938(.A(new_n14374_), .B(new_n14368_), .S0(new_n11885_), .Y(new_n14375_));
  AND2X1   g11939(.A(new_n14303_), .B(new_n12711_), .Y(new_n14376_));
  AOI21X1  g11940(.A0(new_n14375_), .A1(new_n14123_), .B0(new_n14376_), .Y(new_n14377_));
  MX2X1    g11941(.A(new_n14377_), .B(new_n14304_), .S0(new_n12735_), .Y(new_n14378_));
  AOI21X1  g11942(.A0(new_n14303_), .A1(new_n12743_), .B0(pi0715), .Y(new_n14379_));
  OAI21X1  g11943(.A0(new_n14378_), .A1(new_n12743_), .B0(new_n14379_), .Y(new_n14380_));
  NAND3X1  g11944(.A(new_n14380_), .B(new_n14335_), .C(pi1160), .Y(new_n14381_));
  NOR3X1   g11945(.A(new_n12706_), .B(pi0647), .C(new_n12723_), .Y(new_n14382_));
  NOR3X1   g11946(.A(pi1157), .B(new_n12705_), .C(pi0630), .Y(new_n14383_));
  NOR2X1   g11947(.A(new_n14383_), .B(new_n14382_), .Y(new_n14384_));
  INVX1    g11948(.A(new_n14384_), .Y(new_n14385_));
  AND2X1   g11949(.A(pi1157), .B(new_n12723_), .Y(new_n14386_));
  INVX1    g11950(.A(new_n14386_), .Y(new_n14387_));
  AND2X1   g11951(.A(new_n12706_), .B(pi0630), .Y(new_n14388_));
  INVX1    g11952(.A(new_n14388_), .Y(new_n14389_));
  OAI22X1  g11953(.A0(new_n14331_), .A1(new_n14387_), .B0(new_n14330_), .B1(new_n14389_), .Y(new_n14390_));
  AOI21X1  g11954(.A0(new_n14385_), .A1(new_n14377_), .B0(new_n14390_), .Y(new_n14391_));
  AND2X1   g11955(.A(pi0629), .B(new_n12683_), .Y(new_n14392_));
  AND2X1   g11956(.A(new_n12689_), .B(pi0628), .Y(new_n14393_));
  MX2X1    g11957(.A(new_n14393_), .B(new_n14392_), .S0(pi1156), .Y(new_n14394_));
  INVX1    g11958(.A(new_n14394_), .Y(new_n14395_));
  MX2X1    g11959(.A(new_n14327_), .B(new_n14325_), .S0(new_n12689_), .Y(new_n14396_));
  OAI21X1  g11960(.A0(new_n14395_), .A1(new_n14375_), .B0(new_n14396_), .Y(new_n14397_));
  AOI21X1  g11961(.A0(new_n13989_), .A1(pi0145), .B0(new_n14336_), .Y(new_n14398_));
  OAI21X1  g11962(.A0(new_n13986_), .A1(pi0145), .B0(new_n14398_), .Y(new_n14399_));
  OAI21X1  g11963(.A0(new_n12440_), .A1(pi0145), .B0(new_n14336_), .Y(new_n14400_));
  AOI21X1  g11964(.A0(new_n12401_), .A1(pi0145), .B0(new_n14400_), .Y(new_n14401_));
  NOR2X1   g11965(.A(new_n14401_), .B(new_n2959_), .Y(new_n14402_));
  NAND2X1  g11966(.A(new_n12467_), .B(pi0145), .Y(new_n14403_));
  AOI21X1  g11967(.A0(new_n13996_), .A1(new_n5224_), .B0(new_n14336_), .Y(new_n14404_));
  NAND3X1  g11968(.A(new_n12453_), .B(new_n12104_), .C(new_n5224_), .Y(new_n14405_));
  AOI21X1  g11969(.A0(new_n12474_), .A1(pi0145), .B0(pi0767), .Y(new_n14406_));
  AOI22X1  g11970(.A0(new_n14406_), .A1(new_n14405_), .B0(new_n14404_), .B1(new_n14403_), .Y(new_n14407_));
  OAI21X1  g11971(.A0(new_n14407_), .A1(pi0039), .B0(new_n2996_), .Y(new_n14408_));
  AOI21X1  g11972(.A0(new_n14402_), .A1(new_n14399_), .B0(new_n14408_), .Y(new_n14409_));
  OAI21X1  g11973(.A0(new_n12478_), .A1(pi0767), .B0(new_n13669_), .Y(new_n14410_));
  INVX1    g11974(.A(new_n6857_), .Y(new_n14411_));
  AND2X1   g11975(.A(new_n12178_), .B(new_n14336_), .Y(new_n14412_));
  OAI21X1  g11976(.A0(new_n14412_), .A1(new_n13576_), .B0(pi0145), .Y(new_n14413_));
  OAI21X1  g11977(.A0(new_n14413_), .A1(new_n14411_), .B0(pi0038), .Y(new_n14414_));
  AOI21X1  g11978(.A0(new_n14410_), .A1(new_n5224_), .B0(new_n14414_), .Y(new_n14415_));
  OR2X1    g11979(.A(new_n14415_), .B(pi0698), .Y(new_n14416_));
  OAI21X1  g11980(.A0(new_n14416_), .A1(new_n14409_), .B0(new_n3129_), .Y(new_n14417_));
  AOI21X1  g11981(.A0(new_n14345_), .A1(pi0698), .B0(new_n14417_), .Y(new_n14418_));
  AOI21X1  g11982(.A0(new_n3810_), .A1(pi0145), .B0(new_n14418_), .Y(new_n14419_));
  OAI21X1  g11983(.A0(new_n14347_), .A1(new_n12493_), .B0(new_n12494_), .Y(new_n14420_));
  AOI21X1  g11984(.A0(new_n14419_), .A1(new_n12493_), .B0(new_n14420_), .Y(new_n14421_));
  NAND2X1  g11985(.A(new_n14313_), .B(new_n12584_), .Y(new_n14422_));
  OAI21X1  g11986(.A0(new_n14347_), .A1(pi0625), .B0(pi1153), .Y(new_n14423_));
  AOI21X1  g11987(.A0(new_n14419_), .A1(pi0625), .B0(new_n14423_), .Y(new_n14424_));
  NAND2X1  g11988(.A(new_n14315_), .B(pi0608), .Y(new_n14425_));
  OAI22X1  g11989(.A0(new_n14425_), .A1(new_n14424_), .B0(new_n14422_), .B1(new_n14421_), .Y(new_n14426_));
  AND2X1   g11990(.A(new_n14419_), .B(new_n11889_), .Y(new_n14427_));
  AOI21X1  g11991(.A0(new_n14426_), .A1(pi0778), .B0(new_n14427_), .Y(new_n14428_));
  AOI21X1  g11992(.A0(new_n14317_), .A1(pi0609), .B0(pi1155), .Y(new_n14429_));
  OAI21X1  g11993(.A0(new_n14428_), .A1(pi0609), .B0(new_n14429_), .Y(new_n14430_));
  AND2X1   g11994(.A(new_n14351_), .B(new_n12596_), .Y(new_n14431_));
  AOI21X1  g11995(.A0(new_n14317_), .A1(new_n12590_), .B0(new_n12591_), .Y(new_n14432_));
  OAI21X1  g11996(.A0(new_n14428_), .A1(new_n12590_), .B0(new_n14432_), .Y(new_n14433_));
  AND2X1   g11997(.A(new_n14353_), .B(pi0660), .Y(new_n14434_));
  AOI22X1  g11998(.A0(new_n14434_), .A1(new_n14433_), .B0(new_n14431_), .B1(new_n14430_), .Y(new_n14435_));
  MX2X1    g11999(.A(new_n14435_), .B(new_n14428_), .S0(new_n11888_), .Y(new_n14436_));
  AOI21X1  g12000(.A0(new_n14318_), .A1(pi0618), .B0(pi1154), .Y(new_n14437_));
  OAI21X1  g12001(.A0(new_n14436_), .A1(pi0618), .B0(new_n14437_), .Y(new_n14438_));
  AND2X1   g12002(.A(new_n14357_), .B(new_n12622_), .Y(new_n14439_));
  AOI21X1  g12003(.A0(new_n14318_), .A1(new_n12614_), .B0(new_n12615_), .Y(new_n14440_));
  OAI21X1  g12004(.A0(new_n14436_), .A1(new_n12614_), .B0(new_n14440_), .Y(new_n14441_));
  AND2X1   g12005(.A(new_n14359_), .B(pi0627), .Y(new_n14442_));
  AOI22X1  g12006(.A0(new_n14442_), .A1(new_n14441_), .B0(new_n14439_), .B1(new_n14438_), .Y(new_n14443_));
  OR2X1    g12007(.A(new_n14436_), .B(pi0781), .Y(new_n14444_));
  OAI21X1  g12008(.A0(new_n14443_), .A1(new_n11887_), .B0(new_n14444_), .Y(new_n14445_));
  NAND2X1  g12009(.A(new_n14445_), .B(new_n12637_), .Y(new_n14446_));
  AOI21X1  g12010(.A0(new_n14319_), .A1(pi0619), .B0(pi1159), .Y(new_n14447_));
  NAND2X1  g12011(.A(new_n14364_), .B(new_n12645_), .Y(new_n14448_));
  AOI21X1  g12012(.A0(new_n14447_), .A1(new_n14446_), .B0(new_n14448_), .Y(new_n14449_));
  NAND2X1  g12013(.A(new_n14445_), .B(pi0619), .Y(new_n14450_));
  AOI21X1  g12014(.A0(new_n14319_), .A1(new_n12637_), .B0(new_n12638_), .Y(new_n14451_));
  NAND2X1  g12015(.A(new_n14366_), .B(pi0648), .Y(new_n14452_));
  AOI21X1  g12016(.A0(new_n14451_), .A1(new_n14450_), .B0(new_n14452_), .Y(new_n14453_));
  NOR3X1   g12017(.A(new_n14453_), .B(new_n14449_), .C(new_n11886_), .Y(new_n14454_));
  OAI21X1  g12018(.A0(new_n14445_), .A1(pi0789), .B0(new_n12842_), .Y(new_n14455_));
  OR2X1    g12019(.A(new_n14455_), .B(new_n14454_), .Y(new_n14456_));
  NAND3X1  g12020(.A(new_n14373_), .B(new_n14371_), .C(new_n13537_), .Y(new_n14457_));
  OAI21X1  g12021(.A0(new_n14321_), .A1(new_n12770_), .B0(new_n14457_), .Y(new_n14458_));
  AOI21X1  g12022(.A0(new_n14458_), .A1(pi0788), .B0(new_n14273_), .Y(new_n14459_));
  AOI22X1  g12023(.A0(new_n14459_), .A1(new_n14456_), .B0(new_n14397_), .B1(pi0792), .Y(new_n14460_));
  OAI22X1  g12024(.A0(new_n14460_), .A1(new_n14269_), .B0(new_n14391_), .B1(new_n11883_), .Y(new_n14461_));
  NOR2X1   g12025(.A(new_n14461_), .B(pi0644), .Y(new_n14462_));
  OAI21X1  g12026(.A0(new_n14334_), .A1(new_n12743_), .B0(new_n12739_), .Y(new_n14463_));
  AOI21X1  g12027(.A0(new_n14303_), .A1(pi0644), .B0(new_n12739_), .Y(new_n14464_));
  OAI21X1  g12028(.A0(new_n14378_), .A1(pi0644), .B0(new_n14464_), .Y(new_n14465_));
  AND2X1   g12029(.A(new_n14465_), .B(new_n11882_), .Y(new_n14466_));
  OAI21X1  g12030(.A0(new_n14463_), .A1(new_n14462_), .B0(new_n14466_), .Y(new_n14467_));
  AOI21X1  g12031(.A0(new_n14467_), .A1(new_n14381_), .B0(new_n12897_), .Y(new_n14468_));
  NAND3X1  g12032(.A(new_n14380_), .B(pi1160), .C(pi0644), .Y(new_n14469_));
  AOI21X1  g12033(.A0(new_n14469_), .A1(pi0790), .B0(new_n14461_), .Y(new_n14470_));
  OAI21X1  g12034(.A0(new_n14470_), .A1(new_n14468_), .B0(new_n6520_), .Y(new_n14471_));
  AOI21X1  g12035(.A0(po1038), .A1(new_n5224_), .B0(pi0832), .Y(new_n14472_));
  AOI21X1  g12036(.A0(pi1093), .A1(pi1092), .B0(pi0145), .Y(new_n14473_));
  AOI21X1  g12037(.A0(new_n12178_), .A1(new_n14336_), .B0(new_n14473_), .Y(new_n14474_));
  AOI21X1  g12038(.A0(new_n12601_), .A1(new_n2739_), .B0(new_n14474_), .Y(new_n14475_));
  INVX1    g12039(.A(new_n14474_), .Y(new_n14476_));
  AOI21X1  g12040(.A0(new_n14476_), .A1(new_n12776_), .B0(new_n12591_), .Y(new_n14477_));
  AOI21X1  g12041(.A0(new_n14475_), .A1(new_n12779_), .B0(pi1155), .Y(new_n14478_));
  OAI21X1  g12042(.A0(new_n14478_), .A1(new_n14477_), .B0(pi0785), .Y(new_n14479_));
  OAI21X1  g12043(.A0(new_n14475_), .A1(pi0785), .B0(new_n14479_), .Y(new_n14480_));
  INVX1    g12044(.A(new_n14480_), .Y(new_n14481_));
  AOI21X1  g12045(.A0(new_n14481_), .A1(new_n12785_), .B0(new_n12615_), .Y(new_n14482_));
  AOI21X1  g12046(.A0(new_n14481_), .A1(new_n12788_), .B0(pi1154), .Y(new_n14483_));
  OR2X1    g12047(.A(new_n14483_), .B(new_n14482_), .Y(new_n14484_));
  MX2X1    g12048(.A(new_n14484_), .B(new_n14480_), .S0(new_n11887_), .Y(new_n14485_));
  AOI21X1  g12049(.A0(new_n14473_), .A1(new_n12637_), .B0(new_n12638_), .Y(new_n14486_));
  OAI21X1  g12050(.A0(new_n14485_), .A1(new_n12637_), .B0(new_n14486_), .Y(new_n14487_));
  AOI21X1  g12051(.A0(new_n14473_), .A1(pi0619), .B0(pi1159), .Y(new_n14488_));
  OAI21X1  g12052(.A0(new_n14485_), .A1(pi0619), .B0(new_n14488_), .Y(new_n14489_));
  AOI21X1  g12053(.A0(new_n14489_), .A1(new_n14487_), .B0(new_n11886_), .Y(new_n14490_));
  AOI21X1  g12054(.A0(new_n14485_), .A1(new_n11886_), .B0(new_n14490_), .Y(new_n14491_));
  NAND2X1  g12055(.A(new_n14491_), .B(pi0626), .Y(new_n14492_));
  AOI21X1  g12056(.A0(new_n14473_), .A1(new_n12664_), .B0(new_n12676_), .Y(new_n14493_));
  NAND2X1  g12057(.A(new_n14491_), .B(new_n12664_), .Y(new_n14494_));
  AOI21X1  g12058(.A0(new_n14473_), .A1(pi0626), .B0(pi1158), .Y(new_n14495_));
  AOI22X1  g12059(.A0(new_n14495_), .A1(new_n14494_), .B0(new_n14493_), .B1(new_n14492_), .Y(new_n14496_));
  MX2X1    g12060(.A(new_n14496_), .B(new_n14491_), .S0(new_n11885_), .Y(new_n14497_));
  AND2X1   g12061(.A(new_n14473_), .B(new_n12711_), .Y(new_n14498_));
  AOI21X1  g12062(.A0(new_n14497_), .A1(new_n14123_), .B0(new_n14498_), .Y(new_n14499_));
  AOI21X1  g12063(.A0(new_n12566_), .A1(new_n14306_), .B0(new_n14473_), .Y(new_n14500_));
  AND2X1   g12064(.A(new_n12566_), .B(new_n14306_), .Y(new_n14501_));
  AND2X1   g12065(.A(new_n14501_), .B(new_n12493_), .Y(new_n14502_));
  MX2X1    g12066(.A(new_n14473_), .B(pi0625), .S0(new_n14501_), .Y(new_n14503_));
  NOR2X1   g12067(.A(new_n14473_), .B(pi1153), .Y(new_n14504_));
  INVX1    g12068(.A(new_n14504_), .Y(new_n14505_));
  OAI22X1  g12069(.A0(new_n14505_), .A1(new_n14502_), .B0(new_n14503_), .B1(new_n12494_), .Y(new_n14506_));
  MX2X1    g12070(.A(new_n14506_), .B(new_n14500_), .S0(new_n11889_), .Y(new_n14507_));
  NOR3X1   g12071(.A(new_n14507_), .B(new_n12764_), .C(new_n12762_), .Y(new_n14508_));
  INVX1    g12072(.A(new_n14508_), .Y(new_n14509_));
  NOR4X1   g12073(.A(new_n14509_), .B(new_n12870_), .C(new_n12851_), .D(new_n12765_), .Y(new_n14510_));
  INVX1    g12074(.A(new_n14510_), .Y(new_n14511_));
  AOI21X1  g12075(.A0(new_n14473_), .A1(pi0647), .B0(pi1157), .Y(new_n14512_));
  OAI21X1  g12076(.A0(new_n14511_), .A1(pi0647), .B0(new_n14512_), .Y(new_n14513_));
  MX2X1    g12077(.A(new_n14510_), .B(new_n14473_), .S0(new_n12705_), .Y(new_n14514_));
  OAI22X1  g12078(.A0(new_n14514_), .A1(new_n14387_), .B0(new_n14513_), .B1(new_n12723_), .Y(new_n14515_));
  AOI21X1  g12079(.A0(new_n14499_), .A1(new_n14385_), .B0(new_n14515_), .Y(new_n14516_));
  NOR3X1   g12080(.A(new_n14509_), .B(new_n12770_), .C(new_n12765_), .Y(new_n14517_));
  AOI21X1  g12081(.A0(new_n14496_), .A1(new_n13537_), .B0(new_n14517_), .Y(new_n14518_));
  OR2X1    g12082(.A(new_n14518_), .B(new_n11885_), .Y(new_n14519_));
  NOR2X1   g12083(.A(new_n14500_), .B(new_n12120_), .Y(new_n14520_));
  MX2X1    g12084(.A(new_n14474_), .B(pi0625), .S0(new_n14520_), .Y(new_n14521_));
  OAI21X1  g12085(.A0(new_n14503_), .A1(new_n12494_), .B0(new_n12584_), .Y(new_n14522_));
  AOI21X1  g12086(.A0(new_n14521_), .A1(new_n14504_), .B0(new_n14522_), .Y(new_n14523_));
  AOI21X1  g12087(.A0(new_n14501_), .A1(new_n12493_), .B0(new_n14505_), .Y(new_n14524_));
  NOR3X1   g12088(.A(new_n14500_), .B(new_n12120_), .C(new_n12493_), .Y(new_n14525_));
  NOR3X1   g12089(.A(new_n14525_), .B(new_n14476_), .C(new_n12494_), .Y(new_n14526_));
  NOR3X1   g12090(.A(new_n14526_), .B(new_n14524_), .C(new_n12584_), .Y(new_n14527_));
  OAI21X1  g12091(.A0(new_n14527_), .A1(new_n14523_), .B0(pi0778), .Y(new_n14528_));
  OAI21X1  g12092(.A0(new_n14520_), .A1(new_n14476_), .B0(new_n11889_), .Y(new_n14529_));
  NAND2X1  g12093(.A(new_n14529_), .B(new_n14528_), .Y(new_n14530_));
  OAI21X1  g12094(.A0(new_n14507_), .A1(new_n12590_), .B0(new_n12591_), .Y(new_n14531_));
  AOI21X1  g12095(.A0(new_n14530_), .A1(new_n12590_), .B0(new_n14531_), .Y(new_n14532_));
  NOR3X1   g12096(.A(new_n14532_), .B(new_n14477_), .C(pi0660), .Y(new_n14533_));
  OAI21X1  g12097(.A0(new_n14507_), .A1(pi0609), .B0(pi1155), .Y(new_n14534_));
  AOI21X1  g12098(.A0(new_n14530_), .A1(pi0609), .B0(new_n14534_), .Y(new_n14535_));
  NOR3X1   g12099(.A(new_n14535_), .B(new_n14478_), .C(new_n12596_), .Y(new_n14536_));
  OAI21X1  g12100(.A0(new_n14536_), .A1(new_n14533_), .B0(pi0785), .Y(new_n14537_));
  NAND2X1  g12101(.A(new_n14530_), .B(new_n11888_), .Y(new_n14538_));
  AND2X1   g12102(.A(new_n14538_), .B(new_n14537_), .Y(new_n14539_));
  NOR3X1   g12103(.A(new_n14507_), .B(new_n12762_), .C(new_n12614_), .Y(new_n14540_));
  NOR2X1   g12104(.A(new_n14540_), .B(pi1154), .Y(new_n14541_));
  OAI21X1  g12105(.A0(new_n14539_), .A1(pi0618), .B0(new_n14541_), .Y(new_n14542_));
  NOR2X1   g12106(.A(new_n14482_), .B(pi0627), .Y(new_n14543_));
  NOR3X1   g12107(.A(new_n14507_), .B(new_n12762_), .C(pi0618), .Y(new_n14544_));
  NOR2X1   g12108(.A(new_n14544_), .B(new_n12615_), .Y(new_n14545_));
  OAI21X1  g12109(.A0(new_n14539_), .A1(new_n12614_), .B0(new_n14545_), .Y(new_n14546_));
  NOR2X1   g12110(.A(new_n14483_), .B(new_n12622_), .Y(new_n14547_));
  AOI22X1  g12111(.A0(new_n14547_), .A1(new_n14546_), .B0(new_n14543_), .B1(new_n14542_), .Y(new_n14548_));
  MX2X1    g12112(.A(new_n14548_), .B(new_n14539_), .S0(new_n11887_), .Y(new_n14549_));
  AOI21X1  g12113(.A0(new_n14508_), .A1(pi0619), .B0(pi1159), .Y(new_n14550_));
  OAI21X1  g12114(.A0(new_n14549_), .A1(pi0619), .B0(new_n14550_), .Y(new_n14551_));
  AND2X1   g12115(.A(new_n14487_), .B(new_n12645_), .Y(new_n14552_));
  AND2X1   g12116(.A(new_n14552_), .B(new_n14551_), .Y(new_n14553_));
  AOI21X1  g12117(.A0(new_n14508_), .A1(new_n12637_), .B0(new_n12638_), .Y(new_n14554_));
  OAI21X1  g12118(.A0(new_n14549_), .A1(new_n12637_), .B0(new_n14554_), .Y(new_n14555_));
  AND2X1   g12119(.A(new_n14489_), .B(pi0648), .Y(new_n14556_));
  AOI21X1  g12120(.A0(new_n14556_), .A1(new_n14555_), .B0(new_n11886_), .Y(new_n14557_));
  INVX1    g12121(.A(new_n14557_), .Y(new_n14558_));
  AOI21X1  g12122(.A0(new_n14549_), .A1(new_n11886_), .B0(new_n14264_), .Y(new_n14559_));
  OAI21X1  g12123(.A0(new_n14558_), .A1(new_n14553_), .B0(new_n14559_), .Y(new_n14560_));
  AOI21X1  g12124(.A0(new_n14560_), .A1(new_n14519_), .B0(new_n14273_), .Y(new_n14561_));
  INVX1    g12125(.A(new_n14269_), .Y(new_n14562_));
  NOR3X1   g12126(.A(new_n14509_), .B(new_n12851_), .C(new_n12765_), .Y(new_n14563_));
  AOI21X1  g12127(.A0(new_n2739_), .A1(new_n12683_), .B0(new_n12684_), .Y(new_n14564_));
  AOI22X1  g12128(.A0(new_n14564_), .A1(new_n14563_), .B0(new_n14497_), .B1(new_n12867_), .Y(new_n14565_));
  AOI21X1  g12129(.A0(new_n2739_), .A1(pi0628), .B0(pi1156), .Y(new_n14566_));
  AOI22X1  g12130(.A0(new_n14566_), .A1(new_n14563_), .B0(new_n14497_), .B1(new_n12865_), .Y(new_n14567_));
  MX2X1    g12131(.A(new_n14567_), .B(new_n14565_), .S0(new_n12689_), .Y(new_n14568_));
  OAI21X1  g12132(.A0(new_n14568_), .A1(new_n11884_), .B0(new_n14562_), .Y(new_n14569_));
  OAI22X1  g12133(.A0(new_n14569_), .A1(new_n14561_), .B0(new_n14516_), .B1(new_n11883_), .Y(new_n14570_));
  INVX1    g12134(.A(new_n14570_), .Y(new_n14571_));
  OAI21X1  g12135(.A0(new_n14514_), .A1(new_n12706_), .B0(new_n14513_), .Y(new_n14572_));
  MX2X1    g12136(.A(new_n14572_), .B(new_n14511_), .S0(new_n11883_), .Y(new_n14573_));
  OAI21X1  g12137(.A0(new_n14573_), .A1(pi0644), .B0(pi0715), .Y(new_n14574_));
  AOI21X1  g12138(.A0(new_n14571_), .A1(pi0644), .B0(new_n14574_), .Y(new_n14575_));
  INVX1    g12139(.A(new_n14473_), .Y(new_n14576_));
  MX2X1    g12140(.A(new_n14499_), .B(new_n14576_), .S0(new_n12735_), .Y(new_n14577_));
  AOI21X1  g12141(.A0(new_n14473_), .A1(new_n12743_), .B0(pi0715), .Y(new_n14578_));
  OAI21X1  g12142(.A0(new_n14577_), .A1(new_n12743_), .B0(new_n14578_), .Y(new_n14579_));
  NAND2X1  g12143(.A(new_n14579_), .B(pi1160), .Y(new_n14580_));
  OAI21X1  g12144(.A0(new_n14573_), .A1(new_n12743_), .B0(new_n12739_), .Y(new_n14581_));
  AOI21X1  g12145(.A0(new_n14571_), .A1(new_n12743_), .B0(new_n14581_), .Y(new_n14582_));
  AOI21X1  g12146(.A0(new_n14473_), .A1(pi0644), .B0(new_n12739_), .Y(new_n14583_));
  OAI21X1  g12147(.A0(new_n14577_), .A1(pi0644), .B0(new_n14583_), .Y(new_n14584_));
  NAND2X1  g12148(.A(new_n14584_), .B(new_n11882_), .Y(new_n14585_));
  OAI22X1  g12149(.A0(new_n14585_), .A1(new_n14582_), .B0(new_n14580_), .B1(new_n14575_), .Y(new_n14586_));
  OAI21X1  g12150(.A0(new_n14570_), .A1(pi0790), .B0(pi0832), .Y(new_n14587_));
  AOI21X1  g12151(.A0(new_n14586_), .A1(pi0790), .B0(new_n14587_), .Y(new_n14588_));
  AOI21X1  g12152(.A0(new_n14472_), .A1(new_n14471_), .B0(new_n14588_), .Y(po0302));
  INVX1    g12153(.A(pi0947), .Y(new_n14590_));
  AND2X1   g12154(.A(new_n14590_), .B(pi0907), .Y(new_n14591_));
  AOI22X1  g12155(.A0(new_n14591_), .A1(pi0735), .B0(pi0947), .B1(pi0743), .Y(new_n14592_));
  AND2X1   g12156(.A(new_n14592_), .B(new_n2739_), .Y(new_n14593_));
  NOR2X1   g12157(.A(new_n5069_), .B(pi0907), .Y(new_n14594_));
  NOR3X1   g12158(.A(new_n14594_), .B(new_n12063_), .C(new_n2800_), .Y(new_n14595_));
  NAND3X1  g12159(.A(new_n14594_), .B(new_n12073_), .C(pi0146), .Y(new_n14596_));
  OR4X1    g12160(.A(new_n12062_), .B(new_n12058_), .C(new_n5297_), .D(new_n13294_), .Y(new_n14597_));
  AND2X1   g12161(.A(new_n14597_), .B(new_n14590_), .Y(new_n14598_));
  NAND2X1  g12162(.A(new_n12063_), .B(pi0743), .Y(new_n14599_));
  INVX1    g12163(.A(new_n12063_), .Y(new_n14600_));
  AOI21X1  g12164(.A0(new_n14600_), .A1(pi0146), .B0(new_n14590_), .Y(new_n14601_));
  AOI22X1  g12165(.A0(new_n14601_), .A1(new_n14599_), .B0(new_n14598_), .B1(new_n14596_), .Y(new_n14602_));
  OAI21X1  g12166(.A0(new_n14602_), .A1(new_n14595_), .B0(new_n10137_), .Y(new_n14603_));
  INVX1    g12167(.A(new_n14592_), .Y(new_n14604_));
  MX2X1    g12168(.A(new_n14604_), .B(pi0146), .S0(new_n11953_), .Y(new_n14605_));
  AOI21X1  g12169(.A0(new_n14605_), .A1(new_n10136_), .B0(pi0215), .Y(new_n14606_));
  OR2X1    g12170(.A(new_n12086_), .B(new_n2800_), .Y(new_n14607_));
  AOI21X1  g12171(.A0(new_n14604_), .A1(new_n12082_), .B0(new_n2954_), .Y(new_n14608_));
  AOI22X1  g12172(.A0(new_n14608_), .A1(new_n14607_), .B0(new_n14606_), .B1(new_n14603_), .Y(new_n14609_));
  NOR3X1   g12173(.A(new_n14592_), .B(new_n12062_), .C(new_n12058_), .Y(new_n14610_));
  OAI21X1  g12174(.A0(new_n12063_), .A1(new_n2800_), .B0(new_n5051_), .Y(new_n14611_));
  AND2X1   g12175(.A(new_n14604_), .B(new_n12055_), .Y(new_n14612_));
  OAI21X1  g12176(.A0(new_n12055_), .A1(new_n2800_), .B0(new_n5050_), .Y(new_n14613_));
  OAI22X1  g12177(.A0(new_n14613_), .A1(new_n14612_), .B0(new_n14611_), .B1(new_n14610_), .Y(new_n14614_));
  OAI21X1  g12178(.A0(new_n14605_), .A1(new_n2971_), .B0(new_n2964_), .Y(new_n14615_));
  AOI21X1  g12179(.A0(new_n14614_), .A1(new_n2971_), .B0(new_n14615_), .Y(new_n14616_));
  MX2X1    g12180(.A(pi0146), .B(new_n14604_), .S0(new_n12082_), .Y(new_n14617_));
  OAI21X1  g12181(.A0(new_n12008_), .A1(new_n11992_), .B0(new_n2800_), .Y(new_n14618_));
  AOI21X1  g12182(.A0(new_n14592_), .A1(new_n12084_), .B0(new_n5051_), .Y(new_n14619_));
  AOI22X1  g12183(.A0(new_n14619_), .A1(new_n14618_), .B0(new_n14617_), .B1(new_n5051_), .Y(new_n14620_));
  OAI21X1  g12184(.A0(new_n14620_), .A1(new_n2964_), .B0(new_n2953_), .Y(new_n14621_));
  OAI22X1  g12185(.A0(new_n14621_), .A1(new_n14616_), .B0(new_n14609_), .B1(new_n2953_), .Y(new_n14622_));
  OAI21X1  g12186(.A0(new_n14604_), .A1(new_n12091_), .B0(pi0299), .Y(new_n14623_));
  AOI21X1  g12187(.A0(new_n12091_), .A1(new_n2800_), .B0(new_n14623_), .Y(new_n14624_));
  AOI21X1  g12188(.A0(new_n11945_), .A1(new_n11944_), .B0(pi0146), .Y(new_n14625_));
  OAI21X1  g12189(.A0(new_n14604_), .A1(new_n12445_), .B0(new_n2953_), .Y(new_n14626_));
  OAI21X1  g12190(.A0(new_n14626_), .A1(new_n14625_), .B0(new_n2959_), .Y(new_n14627_));
  OAI21X1  g12191(.A0(new_n14627_), .A1(new_n14624_), .B0(new_n2996_), .Y(new_n14628_));
  AOI21X1  g12192(.A0(new_n14622_), .A1(pi0039), .B0(new_n14628_), .Y(new_n14629_));
  OR2X1    g12193(.A(new_n12202_), .B(pi0146), .Y(new_n14630_));
  AOI21X1  g12194(.A0(new_n14593_), .A1(new_n6857_), .B0(new_n2996_), .Y(new_n14631_));
  AND2X1   g12195(.A(new_n14631_), .B(new_n14630_), .Y(new_n14632_));
  NOR3X1   g12196(.A(new_n14632_), .B(new_n14629_), .C(new_n9580_), .Y(new_n14633_));
  OAI21X1  g12197(.A0(new_n7686_), .A1(pi0146), .B0(new_n12898_), .Y(new_n14634_));
  OAI21X1  g12198(.A0(new_n2739_), .A1(pi0146), .B0(pi0832), .Y(new_n14635_));
  OAI22X1  g12199(.A0(new_n14635_), .A1(new_n14593_), .B0(new_n14634_), .B1(new_n14633_), .Y(po0303));
  INVX1    g12200(.A(pi0726), .Y(new_n14637_));
  INVX1    g12201(.A(new_n14591_), .Y(new_n14638_));
  OAI22X1  g12202(.A0(new_n14638_), .A1(new_n14637_), .B0(new_n14590_), .B1(pi0770), .Y(new_n14639_));
  OAI21X1  g12203(.A0(new_n2739_), .A1(pi0147), .B0(pi0832), .Y(new_n14640_));
  AOI21X1  g12204(.A0(new_n14639_), .A1(new_n2739_), .B0(new_n14640_), .Y(new_n14641_));
  AOI21X1  g12205(.A0(new_n11947_), .A1(new_n14590_), .B0(pi0039), .Y(new_n14642_));
  NOR4X1   g12206(.A(new_n12067_), .B(new_n12011_), .C(new_n14590_), .D(pi0299), .Y(new_n14643_));
  INVX1    g12207(.A(new_n14643_), .Y(new_n14644_));
  NOR4X1   g12208(.A(new_n11952_), .B(new_n10137_), .C(new_n2740_), .D(pi0947), .Y(new_n14645_));
  AOI21X1  g12209(.A0(new_n14591_), .A1(new_n12063_), .B0(new_n12075_), .Y(new_n14646_));
  NOR2X1   g12210(.A(new_n14646_), .B(new_n10136_), .Y(new_n14647_));
  NOR3X1   g12211(.A(new_n14647_), .B(new_n14645_), .C(pi0215), .Y(new_n14648_));
  OR2X1    g12212(.A(new_n12085_), .B(new_n12083_), .Y(new_n14649_));
  AND2X1   g12213(.A(new_n14649_), .B(pi0215), .Y(new_n14650_));
  OR4X1    g12214(.A(new_n11990_), .B(new_n11975_), .C(pi0947), .D(new_n5297_), .Y(new_n14651_));
  AND2X1   g12215(.A(new_n14651_), .B(new_n14650_), .Y(new_n14652_));
  OAI21X1  g12216(.A0(new_n14652_), .A1(new_n14648_), .B0(pi0299), .Y(new_n14653_));
  AND2X1   g12217(.A(new_n14653_), .B(new_n12068_), .Y(new_n14654_));
  AOI21X1  g12218(.A0(new_n14654_), .A1(new_n14644_), .B0(new_n2959_), .Y(new_n14655_));
  NOR3X1   g12219(.A(new_n14655_), .B(new_n14642_), .C(pi0038), .Y(new_n14656_));
  NOR4X1   g12220(.A(new_n4996_), .B(new_n2740_), .C(pi0947), .D(new_n2996_), .Y(new_n14657_));
  NOR2X1   g12221(.A(new_n14657_), .B(new_n14656_), .Y(new_n14658_));
  MX2X1    g12222(.A(new_n14658_), .B(new_n12574_), .S0(pi0770), .Y(new_n14659_));
  NOR2X1   g12223(.A(new_n14657_), .B(new_n13402_), .Y(new_n14660_));
  AOI21X1  g12224(.A0(new_n11947_), .A1(pi0947), .B0(pi0039), .Y(new_n14661_));
  NOR3X1   g12225(.A(new_n12067_), .B(new_n12011_), .C(new_n14590_), .Y(new_n14662_));
  NOR2X1   g12226(.A(new_n14662_), .B(pi0299), .Y(new_n14663_));
  INVX1    g12227(.A(new_n14663_), .Y(new_n14664_));
  NOR4X1   g12228(.A(new_n11990_), .B(new_n11975_), .C(new_n14590_), .D(new_n2954_), .Y(new_n14665_));
  INVX1    g12229(.A(new_n14665_), .Y(new_n14666_));
  NOR3X1   g12230(.A(new_n12062_), .B(new_n12058_), .C(new_n14590_), .Y(new_n14667_));
  OR4X1    g12231(.A(new_n11952_), .B(new_n2756_), .C(new_n2755_), .D(new_n14590_), .Y(new_n14668_));
  AOI21X1  g12232(.A0(new_n14668_), .A1(new_n10136_), .B0(pi0215), .Y(new_n14669_));
  OAI21X1  g12233(.A0(new_n14667_), .A1(new_n10136_), .B0(new_n14669_), .Y(new_n14670_));
  NAND3X1  g12234(.A(new_n14670_), .B(new_n14666_), .C(pi0299), .Y(new_n14671_));
  AND2X1   g12235(.A(new_n14671_), .B(new_n14664_), .Y(new_n14672_));
  INVX1    g12236(.A(new_n14672_), .Y(new_n14673_));
  AOI21X1  g12237(.A0(new_n14673_), .A1(pi0039), .B0(new_n14661_), .Y(new_n14674_));
  OAI21X1  g12238(.A0(new_n14674_), .A1(pi0038), .B0(new_n14660_), .Y(new_n14675_));
  OR2X1    g12239(.A(pi0770), .B(new_n8710_), .Y(new_n14676_));
  OAI21X1  g12240(.A0(new_n14676_), .A1(new_n14675_), .B0(new_n14637_), .Y(new_n14677_));
  AOI21X1  g12241(.A0(new_n14659_), .A1(new_n8710_), .B0(new_n14677_), .Y(new_n14678_));
  OR4X1    g12242(.A(new_n14591_), .B(new_n11952_), .C(new_n10137_), .D(new_n2740_), .Y(new_n14679_));
  OR2X1    g12243(.A(new_n14667_), .B(new_n12075_), .Y(new_n14680_));
  AOI21X1  g12244(.A0(new_n14680_), .A1(new_n10137_), .B0(pi0215), .Y(new_n14681_));
  AOI21X1  g12245(.A0(new_n14681_), .A1(new_n14679_), .B0(new_n14650_), .Y(new_n14682_));
  NOR2X1   g12246(.A(new_n14682_), .B(new_n2953_), .Y(new_n14683_));
  AOI22X1  g12247(.A0(new_n12065_), .A1(new_n3630_), .B0(new_n12064_), .B1(new_n2971_), .Y(new_n14684_));
  OAI21X1  g12248(.A0(new_n14684_), .A1(new_n5065_), .B0(new_n2964_), .Y(new_n14685_));
  INVX1    g12249(.A(new_n12010_), .Y(new_n14686_));
  AOI21X1  g12250(.A0(new_n14686_), .A1(new_n14590_), .B0(new_n2964_), .Y(new_n14687_));
  AOI21X1  g12251(.A0(new_n14638_), .A1(new_n14686_), .B0(new_n2964_), .Y(new_n14688_));
  NOR2X1   g12252(.A(new_n14688_), .B(new_n14687_), .Y(new_n14689_));
  AOI21X1  g12253(.A0(new_n14689_), .A1(new_n14685_), .B0(pi0299), .Y(new_n14690_));
  AND2X1   g12254(.A(pi0947), .B(pi0299), .Y(new_n14691_));
  OR2X1    g12255(.A(new_n14691_), .B(new_n14690_), .Y(new_n14692_));
  NOR2X1   g12256(.A(new_n14692_), .B(new_n14683_), .Y(new_n14693_));
  AOI21X1  g12257(.A0(new_n11947_), .A1(new_n5065_), .B0(pi0039), .Y(new_n14694_));
  AOI22X1  g12258(.A0(new_n14694_), .A1(new_n11947_), .B0(new_n14693_), .B1(pi0039), .Y(new_n14695_));
  INVX1    g12259(.A(new_n14695_), .Y(new_n14696_));
  AND2X1   g12260(.A(new_n11947_), .B(new_n5065_), .Y(new_n14697_));
  OR4X1    g12261(.A(new_n12067_), .B(new_n12011_), .C(new_n5064_), .D(pi0299), .Y(new_n14698_));
  AOI21X1  g12262(.A0(new_n12082_), .A1(new_n5065_), .B0(new_n2954_), .Y(new_n14699_));
  OR4X1    g12263(.A(new_n11952_), .B(new_n5064_), .C(new_n2756_), .D(new_n2755_), .Y(new_n14700_));
  OAI21X1  g12264(.A0(new_n14700_), .A1(new_n10137_), .B0(new_n2954_), .Y(new_n14701_));
  OAI21X1  g12265(.A0(new_n14701_), .A1(new_n12076_), .B0(pi0299), .Y(new_n14702_));
  OAI21X1  g12266(.A0(new_n14702_), .A1(new_n14699_), .B0(new_n14698_), .Y(new_n14703_));
  MX2X1    g12267(.A(new_n14703_), .B(new_n14697_), .S0(new_n2959_), .Y(new_n14704_));
  AOI21X1  g12268(.A0(new_n14704_), .A1(pi0147), .B0(pi0038), .Y(new_n14705_));
  OAI21X1  g12269(.A0(new_n14696_), .A1(pi0147), .B0(new_n14705_), .Y(new_n14706_));
  INVX1    g12270(.A(pi0770), .Y(new_n14707_));
  NOR4X1   g12271(.A(new_n5065_), .B(new_n3015_), .C(new_n2740_), .D(pi0039), .Y(new_n14708_));
  AOI21X1  g12272(.A0(new_n12202_), .A1(new_n5065_), .B0(new_n2996_), .Y(new_n14709_));
  OAI21X1  g12273(.A0(new_n14708_), .A1(pi0147), .B0(new_n14709_), .Y(new_n14710_));
  AND2X1   g12274(.A(new_n14710_), .B(new_n14707_), .Y(new_n14711_));
  NOR2X1   g12275(.A(new_n14682_), .B(new_n14665_), .Y(new_n14712_));
  OR4X1    g12276(.A(new_n14591_), .B(new_n12067_), .C(new_n12011_), .D(pi0299), .Y(new_n14713_));
  OAI21X1  g12277(.A0(new_n14712_), .A1(new_n2953_), .B0(new_n14713_), .Y(new_n14714_));
  AND2X1   g12278(.A(new_n14638_), .B(new_n11947_), .Y(new_n14715_));
  MX2X1    g12279(.A(new_n14715_), .B(new_n14714_), .S0(pi0039), .Y(new_n14716_));
  INVX1    g12280(.A(new_n14716_), .Y(new_n14717_));
  NAND2X1  g12281(.A(new_n14651_), .B(pi0215), .Y(new_n14718_));
  AOI21X1  g12282(.A0(new_n14591_), .A1(new_n12063_), .B0(new_n10136_), .Y(new_n14719_));
  NOR4X1   g12283(.A(new_n11952_), .B(new_n2740_), .C(pi0947), .D(new_n5297_), .Y(new_n14720_));
  NOR2X1   g12284(.A(new_n14720_), .B(new_n10137_), .Y(new_n14721_));
  OAI21X1  g12285(.A0(new_n14721_), .A1(new_n14719_), .B0(new_n2954_), .Y(new_n14722_));
  AOI21X1  g12286(.A0(new_n14722_), .A1(new_n14718_), .B0(new_n2953_), .Y(new_n14723_));
  NOR3X1   g12287(.A(new_n14638_), .B(new_n12067_), .C(new_n12011_), .Y(new_n14724_));
  NOR2X1   g12288(.A(new_n14724_), .B(pi0299), .Y(new_n14725_));
  NOR2X1   g12289(.A(new_n14725_), .B(new_n14723_), .Y(new_n14726_));
  AND2X1   g12290(.A(new_n14591_), .B(new_n11947_), .Y(new_n14727_));
  MX2X1    g12291(.A(new_n14727_), .B(new_n14726_), .S0(pi0039), .Y(new_n14728_));
  INVX1    g12292(.A(new_n14728_), .Y(new_n14729_));
  OAI21X1  g12293(.A0(new_n14729_), .A1(new_n8710_), .B0(new_n2996_), .Y(new_n14730_));
  AOI21X1  g12294(.A0(new_n14717_), .A1(new_n8710_), .B0(new_n14730_), .Y(new_n14731_));
  AOI21X1  g12295(.A0(new_n14591_), .A1(new_n12202_), .B0(new_n2996_), .Y(new_n14732_));
  OAI21X1  g12296(.A0(new_n12202_), .A1(pi0147), .B0(new_n14732_), .Y(new_n14733_));
  NAND2X1  g12297(.A(new_n14733_), .B(pi0770), .Y(new_n14734_));
  OAI21X1  g12298(.A0(new_n14734_), .A1(new_n14731_), .B0(pi0726), .Y(new_n14735_));
  AOI21X1  g12299(.A0(new_n14711_), .A1(new_n14706_), .B0(new_n14735_), .Y(new_n14736_));
  OR4X1    g12300(.A(new_n14736_), .B(new_n14678_), .C(po1038), .D(new_n3810_), .Y(new_n14737_));
  AOI21X1  g12301(.A0(new_n9580_), .A1(new_n8710_), .B0(pi0832), .Y(new_n14738_));
  AOI21X1  g12302(.A0(new_n14738_), .A1(new_n14737_), .B0(new_n14641_), .Y(po0304));
  NOR2X1   g12303(.A(new_n12067_), .B(new_n12011_), .Y(new_n14740_));
  INVX1    g12304(.A(new_n14740_), .Y(new_n14741_));
  AOI21X1  g12305(.A0(new_n14741_), .A1(new_n2953_), .B0(new_n14723_), .Y(new_n14742_));
  OAI21X1  g12306(.A0(new_n14742_), .A1(new_n4036_), .B0(new_n12911_), .Y(new_n14743_));
  AOI21X1  g12307(.A0(new_n14714_), .A1(new_n11829_), .B0(new_n14743_), .Y(new_n14744_));
  OAI21X1  g12308(.A0(new_n14703_), .A1(new_n4036_), .B0(pi0749), .Y(new_n14745_));
  AOI21X1  g12309(.A0(new_n14693_), .A1(new_n4036_), .B0(new_n14745_), .Y(new_n14746_));
  NOR3X1   g12310(.A(new_n14746_), .B(new_n14744_), .C(new_n2959_), .Y(new_n14747_));
  AOI21X1  g12311(.A0(new_n11948_), .A1(new_n4036_), .B0(pi0039), .Y(new_n14748_));
  INVX1    g12312(.A(new_n14748_), .Y(new_n14749_));
  AND2X1   g12313(.A(pi0947), .B(new_n12911_), .Y(new_n14750_));
  NOR3X1   g12314(.A(new_n14750_), .B(new_n11948_), .C(new_n5064_), .Y(new_n14751_));
  OAI21X1  g12315(.A0(new_n14751_), .A1(new_n14749_), .B0(new_n2996_), .Y(new_n14752_));
  NAND2X1  g12316(.A(new_n12202_), .B(new_n5065_), .Y(new_n14753_));
  OAI22X1  g12317(.A0(new_n14750_), .A1(new_n14753_), .B0(new_n12202_), .B1(pi0148), .Y(new_n14754_));
  AOI21X1  g12318(.A0(new_n14754_), .A1(pi0038), .B0(new_n12934_), .Y(new_n14755_));
  OAI21X1  g12319(.A0(new_n14752_), .A1(new_n14747_), .B0(new_n14755_), .Y(new_n14756_));
  AND2X1   g12320(.A(new_n5117_), .B(new_n3129_), .Y(new_n14757_));
  INVX1    g12321(.A(new_n14757_), .Y(new_n14758_));
  OR2X1    g12322(.A(new_n14652_), .B(new_n14648_), .Y(new_n14759_));
  AND2X1   g12323(.A(new_n14670_), .B(new_n14666_), .Y(new_n14760_));
  OAI21X1  g12324(.A0(new_n14760_), .A1(new_n4036_), .B0(pi0299), .Y(new_n14761_));
  AOI21X1  g12325(.A0(new_n14759_), .A1(new_n4036_), .B0(new_n14761_), .Y(new_n14762_));
  OAI21X1  g12326(.A0(new_n14740_), .A1(pi0148), .B0(new_n14663_), .Y(new_n14763_));
  NAND2X1  g12327(.A(new_n14763_), .B(pi0749), .Y(new_n14764_));
  NOR2X1   g12328(.A(pi0749), .B(pi0148), .Y(new_n14765_));
  AOI21X1  g12329(.A0(new_n14765_), .A1(new_n12089_), .B0(new_n2959_), .Y(new_n14766_));
  OAI21X1  g12330(.A0(new_n14764_), .A1(new_n14762_), .B0(new_n14766_), .Y(new_n14767_));
  NAND2X1  g12331(.A(pi0947), .B(pi0749), .Y(new_n14768_));
  OAI21X1  g12332(.A0(new_n14768_), .A1(new_n11948_), .B0(new_n14748_), .Y(new_n14769_));
  NAND3X1  g12333(.A(new_n14769_), .B(new_n14767_), .C(new_n2996_), .Y(new_n14770_));
  AOI21X1  g12334(.A0(new_n14768_), .A1(new_n12202_), .B0(new_n2996_), .Y(new_n14771_));
  OAI21X1  g12335(.A0(new_n12572_), .A1(new_n4036_), .B0(new_n14771_), .Y(new_n14772_));
  AND2X1   g12336(.A(new_n14772_), .B(new_n12934_), .Y(new_n14773_));
  AOI21X1  g12337(.A0(new_n14773_), .A1(new_n14770_), .B0(new_n14758_), .Y(new_n14774_));
  OAI21X1  g12338(.A0(new_n14757_), .A1(pi0148), .B0(new_n2436_), .Y(new_n14775_));
  AOI21X1  g12339(.A0(new_n14774_), .A1(new_n14756_), .B0(new_n14775_), .Y(new_n14776_));
  OAI21X1  g12340(.A0(new_n4036_), .A1(new_n2436_), .B0(new_n12898_), .Y(new_n14777_));
  NAND2X1  g12341(.A(new_n14768_), .B(new_n2739_), .Y(new_n14778_));
  AOI21X1  g12342(.A0(new_n14591_), .A1(pi0706), .B0(new_n14778_), .Y(new_n14779_));
  OAI21X1  g12343(.A0(new_n2739_), .A1(new_n4036_), .B0(pi0832), .Y(new_n14780_));
  OAI22X1  g12344(.A0(new_n14780_), .A1(new_n14779_), .B0(new_n14777_), .B1(new_n14776_), .Y(po0305));
  INVX1    g12345(.A(pi0755), .Y(new_n14782_));
  AND2X1   g12346(.A(pi0947), .B(new_n14782_), .Y(new_n14783_));
  INVX1    g12347(.A(new_n14783_), .Y(new_n14784_));
  OAI21X1  g12348(.A0(new_n14638_), .A1(pi0725), .B0(new_n14784_), .Y(new_n14785_));
  OAI21X1  g12349(.A0(new_n2739_), .A1(pi0149), .B0(pi0832), .Y(new_n14786_));
  AOI21X1  g12350(.A0(new_n14785_), .A1(new_n2739_), .B0(new_n14786_), .Y(new_n14787_));
  INVX1    g12351(.A(pi0725), .Y(new_n14788_));
  AOI21X1  g12352(.A0(new_n14784_), .A1(new_n12202_), .B0(new_n2996_), .Y(new_n14789_));
  OAI21X1  g12353(.A0(new_n12572_), .A1(new_n7129_), .B0(new_n14789_), .Y(new_n14790_));
  OR2X1    g12354(.A(new_n2953_), .B(pi0149), .Y(new_n14791_));
  AOI22X1  g12355(.A0(new_n14671_), .A1(new_n14791_), .B0(new_n14759_), .B1(new_n7129_), .Y(new_n14792_));
  OAI21X1  g12356(.A0(new_n14740_), .A1(pi0149), .B0(new_n14663_), .Y(new_n14793_));
  NAND2X1  g12357(.A(new_n14793_), .B(new_n14782_), .Y(new_n14794_));
  AND2X1   g12358(.A(pi0755), .B(new_n7129_), .Y(new_n14795_));
  AOI21X1  g12359(.A0(new_n14795_), .A1(new_n12089_), .B0(new_n2959_), .Y(new_n14796_));
  OAI21X1  g12360(.A0(new_n14794_), .A1(new_n14792_), .B0(new_n14796_), .Y(new_n14797_));
  AOI21X1  g12361(.A0(new_n14783_), .A1(new_n11947_), .B0(pi0039), .Y(new_n14798_));
  OAI21X1  g12362(.A0(new_n11947_), .A1(pi0149), .B0(new_n14798_), .Y(new_n14799_));
  NAND3X1  g12363(.A(new_n14799_), .B(new_n14797_), .C(new_n2996_), .Y(new_n14800_));
  AOI21X1  g12364(.A0(new_n14800_), .A1(new_n14790_), .B0(new_n14788_), .Y(new_n14801_));
  OAI21X1  g12365(.A0(new_n14703_), .A1(new_n7129_), .B0(new_n14782_), .Y(new_n14802_));
  AOI21X1  g12366(.A0(new_n14693_), .A1(new_n7129_), .B0(new_n14802_), .Y(new_n14803_));
  NOR3X1   g12367(.A(new_n14712_), .B(new_n2953_), .C(pi0149), .Y(new_n14804_));
  AND2X1   g12368(.A(new_n14713_), .B(pi0755), .Y(new_n14805_));
  OAI21X1  g12369(.A0(new_n14742_), .A1(new_n7129_), .B0(new_n14805_), .Y(new_n14806_));
  OAI21X1  g12370(.A0(new_n14806_), .A1(new_n14804_), .B0(pi0039), .Y(new_n14807_));
  OAI22X1  g12371(.A0(new_n14807_), .A1(new_n14803_), .B0(new_n14799_), .B1(new_n14727_), .Y(new_n14808_));
  NOR2X1   g12372(.A(new_n12202_), .B(pi0149), .Y(new_n14809_));
  NOR4X1   g12373(.A(new_n5064_), .B(new_n3003_), .C(new_n2740_), .D(new_n2555_), .Y(new_n14810_));
  INVX1    g12374(.A(new_n14810_), .Y(new_n14811_));
  OAI21X1  g12375(.A0(new_n14590_), .A1(new_n14782_), .B0(new_n2959_), .Y(new_n14812_));
  OAI21X1  g12376(.A0(new_n14812_), .A1(new_n14811_), .B0(pi0038), .Y(new_n14813_));
  OAI21X1  g12377(.A0(new_n14813_), .A1(new_n14809_), .B0(new_n14788_), .Y(new_n14814_));
  AOI21X1  g12378(.A0(new_n14808_), .A1(new_n2996_), .B0(new_n14814_), .Y(new_n14815_));
  OAI21X1  g12379(.A0(new_n14815_), .A1(new_n14801_), .B0(new_n7686_), .Y(new_n14816_));
  AOI21X1  g12380(.A0(new_n9580_), .A1(new_n7129_), .B0(pi0832), .Y(new_n14817_));
  AOI21X1  g12381(.A0(new_n14817_), .A1(new_n14816_), .B0(new_n14787_), .Y(po0306));
  AND2X1   g12382(.A(new_n14654_), .B(new_n14644_), .Y(new_n14819_));
  INVX1    g12383(.A(pi0751), .Y(new_n14820_));
  OAI21X1  g12384(.A0(new_n14672_), .A1(new_n9936_), .B0(new_n14820_), .Y(new_n14821_));
  AOI21X1  g12385(.A0(new_n14819_), .A1(new_n9936_), .B0(new_n14821_), .Y(new_n14822_));
  AND2X1   g12386(.A(new_n12088_), .B(new_n12068_), .Y(new_n14823_));
  NOR3X1   g12387(.A(new_n14823_), .B(new_n14820_), .C(pi0150), .Y(new_n14824_));
  OAI21X1  g12388(.A0(new_n14824_), .A1(new_n14822_), .B0(pi0039), .Y(new_n14825_));
  MX2X1    g12389(.A(new_n9936_), .B(new_n14820_), .S0(new_n11947_), .Y(new_n14826_));
  AOI21X1  g12390(.A0(new_n14826_), .A1(new_n14642_), .B0(pi0038), .Y(new_n14827_));
  OR2X1    g12391(.A(new_n14590_), .B(pi0751), .Y(new_n14828_));
  AOI22X1  g12392(.A0(new_n14828_), .A1(new_n12202_), .B0(new_n12573_), .B1(pi0150), .Y(new_n14829_));
  OAI21X1  g12393(.A0(new_n14829_), .A1(new_n2996_), .B0(pi0701), .Y(new_n14830_));
  AOI21X1  g12394(.A0(new_n14827_), .A1(new_n14825_), .B0(new_n14830_), .Y(new_n14831_));
  OAI21X1  g12395(.A0(new_n14726_), .A1(new_n9936_), .B0(pi0751), .Y(new_n14832_));
  AOI21X1  g12396(.A0(new_n14714_), .A1(new_n9936_), .B0(new_n14832_), .Y(new_n14833_));
  OAI21X1  g12397(.A0(new_n14703_), .A1(new_n9936_), .B0(new_n14820_), .Y(new_n14834_));
  AOI21X1  g12398(.A0(new_n14693_), .A1(new_n9936_), .B0(new_n14834_), .Y(new_n14835_));
  OAI21X1  g12399(.A0(new_n14835_), .A1(new_n14833_), .B0(pi0039), .Y(new_n14836_));
  NAND3X1  g12400(.A(new_n14828_), .B(new_n14638_), .C(new_n11947_), .Y(new_n14837_));
  AOI21X1  g12401(.A0(new_n11948_), .A1(pi0150), .B0(pi0039), .Y(new_n14838_));
  AOI21X1  g12402(.A0(new_n14838_), .A1(new_n14837_), .B0(pi0038), .Y(new_n14839_));
  INVX1    g12403(.A(pi0701), .Y(new_n14840_));
  NOR2X1   g12404(.A(new_n12202_), .B(pi0150), .Y(new_n14841_));
  OAI21X1  g12405(.A0(new_n14590_), .A1(new_n14820_), .B0(new_n2959_), .Y(new_n14842_));
  OAI21X1  g12406(.A0(new_n14842_), .A1(new_n14811_), .B0(pi0038), .Y(new_n14843_));
  OAI21X1  g12407(.A0(new_n14843_), .A1(new_n14841_), .B0(new_n14840_), .Y(new_n14844_));
  AOI21X1  g12408(.A0(new_n14839_), .A1(new_n14836_), .B0(new_n14844_), .Y(new_n14845_));
  OAI21X1  g12409(.A0(new_n14845_), .A1(new_n14831_), .B0(new_n7686_), .Y(new_n14846_));
  AOI21X1  g12410(.A0(new_n9580_), .A1(new_n9936_), .B0(pi0832), .Y(new_n14847_));
  OAI21X1  g12411(.A0(new_n14638_), .A1(pi0701), .B0(new_n14828_), .Y(new_n14848_));
  OAI21X1  g12412(.A0(new_n2739_), .A1(pi0150), .B0(pi0832), .Y(new_n14849_));
  AOI21X1  g12413(.A0(new_n14848_), .A1(new_n2739_), .B0(new_n14849_), .Y(new_n14850_));
  AOI21X1  g12414(.A0(new_n14847_), .A1(new_n14846_), .B0(new_n14850_), .Y(po0307));
  OR2X1    g12415(.A(new_n14590_), .B(pi0745), .Y(new_n14852_));
  OAI21X1  g12416(.A0(new_n14638_), .A1(pi0723), .B0(new_n14852_), .Y(new_n14853_));
  OAI21X1  g12417(.A0(new_n2739_), .A1(pi0151), .B0(pi0832), .Y(new_n14854_));
  AOI21X1  g12418(.A0(new_n14853_), .A1(new_n2739_), .B0(new_n14854_), .Y(new_n14855_));
  AOI21X1  g12419(.A0(new_n14591_), .A1(new_n11947_), .B0(pi0039), .Y(new_n14856_));
  INVX1    g12420(.A(new_n14856_), .Y(new_n14857_));
  INVX1    g12421(.A(pi0745), .Y(new_n14858_));
  NAND3X1  g12422(.A(new_n11947_), .B(pi0947), .C(new_n14858_), .Y(new_n14859_));
  OAI21X1  g12423(.A0(new_n11947_), .A1(pi0151), .B0(new_n14859_), .Y(new_n14860_));
  INVX1    g12424(.A(new_n12081_), .Y(new_n14861_));
  AND2X1   g12425(.A(new_n14651_), .B(new_n14649_), .Y(new_n14862_));
  AOI21X1  g12426(.A0(new_n14862_), .A1(new_n3325_), .B0(new_n14861_), .Y(new_n14863_));
  NOR2X1   g12427(.A(new_n14863_), .B(new_n2954_), .Y(new_n14864_));
  NOR3X1   g12428(.A(new_n12062_), .B(new_n12058_), .C(new_n5064_), .Y(new_n14865_));
  INVX1    g12429(.A(new_n14865_), .Y(new_n14866_));
  NOR2X1   g12430(.A(new_n10136_), .B(new_n3325_), .Y(new_n14867_));
  AOI22X1  g12431(.A0(new_n14867_), .A1(new_n14866_), .B0(new_n12075_), .B1(new_n10137_), .Y(new_n14868_));
  OAI21X1  g12432(.A0(new_n11952_), .A1(new_n2740_), .B0(new_n3325_), .Y(new_n14869_));
  AND2X1   g12433(.A(new_n14869_), .B(new_n14721_), .Y(new_n14870_));
  AOI21X1  g12434(.A0(new_n14870_), .A1(new_n14700_), .B0(pi0215), .Y(new_n14871_));
  AOI21X1  g12435(.A0(new_n14871_), .A1(new_n14868_), .B0(new_n14864_), .Y(new_n14872_));
  NOR3X1   g12436(.A(new_n12067_), .B(new_n12011_), .C(new_n5064_), .Y(new_n14873_));
  OAI21X1  g12437(.A0(new_n14873_), .A1(new_n3325_), .B0(new_n14690_), .Y(new_n14874_));
  OAI21X1  g12438(.A0(new_n14872_), .A1(new_n2953_), .B0(new_n14874_), .Y(new_n14875_));
  AND2X1   g12439(.A(new_n14875_), .B(new_n14858_), .Y(new_n14876_));
  AND2X1   g12440(.A(new_n14680_), .B(new_n10137_), .Y(new_n14877_));
  INVX1    g12441(.A(new_n14868_), .Y(new_n14878_));
  NOR4X1   g12442(.A(new_n14870_), .B(new_n14878_), .C(new_n14877_), .D(pi0215), .Y(new_n14879_));
  OAI21X1  g12443(.A0(new_n14879_), .A1(new_n14864_), .B0(new_n14666_), .Y(new_n14880_));
  AND2X1   g12444(.A(new_n14880_), .B(pi0299), .Y(new_n14881_));
  OAI21X1  g12445(.A0(new_n14740_), .A1(pi0151), .B0(new_n14725_), .Y(new_n14882_));
  NAND2X1  g12446(.A(new_n14882_), .B(pi0745), .Y(new_n14883_));
  OAI21X1  g12447(.A0(new_n14883_), .A1(new_n14881_), .B0(pi0039), .Y(new_n14884_));
  OAI22X1  g12448(.A0(new_n14884_), .A1(new_n14876_), .B0(new_n14860_), .B1(new_n14857_), .Y(new_n14885_));
  INVX1    g12449(.A(pi0723), .Y(new_n14886_));
  NOR2X1   g12450(.A(new_n12202_), .B(pi0151), .Y(new_n14887_));
  OAI21X1  g12451(.A0(new_n14590_), .A1(new_n14858_), .B0(new_n2959_), .Y(new_n14888_));
  OAI21X1  g12452(.A0(new_n14888_), .A1(new_n14811_), .B0(pi0038), .Y(new_n14889_));
  OAI21X1  g12453(.A0(new_n14889_), .A1(new_n14887_), .B0(new_n14886_), .Y(new_n14890_));
  AOI21X1  g12454(.A0(new_n14885_), .A1(new_n2996_), .B0(new_n14890_), .Y(new_n14891_));
  AND2X1   g12455(.A(new_n12068_), .B(new_n14858_), .Y(new_n14892_));
  NOR3X1   g12456(.A(new_n14892_), .B(new_n14823_), .C(pi0151), .Y(new_n14893_));
  NOR2X1   g12457(.A(new_n14647_), .B(pi0215), .Y(new_n14894_));
  AND2X1   g12458(.A(new_n14668_), .B(new_n10136_), .Y(new_n14895_));
  AOI21X1  g12459(.A0(new_n14869_), .A1(new_n14895_), .B0(new_n14878_), .Y(new_n14896_));
  OAI21X1  g12460(.A0(new_n14863_), .A1(new_n14718_), .B0(pi0299), .Y(new_n14897_));
  AOI21X1  g12461(.A0(new_n14896_), .A1(new_n14894_), .B0(new_n14897_), .Y(new_n14898_));
  NOR3X1   g12462(.A(new_n14898_), .B(new_n14663_), .C(pi0745), .Y(new_n14899_));
  OAI21X1  g12463(.A0(new_n14899_), .A1(new_n14893_), .B0(pi0039), .Y(new_n14900_));
  AOI21X1  g12464(.A0(new_n14860_), .A1(new_n2959_), .B0(pi0038), .Y(new_n14901_));
  AOI22X1  g12465(.A0(new_n14852_), .A1(new_n12202_), .B0(new_n12573_), .B1(pi0151), .Y(new_n14902_));
  OAI21X1  g12466(.A0(new_n14902_), .A1(new_n2996_), .B0(pi0723), .Y(new_n14903_));
  AOI21X1  g12467(.A0(new_n14901_), .A1(new_n14900_), .B0(new_n14903_), .Y(new_n14904_));
  OAI21X1  g12468(.A0(new_n14904_), .A1(new_n14891_), .B0(new_n7686_), .Y(new_n14905_));
  AOI21X1  g12469(.A0(new_n9580_), .A1(new_n3325_), .B0(pi0832), .Y(new_n14906_));
  AOI21X1  g12470(.A0(new_n14906_), .A1(new_n14905_), .B0(new_n14855_), .Y(po0308));
  INVX1    g12471(.A(pi0759), .Y(new_n14908_));
  MX2X1    g12472(.A(new_n5064_), .B(new_n6900_), .S0(new_n11953_), .Y(new_n14909_));
  AOI21X1  g12473(.A0(new_n14909_), .A1(new_n10136_), .B0(pi0215), .Y(new_n14910_));
  OAI21X1  g12474(.A0(new_n14680_), .A1(new_n6900_), .B0(new_n14719_), .Y(new_n14911_));
  OAI21X1  g12475(.A0(new_n14911_), .A1(new_n14865_), .B0(new_n14910_), .Y(new_n14912_));
  OAI21X1  g12476(.A0(new_n14861_), .A1(pi0152), .B0(new_n14650_), .Y(new_n14913_));
  AND2X1   g12477(.A(new_n14913_), .B(pi0299), .Y(new_n14914_));
  AND2X1   g12478(.A(new_n14914_), .B(new_n14912_), .Y(new_n14915_));
  NOR2X1   g12479(.A(new_n12064_), .B(pi0152), .Y(new_n14916_));
  AOI21X1  g12480(.A0(new_n12064_), .A1(new_n14590_), .B0(new_n2970_), .Y(new_n14917_));
  INVX1    g12481(.A(new_n14917_), .Y(new_n14918_));
  AOI21X1  g12482(.A0(new_n12064_), .A1(new_n5065_), .B0(new_n2970_), .Y(new_n14919_));
  OAI21X1  g12483(.A0(new_n14918_), .A1(new_n14916_), .B0(new_n14919_), .Y(new_n14920_));
  AOI21X1  g12484(.A0(new_n14909_), .A1(new_n2970_), .B0(pi0223), .Y(new_n14921_));
  NAND2X1  g12485(.A(new_n12010_), .B(new_n6900_), .Y(new_n14922_));
  NAND2X1  g12486(.A(new_n14922_), .B(new_n14688_), .Y(new_n14923_));
  AOI21X1  g12487(.A0(new_n14922_), .A1(new_n14687_), .B0(pi0299), .Y(new_n14924_));
  NAND2X1  g12488(.A(new_n14924_), .B(new_n14923_), .Y(new_n14925_));
  AOI21X1  g12489(.A0(new_n14921_), .A1(new_n14920_), .B0(new_n14925_), .Y(new_n14926_));
  NOR3X1   g12490(.A(new_n14926_), .B(new_n14915_), .C(new_n14908_), .Y(new_n14927_));
  AOI21X1  g12491(.A0(new_n11953_), .A1(pi0152), .B0(new_n14720_), .Y(new_n14928_));
  INVX1    g12492(.A(new_n12064_), .Y(new_n14929_));
  OAI21X1  g12493(.A0(new_n14591_), .A1(new_n14929_), .B0(new_n2971_), .Y(new_n14930_));
  OAI22X1  g12494(.A0(new_n14930_), .A1(new_n14916_), .B0(new_n14928_), .B1(new_n2971_), .Y(new_n14931_));
  NAND2X1  g12495(.A(new_n14923_), .B(new_n2953_), .Y(new_n14932_));
  AOI21X1  g12496(.A0(new_n14931_), .A1(new_n2964_), .B0(new_n14932_), .Y(new_n14933_));
  AND2X1   g12497(.A(new_n14910_), .B(new_n14679_), .Y(new_n14934_));
  NOR2X1   g12498(.A(new_n14699_), .B(new_n14591_), .Y(new_n14935_));
  OAI21X1  g12499(.A0(new_n14935_), .A1(new_n14913_), .B0(pi0299), .Y(new_n14936_));
  AOI21X1  g12500(.A0(new_n14934_), .A1(new_n14911_), .B0(new_n14936_), .Y(new_n14937_));
  NOR3X1   g12501(.A(new_n14937_), .B(new_n14933_), .C(pi0759), .Y(new_n14938_));
  NOR3X1   g12502(.A(new_n14938_), .B(new_n14927_), .C(new_n2959_), .Y(new_n14939_));
  NOR2X1   g12503(.A(new_n11947_), .B(pi0039), .Y(new_n14940_));
  AOI21X1  g12504(.A0(pi0947), .A1(pi0759), .B0(pi0039), .Y(new_n14941_));
  OAI22X1  g12505(.A0(new_n14941_), .A1(new_n14940_), .B0(new_n11947_), .B1(new_n6900_), .Y(new_n14942_));
  OAI21X1  g12506(.A0(new_n14942_), .A1(new_n14727_), .B0(new_n2996_), .Y(new_n14943_));
  INVX1    g12507(.A(pi0696), .Y(new_n14944_));
  OR2X1    g12508(.A(new_n12202_), .B(pi0152), .Y(new_n14945_));
  NOR4X1   g12509(.A(new_n14591_), .B(new_n3003_), .C(new_n2740_), .D(new_n2555_), .Y(new_n14946_));
  AOI21X1  g12510(.A0(new_n14946_), .A1(new_n14941_), .B0(new_n2996_), .Y(new_n14947_));
  AOI21X1  g12511(.A0(new_n14947_), .A1(new_n14945_), .B0(new_n14944_), .Y(new_n14948_));
  OAI21X1  g12512(.A0(new_n14943_), .A1(new_n14939_), .B0(new_n14948_), .Y(new_n14949_));
  INVX1    g12513(.A(new_n14647_), .Y(new_n14950_));
  AOI21X1  g12514(.A0(new_n14911_), .A1(new_n14950_), .B0(new_n14667_), .Y(new_n14951_));
  MX2X1    g12515(.A(pi0947), .B(pi0152), .S0(new_n11953_), .Y(new_n14952_));
  OAI21X1  g12516(.A0(new_n14952_), .A1(new_n10137_), .B0(new_n2954_), .Y(new_n14953_));
  OR2X1    g12517(.A(new_n14665_), .B(new_n2953_), .Y(new_n14954_));
  AOI21X1  g12518(.A0(new_n14652_), .A1(pi0152), .B0(new_n14954_), .Y(new_n14955_));
  OAI21X1  g12519(.A0(new_n14953_), .A1(new_n14951_), .B0(new_n14955_), .Y(new_n14956_));
  NOR2X1   g12520(.A(new_n14918_), .B(new_n14916_), .Y(new_n14957_));
  AND2X1   g12521(.A(new_n14952_), .B(new_n2970_), .Y(new_n14958_));
  OAI21X1  g12522(.A0(new_n14958_), .A1(new_n14957_), .B0(new_n2964_), .Y(new_n14959_));
  AOI21X1  g12523(.A0(new_n14959_), .A1(new_n14924_), .B0(new_n14908_), .Y(new_n14960_));
  AOI21X1  g12524(.A0(new_n12088_), .A1(new_n12068_), .B0(pi0759), .Y(new_n14961_));
  AND2X1   g12525(.A(new_n14961_), .B(pi0152), .Y(new_n14962_));
  OR2X1    g12526(.A(new_n14962_), .B(new_n2959_), .Y(new_n14963_));
  AOI21X1  g12527(.A0(new_n14960_), .A1(new_n14956_), .B0(new_n14963_), .Y(new_n14964_));
  NAND2X1  g12528(.A(new_n14942_), .B(new_n2996_), .Y(new_n14965_));
  NAND2X1  g12529(.A(pi0947), .B(pi0759), .Y(new_n14966_));
  AOI21X1  g12530(.A0(new_n14966_), .A1(new_n12202_), .B0(new_n2996_), .Y(new_n14967_));
  OAI21X1  g12531(.A0(new_n12572_), .A1(pi0152), .B0(new_n14967_), .Y(new_n14968_));
  AND2X1   g12532(.A(new_n14968_), .B(new_n14944_), .Y(new_n14969_));
  OAI21X1  g12533(.A0(new_n14965_), .A1(new_n14964_), .B0(new_n14969_), .Y(new_n14970_));
  AOI21X1  g12534(.A0(new_n14970_), .A1(new_n14949_), .B0(new_n9580_), .Y(new_n14971_));
  OAI21X1  g12535(.A0(new_n7686_), .A1(pi0152), .B0(new_n12898_), .Y(new_n14972_));
  NAND2X1  g12536(.A(new_n14966_), .B(new_n2739_), .Y(new_n14973_));
  AOI21X1  g12537(.A0(new_n14591_), .A1(pi0696), .B0(new_n14973_), .Y(new_n14974_));
  OAI21X1  g12538(.A0(new_n2739_), .A1(pi0152), .B0(pi0832), .Y(new_n14975_));
  OAI22X1  g12539(.A0(new_n14975_), .A1(new_n14974_), .B0(new_n14972_), .B1(new_n14971_), .Y(po0309));
  INVX1    g12540(.A(pi0766), .Y(new_n14977_));
  OAI21X1  g12541(.A0(new_n14590_), .A1(new_n14977_), .B0(new_n2739_), .Y(new_n14978_));
  AOI21X1  g12542(.A0(new_n14591_), .A1(pi0700), .B0(new_n14978_), .Y(new_n14979_));
  OAI21X1  g12543(.A0(new_n2739_), .A1(new_n8734_), .B0(pi0832), .Y(new_n14980_));
  INVX1    g12544(.A(new_n14727_), .Y(new_n14981_));
  INVX1    g12545(.A(new_n14661_), .Y(new_n14982_));
  NAND3X1  g12546(.A(new_n11947_), .B(new_n14977_), .C(new_n2959_), .Y(new_n14983_));
  AOI22X1  g12547(.A0(new_n14983_), .A1(new_n14982_), .B0(new_n11948_), .B1(new_n8734_), .Y(new_n14984_));
  INVX1    g12548(.A(new_n14650_), .Y(new_n14985_));
  AOI21X1  g12549(.A0(new_n12082_), .A1(new_n5065_), .B0(new_n8734_), .Y(new_n14986_));
  NOR2X1   g12550(.A(new_n10136_), .B(new_n8734_), .Y(new_n14987_));
  AOI22X1  g12551(.A0(new_n14987_), .A1(new_n14866_), .B0(new_n12075_), .B1(new_n10137_), .Y(new_n14988_));
  INVX1    g12552(.A(new_n14988_), .Y(new_n14989_));
  NOR3X1   g12553(.A(new_n11952_), .B(new_n2740_), .C(new_n5297_), .Y(new_n14990_));
  OAI21X1  g12554(.A0(new_n11952_), .A1(new_n2740_), .B0(new_n8734_), .Y(new_n14991_));
  NAND3X1  g12555(.A(new_n14991_), .B(new_n14668_), .C(new_n10136_), .Y(new_n14992_));
  OAI21X1  g12556(.A0(new_n14992_), .A1(new_n14990_), .B0(new_n2954_), .Y(new_n14993_));
  OAI22X1  g12557(.A0(new_n14993_), .A1(new_n14989_), .B0(new_n14986_), .B1(new_n14985_), .Y(new_n14994_));
  OR2X1    g12558(.A(new_n14873_), .B(new_n8734_), .Y(new_n14995_));
  AOI22X1  g12559(.A0(new_n14995_), .A1(new_n14690_), .B0(new_n14994_), .B1(pi0299), .Y(new_n14996_));
  OR2X1    g12560(.A(new_n14996_), .B(new_n14977_), .Y(new_n14997_));
  AOI22X1  g12561(.A0(new_n14991_), .A1(new_n14721_), .B0(new_n14680_), .B1(new_n10137_), .Y(new_n14998_));
  AOI21X1  g12562(.A0(new_n14998_), .A1(new_n14988_), .B0(pi0215), .Y(new_n14999_));
  INVX1    g12563(.A(new_n14699_), .Y(new_n15000_));
  INVX1    g12564(.A(new_n14986_), .Y(new_n15001_));
  AOI21X1  g12565(.A0(new_n15001_), .A1(new_n14650_), .B0(new_n15000_), .Y(new_n15002_));
  OR2X1    g12566(.A(new_n15002_), .B(new_n14665_), .Y(new_n15003_));
  OAI21X1  g12567(.A0(new_n15003_), .A1(new_n14999_), .B0(pi0299), .Y(new_n15004_));
  OAI21X1  g12568(.A0(new_n14740_), .A1(pi0153), .B0(new_n14725_), .Y(new_n15005_));
  NAND3X1  g12569(.A(new_n15005_), .B(new_n15004_), .C(new_n14977_), .Y(new_n15006_));
  AND2X1   g12570(.A(new_n15006_), .B(pi0039), .Y(new_n15007_));
  AOI22X1  g12571(.A0(new_n15007_), .A1(new_n14997_), .B0(new_n14984_), .B1(new_n14981_), .Y(new_n15008_));
  AOI21X1  g12572(.A0(pi0947), .A1(new_n14977_), .B0(pi0039), .Y(new_n15009_));
  AOI21X1  g12573(.A0(new_n15009_), .A1(new_n14810_), .B0(new_n2996_), .Y(new_n15010_));
  OAI21X1  g12574(.A0(new_n12202_), .A1(pi0153), .B0(new_n15010_), .Y(new_n15011_));
  OAI21X1  g12575(.A0(new_n15008_), .A1(pi0038), .B0(new_n15011_), .Y(new_n15012_));
  OAI21X1  g12576(.A0(new_n14740_), .A1(pi0153), .B0(new_n14663_), .Y(new_n15013_));
  NAND3X1  g12577(.A(new_n14992_), .B(new_n14988_), .C(new_n14894_), .Y(new_n15014_));
  AOI21X1  g12578(.A0(new_n15001_), .A1(new_n14652_), .B0(new_n2953_), .Y(new_n15015_));
  AOI21X1  g12579(.A0(new_n15015_), .A1(new_n15014_), .B0(new_n14977_), .Y(new_n15016_));
  NAND2X1  g12580(.A(new_n15016_), .B(new_n15013_), .Y(new_n15017_));
  NOR2X1   g12581(.A(pi0766), .B(pi0153), .Y(new_n15018_));
  AOI21X1  g12582(.A0(new_n15018_), .A1(new_n12089_), .B0(new_n2959_), .Y(new_n15019_));
  OR2X1    g12583(.A(new_n14984_), .B(pi0038), .Y(new_n15020_));
  AOI21X1  g12584(.A0(new_n15019_), .A1(new_n15017_), .B0(new_n15020_), .Y(new_n15021_));
  INVX1    g12585(.A(pi0700), .Y(new_n15022_));
  AOI21X1  g12586(.A0(new_n4995_), .A1(new_n2739_), .B0(new_n8734_), .Y(new_n15023_));
  OAI21X1  g12587(.A0(new_n14978_), .A1(new_n14411_), .B0(pi0038), .Y(new_n15024_));
  OAI21X1  g12588(.A0(new_n15024_), .A1(new_n15023_), .B0(new_n15022_), .Y(new_n15025_));
  OAI21X1  g12589(.A0(new_n15025_), .A1(new_n15021_), .B0(new_n14757_), .Y(new_n15026_));
  AOI21X1  g12590(.A0(new_n15012_), .A1(pi0700), .B0(new_n15026_), .Y(new_n15027_));
  AOI21X1  g12591(.A0(new_n5117_), .A1(new_n3129_), .B0(pi0153), .Y(new_n15028_));
  NOR3X1   g12592(.A(new_n15028_), .B(new_n15027_), .C(pi0057), .Y(new_n15029_));
  OAI21X1  g12593(.A0(new_n8734_), .A1(new_n2436_), .B0(new_n12898_), .Y(new_n15030_));
  OAI22X1  g12594(.A0(new_n15030_), .A1(new_n15029_), .B0(new_n14980_), .B1(new_n14979_), .Y(po0310));
  OAI22X1  g12595(.A0(new_n14638_), .A1(pi0704), .B0(new_n14590_), .B1(pi0742), .Y(new_n15032_));
  OAI21X1  g12596(.A0(new_n2739_), .A1(pi0154), .B0(pi0832), .Y(new_n15033_));
  AOI21X1  g12597(.A0(new_n15032_), .A1(new_n2739_), .B0(new_n15033_), .Y(new_n15034_));
  OAI21X1  g12598(.A0(new_n11947_), .A1(pi0154), .B0(new_n14856_), .Y(new_n15035_));
  AOI21X1  g12599(.A0(new_n14726_), .A1(pi0154), .B0(new_n2959_), .Y(new_n15036_));
  OAI21X1  g12600(.A0(new_n14714_), .A1(pi0154), .B0(new_n15036_), .Y(new_n15037_));
  AOI21X1  g12601(.A0(new_n15037_), .A1(new_n15035_), .B0(pi0038), .Y(new_n15038_));
  INVX1    g12602(.A(new_n14732_), .Y(new_n15039_));
  NOR2X1   g12603(.A(new_n12202_), .B(pi0154), .Y(new_n15040_));
  OAI21X1  g12604(.A0(new_n15040_), .A1(new_n15039_), .B0(pi0742), .Y(new_n15041_));
  NOR2X1   g12605(.A(new_n15041_), .B(new_n15038_), .Y(new_n15042_));
  AOI21X1  g12606(.A0(new_n14703_), .A1(pi0154), .B0(new_n2959_), .Y(new_n15043_));
  OAI21X1  g12607(.A0(new_n14693_), .A1(pi0154), .B0(new_n15043_), .Y(new_n15044_));
  OAI21X1  g12608(.A0(new_n15035_), .A1(new_n14697_), .B0(new_n15044_), .Y(new_n15045_));
  INVX1    g12609(.A(pi0742), .Y(new_n15046_));
  INVX1    g12610(.A(new_n14709_), .Y(new_n15047_));
  OAI21X1  g12611(.A0(new_n15040_), .A1(new_n15047_), .B0(new_n15046_), .Y(new_n15048_));
  AOI21X1  g12612(.A0(new_n15045_), .A1(new_n2996_), .B0(new_n15048_), .Y(new_n15049_));
  NOR3X1   g12613(.A(new_n15049_), .B(new_n15042_), .C(pi0704), .Y(new_n15050_));
  AOI21X1  g12614(.A0(new_n11948_), .A1(new_n3158_), .B0(new_n14982_), .Y(new_n15051_));
  AOI21X1  g12615(.A0(new_n14654_), .A1(new_n14644_), .B0(pi0154), .Y(new_n15052_));
  AND2X1   g12616(.A(new_n14672_), .B(pi0154), .Y(new_n15053_));
  NOR3X1   g12617(.A(new_n15053_), .B(new_n15052_), .C(new_n2959_), .Y(new_n15054_));
  OAI21X1  g12618(.A0(new_n15054_), .A1(new_n15051_), .B0(new_n2996_), .Y(new_n15055_));
  OAI22X1  g12619(.A0(new_n14657_), .A1(new_n13402_), .B0(new_n12572_), .B1(pi0154), .Y(new_n15056_));
  AND2X1   g12620(.A(new_n15056_), .B(new_n15046_), .Y(new_n15057_));
  OR2X1    g12621(.A(new_n15046_), .B(pi0154), .Y(new_n15058_));
  OAI21X1  g12622(.A0(new_n15058_), .A1(new_n13699_), .B0(pi0704), .Y(new_n15059_));
  AOI21X1  g12623(.A0(new_n15057_), .A1(new_n15055_), .B0(new_n15059_), .Y(new_n15060_));
  OR4X1    g12624(.A(new_n15060_), .B(new_n15050_), .C(po1038), .D(new_n3810_), .Y(new_n15061_));
  AOI21X1  g12625(.A0(new_n9580_), .A1(new_n3158_), .B0(pi0832), .Y(new_n15062_));
  AOI21X1  g12626(.A0(new_n15062_), .A1(new_n15061_), .B0(new_n15034_), .Y(po0311));
  INVX1    g12627(.A(pi0155), .Y(new_n15064_));
  INVX1    g12628(.A(pi0757), .Y(new_n15065_));
  INVX1    g12629(.A(new_n14704_), .Y(new_n15066_));
  AOI21X1  g12630(.A0(new_n15066_), .A1(new_n2996_), .B0(new_n14709_), .Y(new_n15067_));
  NAND2X1  g12631(.A(new_n15067_), .B(new_n15065_), .Y(new_n15068_));
  AOI21X1  g12632(.A0(new_n14729_), .A1(new_n2996_), .B0(new_n14732_), .Y(new_n15069_));
  AOI21X1  g12633(.A0(new_n15069_), .A1(pi0757), .B0(pi0686), .Y(new_n15070_));
  AND2X1   g12634(.A(new_n15070_), .B(new_n15068_), .Y(new_n15071_));
  OR2X1    g12635(.A(new_n14675_), .B(pi0757), .Y(new_n15072_));
  AND2X1   g12636(.A(new_n15072_), .B(pi0686), .Y(new_n15073_));
  NOR3X1   g12637(.A(new_n15073_), .B(new_n15071_), .C(new_n9580_), .Y(new_n15074_));
  MX2X1    g12638(.A(new_n14708_), .B(new_n14696_), .S0(new_n2996_), .Y(new_n15075_));
  OR2X1    g12639(.A(new_n15075_), .B(pi0757), .Y(new_n15076_));
  AOI22X1  g12640(.A0(new_n14732_), .A1(new_n12202_), .B0(new_n14716_), .B1(new_n2996_), .Y(new_n15077_));
  AOI21X1  g12641(.A0(new_n15077_), .A1(pi0757), .B0(pi0686), .Y(new_n15078_));
  OAI21X1  g12642(.A0(new_n13699_), .A1(new_n15065_), .B0(pi0686), .Y(new_n15079_));
  AOI21X1  g12643(.A0(new_n14658_), .A1(new_n15065_), .B0(new_n15079_), .Y(new_n15080_));
  AOI21X1  g12644(.A0(new_n15078_), .A1(new_n15076_), .B0(new_n15080_), .Y(new_n15081_));
  NAND3X1  g12645(.A(new_n6520_), .B(new_n3129_), .C(new_n15064_), .Y(new_n15082_));
  OAI22X1  g12646(.A0(new_n15082_), .A1(new_n15081_), .B0(new_n15074_), .B1(new_n15064_), .Y(new_n15083_));
  OAI22X1  g12647(.A0(new_n14638_), .A1(pi0686), .B0(new_n14590_), .B1(pi0757), .Y(new_n15084_));
  OAI21X1  g12648(.A0(new_n2739_), .A1(pi0155), .B0(pi0832), .Y(new_n15085_));
  AOI21X1  g12649(.A0(new_n15084_), .A1(new_n2739_), .B0(new_n15085_), .Y(new_n15086_));
  AOI21X1  g12650(.A0(new_n15083_), .A1(new_n12898_), .B0(new_n15086_), .Y(po0312));
  OAI22X1  g12651(.A0(new_n14638_), .A1(pi0724), .B0(new_n14590_), .B1(pi0741), .Y(new_n15088_));
  OAI21X1  g12652(.A0(new_n2739_), .A1(pi0156), .B0(pi0832), .Y(new_n15089_));
  AOI21X1  g12653(.A0(new_n15088_), .A1(new_n2739_), .B0(new_n15089_), .Y(new_n15090_));
  INVX1    g12654(.A(pi0741), .Y(new_n15091_));
  INVX1    g12655(.A(pi0724), .Y(new_n15092_));
  OAI21X1  g12656(.A0(new_n15077_), .A1(new_n15091_), .B0(new_n15092_), .Y(new_n15093_));
  AOI21X1  g12657(.A0(new_n15075_), .A1(new_n15091_), .B0(new_n15093_), .Y(new_n15094_));
  AOI21X1  g12658(.A0(new_n13699_), .A1(pi0741), .B0(new_n15092_), .Y(new_n15095_));
  OAI21X1  g12659(.A0(new_n14658_), .A1(pi0741), .B0(new_n15095_), .Y(new_n15096_));
  NAND2X1  g12660(.A(new_n15096_), .B(new_n7686_), .Y(new_n15097_));
  OAI21X1  g12661(.A0(new_n15097_), .A1(new_n15094_), .B0(new_n8876_), .Y(new_n15098_));
  NOR2X1   g12662(.A(new_n15067_), .B(pi0741), .Y(new_n15099_));
  OAI21X1  g12663(.A0(new_n15069_), .A1(new_n15091_), .B0(new_n15092_), .Y(new_n15100_));
  OR2X1    g12664(.A(pi0741), .B(new_n15092_), .Y(new_n15101_));
  OAI22X1  g12665(.A0(new_n15101_), .A1(new_n14675_), .B0(new_n15100_), .B1(new_n15099_), .Y(new_n15102_));
  AND2X1   g12666(.A(new_n7686_), .B(pi0156), .Y(new_n15103_));
  AOI21X1  g12667(.A0(new_n15103_), .A1(new_n15102_), .B0(pi0832), .Y(new_n15104_));
  AOI21X1  g12668(.A0(new_n15104_), .A1(new_n15098_), .B0(new_n15090_), .Y(po0313));
  INVX1    g12669(.A(pi0760), .Y(new_n15106_));
  AND2X1   g12670(.A(pi0947), .B(new_n15106_), .Y(new_n15107_));
  INVX1    g12671(.A(new_n15107_), .Y(new_n15108_));
  OAI21X1  g12672(.A0(new_n14638_), .A1(pi0688), .B0(new_n15108_), .Y(new_n15109_));
  OAI21X1  g12673(.A0(new_n2739_), .A1(pi0157), .B0(pi0832), .Y(new_n15110_));
  AOI21X1  g12674(.A0(new_n15109_), .A1(new_n2739_), .B0(new_n15110_), .Y(new_n15111_));
  INVX1    g12675(.A(pi0688), .Y(new_n15112_));
  AOI21X1  g12676(.A0(new_n15108_), .A1(new_n12202_), .B0(new_n2996_), .Y(new_n15113_));
  OAI21X1  g12677(.A0(new_n12572_), .A1(new_n10060_), .B0(new_n15113_), .Y(new_n15114_));
  OR2X1    g12678(.A(new_n2953_), .B(pi0157), .Y(new_n15115_));
  AOI22X1  g12679(.A0(new_n14671_), .A1(new_n15115_), .B0(new_n14759_), .B1(new_n10060_), .Y(new_n15116_));
  OAI21X1  g12680(.A0(new_n14740_), .A1(pi0157), .B0(new_n14663_), .Y(new_n15117_));
  NAND2X1  g12681(.A(new_n15117_), .B(new_n15106_), .Y(new_n15118_));
  AND2X1   g12682(.A(pi0760), .B(new_n10060_), .Y(new_n15119_));
  AOI21X1  g12683(.A0(new_n15119_), .A1(new_n12089_), .B0(new_n2959_), .Y(new_n15120_));
  OAI21X1  g12684(.A0(new_n15118_), .A1(new_n15116_), .B0(new_n15120_), .Y(new_n15121_));
  AOI21X1  g12685(.A0(new_n15107_), .A1(new_n11947_), .B0(pi0039), .Y(new_n15122_));
  OAI21X1  g12686(.A0(new_n11947_), .A1(pi0157), .B0(new_n15122_), .Y(new_n15123_));
  NAND3X1  g12687(.A(new_n15123_), .B(new_n15121_), .C(new_n2996_), .Y(new_n15124_));
  AOI21X1  g12688(.A0(new_n15124_), .A1(new_n15114_), .B0(new_n15112_), .Y(new_n15125_));
  NOR3X1   g12689(.A(new_n14692_), .B(new_n14683_), .C(pi0760), .Y(new_n15126_));
  OR2X1    g12690(.A(new_n15126_), .B(pi0157), .Y(new_n15127_));
  AOI21X1  g12691(.A0(new_n14714_), .A1(pi0760), .B0(new_n15127_), .Y(new_n15128_));
  NOR2X1   g12692(.A(new_n14703_), .B(pi0760), .Y(new_n15129_));
  OAI21X1  g12693(.A0(new_n14726_), .A1(new_n15106_), .B0(pi0157), .Y(new_n15130_));
  OAI21X1  g12694(.A0(new_n15130_), .A1(new_n15129_), .B0(pi0039), .Y(new_n15131_));
  OAI22X1  g12695(.A0(new_n15131_), .A1(new_n15128_), .B0(new_n15123_), .B1(new_n14727_), .Y(new_n15132_));
  NOR2X1   g12696(.A(new_n12202_), .B(pi0157), .Y(new_n15133_));
  OAI21X1  g12697(.A0(new_n14590_), .A1(new_n15106_), .B0(new_n2959_), .Y(new_n15134_));
  OAI21X1  g12698(.A0(new_n15134_), .A1(new_n14811_), .B0(pi0038), .Y(new_n15135_));
  OAI21X1  g12699(.A0(new_n15135_), .A1(new_n15133_), .B0(new_n15112_), .Y(new_n15136_));
  AOI21X1  g12700(.A0(new_n15132_), .A1(new_n2996_), .B0(new_n15136_), .Y(new_n15137_));
  OAI21X1  g12701(.A0(new_n15137_), .A1(new_n15125_), .B0(new_n7686_), .Y(new_n15138_));
  AOI21X1  g12702(.A0(new_n9580_), .A1(new_n10060_), .B0(pi0832), .Y(new_n15139_));
  AOI21X1  g12703(.A0(new_n15139_), .A1(new_n15138_), .B0(new_n15111_), .Y(po0314));
  INVX1    g12704(.A(pi0753), .Y(new_n15141_));
  OAI21X1  g12705(.A0(new_n14672_), .A1(new_n5128_), .B0(new_n15141_), .Y(new_n15142_));
  AOI21X1  g12706(.A0(new_n14819_), .A1(new_n5128_), .B0(new_n15142_), .Y(new_n15143_));
  NOR3X1   g12707(.A(new_n14823_), .B(new_n15141_), .C(pi0158), .Y(new_n15144_));
  OAI21X1  g12708(.A0(new_n15144_), .A1(new_n15143_), .B0(pi0039), .Y(new_n15145_));
  MX2X1    g12709(.A(new_n5128_), .B(new_n15141_), .S0(new_n11947_), .Y(new_n15146_));
  AOI21X1  g12710(.A0(new_n15146_), .A1(new_n14642_), .B0(pi0038), .Y(new_n15147_));
  OR2X1    g12711(.A(new_n14590_), .B(pi0753), .Y(new_n15148_));
  AOI22X1  g12712(.A0(new_n15148_), .A1(new_n12202_), .B0(new_n12573_), .B1(pi0158), .Y(new_n15149_));
  OAI21X1  g12713(.A0(new_n15149_), .A1(new_n2996_), .B0(pi0702), .Y(new_n15150_));
  AOI21X1  g12714(.A0(new_n15147_), .A1(new_n15145_), .B0(new_n15150_), .Y(new_n15151_));
  OAI21X1  g12715(.A0(new_n14726_), .A1(new_n5128_), .B0(pi0753), .Y(new_n15152_));
  AOI21X1  g12716(.A0(new_n14714_), .A1(new_n5128_), .B0(new_n15152_), .Y(new_n15153_));
  OAI21X1  g12717(.A0(new_n14703_), .A1(new_n5128_), .B0(new_n15141_), .Y(new_n15154_));
  AOI21X1  g12718(.A0(new_n14693_), .A1(new_n5128_), .B0(new_n15154_), .Y(new_n15155_));
  OAI21X1  g12719(.A0(new_n15155_), .A1(new_n15153_), .B0(pi0039), .Y(new_n15156_));
  NAND3X1  g12720(.A(new_n15148_), .B(new_n14638_), .C(new_n11947_), .Y(new_n15157_));
  AOI21X1  g12721(.A0(new_n11948_), .A1(pi0158), .B0(pi0039), .Y(new_n15158_));
  AOI21X1  g12722(.A0(new_n15158_), .A1(new_n15157_), .B0(pi0038), .Y(new_n15159_));
  INVX1    g12723(.A(pi0702), .Y(new_n15160_));
  NOR2X1   g12724(.A(new_n12202_), .B(pi0158), .Y(new_n15161_));
  OAI21X1  g12725(.A0(new_n14590_), .A1(new_n15141_), .B0(new_n2959_), .Y(new_n15162_));
  OAI21X1  g12726(.A0(new_n15162_), .A1(new_n14811_), .B0(pi0038), .Y(new_n15163_));
  OAI21X1  g12727(.A0(new_n15163_), .A1(new_n15161_), .B0(new_n15160_), .Y(new_n15164_));
  AOI21X1  g12728(.A0(new_n15159_), .A1(new_n15156_), .B0(new_n15164_), .Y(new_n15165_));
  OAI21X1  g12729(.A0(new_n15165_), .A1(new_n15151_), .B0(new_n7686_), .Y(new_n15166_));
  AOI21X1  g12730(.A0(new_n9580_), .A1(new_n5128_), .B0(pi0832), .Y(new_n15167_));
  OAI21X1  g12731(.A0(new_n14638_), .A1(pi0702), .B0(new_n15148_), .Y(new_n15168_));
  OAI21X1  g12732(.A0(new_n2739_), .A1(pi0158), .B0(pi0832), .Y(new_n15169_));
  AOI21X1  g12733(.A0(new_n15168_), .A1(new_n2739_), .B0(new_n15169_), .Y(new_n15170_));
  AOI21X1  g12734(.A0(new_n15167_), .A1(new_n15166_), .B0(new_n15170_), .Y(po0315));
  INVX1    g12735(.A(pi0754), .Y(new_n15172_));
  OAI21X1  g12736(.A0(new_n14672_), .A1(new_n5129_), .B0(new_n15172_), .Y(new_n15173_));
  AOI21X1  g12737(.A0(new_n14819_), .A1(new_n5129_), .B0(new_n15173_), .Y(new_n15174_));
  NOR3X1   g12738(.A(new_n14823_), .B(new_n15172_), .C(pi0159), .Y(new_n15175_));
  OAI21X1  g12739(.A0(new_n15175_), .A1(new_n15174_), .B0(pi0039), .Y(new_n15176_));
  MX2X1    g12740(.A(new_n5129_), .B(new_n15172_), .S0(new_n11947_), .Y(new_n15177_));
  AOI21X1  g12741(.A0(new_n15177_), .A1(new_n14642_), .B0(pi0038), .Y(new_n15178_));
  OR2X1    g12742(.A(new_n14590_), .B(pi0754), .Y(new_n15179_));
  AOI22X1  g12743(.A0(new_n15179_), .A1(new_n12202_), .B0(new_n12573_), .B1(pi0159), .Y(new_n15180_));
  OAI21X1  g12744(.A0(new_n15180_), .A1(new_n2996_), .B0(pi0709), .Y(new_n15181_));
  AOI21X1  g12745(.A0(new_n15178_), .A1(new_n15176_), .B0(new_n15181_), .Y(new_n15182_));
  OAI21X1  g12746(.A0(new_n14726_), .A1(new_n5129_), .B0(pi0754), .Y(new_n15183_));
  AOI21X1  g12747(.A0(new_n14714_), .A1(new_n5129_), .B0(new_n15183_), .Y(new_n15184_));
  OAI21X1  g12748(.A0(new_n14703_), .A1(new_n5129_), .B0(new_n15172_), .Y(new_n15185_));
  AOI21X1  g12749(.A0(new_n14693_), .A1(new_n5129_), .B0(new_n15185_), .Y(new_n15186_));
  OAI21X1  g12750(.A0(new_n15186_), .A1(new_n15184_), .B0(pi0039), .Y(new_n15187_));
  NAND3X1  g12751(.A(new_n15179_), .B(new_n14638_), .C(new_n11947_), .Y(new_n15188_));
  AOI21X1  g12752(.A0(new_n11948_), .A1(pi0159), .B0(pi0039), .Y(new_n15189_));
  AOI21X1  g12753(.A0(new_n15189_), .A1(new_n15188_), .B0(pi0038), .Y(new_n15190_));
  INVX1    g12754(.A(pi0709), .Y(new_n15191_));
  NOR2X1   g12755(.A(new_n12202_), .B(pi0159), .Y(new_n15192_));
  OAI21X1  g12756(.A0(new_n14590_), .A1(new_n15172_), .B0(new_n2959_), .Y(new_n15193_));
  OAI21X1  g12757(.A0(new_n15193_), .A1(new_n14811_), .B0(pi0038), .Y(new_n15194_));
  OAI21X1  g12758(.A0(new_n15194_), .A1(new_n15192_), .B0(new_n15191_), .Y(new_n15195_));
  AOI21X1  g12759(.A0(new_n15190_), .A1(new_n15187_), .B0(new_n15195_), .Y(new_n15196_));
  OAI21X1  g12760(.A0(new_n15196_), .A1(new_n15182_), .B0(new_n7686_), .Y(new_n15197_));
  AOI21X1  g12761(.A0(new_n9580_), .A1(new_n5129_), .B0(pi0832), .Y(new_n15198_));
  OAI21X1  g12762(.A0(new_n14638_), .A1(pi0709), .B0(new_n15179_), .Y(new_n15199_));
  OAI21X1  g12763(.A0(new_n2739_), .A1(pi0159), .B0(pi0832), .Y(new_n15200_));
  AOI21X1  g12764(.A0(new_n15199_), .A1(new_n2739_), .B0(new_n15200_), .Y(new_n15201_));
  AOI21X1  g12765(.A0(new_n15198_), .A1(new_n15197_), .B0(new_n15201_), .Y(po0316));
  INVX1    g12766(.A(pi0756), .Y(new_n15203_));
  AND2X1   g12767(.A(pi0947), .B(new_n15203_), .Y(new_n15204_));
  INVX1    g12768(.A(new_n15204_), .Y(new_n15205_));
  OAI21X1  g12769(.A0(new_n14638_), .A1(pi0734), .B0(new_n15205_), .Y(new_n15206_));
  OAI21X1  g12770(.A0(new_n2739_), .A1(pi0160), .B0(pi0832), .Y(new_n15207_));
  AOI21X1  g12771(.A0(new_n15206_), .A1(new_n2739_), .B0(new_n15207_), .Y(new_n15208_));
  INVX1    g12772(.A(pi0734), .Y(new_n15209_));
  AOI21X1  g12773(.A0(new_n15205_), .A1(new_n12202_), .B0(new_n2996_), .Y(new_n15210_));
  OAI21X1  g12774(.A0(new_n12572_), .A1(new_n8747_), .B0(new_n15210_), .Y(new_n15211_));
  OAI21X1  g12775(.A0(new_n14760_), .A1(new_n8747_), .B0(pi0299), .Y(new_n15212_));
  AOI21X1  g12776(.A0(new_n14759_), .A1(new_n8747_), .B0(new_n15212_), .Y(new_n15213_));
  OAI21X1  g12777(.A0(new_n14740_), .A1(pi0160), .B0(new_n14663_), .Y(new_n15214_));
  NAND2X1  g12778(.A(new_n15214_), .B(new_n15203_), .Y(new_n15215_));
  AND2X1   g12779(.A(pi0756), .B(new_n8747_), .Y(new_n15216_));
  AOI21X1  g12780(.A0(new_n15216_), .A1(new_n12089_), .B0(new_n2959_), .Y(new_n15217_));
  OAI21X1  g12781(.A0(new_n15215_), .A1(new_n15213_), .B0(new_n15217_), .Y(new_n15218_));
  AOI21X1  g12782(.A0(new_n15204_), .A1(new_n11947_), .B0(pi0039), .Y(new_n15219_));
  OAI21X1  g12783(.A0(new_n11947_), .A1(pi0160), .B0(new_n15219_), .Y(new_n15220_));
  NAND3X1  g12784(.A(new_n15220_), .B(new_n15218_), .C(new_n2996_), .Y(new_n15221_));
  AOI21X1  g12785(.A0(new_n15221_), .A1(new_n15211_), .B0(new_n15209_), .Y(new_n15222_));
  OAI21X1  g12786(.A0(new_n14703_), .A1(new_n8747_), .B0(new_n15203_), .Y(new_n15223_));
  AOI21X1  g12787(.A0(new_n14693_), .A1(new_n8747_), .B0(new_n15223_), .Y(new_n15224_));
  NOR3X1   g12788(.A(new_n14712_), .B(new_n2953_), .C(pi0160), .Y(new_n15225_));
  AND2X1   g12789(.A(new_n14713_), .B(pi0756), .Y(new_n15226_));
  OAI21X1  g12790(.A0(new_n14742_), .A1(new_n8747_), .B0(new_n15226_), .Y(new_n15227_));
  OAI21X1  g12791(.A0(new_n15227_), .A1(new_n15225_), .B0(pi0039), .Y(new_n15228_));
  OAI22X1  g12792(.A0(new_n15228_), .A1(new_n15224_), .B0(new_n15220_), .B1(new_n14727_), .Y(new_n15229_));
  NOR2X1   g12793(.A(new_n12202_), .B(pi0160), .Y(new_n15230_));
  OAI21X1  g12794(.A0(new_n14590_), .A1(new_n15203_), .B0(new_n2959_), .Y(new_n15231_));
  OAI21X1  g12795(.A0(new_n15231_), .A1(new_n14811_), .B0(pi0038), .Y(new_n15232_));
  OAI21X1  g12796(.A0(new_n15232_), .A1(new_n15230_), .B0(new_n15209_), .Y(new_n15233_));
  AOI21X1  g12797(.A0(new_n15229_), .A1(new_n2996_), .B0(new_n15233_), .Y(new_n15234_));
  OAI21X1  g12798(.A0(new_n15234_), .A1(new_n15222_), .B0(new_n7686_), .Y(new_n15235_));
  AOI21X1  g12799(.A0(new_n9580_), .A1(new_n8747_), .B0(pi0832), .Y(new_n15236_));
  AOI21X1  g12800(.A0(new_n15236_), .A1(new_n15235_), .B0(new_n15208_), .Y(po0317));
  MX2X1    g12801(.A(new_n5064_), .B(new_n4613_), .S0(new_n11953_), .Y(new_n15238_));
  AOI21X1  g12802(.A0(new_n15238_), .A1(new_n10136_), .B0(pi0215), .Y(new_n15239_));
  OAI21X1  g12803(.A0(new_n14680_), .A1(new_n4613_), .B0(new_n14719_), .Y(new_n15240_));
  OAI21X1  g12804(.A0(new_n15240_), .A1(new_n14865_), .B0(new_n15239_), .Y(new_n15241_));
  OAI21X1  g12805(.A0(new_n14861_), .A1(pi0161), .B0(new_n14650_), .Y(new_n15242_));
  AND2X1   g12806(.A(new_n15242_), .B(pi0299), .Y(new_n15243_));
  AND2X1   g12807(.A(new_n15243_), .B(new_n15241_), .Y(new_n15244_));
  NOR2X1   g12808(.A(new_n12064_), .B(pi0161), .Y(new_n15245_));
  OAI21X1  g12809(.A0(new_n15245_), .A1(new_n14918_), .B0(new_n14919_), .Y(new_n15246_));
  AOI21X1  g12810(.A0(new_n15238_), .A1(new_n2970_), .B0(pi0223), .Y(new_n15247_));
  NAND2X1  g12811(.A(new_n12010_), .B(new_n4613_), .Y(new_n15248_));
  NAND2X1  g12812(.A(new_n15248_), .B(new_n14688_), .Y(new_n15249_));
  AOI21X1  g12813(.A0(new_n15248_), .A1(new_n14687_), .B0(pi0299), .Y(new_n15250_));
  NAND2X1  g12814(.A(new_n15250_), .B(new_n15249_), .Y(new_n15251_));
  AOI21X1  g12815(.A0(new_n15247_), .A1(new_n15246_), .B0(new_n15251_), .Y(new_n15252_));
  NOR3X1   g12816(.A(new_n15252_), .B(new_n15244_), .C(new_n13973_), .Y(new_n15253_));
  AOI21X1  g12817(.A0(new_n11953_), .A1(pi0161), .B0(new_n14720_), .Y(new_n15254_));
  OAI22X1  g12818(.A0(new_n15254_), .A1(new_n2971_), .B0(new_n15245_), .B1(new_n14930_), .Y(new_n15255_));
  NAND2X1  g12819(.A(new_n15249_), .B(new_n2953_), .Y(new_n15256_));
  AOI21X1  g12820(.A0(new_n15255_), .A1(new_n2964_), .B0(new_n15256_), .Y(new_n15257_));
  AND2X1   g12821(.A(new_n15239_), .B(new_n14679_), .Y(new_n15258_));
  OAI21X1  g12822(.A0(new_n15242_), .A1(new_n14935_), .B0(pi0299), .Y(new_n15259_));
  AOI21X1  g12823(.A0(new_n15258_), .A1(new_n15240_), .B0(new_n15259_), .Y(new_n15260_));
  NOR3X1   g12824(.A(new_n15260_), .B(new_n15257_), .C(pi0758), .Y(new_n15261_));
  NOR3X1   g12825(.A(new_n15261_), .B(new_n15253_), .C(new_n2959_), .Y(new_n15262_));
  AND2X1   g12826(.A(pi0947), .B(pi0758), .Y(new_n15263_));
  INVX1    g12827(.A(new_n15263_), .Y(new_n15264_));
  AOI21X1  g12828(.A0(new_n11948_), .A1(pi0161), .B0(pi0039), .Y(new_n15265_));
  OAI21X1  g12829(.A0(new_n15264_), .A1(new_n11948_), .B0(new_n15265_), .Y(new_n15266_));
  OAI21X1  g12830(.A0(new_n15266_), .A1(new_n14727_), .B0(new_n2996_), .Y(new_n15267_));
  OR2X1    g12831(.A(new_n12202_), .B(pi0161), .Y(new_n15268_));
  AOI21X1  g12832(.A0(pi0947), .A1(pi0758), .B0(pi0039), .Y(new_n15269_));
  AOI21X1  g12833(.A0(new_n15269_), .A1(new_n14946_), .B0(new_n2996_), .Y(new_n15270_));
  AOI21X1  g12834(.A0(new_n15270_), .A1(new_n15268_), .B0(new_n13969_), .Y(new_n15271_));
  OAI21X1  g12835(.A0(new_n15267_), .A1(new_n15262_), .B0(new_n15271_), .Y(new_n15272_));
  AOI21X1  g12836(.A0(new_n15240_), .A1(new_n14950_), .B0(new_n14667_), .Y(new_n15273_));
  MX2X1    g12837(.A(pi0947), .B(pi0161), .S0(new_n11953_), .Y(new_n15274_));
  OAI21X1  g12838(.A0(new_n15274_), .A1(new_n10137_), .B0(new_n2954_), .Y(new_n15275_));
  AOI21X1  g12839(.A0(new_n14652_), .A1(pi0161), .B0(new_n14954_), .Y(new_n15276_));
  OAI21X1  g12840(.A0(new_n15275_), .A1(new_n15273_), .B0(new_n15276_), .Y(new_n15277_));
  NOR2X1   g12841(.A(new_n15245_), .B(new_n14918_), .Y(new_n15278_));
  AND2X1   g12842(.A(new_n15274_), .B(new_n2970_), .Y(new_n15279_));
  OAI21X1  g12843(.A0(new_n15279_), .A1(new_n15278_), .B0(new_n2964_), .Y(new_n15280_));
  AOI21X1  g12844(.A0(new_n15280_), .A1(new_n15250_), .B0(new_n13973_), .Y(new_n15281_));
  AND2X1   g12845(.A(new_n13970_), .B(pi0161), .Y(new_n15282_));
  OR2X1    g12846(.A(new_n15282_), .B(new_n2959_), .Y(new_n15283_));
  AOI21X1  g12847(.A0(new_n15281_), .A1(new_n15277_), .B0(new_n15283_), .Y(new_n15284_));
  NAND2X1  g12848(.A(new_n15266_), .B(new_n2996_), .Y(new_n15285_));
  AOI21X1  g12849(.A0(new_n15264_), .A1(new_n12202_), .B0(new_n2996_), .Y(new_n15286_));
  OAI21X1  g12850(.A0(new_n12572_), .A1(pi0161), .B0(new_n15286_), .Y(new_n15287_));
  AND2X1   g12851(.A(new_n15287_), .B(new_n13969_), .Y(new_n15288_));
  OAI21X1  g12852(.A0(new_n15285_), .A1(new_n15284_), .B0(new_n15288_), .Y(new_n15289_));
  AOI21X1  g12853(.A0(new_n15289_), .A1(new_n15272_), .B0(new_n9580_), .Y(new_n15290_));
  OAI21X1  g12854(.A0(new_n7686_), .A1(pi0161), .B0(new_n12898_), .Y(new_n15291_));
  OAI21X1  g12855(.A0(new_n14590_), .A1(new_n13973_), .B0(new_n2739_), .Y(new_n15292_));
  AOI21X1  g12856(.A0(new_n14591_), .A1(pi0736), .B0(new_n15292_), .Y(new_n15293_));
  OAI21X1  g12857(.A0(new_n2739_), .A1(pi0161), .B0(pi0832), .Y(new_n15294_));
  OAI22X1  g12858(.A0(new_n15294_), .A1(new_n15293_), .B0(new_n15291_), .B1(new_n15290_), .Y(po0318));
  AND2X1   g12859(.A(pi0947), .B(new_n11890_), .Y(new_n15296_));
  INVX1    g12860(.A(new_n15296_), .Y(new_n15297_));
  AOI21X1  g12861(.A0(new_n15297_), .A1(new_n12202_), .B0(new_n2996_), .Y(new_n15298_));
  OAI21X1  g12862(.A0(new_n12572_), .A1(new_n7349_), .B0(new_n15298_), .Y(new_n15299_));
  OAI21X1  g12863(.A0(new_n12089_), .A1(new_n11890_), .B0(new_n7349_), .Y(new_n15300_));
  AOI21X1  g12864(.A0(new_n14654_), .A1(new_n11890_), .B0(new_n15300_), .Y(new_n15301_));
  AND2X1   g12865(.A(pi0299), .B(pi0162), .Y(new_n15302_));
  INVX1    g12866(.A(new_n15302_), .Y(new_n15303_));
  AOI21X1  g12867(.A0(new_n14670_), .A1(new_n14666_), .B0(new_n15303_), .Y(new_n15304_));
  OAI21X1  g12868(.A0(new_n15304_), .A1(new_n14643_), .B0(new_n11890_), .Y(new_n15305_));
  NAND2X1  g12869(.A(new_n15305_), .B(pi0039), .Y(new_n15306_));
  AOI21X1  g12870(.A0(new_n15296_), .A1(new_n11947_), .B0(pi0039), .Y(new_n15307_));
  OAI21X1  g12871(.A0(new_n11947_), .A1(pi0162), .B0(new_n15307_), .Y(new_n15308_));
  AND2X1   g12872(.A(new_n15308_), .B(new_n2996_), .Y(new_n15309_));
  OAI21X1  g12873(.A0(new_n15306_), .A1(new_n15301_), .B0(new_n15309_), .Y(new_n15310_));
  AOI21X1  g12874(.A0(new_n15310_), .A1(new_n15299_), .B0(new_n12565_), .Y(new_n15311_));
  OAI21X1  g12875(.A0(new_n14742_), .A1(new_n7349_), .B0(pi0761), .Y(new_n15312_));
  AOI21X1  g12876(.A0(new_n14714_), .A1(new_n15303_), .B0(new_n15312_), .Y(new_n15313_));
  NOR3X1   g12877(.A(new_n14692_), .B(new_n14683_), .C(pi0162), .Y(new_n15314_));
  OAI21X1  g12878(.A0(new_n14703_), .A1(new_n7349_), .B0(new_n11890_), .Y(new_n15315_));
  OAI21X1  g12879(.A0(new_n15315_), .A1(new_n15314_), .B0(pi0039), .Y(new_n15316_));
  OAI22X1  g12880(.A0(new_n15316_), .A1(new_n15313_), .B0(new_n15308_), .B1(new_n14727_), .Y(new_n15317_));
  NOR2X1   g12881(.A(new_n12202_), .B(pi0162), .Y(new_n15318_));
  OAI21X1  g12882(.A0(new_n14590_), .A1(new_n11890_), .B0(new_n2959_), .Y(new_n15319_));
  OAI21X1  g12883(.A0(new_n15319_), .A1(new_n14811_), .B0(pi0038), .Y(new_n15320_));
  OAI21X1  g12884(.A0(new_n15320_), .A1(new_n15318_), .B0(new_n12565_), .Y(new_n15321_));
  AOI21X1  g12885(.A0(new_n15317_), .A1(new_n2996_), .B0(new_n15321_), .Y(new_n15322_));
  OAI21X1  g12886(.A0(new_n15322_), .A1(new_n15311_), .B0(new_n7686_), .Y(new_n15323_));
  AOI21X1  g12887(.A0(new_n9580_), .A1(new_n7349_), .B0(pi0832), .Y(new_n15324_));
  OAI21X1  g12888(.A0(new_n14638_), .A1(pi0738), .B0(new_n15297_), .Y(new_n15325_));
  OAI21X1  g12889(.A0(new_n2739_), .A1(pi0162), .B0(pi0832), .Y(new_n15326_));
  AOI21X1  g12890(.A0(new_n15325_), .A1(new_n2739_), .B0(new_n15326_), .Y(new_n15327_));
  AOI21X1  g12891(.A0(new_n15324_), .A1(new_n15323_), .B0(new_n15327_), .Y(po0319));
  INVX1    g12892(.A(pi0777), .Y(new_n15329_));
  AND2X1   g12893(.A(pi0947), .B(new_n15329_), .Y(new_n15330_));
  INVX1    g12894(.A(new_n15330_), .Y(new_n15331_));
  OAI21X1  g12895(.A0(new_n14638_), .A1(pi0737), .B0(new_n15331_), .Y(new_n15332_));
  OAI21X1  g12896(.A0(new_n2739_), .A1(pi0163), .B0(pi0832), .Y(new_n15333_));
  AOI21X1  g12897(.A0(new_n15332_), .A1(new_n2739_), .B0(new_n15333_), .Y(new_n15334_));
  INVX1    g12898(.A(pi0737), .Y(new_n15335_));
  AOI21X1  g12899(.A0(new_n15331_), .A1(new_n12202_), .B0(new_n2996_), .Y(new_n15336_));
  OAI21X1  g12900(.A0(new_n12572_), .A1(new_n8705_), .B0(new_n15336_), .Y(new_n15337_));
  OR2X1    g12901(.A(new_n2953_), .B(pi0163), .Y(new_n15338_));
  AOI22X1  g12902(.A0(new_n14671_), .A1(new_n15338_), .B0(new_n14759_), .B1(new_n8705_), .Y(new_n15339_));
  OAI21X1  g12903(.A0(new_n14740_), .A1(pi0163), .B0(new_n14663_), .Y(new_n15340_));
  NAND2X1  g12904(.A(new_n15340_), .B(new_n15329_), .Y(new_n15341_));
  AND2X1   g12905(.A(pi0777), .B(new_n8705_), .Y(new_n15342_));
  AOI21X1  g12906(.A0(new_n15342_), .A1(new_n12089_), .B0(new_n2959_), .Y(new_n15343_));
  OAI21X1  g12907(.A0(new_n15341_), .A1(new_n15339_), .B0(new_n15343_), .Y(new_n15344_));
  AOI21X1  g12908(.A0(new_n15330_), .A1(new_n11947_), .B0(pi0039), .Y(new_n15345_));
  OAI21X1  g12909(.A0(new_n11947_), .A1(pi0163), .B0(new_n15345_), .Y(new_n15346_));
  NAND3X1  g12910(.A(new_n15346_), .B(new_n15344_), .C(new_n2996_), .Y(new_n15347_));
  AOI21X1  g12911(.A0(new_n15347_), .A1(new_n15337_), .B0(new_n15335_), .Y(new_n15348_));
  OAI21X1  g12912(.A0(new_n14703_), .A1(new_n8705_), .B0(new_n15329_), .Y(new_n15349_));
  AOI21X1  g12913(.A0(new_n14693_), .A1(new_n8705_), .B0(new_n15349_), .Y(new_n15350_));
  NOR3X1   g12914(.A(new_n14712_), .B(new_n2953_), .C(pi0163), .Y(new_n15351_));
  AND2X1   g12915(.A(new_n14713_), .B(pi0777), .Y(new_n15352_));
  OAI21X1  g12916(.A0(new_n14742_), .A1(new_n8705_), .B0(new_n15352_), .Y(new_n15353_));
  OAI21X1  g12917(.A0(new_n15353_), .A1(new_n15351_), .B0(pi0039), .Y(new_n15354_));
  OAI22X1  g12918(.A0(new_n15354_), .A1(new_n15350_), .B0(new_n15346_), .B1(new_n14727_), .Y(new_n15355_));
  NOR2X1   g12919(.A(new_n12202_), .B(pi0163), .Y(new_n15356_));
  OAI21X1  g12920(.A0(new_n14590_), .A1(new_n15329_), .B0(new_n2959_), .Y(new_n15357_));
  OAI21X1  g12921(.A0(new_n15357_), .A1(new_n14811_), .B0(pi0038), .Y(new_n15358_));
  OAI21X1  g12922(.A0(new_n15358_), .A1(new_n15356_), .B0(new_n15335_), .Y(new_n15359_));
  AOI21X1  g12923(.A0(new_n15355_), .A1(new_n2996_), .B0(new_n15359_), .Y(new_n15360_));
  OAI21X1  g12924(.A0(new_n15360_), .A1(new_n15348_), .B0(new_n7686_), .Y(new_n15361_));
  AOI21X1  g12925(.A0(new_n9580_), .A1(new_n8705_), .B0(pi0832), .Y(new_n15362_));
  AOI21X1  g12926(.A0(new_n15362_), .A1(new_n15361_), .B0(new_n15334_), .Y(po0320));
  INVX1    g12927(.A(pi0703), .Y(new_n15364_));
  OAI22X1  g12928(.A0(new_n14638_), .A1(new_n15364_), .B0(new_n14590_), .B1(pi0752), .Y(new_n15365_));
  OAI21X1  g12929(.A0(new_n2739_), .A1(pi0164), .B0(pi0832), .Y(new_n15366_));
  AOI21X1  g12930(.A0(new_n15365_), .A1(new_n2739_), .B0(new_n15366_), .Y(new_n15367_));
  AOI21X1  g12931(.A0(new_n14704_), .A1(pi0164), .B0(pi0038), .Y(new_n15368_));
  OAI21X1  g12932(.A0(new_n14696_), .A1(pi0164), .B0(new_n15368_), .Y(new_n15369_));
  INVX1    g12933(.A(pi0752), .Y(new_n15370_));
  OAI21X1  g12934(.A0(new_n14708_), .A1(pi0164), .B0(new_n14709_), .Y(new_n15371_));
  AND2X1   g12935(.A(new_n15371_), .B(new_n15370_), .Y(new_n15372_));
  AOI21X1  g12936(.A0(new_n14728_), .A1(pi0164), .B0(pi0038), .Y(new_n15373_));
  OAI21X1  g12937(.A0(new_n14716_), .A1(pi0164), .B0(new_n15373_), .Y(new_n15374_));
  OR2X1    g12938(.A(new_n12202_), .B(pi0164), .Y(new_n15375_));
  AOI21X1  g12939(.A0(new_n15375_), .A1(new_n14732_), .B0(new_n15370_), .Y(new_n15376_));
  AOI22X1  g12940(.A0(new_n15376_), .A1(new_n15374_), .B0(new_n15372_), .B1(new_n15369_), .Y(new_n15377_));
  OAI21X1  g12941(.A0(new_n14657_), .A1(new_n7223_), .B0(new_n15370_), .Y(new_n15378_));
  NOR2X1   g12942(.A(new_n15378_), .B(new_n14658_), .Y(new_n15379_));
  OAI21X1  g12943(.A0(new_n14675_), .A1(pi0752), .B0(pi0164), .Y(new_n15380_));
  AOI21X1  g12944(.A0(new_n13699_), .A1(pi0752), .B0(pi0703), .Y(new_n15381_));
  NAND2X1  g12945(.A(new_n15381_), .B(new_n15380_), .Y(new_n15382_));
  OAI22X1  g12946(.A0(new_n15382_), .A1(new_n15379_), .B0(new_n15377_), .B1(new_n15364_), .Y(new_n15383_));
  NAND2X1  g12947(.A(new_n15383_), .B(new_n7686_), .Y(new_n15384_));
  AOI21X1  g12948(.A0(new_n9580_), .A1(new_n7223_), .B0(pi0832), .Y(new_n15385_));
  AOI21X1  g12949(.A0(new_n15385_), .A1(new_n15384_), .B0(new_n15367_), .Y(po0321));
  OAI22X1  g12950(.A0(new_n14638_), .A1(new_n13680_), .B0(new_n14590_), .B1(pi0774), .Y(new_n15387_));
  OAI21X1  g12951(.A0(new_n2739_), .A1(pi0165), .B0(pi0832), .Y(new_n15388_));
  AOI21X1  g12952(.A0(new_n15387_), .A1(new_n2739_), .B0(new_n15388_), .Y(new_n15389_));
  AOI21X1  g12953(.A0(new_n14704_), .A1(pi0165), .B0(pi0038), .Y(new_n15390_));
  OAI21X1  g12954(.A0(new_n14696_), .A1(pi0165), .B0(new_n15390_), .Y(new_n15391_));
  OAI21X1  g12955(.A0(new_n14708_), .A1(pi0165), .B0(new_n14709_), .Y(new_n15392_));
  AND2X1   g12956(.A(new_n15392_), .B(new_n13675_), .Y(new_n15393_));
  AOI21X1  g12957(.A0(new_n14728_), .A1(pi0165), .B0(pi0038), .Y(new_n15394_));
  OAI21X1  g12958(.A0(new_n14716_), .A1(pi0165), .B0(new_n15394_), .Y(new_n15395_));
  OR2X1    g12959(.A(new_n12202_), .B(pi0165), .Y(new_n15396_));
  AOI21X1  g12960(.A0(new_n15396_), .A1(new_n14732_), .B0(new_n13675_), .Y(new_n15397_));
  AOI22X1  g12961(.A0(new_n15397_), .A1(new_n15395_), .B0(new_n15393_), .B1(new_n15391_), .Y(new_n15398_));
  OAI21X1  g12962(.A0(new_n14657_), .A1(new_n9941_), .B0(new_n13675_), .Y(new_n15399_));
  NOR2X1   g12963(.A(new_n15399_), .B(new_n14658_), .Y(new_n15400_));
  OAI21X1  g12964(.A0(new_n14675_), .A1(pi0774), .B0(pi0165), .Y(new_n15401_));
  AOI21X1  g12965(.A0(new_n13699_), .A1(pi0774), .B0(pi0687), .Y(new_n15402_));
  NAND2X1  g12966(.A(new_n15402_), .B(new_n15401_), .Y(new_n15403_));
  OAI22X1  g12967(.A0(new_n15403_), .A1(new_n15400_), .B0(new_n15398_), .B1(new_n13680_), .Y(new_n15404_));
  NAND2X1  g12968(.A(new_n15404_), .B(new_n7686_), .Y(new_n15405_));
  AOI21X1  g12969(.A0(new_n9580_), .A1(new_n9941_), .B0(pi0832), .Y(new_n15406_));
  AOI21X1  g12970(.A0(new_n15406_), .A1(new_n15405_), .B0(new_n15389_), .Y(po0322));
  OAI21X1  g12971(.A0(new_n14680_), .A1(new_n4464_), .B0(new_n14719_), .Y(new_n15408_));
  AOI21X1  g12972(.A0(new_n15408_), .A1(new_n14950_), .B0(new_n14667_), .Y(new_n15409_));
  MX2X1    g12973(.A(pi0947), .B(pi0166), .S0(new_n11953_), .Y(new_n15410_));
  OAI21X1  g12974(.A0(new_n15410_), .A1(new_n10137_), .B0(new_n2954_), .Y(new_n15411_));
  AOI21X1  g12975(.A0(new_n14652_), .A1(pi0166), .B0(new_n14954_), .Y(new_n15412_));
  OAI21X1  g12976(.A0(new_n15411_), .A1(new_n15409_), .B0(new_n15412_), .Y(new_n15413_));
  AND2X1   g12977(.A(new_n12010_), .B(new_n4464_), .Y(new_n15414_));
  INVX1    g12978(.A(new_n15414_), .Y(new_n15415_));
  AOI21X1  g12979(.A0(new_n15415_), .A1(new_n14687_), .B0(pi0299), .Y(new_n15416_));
  OR2X1    g12980(.A(new_n12064_), .B(pi0166), .Y(new_n15417_));
  AOI22X1  g12981(.A0(new_n15417_), .A1(new_n14917_), .B0(new_n15410_), .B1(new_n2970_), .Y(new_n15418_));
  OAI21X1  g12982(.A0(new_n15418_), .A1(pi0223), .B0(new_n15416_), .Y(new_n15419_));
  AND2X1   g12983(.A(new_n15419_), .B(pi0772), .Y(new_n15420_));
  AOI21X1  g12984(.A0(new_n12088_), .A1(new_n12068_), .B0(pi0772), .Y(new_n15421_));
  AND2X1   g12985(.A(new_n15421_), .B(pi0166), .Y(new_n15422_));
  OR2X1    g12986(.A(new_n15422_), .B(new_n2959_), .Y(new_n15423_));
  AOI21X1  g12987(.A0(new_n15420_), .A1(new_n15413_), .B0(new_n15423_), .Y(new_n15424_));
  AOI21X1  g12988(.A0(pi0947), .A1(pi0772), .B0(pi0039), .Y(new_n15425_));
  OAI22X1  g12989(.A0(new_n15425_), .A1(new_n14940_), .B0(new_n11947_), .B1(new_n4464_), .Y(new_n15426_));
  NAND2X1  g12990(.A(new_n15426_), .B(new_n2996_), .Y(new_n15427_));
  INVX1    g12991(.A(pi0727), .Y(new_n15428_));
  AND2X1   g12992(.A(pi0947), .B(pi0772), .Y(new_n15429_));
  INVX1    g12993(.A(new_n15429_), .Y(new_n15430_));
  AOI21X1  g12994(.A0(new_n15430_), .A1(new_n12202_), .B0(new_n2996_), .Y(new_n15431_));
  OAI21X1  g12995(.A0(new_n12572_), .A1(pi0166), .B0(new_n15431_), .Y(new_n15432_));
  AND2X1   g12996(.A(new_n15432_), .B(new_n15428_), .Y(new_n15433_));
  OAI21X1  g12997(.A0(new_n15427_), .A1(new_n15424_), .B0(new_n15433_), .Y(new_n15434_));
  MX2X1    g12998(.A(new_n5064_), .B(new_n4464_), .S0(new_n11953_), .Y(new_n15435_));
  AOI21X1  g12999(.A0(new_n15435_), .A1(new_n10136_), .B0(pi0215), .Y(new_n15436_));
  OAI21X1  g13000(.A0(new_n15408_), .A1(new_n14865_), .B0(new_n15436_), .Y(new_n15437_));
  OAI21X1  g13001(.A0(new_n14861_), .A1(pi0166), .B0(new_n14650_), .Y(new_n15438_));
  AND2X1   g13002(.A(new_n15438_), .B(pi0299), .Y(new_n15439_));
  AOI21X1  g13003(.A0(new_n15435_), .A1(new_n2970_), .B0(pi0223), .Y(new_n15440_));
  INVX1    g13004(.A(new_n15440_), .Y(new_n15441_));
  MX2X1    g13005(.A(new_n4464_), .B(new_n14638_), .S0(new_n12064_), .Y(new_n15442_));
  AOI21X1  g13006(.A0(new_n15442_), .A1(new_n14919_), .B0(new_n15441_), .Y(new_n15443_));
  OAI21X1  g13007(.A0(new_n12010_), .A1(new_n5064_), .B0(new_n4464_), .Y(new_n15444_));
  AND2X1   g13008(.A(new_n15444_), .B(new_n14688_), .Y(new_n15445_));
  INVX1    g13009(.A(new_n15445_), .Y(new_n15446_));
  NAND2X1  g13010(.A(new_n15446_), .B(new_n15416_), .Y(new_n15447_));
  OAI21X1  g13011(.A0(new_n15447_), .A1(new_n15443_), .B0(pi0772), .Y(new_n15448_));
  AOI21X1  g13012(.A0(new_n15439_), .A1(new_n15437_), .B0(new_n15448_), .Y(new_n15449_));
  OAI21X1  g13013(.A0(new_n14668_), .A1(new_n2971_), .B0(new_n15440_), .Y(new_n15450_));
  AOI21X1  g13014(.A0(new_n15442_), .A1(new_n2971_), .B0(new_n15450_), .Y(new_n15451_));
  NOR3X1   g13015(.A(new_n15451_), .B(new_n15445_), .C(pi0299), .Y(new_n15452_));
  AND2X1   g13016(.A(new_n15436_), .B(new_n14679_), .Y(new_n15453_));
  OAI21X1  g13017(.A0(new_n15438_), .A1(new_n14935_), .B0(pi0299), .Y(new_n15454_));
  AOI21X1  g13018(.A0(new_n15453_), .A1(new_n15408_), .B0(new_n15454_), .Y(new_n15455_));
  NOR3X1   g13019(.A(new_n15455_), .B(new_n15452_), .C(pi0772), .Y(new_n15456_));
  NOR3X1   g13020(.A(new_n15456_), .B(new_n15449_), .C(new_n2959_), .Y(new_n15457_));
  OAI21X1  g13021(.A0(new_n15426_), .A1(new_n14727_), .B0(new_n2996_), .Y(new_n15458_));
  NAND2X1  g13022(.A(new_n15425_), .B(new_n14946_), .Y(new_n15459_));
  AOI21X1  g13023(.A0(new_n12901_), .A1(new_n4464_), .B0(new_n2996_), .Y(new_n15460_));
  AOI21X1  g13024(.A0(new_n15460_), .A1(new_n15459_), .B0(new_n15428_), .Y(new_n15461_));
  OAI21X1  g13025(.A0(new_n15458_), .A1(new_n15457_), .B0(new_n15461_), .Y(new_n15462_));
  AOI21X1  g13026(.A0(new_n15462_), .A1(new_n15434_), .B0(new_n9580_), .Y(new_n15463_));
  OAI21X1  g13027(.A0(new_n7686_), .A1(pi0166), .B0(new_n12898_), .Y(new_n15464_));
  INVX1    g13028(.A(pi0772), .Y(new_n15465_));
  OAI21X1  g13029(.A0(new_n14590_), .A1(new_n15465_), .B0(new_n2739_), .Y(new_n15466_));
  AOI21X1  g13030(.A0(new_n14591_), .A1(pi0727), .B0(new_n15466_), .Y(new_n15467_));
  OAI21X1  g13031(.A0(new_n2739_), .A1(pi0166), .B0(pi0832), .Y(new_n15468_));
  OAI22X1  g13032(.A0(new_n15468_), .A1(new_n15467_), .B0(new_n15464_), .B1(new_n15463_), .Y(po0323));
  INVX1    g13033(.A(pi0705), .Y(new_n15470_));
  OAI22X1  g13034(.A0(new_n14638_), .A1(new_n15470_), .B0(new_n14590_), .B1(pi0768), .Y(new_n15471_));
  OAI21X1  g13035(.A0(new_n2739_), .A1(pi0167), .B0(pi0832), .Y(new_n15472_));
  AOI21X1  g13036(.A0(new_n15471_), .A1(new_n2739_), .B0(new_n15472_), .Y(new_n15473_));
  INVX1    g13037(.A(pi0768), .Y(new_n15474_));
  OAI21X1  g13038(.A0(new_n14729_), .A1(new_n7354_), .B0(new_n2996_), .Y(new_n15475_));
  AOI21X1  g13039(.A0(new_n14717_), .A1(new_n7354_), .B0(new_n15475_), .Y(new_n15476_));
  AOI21X1  g13040(.A0(new_n12901_), .A1(new_n7354_), .B0(new_n15039_), .Y(new_n15477_));
  NOR3X1   g13041(.A(new_n15477_), .B(new_n15476_), .C(new_n15474_), .Y(new_n15478_));
  OAI21X1  g13042(.A0(new_n15066_), .A1(new_n7354_), .B0(new_n2996_), .Y(new_n15479_));
  AOI21X1  g13043(.A0(new_n14695_), .A1(new_n7354_), .B0(new_n15479_), .Y(new_n15480_));
  OAI21X1  g13044(.A0(new_n14708_), .A1(pi0167), .B0(new_n14709_), .Y(new_n15481_));
  NAND2X1  g13045(.A(new_n15481_), .B(new_n15474_), .Y(new_n15482_));
  OAI21X1  g13046(.A0(new_n15482_), .A1(new_n15480_), .B0(pi0705), .Y(new_n15483_));
  OAI21X1  g13047(.A0(new_n14655_), .A1(new_n14642_), .B0(new_n7354_), .Y(new_n15484_));
  AOI21X1  g13048(.A0(new_n14674_), .A1(pi0167), .B0(pi0038), .Y(new_n15485_));
  NAND2X1  g13049(.A(new_n15485_), .B(new_n15484_), .Y(new_n15486_));
  OAI22X1  g13050(.A0(new_n14657_), .A1(new_n13402_), .B0(new_n12572_), .B1(pi0167), .Y(new_n15487_));
  NAND3X1  g13051(.A(new_n15487_), .B(new_n15486_), .C(new_n15474_), .Y(new_n15488_));
  NAND3X1  g13052(.A(new_n12574_), .B(pi0768), .C(new_n7354_), .Y(new_n15489_));
  AND2X1   g13053(.A(new_n15489_), .B(new_n15470_), .Y(new_n15490_));
  AOI21X1  g13054(.A0(new_n15490_), .A1(new_n15488_), .B0(new_n9580_), .Y(new_n15491_));
  OAI21X1  g13055(.A0(new_n15483_), .A1(new_n15478_), .B0(new_n15491_), .Y(new_n15492_));
  AOI21X1  g13056(.A0(new_n9580_), .A1(new_n7354_), .B0(pi0832), .Y(new_n15493_));
  AOI21X1  g13057(.A0(new_n15493_), .A1(new_n15492_), .B0(new_n15473_), .Y(po0324));
  INVX1    g13058(.A(pi0763), .Y(new_n15495_));
  OAI21X1  g13059(.A0(new_n14590_), .A1(new_n15495_), .B0(new_n2739_), .Y(new_n15496_));
  AOI21X1  g13060(.A0(new_n14591_), .A1(pi0699), .B0(new_n15496_), .Y(new_n15497_));
  OAI21X1  g13061(.A0(new_n2739_), .A1(new_n4351_), .B0(pi0832), .Y(new_n15498_));
  NAND3X1  g13062(.A(new_n11947_), .B(new_n15495_), .C(new_n2959_), .Y(new_n15499_));
  AOI22X1  g13063(.A0(new_n15499_), .A1(new_n14982_), .B0(new_n11948_), .B1(new_n4351_), .Y(new_n15500_));
  AOI21X1  g13064(.A0(new_n12082_), .A1(new_n5065_), .B0(new_n4351_), .Y(new_n15501_));
  NOR2X1   g13065(.A(new_n10136_), .B(new_n4351_), .Y(new_n15502_));
  AOI22X1  g13066(.A0(new_n15502_), .A1(new_n14866_), .B0(new_n12075_), .B1(new_n10137_), .Y(new_n15503_));
  INVX1    g13067(.A(new_n15503_), .Y(new_n15504_));
  OAI21X1  g13068(.A0(new_n11952_), .A1(new_n2740_), .B0(new_n4351_), .Y(new_n15505_));
  NAND3X1  g13069(.A(new_n15505_), .B(new_n14668_), .C(new_n10136_), .Y(new_n15506_));
  OAI21X1  g13070(.A0(new_n15506_), .A1(new_n14990_), .B0(new_n2954_), .Y(new_n15507_));
  OAI22X1  g13071(.A0(new_n15507_), .A1(new_n15504_), .B0(new_n15501_), .B1(new_n14985_), .Y(new_n15508_));
  OR2X1    g13072(.A(new_n14873_), .B(new_n4351_), .Y(new_n15509_));
  AOI22X1  g13073(.A0(new_n15509_), .A1(new_n14690_), .B0(new_n15508_), .B1(pi0299), .Y(new_n15510_));
  OR2X1    g13074(.A(new_n15510_), .B(new_n15495_), .Y(new_n15511_));
  AOI22X1  g13075(.A0(new_n15505_), .A1(new_n14721_), .B0(new_n14680_), .B1(new_n10137_), .Y(new_n15512_));
  AOI21X1  g13076(.A0(new_n15512_), .A1(new_n15503_), .B0(pi0215), .Y(new_n15513_));
  INVX1    g13077(.A(new_n15501_), .Y(new_n15514_));
  AOI21X1  g13078(.A0(new_n15514_), .A1(new_n14650_), .B0(new_n15000_), .Y(new_n15515_));
  OR2X1    g13079(.A(new_n15515_), .B(new_n14665_), .Y(new_n15516_));
  OAI21X1  g13080(.A0(new_n15516_), .A1(new_n15513_), .B0(pi0299), .Y(new_n15517_));
  OAI21X1  g13081(.A0(new_n14740_), .A1(pi0168), .B0(new_n14725_), .Y(new_n15518_));
  NAND3X1  g13082(.A(new_n15518_), .B(new_n15517_), .C(new_n15495_), .Y(new_n15519_));
  AND2X1   g13083(.A(new_n15519_), .B(pi0039), .Y(new_n15520_));
  AOI22X1  g13084(.A0(new_n15520_), .A1(new_n15511_), .B0(new_n15500_), .B1(new_n14981_), .Y(new_n15521_));
  AOI21X1  g13085(.A0(pi0947), .A1(new_n15495_), .B0(pi0039), .Y(new_n15522_));
  AOI21X1  g13086(.A0(new_n15522_), .A1(new_n14810_), .B0(new_n2996_), .Y(new_n15523_));
  OAI21X1  g13087(.A0(new_n12202_), .A1(pi0168), .B0(new_n15523_), .Y(new_n15524_));
  OAI21X1  g13088(.A0(new_n15521_), .A1(pi0038), .B0(new_n15524_), .Y(new_n15525_));
  OAI21X1  g13089(.A0(new_n14740_), .A1(pi0168), .B0(new_n14663_), .Y(new_n15526_));
  NAND3X1  g13090(.A(new_n15506_), .B(new_n15503_), .C(new_n14894_), .Y(new_n15527_));
  AOI21X1  g13091(.A0(new_n15514_), .A1(new_n14652_), .B0(new_n2953_), .Y(new_n15528_));
  AOI21X1  g13092(.A0(new_n15528_), .A1(new_n15527_), .B0(new_n15495_), .Y(new_n15529_));
  NAND2X1  g13093(.A(new_n15529_), .B(new_n15526_), .Y(new_n15530_));
  NOR2X1   g13094(.A(pi0763), .B(pi0168), .Y(new_n15531_));
  AOI21X1  g13095(.A0(new_n15531_), .A1(new_n12089_), .B0(new_n2959_), .Y(new_n15532_));
  OR2X1    g13096(.A(new_n15500_), .B(pi0038), .Y(new_n15533_));
  AOI21X1  g13097(.A0(new_n15532_), .A1(new_n15530_), .B0(new_n15533_), .Y(new_n15534_));
  INVX1    g13098(.A(pi0699), .Y(new_n15535_));
  AOI21X1  g13099(.A0(new_n4995_), .A1(new_n2739_), .B0(new_n4351_), .Y(new_n15536_));
  OAI21X1  g13100(.A0(new_n15496_), .A1(new_n14411_), .B0(pi0038), .Y(new_n15537_));
  OAI21X1  g13101(.A0(new_n15537_), .A1(new_n15536_), .B0(new_n15535_), .Y(new_n15538_));
  OAI21X1  g13102(.A0(new_n15538_), .A1(new_n15534_), .B0(new_n14757_), .Y(new_n15539_));
  AOI21X1  g13103(.A0(new_n15525_), .A1(pi0699), .B0(new_n15539_), .Y(new_n15540_));
  AOI21X1  g13104(.A0(new_n5117_), .A1(new_n3129_), .B0(pi0168), .Y(new_n15541_));
  NOR3X1   g13105(.A(new_n15541_), .B(new_n15540_), .C(pi0057), .Y(new_n15542_));
  OAI21X1  g13106(.A0(new_n4351_), .A1(new_n2436_), .B0(new_n12898_), .Y(new_n15543_));
  OAI22X1  g13107(.A0(new_n15543_), .A1(new_n15542_), .B0(new_n15498_), .B1(new_n15497_), .Y(po0325));
  INVX1    g13108(.A(pi0746), .Y(new_n15545_));
  OAI21X1  g13109(.A0(new_n14590_), .A1(new_n15545_), .B0(new_n2739_), .Y(new_n15546_));
  AOI21X1  g13110(.A0(new_n14591_), .A1(pi0729), .B0(new_n15546_), .Y(new_n15547_));
  OAI21X1  g13111(.A0(new_n2739_), .A1(new_n4210_), .B0(pi0832), .Y(new_n15548_));
  NAND3X1  g13112(.A(new_n11947_), .B(new_n15545_), .C(new_n2959_), .Y(new_n15549_));
  AOI22X1  g13113(.A0(new_n15549_), .A1(new_n14982_), .B0(new_n11948_), .B1(new_n4210_), .Y(new_n15550_));
  AOI21X1  g13114(.A0(new_n12082_), .A1(new_n5065_), .B0(new_n4210_), .Y(new_n15551_));
  NOR2X1   g13115(.A(new_n10136_), .B(new_n4210_), .Y(new_n15552_));
  AOI22X1  g13116(.A0(new_n15552_), .A1(new_n14866_), .B0(new_n12075_), .B1(new_n10137_), .Y(new_n15553_));
  INVX1    g13117(.A(new_n15553_), .Y(new_n15554_));
  OAI21X1  g13118(.A0(new_n11952_), .A1(new_n2740_), .B0(new_n4210_), .Y(new_n15555_));
  NAND3X1  g13119(.A(new_n15555_), .B(new_n14668_), .C(new_n10136_), .Y(new_n15556_));
  OAI21X1  g13120(.A0(new_n15556_), .A1(new_n14990_), .B0(new_n2954_), .Y(new_n15557_));
  OAI22X1  g13121(.A0(new_n15557_), .A1(new_n15554_), .B0(new_n15551_), .B1(new_n14985_), .Y(new_n15558_));
  OR2X1    g13122(.A(new_n14873_), .B(new_n4210_), .Y(new_n15559_));
  AOI22X1  g13123(.A0(new_n15559_), .A1(new_n14690_), .B0(new_n15558_), .B1(pi0299), .Y(new_n15560_));
  OR2X1    g13124(.A(new_n15560_), .B(new_n15545_), .Y(new_n15561_));
  AOI22X1  g13125(.A0(new_n15555_), .A1(new_n14721_), .B0(new_n14680_), .B1(new_n10137_), .Y(new_n15562_));
  AOI21X1  g13126(.A0(new_n15562_), .A1(new_n15553_), .B0(pi0215), .Y(new_n15563_));
  INVX1    g13127(.A(new_n15551_), .Y(new_n15564_));
  AOI21X1  g13128(.A0(new_n15564_), .A1(new_n14650_), .B0(new_n15000_), .Y(new_n15565_));
  OR2X1    g13129(.A(new_n15565_), .B(new_n14665_), .Y(new_n15566_));
  OAI21X1  g13130(.A0(new_n15566_), .A1(new_n15563_), .B0(pi0299), .Y(new_n15567_));
  OAI21X1  g13131(.A0(new_n14740_), .A1(pi0169), .B0(new_n14725_), .Y(new_n15568_));
  NAND3X1  g13132(.A(new_n15568_), .B(new_n15567_), .C(new_n15545_), .Y(new_n15569_));
  AND2X1   g13133(.A(new_n15569_), .B(pi0039), .Y(new_n15570_));
  AOI22X1  g13134(.A0(new_n15570_), .A1(new_n15561_), .B0(new_n15550_), .B1(new_n14981_), .Y(new_n15571_));
  AOI21X1  g13135(.A0(pi0947), .A1(new_n15545_), .B0(pi0039), .Y(new_n15572_));
  AOI21X1  g13136(.A0(new_n15572_), .A1(new_n14810_), .B0(new_n2996_), .Y(new_n15573_));
  OAI21X1  g13137(.A0(new_n12202_), .A1(pi0169), .B0(new_n15573_), .Y(new_n15574_));
  OAI21X1  g13138(.A0(new_n15571_), .A1(pi0038), .B0(new_n15574_), .Y(new_n15575_));
  OAI21X1  g13139(.A0(new_n14740_), .A1(pi0169), .B0(new_n14663_), .Y(new_n15576_));
  NAND3X1  g13140(.A(new_n15556_), .B(new_n15553_), .C(new_n14894_), .Y(new_n15577_));
  AOI21X1  g13141(.A0(new_n15564_), .A1(new_n14652_), .B0(new_n2953_), .Y(new_n15578_));
  AOI21X1  g13142(.A0(new_n15578_), .A1(new_n15577_), .B0(new_n15545_), .Y(new_n15579_));
  NAND2X1  g13143(.A(new_n15579_), .B(new_n15576_), .Y(new_n15580_));
  NOR2X1   g13144(.A(pi0746), .B(pi0169), .Y(new_n15581_));
  AOI21X1  g13145(.A0(new_n15581_), .A1(new_n12089_), .B0(new_n2959_), .Y(new_n15582_));
  OR2X1    g13146(.A(new_n15550_), .B(pi0038), .Y(new_n15583_));
  AOI21X1  g13147(.A0(new_n15582_), .A1(new_n15580_), .B0(new_n15583_), .Y(new_n15584_));
  INVX1    g13148(.A(pi0729), .Y(new_n15585_));
  AOI21X1  g13149(.A0(new_n4995_), .A1(new_n2739_), .B0(new_n4210_), .Y(new_n15586_));
  OAI21X1  g13150(.A0(new_n15546_), .A1(new_n14411_), .B0(pi0038), .Y(new_n15587_));
  OAI21X1  g13151(.A0(new_n15587_), .A1(new_n15586_), .B0(new_n15585_), .Y(new_n15588_));
  OAI21X1  g13152(.A0(new_n15588_), .A1(new_n15584_), .B0(new_n14757_), .Y(new_n15589_));
  AOI21X1  g13153(.A0(new_n15575_), .A1(pi0729), .B0(new_n15589_), .Y(new_n15590_));
  AOI21X1  g13154(.A0(new_n5117_), .A1(new_n3129_), .B0(pi0169), .Y(new_n15591_));
  NOR3X1   g13155(.A(new_n15591_), .B(new_n15590_), .C(pi0057), .Y(new_n15592_));
  OAI21X1  g13156(.A0(new_n4210_), .A1(new_n2436_), .B0(new_n12898_), .Y(new_n15593_));
  OAI22X1  g13157(.A0(new_n15593_), .A1(new_n15592_), .B0(new_n15548_), .B1(new_n15547_), .Y(po0326));
  INVX1    g13158(.A(pi0748), .Y(new_n15595_));
  OAI21X1  g13159(.A0(new_n14590_), .A1(new_n15595_), .B0(new_n2739_), .Y(new_n15596_));
  AOI21X1  g13160(.A0(new_n14591_), .A1(pi0730), .B0(new_n15596_), .Y(new_n15597_));
  OAI21X1  g13161(.A0(new_n2739_), .A1(new_n3917_), .B0(pi0832), .Y(new_n15598_));
  INVX1    g13162(.A(new_n14877_), .Y(new_n15599_));
  NOR2X1   g13163(.A(new_n10136_), .B(new_n3917_), .Y(new_n15600_));
  AOI22X1  g13164(.A0(new_n15600_), .A1(new_n14866_), .B0(new_n12075_), .B1(new_n10137_), .Y(new_n15601_));
  OAI21X1  g13165(.A0(new_n12012_), .A1(pi0170), .B0(new_n14721_), .Y(new_n15602_));
  NAND3X1  g13166(.A(new_n15602_), .B(new_n15601_), .C(new_n15599_), .Y(new_n15603_));
  AOI21X1  g13167(.A0(new_n12082_), .A1(new_n5065_), .B0(new_n3917_), .Y(new_n15604_));
  OAI21X1  g13168(.A0(new_n15604_), .A1(new_n14985_), .B0(new_n14699_), .Y(new_n15605_));
  NAND2X1  g13169(.A(new_n15605_), .B(new_n14666_), .Y(new_n15606_));
  AOI21X1  g13170(.A0(new_n15603_), .A1(new_n2954_), .B0(new_n15606_), .Y(new_n15607_));
  OAI21X1  g13171(.A0(new_n14740_), .A1(pi0170), .B0(new_n2953_), .Y(new_n15608_));
  OAI22X1  g13172(.A0(new_n15608_), .A1(new_n14724_), .B0(new_n15607_), .B1(new_n2953_), .Y(new_n15609_));
  OR2X1    g13173(.A(new_n11947_), .B(pi0170), .Y(new_n15610_));
  AOI22X1  g13174(.A0(new_n15610_), .A1(new_n14856_), .B0(new_n15609_), .B1(pi0039), .Y(new_n15611_));
  OR2X1    g13175(.A(new_n12202_), .B(pi0170), .Y(new_n15612_));
  AOI21X1  g13176(.A0(new_n15612_), .A1(new_n14732_), .B0(pi0748), .Y(new_n15613_));
  OAI21X1  g13177(.A0(new_n15611_), .A1(pi0038), .B0(new_n15613_), .Y(new_n15614_));
  OAI21X1  g13178(.A0(new_n14873_), .A1(new_n3917_), .B0(new_n14690_), .Y(new_n15615_));
  INVX1    g13179(.A(new_n15601_), .Y(new_n15616_));
  OAI21X1  g13180(.A0(new_n12012_), .A1(pi0170), .B0(new_n14895_), .Y(new_n15617_));
  OAI21X1  g13181(.A0(new_n15617_), .A1(new_n14990_), .B0(new_n2954_), .Y(new_n15618_));
  OAI22X1  g13182(.A0(new_n15618_), .A1(new_n15616_), .B0(new_n15604_), .B1(new_n14985_), .Y(new_n15619_));
  AOI21X1  g13183(.A0(new_n15619_), .A1(pi0299), .B0(new_n2959_), .Y(new_n15620_));
  AOI22X1  g13184(.A0(new_n15620_), .A1(new_n15615_), .B0(new_n15610_), .B1(new_n14694_), .Y(new_n15621_));
  AOI21X1  g13185(.A0(new_n15612_), .A1(new_n14709_), .B0(new_n15595_), .Y(new_n15622_));
  OAI21X1  g13186(.A0(new_n15621_), .A1(pi0038), .B0(new_n15622_), .Y(new_n15623_));
  NAND3X1  g13187(.A(new_n15623_), .B(new_n15614_), .C(pi0730), .Y(new_n15624_));
  NAND2X1  g13188(.A(new_n15617_), .B(new_n15601_), .Y(new_n15625_));
  NOR3X1   g13189(.A(new_n15625_), .B(new_n14647_), .C(pi0215), .Y(new_n15626_));
  OAI21X1  g13190(.A0(new_n14861_), .A1(new_n3917_), .B0(new_n14652_), .Y(new_n15627_));
  NAND2X1  g13191(.A(new_n15627_), .B(pi0299), .Y(new_n15628_));
  OAI22X1  g13192(.A0(new_n15628_), .A1(new_n15626_), .B0(new_n15608_), .B1(new_n14662_), .Y(new_n15629_));
  AOI22X1  g13193(.A0(new_n15629_), .A1(pi0039), .B0(new_n15610_), .B1(new_n14661_), .Y(new_n15630_));
  OAI22X1  g13194(.A0(new_n14657_), .A1(new_n13402_), .B0(new_n12572_), .B1(pi0170), .Y(new_n15631_));
  AND2X1   g13195(.A(new_n15631_), .B(pi0748), .Y(new_n15632_));
  OAI21X1  g13196(.A0(new_n15630_), .A1(pi0038), .B0(new_n15632_), .Y(new_n15633_));
  NOR2X1   g13197(.A(pi0748), .B(pi0170), .Y(new_n15634_));
  AOI21X1  g13198(.A0(new_n15634_), .A1(new_n12574_), .B0(pi0730), .Y(new_n15635_));
  AOI21X1  g13199(.A0(new_n15635_), .A1(new_n15633_), .B0(new_n14758_), .Y(new_n15636_));
  OAI21X1  g13200(.A0(new_n14757_), .A1(pi0170), .B0(new_n2436_), .Y(new_n15637_));
  AOI21X1  g13201(.A0(new_n15636_), .A1(new_n15624_), .B0(new_n15637_), .Y(new_n15638_));
  OAI21X1  g13202(.A0(new_n3917_), .A1(new_n2436_), .B0(new_n12898_), .Y(new_n15639_));
  OAI22X1  g13203(.A0(new_n15639_), .A1(new_n15638_), .B0(new_n15598_), .B1(new_n15597_), .Y(po0327));
  INVX1    g13204(.A(pi0764), .Y(new_n15641_));
  OAI21X1  g13205(.A0(new_n14590_), .A1(new_n15641_), .B0(new_n2739_), .Y(new_n15642_));
  AOI21X1  g13206(.A0(new_n14591_), .A1(pi0691), .B0(new_n15642_), .Y(new_n15643_));
  OAI21X1  g13207(.A0(new_n2739_), .A1(new_n3774_), .B0(pi0832), .Y(new_n15644_));
  NAND3X1  g13208(.A(new_n11947_), .B(new_n15641_), .C(new_n2959_), .Y(new_n15645_));
  AOI22X1  g13209(.A0(new_n15645_), .A1(new_n14982_), .B0(new_n11948_), .B1(new_n3774_), .Y(new_n15646_));
  AOI21X1  g13210(.A0(new_n12082_), .A1(new_n5065_), .B0(new_n3774_), .Y(new_n15647_));
  NOR2X1   g13211(.A(new_n10136_), .B(new_n3774_), .Y(new_n15648_));
  AOI22X1  g13212(.A0(new_n15648_), .A1(new_n14866_), .B0(new_n12075_), .B1(new_n10137_), .Y(new_n15649_));
  INVX1    g13213(.A(new_n15649_), .Y(new_n15650_));
  OAI21X1  g13214(.A0(new_n11952_), .A1(new_n2740_), .B0(new_n3774_), .Y(new_n15651_));
  NAND3X1  g13215(.A(new_n15651_), .B(new_n14668_), .C(new_n10136_), .Y(new_n15652_));
  OAI21X1  g13216(.A0(new_n15652_), .A1(new_n14990_), .B0(new_n2954_), .Y(new_n15653_));
  OAI22X1  g13217(.A0(new_n15653_), .A1(new_n15650_), .B0(new_n15647_), .B1(new_n14985_), .Y(new_n15654_));
  OR2X1    g13218(.A(new_n14873_), .B(new_n3774_), .Y(new_n15655_));
  AOI22X1  g13219(.A0(new_n15655_), .A1(new_n14690_), .B0(new_n15654_), .B1(pi0299), .Y(new_n15656_));
  OR2X1    g13220(.A(new_n15656_), .B(new_n15641_), .Y(new_n15657_));
  AOI22X1  g13221(.A0(new_n15651_), .A1(new_n14721_), .B0(new_n14680_), .B1(new_n10137_), .Y(new_n15658_));
  AOI21X1  g13222(.A0(new_n15658_), .A1(new_n15649_), .B0(pi0215), .Y(new_n15659_));
  INVX1    g13223(.A(new_n15647_), .Y(new_n15660_));
  AOI21X1  g13224(.A0(new_n15660_), .A1(new_n14650_), .B0(new_n15000_), .Y(new_n15661_));
  OR2X1    g13225(.A(new_n15661_), .B(new_n14665_), .Y(new_n15662_));
  OAI21X1  g13226(.A0(new_n15662_), .A1(new_n15659_), .B0(pi0299), .Y(new_n15663_));
  OAI21X1  g13227(.A0(new_n14740_), .A1(pi0171), .B0(new_n14725_), .Y(new_n15664_));
  NAND3X1  g13228(.A(new_n15664_), .B(new_n15663_), .C(new_n15641_), .Y(new_n15665_));
  AND2X1   g13229(.A(new_n15665_), .B(pi0039), .Y(new_n15666_));
  AOI22X1  g13230(.A0(new_n15666_), .A1(new_n15657_), .B0(new_n15646_), .B1(new_n14981_), .Y(new_n15667_));
  AOI21X1  g13231(.A0(pi0947), .A1(new_n15641_), .B0(pi0039), .Y(new_n15668_));
  AOI21X1  g13232(.A0(new_n15668_), .A1(new_n14810_), .B0(new_n2996_), .Y(new_n15669_));
  OAI21X1  g13233(.A0(new_n12202_), .A1(pi0171), .B0(new_n15669_), .Y(new_n15670_));
  OAI21X1  g13234(.A0(new_n15667_), .A1(pi0038), .B0(new_n15670_), .Y(new_n15671_));
  OAI21X1  g13235(.A0(new_n14740_), .A1(pi0171), .B0(new_n14663_), .Y(new_n15672_));
  NAND3X1  g13236(.A(new_n15652_), .B(new_n15649_), .C(new_n14894_), .Y(new_n15673_));
  AOI21X1  g13237(.A0(new_n15660_), .A1(new_n14652_), .B0(new_n2953_), .Y(new_n15674_));
  AOI21X1  g13238(.A0(new_n15674_), .A1(new_n15673_), .B0(new_n15641_), .Y(new_n15675_));
  NAND2X1  g13239(.A(new_n15675_), .B(new_n15672_), .Y(new_n15676_));
  NOR2X1   g13240(.A(pi0764), .B(pi0171), .Y(new_n15677_));
  AOI21X1  g13241(.A0(new_n15677_), .A1(new_n12089_), .B0(new_n2959_), .Y(new_n15678_));
  OR2X1    g13242(.A(new_n15646_), .B(pi0038), .Y(new_n15679_));
  AOI21X1  g13243(.A0(new_n15678_), .A1(new_n15676_), .B0(new_n15679_), .Y(new_n15680_));
  INVX1    g13244(.A(pi0691), .Y(new_n15681_));
  AOI21X1  g13245(.A0(new_n4995_), .A1(new_n2739_), .B0(new_n3774_), .Y(new_n15682_));
  OAI21X1  g13246(.A0(new_n15642_), .A1(new_n14411_), .B0(pi0038), .Y(new_n15683_));
  OAI21X1  g13247(.A0(new_n15683_), .A1(new_n15682_), .B0(new_n15681_), .Y(new_n15684_));
  OAI21X1  g13248(.A0(new_n15684_), .A1(new_n15680_), .B0(new_n14757_), .Y(new_n15685_));
  AOI21X1  g13249(.A0(new_n15671_), .A1(pi0691), .B0(new_n15685_), .Y(new_n15686_));
  AOI21X1  g13250(.A0(new_n5117_), .A1(new_n3129_), .B0(pi0171), .Y(new_n15687_));
  NOR3X1   g13251(.A(new_n15687_), .B(new_n15686_), .C(pi0057), .Y(new_n15688_));
  OAI21X1  g13252(.A0(new_n3774_), .A1(new_n2436_), .B0(new_n12898_), .Y(new_n15689_));
  OAI22X1  g13253(.A0(new_n15689_), .A1(new_n15688_), .B0(new_n15644_), .B1(new_n15643_), .Y(po0328));
  NAND2X1  g13254(.A(pi0947), .B(pi0739), .Y(new_n15691_));
  NAND2X1  g13255(.A(new_n15691_), .B(new_n2739_), .Y(new_n15692_));
  AOI21X1  g13256(.A0(new_n14591_), .A1(pi0690), .B0(new_n15692_), .Y(new_n15693_));
  OAI21X1  g13257(.A0(new_n2739_), .A1(new_n3601_), .B0(pi0832), .Y(new_n15694_));
  OAI21X1  g13258(.A0(new_n15691_), .A1(new_n11948_), .B0(new_n2959_), .Y(new_n15695_));
  AOI21X1  g13259(.A0(new_n11948_), .A1(new_n3601_), .B0(new_n15695_), .Y(new_n15696_));
  INVX1    g13260(.A(pi0739), .Y(new_n15697_));
  AOI21X1  g13261(.A0(new_n12082_), .A1(new_n5065_), .B0(new_n3601_), .Y(new_n15698_));
  NOR2X1   g13262(.A(new_n10136_), .B(new_n3601_), .Y(new_n15699_));
  AOI22X1  g13263(.A0(new_n15699_), .A1(new_n14866_), .B0(new_n12075_), .B1(new_n10137_), .Y(new_n15700_));
  INVX1    g13264(.A(new_n15700_), .Y(new_n15701_));
  OAI21X1  g13265(.A0(new_n11952_), .A1(new_n2740_), .B0(new_n3601_), .Y(new_n15702_));
  NAND3X1  g13266(.A(new_n15702_), .B(new_n14668_), .C(new_n10136_), .Y(new_n15703_));
  OAI21X1  g13267(.A0(new_n15703_), .A1(new_n14990_), .B0(new_n2954_), .Y(new_n15704_));
  OAI22X1  g13268(.A0(new_n15704_), .A1(new_n15701_), .B0(new_n15698_), .B1(new_n14985_), .Y(new_n15705_));
  OR2X1    g13269(.A(new_n14873_), .B(new_n3601_), .Y(new_n15706_));
  AOI22X1  g13270(.A0(new_n15706_), .A1(new_n14690_), .B0(new_n15705_), .B1(pi0299), .Y(new_n15707_));
  OR2X1    g13271(.A(new_n15707_), .B(new_n15697_), .Y(new_n15708_));
  AOI22X1  g13272(.A0(new_n15702_), .A1(new_n14721_), .B0(new_n14680_), .B1(new_n10137_), .Y(new_n15709_));
  AOI21X1  g13273(.A0(new_n15709_), .A1(new_n15700_), .B0(pi0215), .Y(new_n15710_));
  INVX1    g13274(.A(new_n15698_), .Y(new_n15711_));
  AOI21X1  g13275(.A0(new_n15711_), .A1(new_n14650_), .B0(new_n15000_), .Y(new_n15712_));
  OR2X1    g13276(.A(new_n15712_), .B(new_n14665_), .Y(new_n15713_));
  OAI21X1  g13277(.A0(new_n15713_), .A1(new_n15710_), .B0(pi0299), .Y(new_n15714_));
  OAI21X1  g13278(.A0(new_n14740_), .A1(pi0172), .B0(new_n14725_), .Y(new_n15715_));
  NAND3X1  g13279(.A(new_n15715_), .B(new_n15714_), .C(new_n15697_), .Y(new_n15716_));
  AND2X1   g13280(.A(new_n15716_), .B(pi0039), .Y(new_n15717_));
  AOI22X1  g13281(.A0(new_n15717_), .A1(new_n15708_), .B0(new_n15696_), .B1(new_n14981_), .Y(new_n15718_));
  AOI21X1  g13282(.A0(pi0947), .A1(new_n15697_), .B0(pi0039), .Y(new_n15719_));
  AOI21X1  g13283(.A0(new_n15719_), .A1(new_n14810_), .B0(new_n2996_), .Y(new_n15720_));
  OAI21X1  g13284(.A0(new_n12202_), .A1(pi0172), .B0(new_n15720_), .Y(new_n15721_));
  OAI21X1  g13285(.A0(new_n15718_), .A1(pi0038), .B0(new_n15721_), .Y(new_n15722_));
  OAI21X1  g13286(.A0(new_n14740_), .A1(pi0172), .B0(new_n14663_), .Y(new_n15723_));
  NAND3X1  g13287(.A(new_n15703_), .B(new_n15700_), .C(new_n14894_), .Y(new_n15724_));
  AOI21X1  g13288(.A0(new_n15711_), .A1(new_n14652_), .B0(new_n2953_), .Y(new_n15725_));
  AOI21X1  g13289(.A0(new_n15725_), .A1(new_n15724_), .B0(new_n15697_), .Y(new_n15726_));
  NAND2X1  g13290(.A(new_n15726_), .B(new_n15723_), .Y(new_n15727_));
  NOR2X1   g13291(.A(pi0739), .B(pi0172), .Y(new_n15728_));
  AOI21X1  g13292(.A0(new_n15728_), .A1(new_n12089_), .B0(new_n2959_), .Y(new_n15729_));
  OR2X1    g13293(.A(new_n15696_), .B(pi0038), .Y(new_n15730_));
  AOI21X1  g13294(.A0(new_n15729_), .A1(new_n15727_), .B0(new_n15730_), .Y(new_n15731_));
  INVX1    g13295(.A(pi0690), .Y(new_n15732_));
  AOI21X1  g13296(.A0(new_n4995_), .A1(new_n2739_), .B0(new_n3601_), .Y(new_n15733_));
  OAI21X1  g13297(.A0(new_n15692_), .A1(new_n14411_), .B0(pi0038), .Y(new_n15734_));
  OAI21X1  g13298(.A0(new_n15734_), .A1(new_n15733_), .B0(new_n15732_), .Y(new_n15735_));
  OAI21X1  g13299(.A0(new_n15735_), .A1(new_n15731_), .B0(new_n14757_), .Y(new_n15736_));
  AOI21X1  g13300(.A0(new_n15722_), .A1(pi0690), .B0(new_n15736_), .Y(new_n15737_));
  AOI21X1  g13301(.A0(new_n5117_), .A1(new_n3129_), .B0(pi0172), .Y(new_n15738_));
  NOR3X1   g13302(.A(new_n15738_), .B(new_n15737_), .C(pi0057), .Y(new_n15739_));
  OAI21X1  g13303(.A0(new_n3601_), .A1(new_n2436_), .B0(new_n12898_), .Y(new_n15740_));
  OAI22X1  g13304(.A0(new_n15740_), .A1(new_n15739_), .B0(new_n15694_), .B1(new_n15693_), .Y(po0329));
  AOI21X1  g13305(.A0(new_n13699_), .A1(new_n3129_), .B0(pi0173), .Y(new_n15742_));
  INVX1    g13306(.A(new_n15742_), .Y(new_n15743_));
  OAI21X1  g13307(.A0(new_n3810_), .A1(pi0723), .B0(new_n15742_), .Y(new_n15744_));
  AOI21X1  g13308(.A0(new_n12955_), .A1(pi0173), .B0(pi0038), .Y(new_n15745_));
  OAI22X1  g13309(.A0(new_n15745_), .A1(new_n3810_), .B0(new_n12953_), .B1(pi0173), .Y(new_n15746_));
  OAI21X1  g13310(.A0(new_n12202_), .A1(pi0173), .B0(new_n12567_), .Y(new_n15747_));
  NAND3X1  g13311(.A(new_n15747_), .B(new_n15746_), .C(new_n14886_), .Y(new_n15748_));
  AND2X1   g13312(.A(new_n15748_), .B(new_n15744_), .Y(new_n15749_));
  AOI21X1  g13313(.A0(new_n15742_), .A1(new_n12493_), .B0(new_n12494_), .Y(new_n15750_));
  OAI21X1  g13314(.A0(new_n15749_), .A1(new_n12493_), .B0(new_n15750_), .Y(new_n15751_));
  AOI21X1  g13315(.A0(new_n15742_), .A1(pi0625), .B0(pi1153), .Y(new_n15752_));
  OAI21X1  g13316(.A0(new_n15749_), .A1(pi0625), .B0(new_n15752_), .Y(new_n15753_));
  AOI21X1  g13317(.A0(new_n15753_), .A1(new_n15751_), .B0(new_n11889_), .Y(new_n15754_));
  AOI21X1  g13318(.A0(new_n15749_), .A1(new_n11889_), .B0(new_n15754_), .Y(new_n15755_));
  MX2X1    g13319(.A(new_n15755_), .B(new_n15742_), .S0(new_n12618_), .Y(new_n15756_));
  MX2X1    g13320(.A(new_n15756_), .B(new_n15742_), .S0(new_n12641_), .Y(new_n15757_));
  MX2X1    g13321(.A(new_n15757_), .B(new_n15742_), .S0(new_n12659_), .Y(new_n15758_));
  INVX1    g13322(.A(new_n15758_), .Y(new_n15759_));
  MX2X1    g13323(.A(new_n15759_), .B(new_n15743_), .S0(new_n12691_), .Y(new_n15760_));
  AND2X1   g13324(.A(new_n15760_), .B(new_n11884_), .Y(new_n15761_));
  AOI21X1  g13325(.A0(new_n15742_), .A1(new_n12683_), .B0(new_n12684_), .Y(new_n15762_));
  OAI21X1  g13326(.A0(new_n15760_), .A1(new_n12683_), .B0(new_n15762_), .Y(new_n15763_));
  AOI21X1  g13327(.A0(new_n15742_), .A1(pi0628), .B0(pi1156), .Y(new_n15764_));
  OAI21X1  g13328(.A0(new_n15760_), .A1(pi0628), .B0(new_n15764_), .Y(new_n15765_));
  AOI21X1  g13329(.A0(new_n15765_), .A1(new_n15763_), .B0(new_n11884_), .Y(new_n15766_));
  NOR2X1   g13330(.A(new_n15766_), .B(new_n15761_), .Y(new_n15767_));
  MX2X1    g13331(.A(new_n15767_), .B(new_n15742_), .S0(pi0647), .Y(new_n15768_));
  MX2X1    g13332(.A(new_n15767_), .B(new_n15742_), .S0(new_n12705_), .Y(new_n15769_));
  MX2X1    g13333(.A(new_n15769_), .B(new_n15768_), .S0(new_n12706_), .Y(new_n15770_));
  NOR3X1   g13334(.A(new_n15766_), .B(new_n15761_), .C(pi0787), .Y(new_n15771_));
  AOI21X1  g13335(.A0(new_n15770_), .A1(pi0787), .B0(new_n15771_), .Y(new_n15772_));
  OAI21X1  g13336(.A0(new_n15772_), .A1(pi0644), .B0(pi0715), .Y(new_n15773_));
  AOI21X1  g13337(.A0(new_n12090_), .A1(new_n9989_), .B0(new_n14858_), .Y(new_n15774_));
  NOR2X1   g13338(.A(pi0745), .B(pi0173), .Y(new_n15775_));
  INVX1    g13339(.A(new_n15775_), .Y(new_n15776_));
  OAI22X1  g13340(.A0(new_n15776_), .A1(new_n12910_), .B0(new_n12199_), .B1(new_n9989_), .Y(new_n15777_));
  OAI21X1  g13341(.A0(new_n15777_), .A1(new_n15774_), .B0(new_n2996_), .Y(new_n15778_));
  AOI21X1  g13342(.A0(new_n12901_), .A1(new_n9989_), .B0(new_n2996_), .Y(new_n15779_));
  OAI21X1  g13343(.A0(new_n14342_), .A1(pi0745), .B0(new_n15779_), .Y(new_n15780_));
  AND2X1   g13344(.A(new_n15780_), .B(new_n15778_), .Y(new_n15781_));
  MX2X1    g13345(.A(new_n15781_), .B(new_n9989_), .S0(new_n3810_), .Y(new_n15782_));
  INVX1    g13346(.A(new_n15782_), .Y(new_n15783_));
  MX2X1    g13347(.A(new_n15783_), .B(new_n15743_), .S0(new_n12601_), .Y(new_n15784_));
  NOR2X1   g13348(.A(new_n15782_), .B(new_n12601_), .Y(new_n15785_));
  AOI22X1  g13349(.A0(new_n15785_), .A1(pi0609), .B0(new_n15743_), .B1(new_n13430_), .Y(new_n15786_));
  OR2X1    g13350(.A(new_n15786_), .B(new_n12591_), .Y(new_n15787_));
  AOI22X1  g13351(.A0(new_n15785_), .A1(new_n12590_), .B0(new_n15743_), .B1(new_n13436_), .Y(new_n15788_));
  OR2X1    g13352(.A(new_n15788_), .B(pi1155), .Y(new_n15789_));
  NAND2X1  g13353(.A(new_n15789_), .B(new_n15787_), .Y(new_n15790_));
  MX2X1    g13354(.A(new_n15790_), .B(new_n15784_), .S0(new_n11888_), .Y(new_n15791_));
  AOI21X1  g13355(.A0(new_n15742_), .A1(new_n12614_), .B0(new_n12615_), .Y(new_n15792_));
  OAI21X1  g13356(.A0(new_n15791_), .A1(new_n12614_), .B0(new_n15792_), .Y(new_n15793_));
  AOI21X1  g13357(.A0(new_n15742_), .A1(pi0618), .B0(pi1154), .Y(new_n15794_));
  OAI21X1  g13358(.A0(new_n15791_), .A1(pi0618), .B0(new_n15794_), .Y(new_n15795_));
  NAND2X1  g13359(.A(new_n15795_), .B(new_n15793_), .Y(new_n15796_));
  MX2X1    g13360(.A(new_n15796_), .B(new_n15791_), .S0(new_n11887_), .Y(new_n15797_));
  AND2X1   g13361(.A(new_n15797_), .B(new_n11886_), .Y(new_n15798_));
  AOI21X1  g13362(.A0(new_n15742_), .A1(new_n12637_), .B0(new_n12638_), .Y(new_n15799_));
  OAI21X1  g13363(.A0(new_n15797_), .A1(new_n12637_), .B0(new_n15799_), .Y(new_n15800_));
  AOI21X1  g13364(.A0(new_n15742_), .A1(pi0619), .B0(pi1159), .Y(new_n15801_));
  OAI21X1  g13365(.A0(new_n15797_), .A1(pi0619), .B0(new_n15801_), .Y(new_n15802_));
  AOI21X1  g13366(.A0(new_n15802_), .A1(new_n15800_), .B0(new_n11886_), .Y(new_n15803_));
  NOR2X1   g13367(.A(new_n15803_), .B(new_n15798_), .Y(new_n15804_));
  INVX1    g13368(.A(new_n15804_), .Y(new_n15805_));
  AOI21X1  g13369(.A0(new_n15742_), .A1(new_n12664_), .B0(new_n12676_), .Y(new_n15806_));
  OAI21X1  g13370(.A0(new_n15805_), .A1(new_n12664_), .B0(new_n15806_), .Y(new_n15807_));
  AOI21X1  g13371(.A0(new_n15742_), .A1(pi0626), .B0(pi1158), .Y(new_n15808_));
  OAI21X1  g13372(.A0(new_n15805_), .A1(pi0626), .B0(new_n15808_), .Y(new_n15809_));
  AND2X1   g13373(.A(new_n15809_), .B(new_n15807_), .Y(new_n15810_));
  MX2X1    g13374(.A(new_n15810_), .B(new_n15804_), .S0(new_n11885_), .Y(new_n15811_));
  AND2X1   g13375(.A(new_n15742_), .B(new_n12711_), .Y(new_n15812_));
  AOI21X1  g13376(.A0(new_n15811_), .A1(new_n14123_), .B0(new_n15812_), .Y(new_n15813_));
  MX2X1    g13377(.A(new_n15813_), .B(new_n15743_), .S0(new_n12735_), .Y(new_n15814_));
  AOI21X1  g13378(.A0(new_n15742_), .A1(new_n12743_), .B0(pi0715), .Y(new_n15815_));
  OAI21X1  g13379(.A0(new_n15814_), .A1(new_n12743_), .B0(new_n15815_), .Y(new_n15816_));
  NAND3X1  g13380(.A(new_n15816_), .B(new_n15773_), .C(pi1160), .Y(new_n15817_));
  OAI22X1  g13381(.A0(new_n15769_), .A1(new_n14387_), .B0(new_n15768_), .B1(new_n14389_), .Y(new_n15818_));
  AOI21X1  g13382(.A0(new_n15813_), .A1(new_n14385_), .B0(new_n15818_), .Y(new_n15819_));
  MX2X1    g13383(.A(new_n15765_), .B(new_n15763_), .S0(new_n12689_), .Y(new_n15820_));
  OAI21X1  g13384(.A0(new_n15811_), .A1(new_n14395_), .B0(new_n15820_), .Y(new_n15821_));
  AOI21X1  g13385(.A0(new_n13989_), .A1(pi0173), .B0(new_n14858_), .Y(new_n15822_));
  OAI21X1  g13386(.A0(new_n13986_), .A1(pi0173), .B0(new_n15822_), .Y(new_n15823_));
  OAI21X1  g13387(.A0(new_n12440_), .A1(pi0173), .B0(new_n14858_), .Y(new_n15824_));
  AOI21X1  g13388(.A0(new_n12401_), .A1(pi0173), .B0(new_n15824_), .Y(new_n15825_));
  NOR2X1   g13389(.A(new_n15825_), .B(new_n2959_), .Y(new_n15826_));
  NAND2X1  g13390(.A(new_n12467_), .B(pi0173), .Y(new_n15827_));
  AOI21X1  g13391(.A0(new_n13996_), .A1(new_n9989_), .B0(new_n14858_), .Y(new_n15828_));
  NAND3X1  g13392(.A(new_n12453_), .B(new_n12104_), .C(new_n9989_), .Y(new_n15829_));
  AOI21X1  g13393(.A0(new_n12474_), .A1(pi0173), .B0(pi0745), .Y(new_n15830_));
  AOI22X1  g13394(.A0(new_n15830_), .A1(new_n15829_), .B0(new_n15828_), .B1(new_n15827_), .Y(new_n15831_));
  OAI21X1  g13395(.A0(new_n15831_), .A1(pi0039), .B0(new_n2996_), .Y(new_n15832_));
  AOI21X1  g13396(.A0(new_n15826_), .A1(new_n15823_), .B0(new_n15832_), .Y(new_n15833_));
  OAI21X1  g13397(.A0(new_n12478_), .A1(pi0745), .B0(new_n13669_), .Y(new_n15834_));
  AND2X1   g13398(.A(new_n12178_), .B(new_n14858_), .Y(new_n15835_));
  OAI21X1  g13399(.A0(new_n15835_), .A1(new_n13576_), .B0(pi0173), .Y(new_n15836_));
  OAI21X1  g13400(.A0(new_n15836_), .A1(new_n14411_), .B0(pi0038), .Y(new_n15837_));
  AOI21X1  g13401(.A0(new_n15834_), .A1(new_n9989_), .B0(new_n15837_), .Y(new_n15838_));
  OR2X1    g13402(.A(new_n15838_), .B(pi0723), .Y(new_n15839_));
  OAI21X1  g13403(.A0(new_n15839_), .A1(new_n15833_), .B0(new_n3129_), .Y(new_n15840_));
  AOI21X1  g13404(.A0(new_n15781_), .A1(pi0723), .B0(new_n15840_), .Y(new_n15841_));
  AOI21X1  g13405(.A0(new_n3810_), .A1(pi0173), .B0(new_n15841_), .Y(new_n15842_));
  OAI21X1  g13406(.A0(new_n15783_), .A1(new_n12493_), .B0(new_n12494_), .Y(new_n15843_));
  AOI21X1  g13407(.A0(new_n15842_), .A1(new_n12493_), .B0(new_n15843_), .Y(new_n15844_));
  NAND2X1  g13408(.A(new_n15751_), .B(new_n12584_), .Y(new_n15845_));
  OAI21X1  g13409(.A0(new_n15783_), .A1(pi0625), .B0(pi1153), .Y(new_n15846_));
  AOI21X1  g13410(.A0(new_n15842_), .A1(pi0625), .B0(new_n15846_), .Y(new_n15847_));
  NAND2X1  g13411(.A(new_n15753_), .B(pi0608), .Y(new_n15848_));
  OAI22X1  g13412(.A0(new_n15848_), .A1(new_n15847_), .B0(new_n15845_), .B1(new_n15844_), .Y(new_n15849_));
  AND2X1   g13413(.A(new_n15842_), .B(new_n11889_), .Y(new_n15850_));
  AOI21X1  g13414(.A0(new_n15849_), .A1(pi0778), .B0(new_n15850_), .Y(new_n15851_));
  AOI21X1  g13415(.A0(new_n15755_), .A1(pi0609), .B0(pi1155), .Y(new_n15852_));
  OAI21X1  g13416(.A0(new_n15851_), .A1(pi0609), .B0(new_n15852_), .Y(new_n15853_));
  AND2X1   g13417(.A(new_n15787_), .B(new_n12596_), .Y(new_n15854_));
  AOI21X1  g13418(.A0(new_n15755_), .A1(new_n12590_), .B0(new_n12591_), .Y(new_n15855_));
  OAI21X1  g13419(.A0(new_n15851_), .A1(new_n12590_), .B0(new_n15855_), .Y(new_n15856_));
  AND2X1   g13420(.A(new_n15789_), .B(pi0660), .Y(new_n15857_));
  AOI22X1  g13421(.A0(new_n15857_), .A1(new_n15856_), .B0(new_n15854_), .B1(new_n15853_), .Y(new_n15858_));
  MX2X1    g13422(.A(new_n15858_), .B(new_n15851_), .S0(new_n11888_), .Y(new_n15859_));
  AOI21X1  g13423(.A0(new_n15756_), .A1(pi0618), .B0(pi1154), .Y(new_n15860_));
  OAI21X1  g13424(.A0(new_n15859_), .A1(pi0618), .B0(new_n15860_), .Y(new_n15861_));
  AND2X1   g13425(.A(new_n15793_), .B(new_n12622_), .Y(new_n15862_));
  AOI21X1  g13426(.A0(new_n15756_), .A1(new_n12614_), .B0(new_n12615_), .Y(new_n15863_));
  OAI21X1  g13427(.A0(new_n15859_), .A1(new_n12614_), .B0(new_n15863_), .Y(new_n15864_));
  AND2X1   g13428(.A(new_n15795_), .B(pi0627), .Y(new_n15865_));
  AOI22X1  g13429(.A0(new_n15865_), .A1(new_n15864_), .B0(new_n15862_), .B1(new_n15861_), .Y(new_n15866_));
  OR2X1    g13430(.A(new_n15859_), .B(pi0781), .Y(new_n15867_));
  OAI21X1  g13431(.A0(new_n15866_), .A1(new_n11887_), .B0(new_n15867_), .Y(new_n15868_));
  NAND2X1  g13432(.A(new_n15868_), .B(new_n12637_), .Y(new_n15869_));
  AOI21X1  g13433(.A0(new_n15757_), .A1(pi0619), .B0(pi1159), .Y(new_n15870_));
  NAND2X1  g13434(.A(new_n15800_), .B(new_n12645_), .Y(new_n15871_));
  AOI21X1  g13435(.A0(new_n15870_), .A1(new_n15869_), .B0(new_n15871_), .Y(new_n15872_));
  NAND2X1  g13436(.A(new_n15868_), .B(pi0619), .Y(new_n15873_));
  AOI21X1  g13437(.A0(new_n15757_), .A1(new_n12637_), .B0(new_n12638_), .Y(new_n15874_));
  NAND2X1  g13438(.A(new_n15802_), .B(pi0648), .Y(new_n15875_));
  AOI21X1  g13439(.A0(new_n15874_), .A1(new_n15873_), .B0(new_n15875_), .Y(new_n15876_));
  NOR3X1   g13440(.A(new_n15876_), .B(new_n15872_), .C(new_n11886_), .Y(new_n15877_));
  OAI21X1  g13441(.A0(new_n15868_), .A1(pi0789), .B0(new_n12842_), .Y(new_n15878_));
  OR2X1    g13442(.A(new_n15878_), .B(new_n15877_), .Y(new_n15879_));
  NAND3X1  g13443(.A(new_n15809_), .B(new_n15807_), .C(new_n13537_), .Y(new_n15880_));
  OAI21X1  g13444(.A0(new_n15759_), .A1(new_n12770_), .B0(new_n15880_), .Y(new_n15881_));
  AOI21X1  g13445(.A0(new_n15881_), .A1(pi0788), .B0(new_n14273_), .Y(new_n15882_));
  AOI22X1  g13446(.A0(new_n15882_), .A1(new_n15879_), .B0(new_n15821_), .B1(pi0792), .Y(new_n15883_));
  OAI22X1  g13447(.A0(new_n15883_), .A1(new_n14269_), .B0(new_n15819_), .B1(new_n11883_), .Y(new_n15884_));
  NOR2X1   g13448(.A(new_n15884_), .B(pi0644), .Y(new_n15885_));
  OAI21X1  g13449(.A0(new_n15772_), .A1(new_n12743_), .B0(new_n12739_), .Y(new_n15886_));
  AOI21X1  g13450(.A0(new_n15742_), .A1(pi0644), .B0(new_n12739_), .Y(new_n15887_));
  OAI21X1  g13451(.A0(new_n15814_), .A1(pi0644), .B0(new_n15887_), .Y(new_n15888_));
  AND2X1   g13452(.A(new_n15888_), .B(new_n11882_), .Y(new_n15889_));
  OAI21X1  g13453(.A0(new_n15886_), .A1(new_n15885_), .B0(new_n15889_), .Y(new_n15890_));
  AOI21X1  g13454(.A0(new_n15890_), .A1(new_n15817_), .B0(new_n12897_), .Y(new_n15891_));
  NAND3X1  g13455(.A(new_n15816_), .B(pi1160), .C(pi0644), .Y(new_n15892_));
  AOI21X1  g13456(.A0(new_n15892_), .A1(pi0790), .B0(new_n15884_), .Y(new_n15893_));
  OAI21X1  g13457(.A0(new_n15893_), .A1(new_n15891_), .B0(new_n6520_), .Y(new_n15894_));
  AOI21X1  g13458(.A0(po1038), .A1(new_n9989_), .B0(pi0832), .Y(new_n15895_));
  AOI21X1  g13459(.A0(pi1093), .A1(pi1092), .B0(pi0173), .Y(new_n15896_));
  AOI21X1  g13460(.A0(new_n12178_), .A1(new_n14858_), .B0(new_n15896_), .Y(new_n15897_));
  AOI21X1  g13461(.A0(new_n12601_), .A1(new_n2739_), .B0(new_n15897_), .Y(new_n15898_));
  AND2X1   g13462(.A(new_n15835_), .B(new_n12608_), .Y(new_n15899_));
  INVX1    g13463(.A(new_n15899_), .Y(new_n15900_));
  AOI21X1  g13464(.A0(new_n15900_), .A1(new_n15898_), .B0(new_n12591_), .Y(new_n15901_));
  NOR3X1   g13465(.A(new_n15899_), .B(new_n15896_), .C(pi1155), .Y(new_n15902_));
  NOR2X1   g13466(.A(new_n15902_), .B(new_n15901_), .Y(new_n15903_));
  MX2X1    g13467(.A(new_n15903_), .B(new_n15898_), .S0(new_n11888_), .Y(new_n15904_));
  AOI21X1  g13468(.A0(new_n15904_), .A1(new_n12785_), .B0(new_n12615_), .Y(new_n15905_));
  AOI21X1  g13469(.A0(new_n15904_), .A1(new_n12788_), .B0(pi1154), .Y(new_n15906_));
  NOR2X1   g13470(.A(new_n15906_), .B(new_n15905_), .Y(new_n15907_));
  MX2X1    g13471(.A(new_n15907_), .B(new_n15904_), .S0(new_n11887_), .Y(new_n15908_));
  OR2X1    g13472(.A(new_n15908_), .B(pi0789), .Y(new_n15909_));
  NAND2X1  g13473(.A(new_n2739_), .B(new_n12637_), .Y(new_n15910_));
  AOI21X1  g13474(.A0(new_n15910_), .A1(new_n15908_), .B0(new_n12638_), .Y(new_n15911_));
  NAND3X1  g13475(.A(pi1093), .B(pi1092), .C(pi0619), .Y(new_n15912_));
  AOI21X1  g13476(.A0(new_n15912_), .A1(new_n15908_), .B0(pi1159), .Y(new_n15913_));
  OAI21X1  g13477(.A0(new_n15913_), .A1(new_n15911_), .B0(pi0789), .Y(new_n15914_));
  AND2X1   g13478(.A(new_n15914_), .B(new_n15909_), .Y(new_n15915_));
  NAND3X1  g13479(.A(new_n15914_), .B(new_n15909_), .C(pi0626), .Y(new_n15916_));
  AOI21X1  g13480(.A0(new_n15896_), .A1(new_n12664_), .B0(new_n12676_), .Y(new_n15917_));
  NAND3X1  g13481(.A(new_n15914_), .B(new_n15909_), .C(new_n12664_), .Y(new_n15918_));
  AOI21X1  g13482(.A0(new_n15896_), .A1(pi0626), .B0(pi1158), .Y(new_n15919_));
  AOI22X1  g13483(.A0(new_n15919_), .A1(new_n15918_), .B0(new_n15917_), .B1(new_n15916_), .Y(new_n15920_));
  MX2X1    g13484(.A(new_n15920_), .B(new_n15915_), .S0(new_n11885_), .Y(new_n15921_));
  AND2X1   g13485(.A(new_n15896_), .B(new_n12711_), .Y(new_n15922_));
  AOI21X1  g13486(.A0(new_n15921_), .A1(new_n14123_), .B0(new_n15922_), .Y(new_n15923_));
  AOI21X1  g13487(.A0(new_n12566_), .A1(new_n14886_), .B0(new_n15896_), .Y(new_n15924_));
  INVX1    g13488(.A(new_n15924_), .Y(new_n15925_));
  NOR3X1   g13489(.A(new_n13585_), .B(pi0723), .C(pi0625), .Y(new_n15926_));
  INVX1    g13490(.A(new_n15926_), .Y(new_n15927_));
  AOI21X1  g13491(.A0(new_n15927_), .A1(new_n15925_), .B0(new_n12494_), .Y(new_n15928_));
  INVX1    g13492(.A(new_n15928_), .Y(new_n15929_));
  NOR2X1   g13493(.A(new_n15896_), .B(pi1153), .Y(new_n15930_));
  AOI21X1  g13494(.A0(new_n15930_), .A1(new_n15927_), .B0(new_n11889_), .Y(new_n15931_));
  AOI22X1  g13495(.A0(new_n15931_), .A1(new_n15929_), .B0(new_n15925_), .B1(new_n11889_), .Y(new_n15932_));
  NOR3X1   g13496(.A(new_n15932_), .B(new_n12764_), .C(new_n12762_), .Y(new_n15933_));
  INVX1    g13497(.A(new_n15933_), .Y(new_n15934_));
  NOR4X1   g13498(.A(new_n15934_), .B(new_n12870_), .C(new_n12851_), .D(new_n12765_), .Y(new_n15935_));
  INVX1    g13499(.A(new_n15935_), .Y(new_n15936_));
  AOI21X1  g13500(.A0(new_n15896_), .A1(pi0647), .B0(pi1157), .Y(new_n15937_));
  OAI21X1  g13501(.A0(new_n15936_), .A1(pi0647), .B0(new_n15937_), .Y(new_n15938_));
  MX2X1    g13502(.A(new_n15935_), .B(new_n15896_), .S0(new_n12705_), .Y(new_n15939_));
  OAI22X1  g13503(.A0(new_n15939_), .A1(new_n14387_), .B0(new_n15938_), .B1(new_n12723_), .Y(new_n15940_));
  AOI21X1  g13504(.A0(new_n15923_), .A1(new_n14385_), .B0(new_n15940_), .Y(new_n15941_));
  NOR3X1   g13505(.A(new_n15934_), .B(new_n12770_), .C(new_n12765_), .Y(new_n15942_));
  AND2X1   g13506(.A(new_n15920_), .B(new_n13537_), .Y(new_n15943_));
  OR2X1    g13507(.A(new_n15943_), .B(new_n15942_), .Y(new_n15944_));
  INVX1    g13508(.A(new_n15897_), .Y(new_n15945_));
  AOI21X1  g13509(.A0(new_n15925_), .A1(new_n12171_), .B0(new_n15945_), .Y(new_n15946_));
  NOR3X1   g13510(.A(new_n15924_), .B(new_n12120_), .C(new_n12493_), .Y(new_n15947_));
  OR2X1    g13511(.A(new_n15946_), .B(new_n15947_), .Y(new_n15948_));
  OR2X1    g13512(.A(new_n15928_), .B(pi0608), .Y(new_n15949_));
  AOI21X1  g13513(.A0(new_n15948_), .A1(new_n15930_), .B0(new_n15949_), .Y(new_n15950_));
  NOR3X1   g13514(.A(new_n15947_), .B(new_n15945_), .C(new_n12494_), .Y(new_n15951_));
  INVX1    g13515(.A(new_n15930_), .Y(new_n15952_));
  OAI21X1  g13516(.A0(new_n15952_), .A1(new_n15926_), .B0(pi0608), .Y(new_n15953_));
  NOR2X1   g13517(.A(new_n15953_), .B(new_n15951_), .Y(new_n15954_));
  OAI21X1  g13518(.A0(new_n15954_), .A1(new_n15950_), .B0(pi0778), .Y(new_n15955_));
  OAI21X1  g13519(.A0(new_n15946_), .A1(pi0778), .B0(new_n15955_), .Y(new_n15956_));
  OAI21X1  g13520(.A0(new_n15932_), .A1(new_n12590_), .B0(new_n12591_), .Y(new_n15957_));
  AOI21X1  g13521(.A0(new_n15956_), .A1(new_n12590_), .B0(new_n15957_), .Y(new_n15958_));
  OR2X1    g13522(.A(new_n15901_), .B(pi0660), .Y(new_n15959_));
  OAI21X1  g13523(.A0(new_n15932_), .A1(pi0609), .B0(pi1155), .Y(new_n15960_));
  AOI21X1  g13524(.A0(new_n15956_), .A1(pi0609), .B0(new_n15960_), .Y(new_n15961_));
  OR2X1    g13525(.A(new_n15902_), .B(new_n12596_), .Y(new_n15962_));
  OAI22X1  g13526(.A0(new_n15962_), .A1(new_n15961_), .B0(new_n15959_), .B1(new_n15958_), .Y(new_n15963_));
  MX2X1    g13527(.A(new_n15963_), .B(new_n15956_), .S0(new_n11888_), .Y(new_n15964_));
  INVX1    g13528(.A(new_n15964_), .Y(new_n15965_));
  NOR3X1   g13529(.A(new_n15932_), .B(new_n12762_), .C(new_n12614_), .Y(new_n15966_));
  NOR2X1   g13530(.A(new_n15966_), .B(pi1154), .Y(new_n15967_));
  OAI21X1  g13531(.A0(new_n15965_), .A1(pi0618), .B0(new_n15967_), .Y(new_n15968_));
  NOR2X1   g13532(.A(new_n15905_), .B(pi0627), .Y(new_n15969_));
  NOR3X1   g13533(.A(new_n15932_), .B(new_n12762_), .C(pi0618), .Y(new_n15970_));
  NOR2X1   g13534(.A(new_n15970_), .B(new_n12615_), .Y(new_n15971_));
  OAI21X1  g13535(.A0(new_n15965_), .A1(new_n12614_), .B0(new_n15971_), .Y(new_n15972_));
  NOR2X1   g13536(.A(new_n15906_), .B(new_n12622_), .Y(new_n15973_));
  AOI22X1  g13537(.A0(new_n15973_), .A1(new_n15972_), .B0(new_n15969_), .B1(new_n15968_), .Y(new_n15974_));
  MX2X1    g13538(.A(new_n15974_), .B(new_n15965_), .S0(new_n11887_), .Y(new_n15975_));
  AOI21X1  g13539(.A0(new_n15933_), .A1(pi0619), .B0(pi1159), .Y(new_n15976_));
  OAI21X1  g13540(.A0(new_n15975_), .A1(pi0619), .B0(new_n15976_), .Y(new_n15977_));
  NOR2X1   g13541(.A(new_n15911_), .B(pi0648), .Y(new_n15978_));
  AND2X1   g13542(.A(new_n15978_), .B(new_n15977_), .Y(new_n15979_));
  AOI21X1  g13543(.A0(new_n15933_), .A1(new_n12637_), .B0(new_n12638_), .Y(new_n15980_));
  OAI21X1  g13544(.A0(new_n15975_), .A1(new_n12637_), .B0(new_n15980_), .Y(new_n15981_));
  NOR2X1   g13545(.A(new_n15913_), .B(new_n12645_), .Y(new_n15982_));
  AOI21X1  g13546(.A0(new_n15982_), .A1(new_n15981_), .B0(new_n11886_), .Y(new_n15983_));
  INVX1    g13547(.A(new_n15983_), .Y(new_n15984_));
  OR2X1    g13548(.A(new_n15984_), .B(new_n15979_), .Y(new_n15985_));
  AOI21X1  g13549(.A0(new_n15975_), .A1(new_n11886_), .B0(new_n14264_), .Y(new_n15986_));
  AOI22X1  g13550(.A0(new_n15986_), .A1(new_n15985_), .B0(new_n15944_), .B1(pi0788), .Y(new_n15987_));
  NOR2X1   g13551(.A(new_n15987_), .B(new_n14273_), .Y(new_n15988_));
  NOR3X1   g13552(.A(new_n15934_), .B(new_n12851_), .C(new_n12765_), .Y(new_n15989_));
  AOI22X1  g13553(.A0(new_n15989_), .A1(new_n14564_), .B0(new_n15921_), .B1(new_n12867_), .Y(new_n15990_));
  AOI22X1  g13554(.A0(new_n15989_), .A1(new_n14566_), .B0(new_n15921_), .B1(new_n12865_), .Y(new_n15991_));
  MX2X1    g13555(.A(new_n15991_), .B(new_n15990_), .S0(new_n12689_), .Y(new_n15992_));
  OAI21X1  g13556(.A0(new_n15992_), .A1(new_n11884_), .B0(new_n14562_), .Y(new_n15993_));
  OAI22X1  g13557(.A0(new_n15993_), .A1(new_n15988_), .B0(new_n15941_), .B1(new_n11883_), .Y(new_n15994_));
  INVX1    g13558(.A(new_n15994_), .Y(new_n15995_));
  OAI21X1  g13559(.A0(new_n15939_), .A1(new_n12706_), .B0(new_n15938_), .Y(new_n15996_));
  MX2X1    g13560(.A(new_n15996_), .B(new_n15936_), .S0(new_n11883_), .Y(new_n15997_));
  OAI21X1  g13561(.A0(new_n15997_), .A1(pi0644), .B0(pi0715), .Y(new_n15998_));
  AOI21X1  g13562(.A0(new_n15995_), .A1(pi0644), .B0(new_n15998_), .Y(new_n15999_));
  OR4X1    g13563(.A(new_n12734_), .B(new_n2739_), .C(new_n11883_), .D(pi0173), .Y(new_n16000_));
  OAI21X1  g13564(.A0(new_n15923_), .A1(new_n12735_), .B0(new_n16000_), .Y(new_n16001_));
  INVX1    g13565(.A(new_n15896_), .Y(new_n16002_));
  OAI21X1  g13566(.A0(new_n16002_), .A1(pi0644), .B0(new_n12739_), .Y(new_n16003_));
  AOI21X1  g13567(.A0(new_n16001_), .A1(pi0644), .B0(new_n16003_), .Y(new_n16004_));
  OR2X1    g13568(.A(new_n16004_), .B(new_n11882_), .Y(new_n16005_));
  OAI21X1  g13569(.A0(new_n15997_), .A1(new_n12743_), .B0(new_n12739_), .Y(new_n16006_));
  AOI21X1  g13570(.A0(new_n15995_), .A1(new_n12743_), .B0(new_n16006_), .Y(new_n16007_));
  OAI21X1  g13571(.A0(new_n16002_), .A1(new_n12743_), .B0(pi0715), .Y(new_n16008_));
  AOI21X1  g13572(.A0(new_n16001_), .A1(new_n12743_), .B0(new_n16008_), .Y(new_n16009_));
  OR2X1    g13573(.A(new_n16009_), .B(pi1160), .Y(new_n16010_));
  OAI22X1  g13574(.A0(new_n16010_), .A1(new_n16007_), .B0(new_n16005_), .B1(new_n15999_), .Y(new_n16011_));
  OAI21X1  g13575(.A0(new_n15994_), .A1(pi0790), .B0(pi0832), .Y(new_n16012_));
  AOI21X1  g13576(.A0(new_n16011_), .A1(pi0790), .B0(new_n16012_), .Y(new_n16013_));
  AOI21X1  g13577(.A0(new_n15895_), .A1(new_n15894_), .B0(new_n16013_), .Y(po0330));
  AND2X1   g13578(.A(new_n12161_), .B(pi0759), .Y(new_n16015_));
  OAI21X1  g13579(.A0(new_n16015_), .A1(new_n14961_), .B0(pi0039), .Y(new_n16016_));
  AOI21X1  g13580(.A0(new_n11947_), .A1(new_n14908_), .B0(pi0039), .Y(new_n16017_));
  OAI21X1  g13581(.A0(new_n12909_), .A1(new_n14908_), .B0(new_n16017_), .Y(new_n16018_));
  AOI21X1  g13582(.A0(new_n16018_), .A1(new_n16016_), .B0(new_n7008_), .Y(new_n16019_));
  NOR3X1   g13583(.A(new_n13977_), .B(new_n14908_), .C(pi0174), .Y(new_n16020_));
  OAI21X1  g13584(.A0(new_n16020_), .A1(new_n16019_), .B0(new_n2996_), .Y(new_n16021_));
  NOR2X1   g13585(.A(new_n12202_), .B(pi0174), .Y(new_n16022_));
  AOI21X1  g13586(.A0(new_n12120_), .A1(pi0759), .B0(new_n12901_), .Y(new_n16023_));
  NOR3X1   g13587(.A(new_n16023_), .B(new_n16022_), .C(new_n2996_), .Y(new_n16024_));
  INVX1    g13588(.A(new_n16024_), .Y(new_n16025_));
  NAND3X1  g13589(.A(new_n16025_), .B(new_n16021_), .C(new_n14944_), .Y(new_n16026_));
  OAI21X1  g13590(.A0(new_n13989_), .A1(pi0174), .B0(new_n14908_), .Y(new_n16027_));
  AOI21X1  g13591(.A0(new_n13986_), .A1(pi0174), .B0(new_n16027_), .Y(new_n16028_));
  AOI21X1  g13592(.A0(new_n12440_), .A1(pi0174), .B0(new_n14908_), .Y(new_n16029_));
  OAI21X1  g13593(.A0(new_n12401_), .A1(pi0174), .B0(new_n16029_), .Y(new_n16030_));
  NAND2X1  g13594(.A(new_n16030_), .B(pi0039), .Y(new_n16031_));
  AOI21X1  g13595(.A0(new_n13996_), .A1(pi0174), .B0(pi0759), .Y(new_n16032_));
  OAI21X1  g13596(.A0(new_n13995_), .A1(pi0174), .B0(new_n16032_), .Y(new_n16033_));
  NAND3X1  g13597(.A(new_n12453_), .B(new_n12104_), .C(pi0174), .Y(new_n16034_));
  AOI21X1  g13598(.A0(new_n12474_), .A1(new_n7008_), .B0(new_n14908_), .Y(new_n16035_));
  AOI21X1  g13599(.A0(new_n16035_), .A1(new_n16034_), .B0(pi0039), .Y(new_n16036_));
  AOI21X1  g13600(.A0(new_n16036_), .A1(new_n16033_), .B0(pi0038), .Y(new_n16037_));
  OAI21X1  g13601(.A0(new_n16031_), .A1(new_n16028_), .B0(new_n16037_), .Y(new_n16038_));
  NOR3X1   g13602(.A(new_n16024_), .B(new_n13676_), .C(new_n14944_), .Y(new_n16039_));
  AOI21X1  g13603(.A0(new_n16039_), .A1(new_n16038_), .B0(new_n3810_), .Y(new_n16040_));
  AOI22X1  g13604(.A0(new_n16040_), .A1(new_n16026_), .B0(new_n3810_), .B1(pi0174), .Y(new_n16041_));
  AND2X1   g13605(.A(new_n16041_), .B(new_n12493_), .Y(new_n16042_));
  NAND2X1  g13606(.A(new_n16025_), .B(new_n16021_), .Y(new_n16043_));
  MX2X1    g13607(.A(new_n16043_), .B(pi0174), .S0(new_n3810_), .Y(new_n16044_));
  OAI21X1  g13608(.A0(new_n16044_), .A1(new_n12493_), .B0(new_n12494_), .Y(new_n16045_));
  OAI21X1  g13609(.A0(new_n12574_), .A1(new_n3810_), .B0(pi0174), .Y(new_n16046_));
  NOR4X1   g13610(.A(new_n3125_), .B(new_n14944_), .C(pi0100), .D(pi0087), .Y(new_n16047_));
  INVX1    g13611(.A(new_n16047_), .Y(new_n16048_));
  OAI21X1  g13612(.A0(new_n12955_), .A1(pi0174), .B0(new_n2996_), .Y(new_n16049_));
  AOI21X1  g13613(.A0(new_n12953_), .A1(pi0174), .B0(new_n16049_), .Y(new_n16050_));
  OAI21X1  g13614(.A0(new_n16022_), .A1(new_n14017_), .B0(new_n16047_), .Y(new_n16051_));
  NOR2X1   g13615(.A(new_n16051_), .B(new_n16050_), .Y(new_n16052_));
  AOI21X1  g13616(.A0(new_n16048_), .A1(new_n16046_), .B0(new_n16052_), .Y(new_n16053_));
  AOI21X1  g13617(.A0(new_n16046_), .A1(new_n12493_), .B0(new_n12494_), .Y(new_n16054_));
  OAI21X1  g13618(.A0(new_n16053_), .A1(new_n12493_), .B0(new_n16054_), .Y(new_n16055_));
  AND2X1   g13619(.A(new_n16055_), .B(new_n12584_), .Y(new_n16056_));
  OAI21X1  g13620(.A0(new_n16045_), .A1(new_n16042_), .B0(new_n16056_), .Y(new_n16057_));
  AND2X1   g13621(.A(new_n16041_), .B(pi0625), .Y(new_n16058_));
  OAI21X1  g13622(.A0(new_n16044_), .A1(pi0625), .B0(pi1153), .Y(new_n16059_));
  AOI21X1  g13623(.A0(new_n16046_), .A1(pi0625), .B0(pi1153), .Y(new_n16060_));
  OAI21X1  g13624(.A0(new_n16053_), .A1(pi0625), .B0(new_n16060_), .Y(new_n16061_));
  AND2X1   g13625(.A(new_n16061_), .B(pi0608), .Y(new_n16062_));
  OAI21X1  g13626(.A0(new_n16059_), .A1(new_n16058_), .B0(new_n16062_), .Y(new_n16063_));
  AOI21X1  g13627(.A0(new_n16063_), .A1(new_n16057_), .B0(new_n11889_), .Y(new_n16064_));
  AND2X1   g13628(.A(new_n16041_), .B(new_n11889_), .Y(new_n16065_));
  OAI21X1  g13629(.A0(new_n16065_), .A1(new_n16064_), .B0(new_n12590_), .Y(new_n16066_));
  AND2X1   g13630(.A(new_n16053_), .B(new_n11889_), .Y(new_n16067_));
  NAND2X1  g13631(.A(new_n16061_), .B(new_n16055_), .Y(new_n16068_));
  AOI21X1  g13632(.A0(new_n16068_), .A1(pi0778), .B0(new_n16067_), .Y(new_n16069_));
  AOI21X1  g13633(.A0(new_n16069_), .A1(pi0609), .B0(pi1155), .Y(new_n16070_));
  NAND2X1  g13634(.A(new_n16046_), .B(new_n12601_), .Y(new_n16071_));
  OAI21X1  g13635(.A0(new_n16044_), .A1(new_n12601_), .B0(new_n16071_), .Y(new_n16072_));
  INVX1    g13636(.A(new_n16046_), .Y(new_n16073_));
  OAI21X1  g13637(.A0(new_n16073_), .A1(pi0609), .B0(pi1155), .Y(new_n16074_));
  AOI21X1  g13638(.A0(new_n16072_), .A1(pi0609), .B0(new_n16074_), .Y(new_n16075_));
  OR2X1    g13639(.A(new_n16075_), .B(pi0660), .Y(new_n16076_));
  AOI21X1  g13640(.A0(new_n16070_), .A1(new_n16066_), .B0(new_n16076_), .Y(new_n16077_));
  OAI21X1  g13641(.A0(new_n16065_), .A1(new_n16064_), .B0(pi0609), .Y(new_n16078_));
  AOI21X1  g13642(.A0(new_n16069_), .A1(new_n12590_), .B0(new_n12591_), .Y(new_n16079_));
  OAI21X1  g13643(.A0(new_n16073_), .A1(new_n12590_), .B0(new_n12591_), .Y(new_n16080_));
  AOI21X1  g13644(.A0(new_n16072_), .A1(new_n12590_), .B0(new_n16080_), .Y(new_n16081_));
  OR2X1    g13645(.A(new_n16081_), .B(new_n12596_), .Y(new_n16082_));
  AOI21X1  g13646(.A0(new_n16079_), .A1(new_n16078_), .B0(new_n16082_), .Y(new_n16083_));
  OAI21X1  g13647(.A0(new_n16083_), .A1(new_n16077_), .B0(pi0785), .Y(new_n16084_));
  OAI21X1  g13648(.A0(new_n16065_), .A1(new_n16064_), .B0(new_n11888_), .Y(new_n16085_));
  AOI21X1  g13649(.A0(new_n16085_), .A1(new_n16084_), .B0(pi0618), .Y(new_n16086_));
  AND2X1   g13650(.A(new_n16046_), .B(new_n12618_), .Y(new_n16087_));
  AOI21X1  g13651(.A0(new_n16069_), .A1(new_n13598_), .B0(new_n16087_), .Y(new_n16088_));
  OAI21X1  g13652(.A0(new_n16088_), .A1(new_n12614_), .B0(new_n12615_), .Y(new_n16089_));
  OAI21X1  g13653(.A0(new_n16081_), .A1(new_n16075_), .B0(pi0785), .Y(new_n16090_));
  OAI21X1  g13654(.A0(new_n16072_), .A1(pi0785), .B0(new_n16090_), .Y(new_n16091_));
  AOI21X1  g13655(.A0(new_n16046_), .A1(new_n12614_), .B0(new_n12615_), .Y(new_n16092_));
  OAI21X1  g13656(.A0(new_n16091_), .A1(new_n12614_), .B0(new_n16092_), .Y(new_n16093_));
  AND2X1   g13657(.A(new_n16093_), .B(new_n12622_), .Y(new_n16094_));
  OAI21X1  g13658(.A0(new_n16089_), .A1(new_n16086_), .B0(new_n16094_), .Y(new_n16095_));
  AOI21X1  g13659(.A0(new_n16085_), .A1(new_n16084_), .B0(new_n12614_), .Y(new_n16096_));
  OAI21X1  g13660(.A0(new_n16088_), .A1(pi0618), .B0(pi1154), .Y(new_n16097_));
  AOI21X1  g13661(.A0(new_n16046_), .A1(pi0618), .B0(pi1154), .Y(new_n16098_));
  OAI21X1  g13662(.A0(new_n16091_), .A1(pi0618), .B0(new_n16098_), .Y(new_n16099_));
  AND2X1   g13663(.A(new_n16099_), .B(pi0627), .Y(new_n16100_));
  OAI21X1  g13664(.A0(new_n16097_), .A1(new_n16096_), .B0(new_n16100_), .Y(new_n16101_));
  AOI21X1  g13665(.A0(new_n16101_), .A1(new_n16095_), .B0(new_n11887_), .Y(new_n16102_));
  AOI21X1  g13666(.A0(new_n16085_), .A1(new_n16084_), .B0(pi0781), .Y(new_n16103_));
  OAI21X1  g13667(.A0(new_n16103_), .A1(new_n16102_), .B0(new_n12637_), .Y(new_n16104_));
  MX2X1    g13668(.A(new_n16088_), .B(new_n16073_), .S0(new_n12641_), .Y(new_n16105_));
  INVX1    g13669(.A(new_n16105_), .Y(new_n16106_));
  AOI21X1  g13670(.A0(new_n16106_), .A1(pi0619), .B0(pi1159), .Y(new_n16107_));
  AOI21X1  g13671(.A0(new_n16099_), .A1(new_n16093_), .B0(new_n11887_), .Y(new_n16108_));
  AOI21X1  g13672(.A0(new_n16091_), .A1(new_n11887_), .B0(new_n16108_), .Y(new_n16109_));
  OAI21X1  g13673(.A0(new_n16073_), .A1(pi0619), .B0(pi1159), .Y(new_n16110_));
  AOI21X1  g13674(.A0(new_n16109_), .A1(pi0619), .B0(new_n16110_), .Y(new_n16111_));
  OR2X1    g13675(.A(new_n16111_), .B(pi0648), .Y(new_n16112_));
  AOI21X1  g13676(.A0(new_n16107_), .A1(new_n16104_), .B0(new_n16112_), .Y(new_n16113_));
  OAI21X1  g13677(.A0(new_n16103_), .A1(new_n16102_), .B0(pi0619), .Y(new_n16114_));
  AOI21X1  g13678(.A0(new_n16106_), .A1(new_n12637_), .B0(new_n12638_), .Y(new_n16115_));
  OAI21X1  g13679(.A0(new_n16073_), .A1(new_n12637_), .B0(new_n12638_), .Y(new_n16116_));
  AOI21X1  g13680(.A0(new_n16109_), .A1(new_n12637_), .B0(new_n16116_), .Y(new_n16117_));
  OR2X1    g13681(.A(new_n16117_), .B(new_n12645_), .Y(new_n16118_));
  AOI21X1  g13682(.A0(new_n16115_), .A1(new_n16114_), .B0(new_n16118_), .Y(new_n16119_));
  OAI21X1  g13683(.A0(new_n16119_), .A1(new_n16113_), .B0(pi0789), .Y(new_n16120_));
  OAI21X1  g13684(.A0(new_n16103_), .A1(new_n16102_), .B0(new_n11886_), .Y(new_n16121_));
  NAND3X1  g13685(.A(new_n16121_), .B(new_n16120_), .C(new_n11885_), .Y(new_n16122_));
  NAND3X1  g13686(.A(new_n16121_), .B(new_n16120_), .C(new_n12664_), .Y(new_n16123_));
  MX2X1    g13687(.A(new_n16105_), .B(new_n16073_), .S0(new_n12659_), .Y(new_n16124_));
  AOI21X1  g13688(.A0(new_n16124_), .A1(pi0626), .B0(pi0641), .Y(new_n16125_));
  NOR2X1   g13689(.A(new_n16117_), .B(new_n16111_), .Y(new_n16126_));
  MX2X1    g13690(.A(new_n16126_), .B(new_n16109_), .S0(new_n11886_), .Y(new_n16127_));
  AOI21X1  g13691(.A0(new_n16073_), .A1(pi0626), .B0(new_n12672_), .Y(new_n16128_));
  OAI21X1  g13692(.A0(new_n16127_), .A1(pi0626), .B0(new_n16128_), .Y(new_n16129_));
  NAND2X1  g13693(.A(new_n16129_), .B(new_n12676_), .Y(new_n16130_));
  AOI21X1  g13694(.A0(new_n16125_), .A1(new_n16123_), .B0(new_n16130_), .Y(new_n16131_));
  NAND3X1  g13695(.A(new_n16121_), .B(new_n16120_), .C(pi0626), .Y(new_n16132_));
  AOI21X1  g13696(.A0(new_n16124_), .A1(new_n12664_), .B0(new_n12672_), .Y(new_n16133_));
  AOI21X1  g13697(.A0(new_n16073_), .A1(new_n12664_), .B0(pi0641), .Y(new_n16134_));
  OAI21X1  g13698(.A0(new_n16127_), .A1(new_n12664_), .B0(new_n16134_), .Y(new_n16135_));
  NAND2X1  g13699(.A(new_n16135_), .B(pi1158), .Y(new_n16136_));
  AOI21X1  g13700(.A0(new_n16133_), .A1(new_n16132_), .B0(new_n16136_), .Y(new_n16137_));
  OAI21X1  g13701(.A0(new_n16137_), .A1(new_n16131_), .B0(pi0788), .Y(new_n16138_));
  NAND3X1  g13702(.A(new_n16138_), .B(new_n16122_), .C(new_n12683_), .Y(new_n16139_));
  MX2X1    g13703(.A(new_n16127_), .B(new_n16046_), .S0(new_n12841_), .Y(new_n16140_));
  AOI21X1  g13704(.A0(new_n16140_), .A1(pi0628), .B0(pi1156), .Y(new_n16141_));
  MX2X1    g13705(.A(new_n16124_), .B(new_n16073_), .S0(new_n12691_), .Y(new_n16142_));
  AOI21X1  g13706(.A0(new_n16046_), .A1(new_n12683_), .B0(new_n12684_), .Y(new_n16143_));
  OAI21X1  g13707(.A0(new_n16142_), .A1(new_n12683_), .B0(new_n16143_), .Y(new_n16144_));
  NAND2X1  g13708(.A(new_n16144_), .B(new_n12689_), .Y(new_n16145_));
  AOI21X1  g13709(.A0(new_n16141_), .A1(new_n16139_), .B0(new_n16145_), .Y(new_n16146_));
  NAND3X1  g13710(.A(new_n16138_), .B(new_n16122_), .C(pi0628), .Y(new_n16147_));
  AOI21X1  g13711(.A0(new_n16140_), .A1(new_n12683_), .B0(new_n12684_), .Y(new_n16148_));
  AOI21X1  g13712(.A0(new_n16046_), .A1(pi0628), .B0(pi1156), .Y(new_n16149_));
  OAI21X1  g13713(.A0(new_n16142_), .A1(pi0628), .B0(new_n16149_), .Y(new_n16150_));
  NAND2X1  g13714(.A(new_n16150_), .B(pi0629), .Y(new_n16151_));
  AOI21X1  g13715(.A0(new_n16148_), .A1(new_n16147_), .B0(new_n16151_), .Y(new_n16152_));
  OAI21X1  g13716(.A0(new_n16152_), .A1(new_n16146_), .B0(pi0792), .Y(new_n16153_));
  NAND3X1  g13717(.A(new_n16138_), .B(new_n16122_), .C(new_n11884_), .Y(new_n16154_));
  AOI21X1  g13718(.A0(new_n16154_), .A1(new_n16153_), .B0(pi0647), .Y(new_n16155_));
  MX2X1    g13719(.A(new_n16140_), .B(new_n16046_), .S0(new_n12711_), .Y(new_n16156_));
  INVX1    g13720(.A(new_n16156_), .Y(new_n16157_));
  OAI21X1  g13721(.A0(new_n16157_), .A1(new_n12705_), .B0(new_n12706_), .Y(new_n16158_));
  AND2X1   g13722(.A(new_n16142_), .B(new_n11884_), .Y(new_n16159_));
  AOI21X1  g13723(.A0(new_n16150_), .A1(new_n16144_), .B0(new_n11884_), .Y(new_n16160_));
  NOR2X1   g13724(.A(new_n16160_), .B(new_n16159_), .Y(new_n16161_));
  INVX1    g13725(.A(new_n16161_), .Y(new_n16162_));
  AOI21X1  g13726(.A0(new_n16046_), .A1(new_n12705_), .B0(new_n12706_), .Y(new_n16163_));
  OAI21X1  g13727(.A0(new_n16162_), .A1(new_n12705_), .B0(new_n16163_), .Y(new_n16164_));
  AND2X1   g13728(.A(new_n16164_), .B(new_n12723_), .Y(new_n16165_));
  OAI21X1  g13729(.A0(new_n16158_), .A1(new_n16155_), .B0(new_n16165_), .Y(new_n16166_));
  AOI21X1  g13730(.A0(new_n16154_), .A1(new_n16153_), .B0(new_n12705_), .Y(new_n16167_));
  OAI21X1  g13731(.A0(new_n16157_), .A1(pi0647), .B0(pi1157), .Y(new_n16168_));
  AOI21X1  g13732(.A0(new_n16046_), .A1(pi0647), .B0(pi1157), .Y(new_n16169_));
  OAI21X1  g13733(.A0(new_n16162_), .A1(pi0647), .B0(new_n16169_), .Y(new_n16170_));
  AND2X1   g13734(.A(new_n16170_), .B(pi0630), .Y(new_n16171_));
  OAI21X1  g13735(.A0(new_n16168_), .A1(new_n16167_), .B0(new_n16171_), .Y(new_n16172_));
  AOI21X1  g13736(.A0(new_n16172_), .A1(new_n16166_), .B0(new_n11883_), .Y(new_n16173_));
  AOI21X1  g13737(.A0(new_n16154_), .A1(new_n16153_), .B0(pi0787), .Y(new_n16174_));
  OAI21X1  g13738(.A0(new_n16174_), .A1(new_n16173_), .B0(pi0644), .Y(new_n16175_));
  AND2X1   g13739(.A(new_n16170_), .B(new_n16164_), .Y(new_n16176_));
  MX2X1    g13740(.A(new_n16176_), .B(new_n16161_), .S0(new_n11883_), .Y(new_n16177_));
  AOI21X1  g13741(.A0(new_n16177_), .A1(new_n12743_), .B0(new_n12739_), .Y(new_n16178_));
  MX2X1    g13742(.A(new_n16156_), .B(new_n16046_), .S0(new_n12735_), .Y(new_n16179_));
  OAI21X1  g13743(.A0(new_n16073_), .A1(pi0644), .B0(new_n12739_), .Y(new_n16180_));
  AOI21X1  g13744(.A0(new_n16179_), .A1(pi0644), .B0(new_n16180_), .Y(new_n16181_));
  OR2X1    g13745(.A(new_n16181_), .B(new_n11882_), .Y(new_n16182_));
  AOI21X1  g13746(.A0(new_n16178_), .A1(new_n16175_), .B0(new_n16182_), .Y(new_n16183_));
  OAI21X1  g13747(.A0(new_n16174_), .A1(new_n16173_), .B0(new_n12743_), .Y(new_n16184_));
  AOI21X1  g13748(.A0(new_n16177_), .A1(pi0644), .B0(pi0715), .Y(new_n16185_));
  OAI21X1  g13749(.A0(new_n16073_), .A1(new_n12743_), .B0(pi0715), .Y(new_n16186_));
  AOI21X1  g13750(.A0(new_n16179_), .A1(new_n12743_), .B0(new_n16186_), .Y(new_n16187_));
  OR2X1    g13751(.A(new_n16187_), .B(pi1160), .Y(new_n16188_));
  AOI21X1  g13752(.A0(new_n16185_), .A1(new_n16184_), .B0(new_n16188_), .Y(new_n16189_));
  NOR3X1   g13753(.A(new_n16189_), .B(new_n16183_), .C(new_n12897_), .Y(new_n16190_));
  NOR3X1   g13754(.A(new_n16174_), .B(new_n16173_), .C(pi0790), .Y(new_n16191_));
  OR2X1    g13755(.A(new_n16191_), .B(new_n5118_), .Y(new_n16192_));
  AOI21X1  g13756(.A0(new_n5118_), .A1(new_n7008_), .B0(pi0057), .Y(new_n16193_));
  OAI21X1  g13757(.A0(new_n16192_), .A1(new_n16190_), .B0(new_n16193_), .Y(new_n16194_));
  AOI21X1  g13758(.A0(pi0174), .A1(pi0057), .B0(pi0832), .Y(new_n16195_));
  NOR2X1   g13759(.A(new_n2739_), .B(new_n7008_), .Y(new_n16196_));
  AOI21X1  g13760(.A0(new_n12178_), .A1(pi0759), .B0(new_n16196_), .Y(new_n16197_));
  OAI21X1  g13761(.A0(new_n14209_), .A1(new_n14944_), .B0(new_n16197_), .Y(new_n16198_));
  NOR4X1   g13762(.A(new_n13585_), .B(new_n12120_), .C(new_n14944_), .D(new_n12493_), .Y(new_n16199_));
  INVX1    g13763(.A(new_n16199_), .Y(new_n16200_));
  AOI21X1  g13764(.A0(new_n16200_), .A1(new_n16198_), .B0(pi1153), .Y(new_n16201_));
  NOR3X1   g13765(.A(new_n13585_), .B(new_n14944_), .C(new_n12493_), .Y(new_n16202_));
  NOR3X1   g13766(.A(new_n16202_), .B(new_n16196_), .C(new_n12494_), .Y(new_n16203_));
  OR2X1    g13767(.A(new_n16203_), .B(pi0608), .Y(new_n16204_));
  AOI21X1  g13768(.A0(new_n12566_), .A1(pi0696), .B0(new_n16196_), .Y(new_n16205_));
  OR2X1    g13769(.A(new_n16205_), .B(new_n16202_), .Y(new_n16206_));
  AND2X1   g13770(.A(new_n16206_), .B(new_n12494_), .Y(new_n16207_));
  NAND2X1  g13771(.A(new_n16197_), .B(pi1153), .Y(new_n16208_));
  OAI21X1  g13772(.A0(new_n16208_), .A1(new_n16199_), .B0(pi0608), .Y(new_n16209_));
  OAI22X1  g13773(.A0(new_n16209_), .A1(new_n16207_), .B0(new_n16204_), .B1(new_n16201_), .Y(new_n16210_));
  MX2X1    g13774(.A(new_n16210_), .B(new_n16198_), .S0(new_n11889_), .Y(new_n16211_));
  INVX1    g13775(.A(new_n16205_), .Y(new_n16212_));
  AOI21X1  g13776(.A0(new_n16206_), .A1(new_n12494_), .B0(new_n16203_), .Y(new_n16213_));
  MX2X1    g13777(.A(new_n16213_), .B(new_n16212_), .S0(new_n11889_), .Y(new_n16214_));
  INVX1    g13778(.A(new_n16214_), .Y(new_n16215_));
  OAI21X1  g13779(.A0(new_n16215_), .A1(new_n12590_), .B0(new_n12591_), .Y(new_n16216_));
  AOI21X1  g13780(.A0(new_n16211_), .A1(new_n12590_), .B0(new_n16216_), .Y(new_n16217_));
  NOR3X1   g13781(.A(new_n13430_), .B(new_n12204_), .C(new_n14908_), .Y(new_n16218_));
  OAI21X1  g13782(.A0(new_n2739_), .A1(new_n7008_), .B0(pi1155), .Y(new_n16219_));
  OAI21X1  g13783(.A0(new_n16219_), .A1(new_n16218_), .B0(new_n12596_), .Y(new_n16220_));
  OAI21X1  g13784(.A0(new_n16215_), .A1(pi0609), .B0(pi1155), .Y(new_n16221_));
  AOI21X1  g13785(.A0(new_n16211_), .A1(pi0609), .B0(new_n16221_), .Y(new_n16222_));
  NOR3X1   g13786(.A(new_n13436_), .B(new_n12204_), .C(new_n14908_), .Y(new_n16223_));
  OAI21X1  g13787(.A0(new_n2739_), .A1(new_n7008_), .B0(new_n12591_), .Y(new_n16224_));
  OAI21X1  g13788(.A0(new_n16224_), .A1(new_n16223_), .B0(pi0660), .Y(new_n16225_));
  OAI22X1  g13789(.A0(new_n16225_), .A1(new_n16222_), .B0(new_n16220_), .B1(new_n16217_), .Y(new_n16226_));
  MX2X1    g13790(.A(new_n16226_), .B(new_n16211_), .S0(new_n11888_), .Y(new_n16227_));
  NAND2X1  g13791(.A(new_n16227_), .B(new_n12614_), .Y(new_n16228_));
  OAI22X1  g13792(.A0(new_n16215_), .A1(new_n12618_), .B0(new_n2739_), .B1(new_n7008_), .Y(new_n16229_));
  AOI21X1  g13793(.A0(new_n16229_), .A1(pi0618), .B0(pi1154), .Y(new_n16230_));
  OR4X1    g13794(.A(new_n14178_), .B(new_n12171_), .C(new_n2740_), .D(new_n14908_), .Y(new_n16231_));
  NOR3X1   g13795(.A(new_n16231_), .B(new_n12601_), .C(new_n12614_), .Y(new_n16232_));
  OAI21X1  g13796(.A0(new_n2739_), .A1(new_n7008_), .B0(pi1154), .Y(new_n16233_));
  OAI21X1  g13797(.A0(new_n16233_), .A1(new_n16232_), .B0(new_n12622_), .Y(new_n16234_));
  AOI21X1  g13798(.A0(new_n16230_), .A1(new_n16228_), .B0(new_n16234_), .Y(new_n16235_));
  NAND2X1  g13799(.A(new_n16227_), .B(pi0618), .Y(new_n16236_));
  AOI21X1  g13800(.A0(new_n16229_), .A1(new_n12614_), .B0(new_n12615_), .Y(new_n16237_));
  NOR3X1   g13801(.A(new_n16231_), .B(new_n12601_), .C(pi0618), .Y(new_n16238_));
  OAI21X1  g13802(.A0(new_n2739_), .A1(new_n7008_), .B0(new_n12615_), .Y(new_n16239_));
  OAI21X1  g13803(.A0(new_n16239_), .A1(new_n16238_), .B0(pi0627), .Y(new_n16240_));
  AOI21X1  g13804(.A0(new_n16237_), .A1(new_n16236_), .B0(new_n16240_), .Y(new_n16241_));
  OAI21X1  g13805(.A0(new_n16241_), .A1(new_n16235_), .B0(pi0781), .Y(new_n16242_));
  INVX1    g13806(.A(new_n12658_), .Y(new_n16243_));
  NOR3X1   g13807(.A(new_n12638_), .B(new_n12645_), .C(pi0619), .Y(new_n16244_));
  NOR3X1   g13808(.A(pi1159), .B(pi0648), .C(new_n12637_), .Y(new_n16245_));
  OR2X1    g13809(.A(new_n16245_), .B(new_n16244_), .Y(new_n16246_));
  NOR2X1   g13810(.A(new_n16246_), .B(new_n16243_), .Y(new_n16247_));
  NOR2X1   g13811(.A(new_n16247_), .B(new_n11886_), .Y(new_n16248_));
  AOI21X1  g13812(.A0(new_n16227_), .A1(new_n11887_), .B0(new_n16248_), .Y(new_n16249_));
  NAND3X1  g13813(.A(new_n16214_), .B(new_n14198_), .C(new_n13598_), .Y(new_n16250_));
  OR2X1    g13814(.A(new_n12638_), .B(pi0648), .Y(new_n16251_));
  OR2X1    g13815(.A(pi1159), .B(new_n12645_), .Y(new_n16252_));
  NOR4X1   g13816(.A(new_n16231_), .B(new_n14183_), .C(new_n12601_), .D(pi0619), .Y(new_n16253_));
  NOR4X1   g13817(.A(new_n16231_), .B(new_n14183_), .C(new_n12601_), .D(new_n12637_), .Y(new_n16254_));
  OAI22X1  g13818(.A0(new_n16254_), .A1(new_n16251_), .B0(new_n16253_), .B1(new_n16252_), .Y(new_n16255_));
  AOI21X1  g13819(.A0(new_n16250_), .A1(new_n16246_), .B0(new_n16255_), .Y(new_n16256_));
  OAI21X1  g13820(.A0(new_n2739_), .A1(new_n7008_), .B0(pi0789), .Y(new_n16257_));
  OAI21X1  g13821(.A0(new_n16257_), .A1(new_n16256_), .B0(new_n12842_), .Y(new_n16258_));
  AOI21X1  g13822(.A0(new_n16249_), .A1(new_n16242_), .B0(new_n16258_), .Y(new_n16259_));
  OAI22X1  g13823(.A0(new_n16250_), .A1(new_n12659_), .B0(new_n2739_), .B1(new_n7008_), .Y(new_n16260_));
  NOR2X1   g13824(.A(new_n16231_), .B(new_n14185_), .Y(new_n16261_));
  AOI21X1  g13825(.A0(new_n16261_), .A1(new_n12664_), .B0(new_n16196_), .Y(new_n16262_));
  OAI21X1  g13826(.A0(new_n16262_), .A1(pi1158), .B0(pi0641), .Y(new_n16263_));
  AOI21X1  g13827(.A0(new_n16260_), .A1(new_n14196_), .B0(new_n16263_), .Y(new_n16264_));
  AOI21X1  g13828(.A0(new_n16261_), .A1(pi0626), .B0(new_n16196_), .Y(new_n16265_));
  OAI21X1  g13829(.A0(new_n16265_), .A1(new_n12676_), .B0(new_n12672_), .Y(new_n16266_));
  AOI21X1  g13830(.A0(new_n16260_), .A1(new_n14204_), .B0(new_n16266_), .Y(new_n16267_));
  NOR3X1   g13831(.A(new_n16267_), .B(new_n16264_), .C(new_n11885_), .Y(new_n16268_));
  OR2X1    g13832(.A(new_n16268_), .B(new_n14273_), .Y(new_n16269_));
  NOR3X1   g13833(.A(new_n16231_), .B(new_n14185_), .C(new_n12841_), .Y(new_n16270_));
  INVX1    g13834(.A(new_n16270_), .Y(new_n16271_));
  OAI21X1  g13835(.A0(new_n16271_), .A1(pi0629), .B0(pi0628), .Y(new_n16272_));
  NOR2X1   g13836(.A(new_n16215_), .B(new_n13624_), .Y(new_n16273_));
  OAI21X1  g13837(.A0(new_n16273_), .A1(new_n12689_), .B0(new_n16272_), .Y(new_n16274_));
  OAI21X1  g13838(.A0(new_n16270_), .A1(pi0628), .B0(pi0629), .Y(new_n16275_));
  NAND2X1  g13839(.A(new_n16275_), .B(pi1156), .Y(new_n16276_));
  AOI21X1  g13840(.A0(new_n16273_), .A1(pi0628), .B0(new_n16276_), .Y(new_n16277_));
  AOI21X1  g13841(.A0(new_n16274_), .A1(new_n12684_), .B0(new_n16277_), .Y(new_n16278_));
  OAI21X1  g13842(.A0(new_n2739_), .A1(new_n7008_), .B0(pi0792), .Y(new_n16279_));
  OAI22X1  g13843(.A0(new_n16279_), .A1(new_n16278_), .B0(new_n16269_), .B1(new_n16259_), .Y(new_n16280_));
  OR4X1    g13844(.A(new_n16231_), .B(new_n14185_), .C(new_n12841_), .D(new_n12711_), .Y(new_n16281_));
  OR2X1    g13845(.A(new_n16281_), .B(pi0630), .Y(new_n16282_));
  NOR3X1   g13846(.A(new_n16215_), .B(new_n13639_), .C(new_n13624_), .Y(new_n16283_));
  INVX1    g13847(.A(new_n16283_), .Y(new_n16284_));
  AOI22X1  g13848(.A0(new_n16284_), .A1(pi0630), .B0(new_n16282_), .B1(pi0647), .Y(new_n16285_));
  AOI21X1  g13849(.A0(new_n16284_), .A1(new_n12723_), .B0(new_n12705_), .Y(new_n16286_));
  OAI21X1  g13850(.A0(new_n16281_), .A1(new_n12723_), .B0(pi1157), .Y(new_n16287_));
  OAI22X1  g13851(.A0(new_n16287_), .A1(new_n16286_), .B0(new_n16285_), .B1(pi1157), .Y(new_n16288_));
  NOR2X1   g13852(.A(new_n16196_), .B(new_n11883_), .Y(new_n16289_));
  AOI22X1  g13853(.A0(new_n16289_), .A1(new_n16288_), .B0(new_n16280_), .B1(new_n14562_), .Y(new_n16290_));
  AOI21X1  g13854(.A0(new_n16283_), .A1(new_n14286_), .B0(new_n16196_), .Y(new_n16291_));
  OAI21X1  g13855(.A0(new_n16291_), .A1(pi0644), .B0(pi0715), .Y(new_n16292_));
  AOI21X1  g13856(.A0(new_n16290_), .A1(pi0644), .B0(new_n16292_), .Y(new_n16293_));
  OR2X1    g13857(.A(new_n12735_), .B(new_n12711_), .Y(new_n16294_));
  NOR3X1   g13858(.A(new_n16294_), .B(new_n16271_), .C(new_n12743_), .Y(new_n16295_));
  OAI21X1  g13859(.A0(new_n2739_), .A1(new_n7008_), .B0(new_n12739_), .Y(new_n16296_));
  OAI21X1  g13860(.A0(new_n16296_), .A1(new_n16295_), .B0(pi1160), .Y(new_n16297_));
  OAI21X1  g13861(.A0(new_n16291_), .A1(new_n12743_), .B0(new_n12739_), .Y(new_n16298_));
  AOI21X1  g13862(.A0(new_n16290_), .A1(new_n12743_), .B0(new_n16298_), .Y(new_n16299_));
  NOR3X1   g13863(.A(new_n16294_), .B(new_n16271_), .C(pi0644), .Y(new_n16300_));
  OAI21X1  g13864(.A0(new_n2739_), .A1(new_n7008_), .B0(pi0715), .Y(new_n16301_));
  OAI21X1  g13865(.A0(new_n16301_), .A1(new_n16300_), .B0(new_n11882_), .Y(new_n16302_));
  OAI22X1  g13866(.A0(new_n16302_), .A1(new_n16299_), .B0(new_n16297_), .B1(new_n16293_), .Y(new_n16303_));
  NAND2X1  g13867(.A(new_n16303_), .B(pi0790), .Y(new_n16304_));
  AOI21X1  g13868(.A0(new_n16290_), .A1(new_n12897_), .B0(new_n12898_), .Y(new_n16305_));
  AOI22X1  g13869(.A0(new_n16305_), .A1(new_n16304_), .B0(new_n16195_), .B1(new_n16194_), .Y(po0331));
  AOI21X1  g13870(.A0(pi1093), .A1(pi1092), .B0(pi0175), .Y(new_n16307_));
  INVX1    g13871(.A(new_n16307_), .Y(new_n16308_));
  AOI21X1  g13872(.A0(new_n12178_), .A1(pi0766), .B0(new_n16307_), .Y(new_n16309_));
  AOI21X1  g13873(.A0(new_n12601_), .A1(new_n2739_), .B0(new_n16309_), .Y(new_n16310_));
  AND2X1   g13874(.A(new_n12178_), .B(pi0766), .Y(new_n16311_));
  AND2X1   g13875(.A(new_n16311_), .B(new_n12608_), .Y(new_n16312_));
  INVX1    g13876(.A(new_n16312_), .Y(new_n16313_));
  AOI21X1  g13877(.A0(new_n16313_), .A1(new_n16310_), .B0(new_n12591_), .Y(new_n16314_));
  NOR3X1   g13878(.A(new_n16312_), .B(new_n16307_), .C(pi1155), .Y(new_n16315_));
  OAI21X1  g13879(.A0(new_n16315_), .A1(new_n16314_), .B0(pi0785), .Y(new_n16316_));
  OAI21X1  g13880(.A0(new_n16310_), .A1(pi0785), .B0(new_n16316_), .Y(new_n16317_));
  INVX1    g13881(.A(new_n16317_), .Y(new_n16318_));
  AOI21X1  g13882(.A0(new_n16318_), .A1(new_n12785_), .B0(new_n12615_), .Y(new_n16319_));
  AOI21X1  g13883(.A0(new_n16318_), .A1(new_n12788_), .B0(pi1154), .Y(new_n16320_));
  NOR2X1   g13884(.A(new_n16320_), .B(new_n16319_), .Y(new_n16321_));
  MX2X1    g13885(.A(new_n16321_), .B(new_n16318_), .S0(new_n11887_), .Y(new_n16322_));
  OR2X1    g13886(.A(new_n16322_), .B(pi0789), .Y(new_n16323_));
  AOI21X1  g13887(.A0(new_n16322_), .A1(new_n15910_), .B0(new_n12638_), .Y(new_n16324_));
  AOI21X1  g13888(.A0(new_n16322_), .A1(new_n15912_), .B0(pi1159), .Y(new_n16325_));
  OAI21X1  g13889(.A0(new_n16325_), .A1(new_n16324_), .B0(pi0789), .Y(new_n16326_));
  AND2X1   g13890(.A(new_n16326_), .B(new_n16323_), .Y(new_n16327_));
  INVX1    g13891(.A(new_n16327_), .Y(new_n16328_));
  MX2X1    g13892(.A(new_n16328_), .B(new_n16308_), .S0(new_n12841_), .Y(new_n16329_));
  MX2X1    g13893(.A(new_n16329_), .B(new_n16308_), .S0(new_n12711_), .Y(new_n16330_));
  AOI21X1  g13894(.A0(new_n12566_), .A1(pi0700), .B0(new_n16307_), .Y(new_n16331_));
  INVX1    g13895(.A(new_n16331_), .Y(new_n16332_));
  NOR3X1   g13896(.A(new_n13585_), .B(new_n15022_), .C(pi0625), .Y(new_n16333_));
  OR2X1    g13897(.A(new_n16333_), .B(new_n16331_), .Y(new_n16334_));
  NOR2X1   g13898(.A(new_n16307_), .B(pi1153), .Y(new_n16335_));
  INVX1    g13899(.A(new_n16335_), .Y(new_n16336_));
  OAI21X1  g13900(.A0(new_n16336_), .A1(new_n16333_), .B0(pi0778), .Y(new_n16337_));
  AOI21X1  g13901(.A0(new_n16334_), .A1(pi1153), .B0(new_n16337_), .Y(new_n16338_));
  AOI21X1  g13902(.A0(new_n16332_), .A1(new_n11889_), .B0(new_n16338_), .Y(new_n16339_));
  NOR4X1   g13903(.A(new_n16339_), .B(new_n12765_), .C(new_n12764_), .D(new_n12762_), .Y(new_n16340_));
  INVX1    g13904(.A(new_n16340_), .Y(new_n16341_));
  NOR3X1   g13905(.A(new_n16341_), .B(new_n12870_), .C(new_n12851_), .Y(new_n16342_));
  INVX1    g13906(.A(new_n16342_), .Y(new_n16343_));
  AOI21X1  g13907(.A0(new_n16307_), .A1(pi0647), .B0(pi1157), .Y(new_n16344_));
  OAI21X1  g13908(.A0(new_n16343_), .A1(pi0647), .B0(new_n16344_), .Y(new_n16345_));
  MX2X1    g13909(.A(new_n16342_), .B(new_n16307_), .S0(new_n12705_), .Y(new_n16346_));
  OAI22X1  g13910(.A0(new_n16346_), .A1(new_n14387_), .B0(new_n16345_), .B1(new_n12723_), .Y(new_n16347_));
  AOI21X1  g13911(.A0(new_n16330_), .A1(new_n14385_), .B0(new_n16347_), .Y(new_n16348_));
  NOR2X1   g13912(.A(new_n16348_), .B(new_n11883_), .Y(new_n16349_));
  INVX1    g13913(.A(new_n14273_), .Y(new_n16350_));
  AND2X1   g13914(.A(new_n12676_), .B(pi0641), .Y(new_n16351_));
  INVX1    g13915(.A(new_n16351_), .Y(new_n16352_));
  AOI21X1  g13916(.A0(new_n16308_), .A1(pi0626), .B0(new_n16352_), .Y(new_n16353_));
  OAI21X1  g13917(.A0(new_n16327_), .A1(pi0626), .B0(new_n16353_), .Y(new_n16354_));
  AND2X1   g13918(.A(pi1158), .B(new_n12672_), .Y(new_n16355_));
  INVX1    g13919(.A(new_n16355_), .Y(new_n16356_));
  AOI21X1  g13920(.A0(new_n16326_), .A1(new_n16323_), .B0(new_n12664_), .Y(new_n16357_));
  NOR2X1   g13921(.A(new_n16307_), .B(pi0626), .Y(new_n16358_));
  NOR3X1   g13922(.A(new_n16358_), .B(new_n16357_), .C(new_n16356_), .Y(new_n16359_));
  AOI21X1  g13923(.A0(new_n16340_), .A1(new_n12769_), .B0(new_n16359_), .Y(new_n16360_));
  AOI21X1  g13924(.A0(new_n16360_), .A1(new_n16354_), .B0(new_n11885_), .Y(new_n16361_));
  INVX1    g13925(.A(new_n16309_), .Y(new_n16362_));
  AOI21X1  g13926(.A0(new_n16332_), .A1(new_n12171_), .B0(new_n16362_), .Y(new_n16363_));
  NOR3X1   g13927(.A(new_n16331_), .B(new_n12120_), .C(new_n12493_), .Y(new_n16364_));
  OR2X1    g13928(.A(new_n16363_), .B(new_n16364_), .Y(new_n16365_));
  NOR2X1   g13929(.A(new_n16333_), .B(new_n16331_), .Y(new_n16366_));
  OAI21X1  g13930(.A0(new_n16366_), .A1(new_n12494_), .B0(new_n12584_), .Y(new_n16367_));
  AOI21X1  g13931(.A0(new_n16365_), .A1(new_n16335_), .B0(new_n16367_), .Y(new_n16368_));
  NOR3X1   g13932(.A(new_n16364_), .B(new_n16362_), .C(new_n12494_), .Y(new_n16369_));
  OAI21X1  g13933(.A0(new_n16336_), .A1(new_n16333_), .B0(pi0608), .Y(new_n16370_));
  NOR2X1   g13934(.A(new_n16370_), .B(new_n16369_), .Y(new_n16371_));
  OAI21X1  g13935(.A0(new_n16371_), .A1(new_n16368_), .B0(pi0778), .Y(new_n16372_));
  OAI21X1  g13936(.A0(new_n16363_), .A1(pi0778), .B0(new_n16372_), .Y(new_n16373_));
  OAI21X1  g13937(.A0(new_n16339_), .A1(new_n12590_), .B0(new_n12591_), .Y(new_n16374_));
  AOI21X1  g13938(.A0(new_n16373_), .A1(new_n12590_), .B0(new_n16374_), .Y(new_n16375_));
  NOR3X1   g13939(.A(new_n16375_), .B(new_n16314_), .C(pi0660), .Y(new_n16376_));
  OAI21X1  g13940(.A0(new_n16339_), .A1(pi0609), .B0(pi1155), .Y(new_n16377_));
  AOI21X1  g13941(.A0(new_n16373_), .A1(pi0609), .B0(new_n16377_), .Y(new_n16378_));
  NOR3X1   g13942(.A(new_n16378_), .B(new_n16315_), .C(new_n12596_), .Y(new_n16379_));
  OAI21X1  g13943(.A0(new_n16379_), .A1(new_n16376_), .B0(pi0785), .Y(new_n16380_));
  NAND2X1  g13944(.A(new_n16373_), .B(new_n11888_), .Y(new_n16381_));
  AND2X1   g13945(.A(new_n16381_), .B(new_n16380_), .Y(new_n16382_));
  NOR3X1   g13946(.A(new_n16339_), .B(new_n12762_), .C(new_n12614_), .Y(new_n16383_));
  NOR2X1   g13947(.A(new_n16383_), .B(pi1154), .Y(new_n16384_));
  OAI21X1  g13948(.A0(new_n16382_), .A1(pi0618), .B0(new_n16384_), .Y(new_n16385_));
  NOR2X1   g13949(.A(new_n16319_), .B(pi0627), .Y(new_n16386_));
  NOR3X1   g13950(.A(new_n16339_), .B(new_n12762_), .C(pi0618), .Y(new_n16387_));
  NOR2X1   g13951(.A(new_n16387_), .B(new_n12615_), .Y(new_n16388_));
  OAI21X1  g13952(.A0(new_n16382_), .A1(new_n12614_), .B0(new_n16388_), .Y(new_n16389_));
  NOR2X1   g13953(.A(new_n16320_), .B(new_n12622_), .Y(new_n16390_));
  AOI22X1  g13954(.A0(new_n16390_), .A1(new_n16389_), .B0(new_n16386_), .B1(new_n16385_), .Y(new_n16391_));
  MX2X1    g13955(.A(new_n16391_), .B(new_n16382_), .S0(new_n11887_), .Y(new_n16392_));
  OR4X1    g13956(.A(new_n16339_), .B(new_n12764_), .C(new_n12762_), .D(new_n12637_), .Y(new_n16393_));
  AND2X1   g13957(.A(new_n16393_), .B(new_n12638_), .Y(new_n16394_));
  OAI21X1  g13958(.A0(new_n16392_), .A1(pi0619), .B0(new_n16394_), .Y(new_n16395_));
  NOR2X1   g13959(.A(new_n16324_), .B(pi0648), .Y(new_n16396_));
  AND2X1   g13960(.A(new_n16396_), .B(new_n16395_), .Y(new_n16397_));
  INVX1    g13961(.A(new_n16397_), .Y(new_n16398_));
  NOR4X1   g13962(.A(new_n16339_), .B(new_n12764_), .C(new_n12762_), .D(pi0619), .Y(new_n16399_));
  NOR2X1   g13963(.A(new_n16399_), .B(new_n12638_), .Y(new_n16400_));
  OAI21X1  g13964(.A0(new_n16392_), .A1(new_n12637_), .B0(new_n16400_), .Y(new_n16401_));
  NOR2X1   g13965(.A(new_n16325_), .B(new_n12645_), .Y(new_n16402_));
  AOI21X1  g13966(.A0(new_n16402_), .A1(new_n16401_), .B0(new_n11886_), .Y(new_n16403_));
  AOI21X1  g13967(.A0(new_n16392_), .A1(new_n11886_), .B0(new_n14264_), .Y(new_n16404_));
  INVX1    g13968(.A(new_n16404_), .Y(new_n16405_));
  AOI21X1  g13969(.A0(new_n16403_), .A1(new_n16398_), .B0(new_n16405_), .Y(new_n16406_));
  OAI21X1  g13970(.A0(new_n16406_), .A1(new_n16361_), .B0(new_n16350_), .Y(new_n16407_));
  INVX1    g13971(.A(new_n16329_), .Y(new_n16408_));
  AND2X1   g13972(.A(new_n16340_), .B(new_n12852_), .Y(new_n16409_));
  AOI22X1  g13973(.A0(new_n16409_), .A1(new_n14564_), .B0(new_n16408_), .B1(new_n12867_), .Y(new_n16410_));
  AOI22X1  g13974(.A0(new_n16409_), .A1(new_n14566_), .B0(new_n16408_), .B1(new_n12865_), .Y(new_n16411_));
  MX2X1    g13975(.A(new_n16411_), .B(new_n16410_), .S0(new_n12689_), .Y(new_n16412_));
  OAI21X1  g13976(.A0(new_n16412_), .A1(new_n11884_), .B0(new_n14562_), .Y(new_n16413_));
  INVX1    g13977(.A(new_n16413_), .Y(new_n16414_));
  AOI21X1  g13978(.A0(new_n16414_), .A1(new_n16407_), .B0(new_n16349_), .Y(new_n16415_));
  OAI21X1  g13979(.A0(new_n16346_), .A1(new_n12706_), .B0(new_n16345_), .Y(new_n16416_));
  MX2X1    g13980(.A(new_n16416_), .B(new_n16343_), .S0(new_n11883_), .Y(new_n16417_));
  OAI21X1  g13981(.A0(new_n16417_), .A1(pi0644), .B0(pi0715), .Y(new_n16418_));
  AOI21X1  g13982(.A0(new_n16415_), .A1(pi0644), .B0(new_n16418_), .Y(new_n16419_));
  OR4X1    g13983(.A(new_n12734_), .B(new_n2739_), .C(new_n11883_), .D(pi0175), .Y(new_n16420_));
  OAI21X1  g13984(.A0(new_n16330_), .A1(new_n12735_), .B0(new_n16420_), .Y(new_n16421_));
  OAI21X1  g13985(.A0(new_n16308_), .A1(pi0644), .B0(new_n12739_), .Y(new_n16422_));
  AOI21X1  g13986(.A0(new_n16421_), .A1(pi0644), .B0(new_n16422_), .Y(new_n16423_));
  OR2X1    g13987(.A(new_n16423_), .B(new_n11882_), .Y(new_n16424_));
  OAI21X1  g13988(.A0(new_n16417_), .A1(new_n12743_), .B0(new_n12739_), .Y(new_n16425_));
  AOI21X1  g13989(.A0(new_n16415_), .A1(new_n12743_), .B0(new_n16425_), .Y(new_n16426_));
  OAI21X1  g13990(.A0(new_n16308_), .A1(new_n12743_), .B0(pi0715), .Y(new_n16427_));
  AOI21X1  g13991(.A0(new_n16421_), .A1(new_n12743_), .B0(new_n16427_), .Y(new_n16428_));
  OR2X1    g13992(.A(new_n16428_), .B(pi1160), .Y(new_n16429_));
  OAI22X1  g13993(.A0(new_n16429_), .A1(new_n16426_), .B0(new_n16424_), .B1(new_n16419_), .Y(new_n16430_));
  NAND2X1  g13994(.A(new_n16430_), .B(pi0790), .Y(new_n16431_));
  AOI21X1  g13995(.A0(new_n16415_), .A1(new_n12897_), .B0(new_n12898_), .Y(new_n16432_));
  AOI21X1  g13996(.A0(new_n13699_), .A1(new_n3129_), .B0(pi0175), .Y(new_n16433_));
  INVX1    g13997(.A(new_n16433_), .Y(new_n16434_));
  MX2X1    g13998(.A(new_n12560_), .B(new_n13391_), .S0(new_n2959_), .Y(new_n16435_));
  MX2X1    g13999(.A(new_n12522_), .B(new_n13685_), .S0(new_n2959_), .Y(new_n16436_));
  OAI21X1  g14000(.A0(new_n16436_), .A1(new_n11203_), .B0(new_n2996_), .Y(new_n16437_));
  AOI21X1  g14001(.A0(new_n16435_), .A1(new_n11203_), .B0(new_n16437_), .Y(new_n16438_));
  AOI21X1  g14002(.A0(new_n12901_), .A1(new_n11203_), .B0(new_n12568_), .Y(new_n16439_));
  NOR3X1   g14003(.A(new_n16439_), .B(new_n16438_), .C(new_n15022_), .Y(new_n16440_));
  OR2X1    g14004(.A(pi0700), .B(pi0175), .Y(new_n16441_));
  OAI21X1  g14005(.A0(new_n16441_), .A1(new_n13699_), .B0(new_n3129_), .Y(new_n16442_));
  OAI22X1  g14006(.A0(new_n16442_), .A1(new_n16440_), .B0(new_n3129_), .B1(new_n11203_), .Y(new_n16443_));
  AND2X1   g14007(.A(new_n16443_), .B(new_n11889_), .Y(new_n16444_));
  AOI21X1  g14008(.A0(new_n16433_), .A1(new_n12493_), .B0(new_n12494_), .Y(new_n16445_));
  OAI21X1  g14009(.A0(new_n16443_), .A1(new_n12493_), .B0(new_n16445_), .Y(new_n16446_));
  AOI21X1  g14010(.A0(new_n16433_), .A1(pi0625), .B0(pi1153), .Y(new_n16447_));
  OAI21X1  g14011(.A0(new_n16443_), .A1(pi0625), .B0(new_n16447_), .Y(new_n16448_));
  AOI21X1  g14012(.A0(new_n16448_), .A1(new_n16446_), .B0(new_n11889_), .Y(new_n16449_));
  NOR2X1   g14013(.A(new_n16449_), .B(new_n16444_), .Y(new_n16450_));
  MX2X1    g14014(.A(new_n16450_), .B(new_n16433_), .S0(new_n12618_), .Y(new_n16451_));
  AND2X1   g14015(.A(new_n16433_), .B(new_n12641_), .Y(new_n16452_));
  AOI21X1  g14016(.A0(new_n16451_), .A1(new_n14198_), .B0(new_n16452_), .Y(new_n16453_));
  MX2X1    g14017(.A(new_n16453_), .B(new_n16434_), .S0(new_n12659_), .Y(new_n16454_));
  MX2X1    g14018(.A(new_n16454_), .B(new_n16434_), .S0(new_n12691_), .Y(new_n16455_));
  MX2X1    g14019(.A(new_n16455_), .B(new_n16434_), .S0(pi0628), .Y(new_n16456_));
  MX2X1    g14020(.A(new_n16455_), .B(new_n16434_), .S0(new_n12683_), .Y(new_n16457_));
  MX2X1    g14021(.A(new_n16457_), .B(new_n16456_), .S0(new_n12684_), .Y(new_n16458_));
  MX2X1    g14022(.A(new_n16458_), .B(new_n16455_), .S0(new_n11884_), .Y(new_n16459_));
  MX2X1    g14023(.A(new_n16459_), .B(new_n16434_), .S0(pi0647), .Y(new_n16460_));
  MX2X1    g14024(.A(new_n16459_), .B(new_n16434_), .S0(new_n12705_), .Y(new_n16461_));
  MX2X1    g14025(.A(new_n16461_), .B(new_n16460_), .S0(new_n12706_), .Y(new_n16462_));
  MX2X1    g14026(.A(new_n16462_), .B(new_n16459_), .S0(new_n11883_), .Y(new_n16463_));
  OAI21X1  g14027(.A0(new_n16463_), .A1(pi0644), .B0(pi0715), .Y(new_n16464_));
  OAI22X1  g14028(.A0(new_n12904_), .A1(new_n11203_), .B0(new_n12089_), .B1(pi0766), .Y(new_n16465_));
  NAND2X1  g14029(.A(new_n16465_), .B(pi0039), .Y(new_n16466_));
  AND2X1   g14030(.A(pi0766), .B(new_n11203_), .Y(new_n16467_));
  AOI21X1  g14031(.A0(new_n13683_), .A1(new_n2959_), .B0(new_n14977_), .Y(new_n16468_));
  OAI21X1  g14032(.A0(new_n16468_), .A1(new_n11203_), .B0(new_n14983_), .Y(new_n16469_));
  AOI21X1  g14033(.A0(new_n16467_), .A1(new_n12162_), .B0(new_n16469_), .Y(new_n16470_));
  AOI21X1  g14034(.A0(new_n16470_), .A1(new_n16466_), .B0(pi0038), .Y(new_n16471_));
  OAI21X1  g14035(.A0(new_n12202_), .A1(pi0175), .B0(pi0038), .Y(new_n16472_));
  AOI21X1  g14036(.A0(new_n12205_), .A1(pi0766), .B0(new_n16472_), .Y(new_n16473_));
  NOR2X1   g14037(.A(new_n16473_), .B(new_n16471_), .Y(new_n16474_));
  MX2X1    g14038(.A(new_n16474_), .B(new_n11203_), .S0(new_n3810_), .Y(new_n16475_));
  MX2X1    g14039(.A(new_n16475_), .B(new_n16433_), .S0(new_n12601_), .Y(new_n16476_));
  NOR2X1   g14040(.A(new_n16475_), .B(new_n12601_), .Y(new_n16477_));
  AOI22X1  g14041(.A0(new_n16477_), .A1(pi0609), .B0(new_n16434_), .B1(new_n13430_), .Y(new_n16478_));
  AOI22X1  g14042(.A0(new_n16477_), .A1(new_n12590_), .B0(new_n16434_), .B1(new_n13436_), .Y(new_n16479_));
  MX2X1    g14043(.A(new_n16479_), .B(new_n16478_), .S0(pi1155), .Y(new_n16480_));
  MX2X1    g14044(.A(new_n16480_), .B(new_n16476_), .S0(new_n11888_), .Y(new_n16481_));
  OAI21X1  g14045(.A0(new_n16434_), .A1(pi0618), .B0(pi1154), .Y(new_n16482_));
  AOI21X1  g14046(.A0(new_n16481_), .A1(pi0618), .B0(new_n16482_), .Y(new_n16483_));
  OAI21X1  g14047(.A0(new_n16434_), .A1(new_n12614_), .B0(new_n12615_), .Y(new_n16484_));
  AOI21X1  g14048(.A0(new_n16481_), .A1(new_n12614_), .B0(new_n16484_), .Y(new_n16485_));
  NOR2X1   g14049(.A(new_n16485_), .B(new_n16483_), .Y(new_n16486_));
  MX2X1    g14050(.A(new_n16486_), .B(new_n16481_), .S0(new_n11887_), .Y(new_n16487_));
  OAI21X1  g14051(.A0(new_n16434_), .A1(pi0619), .B0(pi1159), .Y(new_n16488_));
  AOI21X1  g14052(.A0(new_n16487_), .A1(pi0619), .B0(new_n16488_), .Y(new_n16489_));
  OAI21X1  g14053(.A0(new_n16434_), .A1(new_n12637_), .B0(new_n12638_), .Y(new_n16490_));
  AOI21X1  g14054(.A0(new_n16487_), .A1(new_n12637_), .B0(new_n16490_), .Y(new_n16491_));
  NOR2X1   g14055(.A(new_n16491_), .B(new_n16489_), .Y(new_n16492_));
  MX2X1    g14056(.A(new_n16492_), .B(new_n16487_), .S0(new_n11886_), .Y(new_n16493_));
  MX2X1    g14057(.A(new_n16493_), .B(new_n16433_), .S0(new_n12841_), .Y(new_n16494_));
  MX2X1    g14058(.A(new_n16494_), .B(new_n16433_), .S0(new_n12711_), .Y(new_n16495_));
  MX2X1    g14059(.A(new_n16495_), .B(new_n16433_), .S0(new_n12735_), .Y(new_n16496_));
  OAI21X1  g14060(.A0(new_n16434_), .A1(pi0644), .B0(new_n12739_), .Y(new_n16497_));
  AOI21X1  g14061(.A0(new_n16496_), .A1(pi0644), .B0(new_n16497_), .Y(new_n16498_));
  NOR2X1   g14062(.A(new_n16498_), .B(new_n11882_), .Y(new_n16499_));
  OAI21X1  g14063(.A0(new_n16463_), .A1(new_n12743_), .B0(new_n12739_), .Y(new_n16500_));
  OAI21X1  g14064(.A0(new_n16434_), .A1(new_n12743_), .B0(pi0715), .Y(new_n16501_));
  AOI21X1  g14065(.A0(new_n16496_), .A1(new_n12743_), .B0(new_n16501_), .Y(new_n16502_));
  NOR2X1   g14066(.A(new_n16502_), .B(pi1160), .Y(new_n16503_));
  AOI22X1  g14067(.A0(new_n16503_), .A1(new_n16500_), .B0(new_n16499_), .B1(new_n16464_), .Y(new_n16504_));
  NOR3X1   g14068(.A(new_n16502_), .B(pi1160), .C(pi0644), .Y(new_n16505_));
  NOR3X1   g14069(.A(new_n16498_), .B(new_n11882_), .C(new_n12743_), .Y(new_n16506_));
  NOR3X1   g14070(.A(new_n16506_), .B(new_n16505_), .C(new_n12897_), .Y(new_n16507_));
  AOI22X1  g14071(.A0(new_n16457_), .A1(new_n12707_), .B0(new_n16456_), .B1(new_n12709_), .Y(new_n16508_));
  OAI21X1  g14072(.A0(new_n16494_), .A1(new_n14395_), .B0(new_n16508_), .Y(new_n16509_));
  NOR3X1   g14073(.A(new_n16473_), .B(new_n16471_), .C(pi0700), .Y(new_n16510_));
  INVX1    g14074(.A(new_n16510_), .Y(new_n16511_));
  AOI21X1  g14075(.A0(new_n13989_), .A1(pi0175), .B0(pi0766), .Y(new_n16512_));
  OAI21X1  g14076(.A0(new_n13986_), .A1(pi0175), .B0(new_n16512_), .Y(new_n16513_));
  OAI21X1  g14077(.A0(new_n12440_), .A1(pi0175), .B0(pi0766), .Y(new_n16514_));
  AOI21X1  g14078(.A0(new_n12401_), .A1(pi0175), .B0(new_n16514_), .Y(new_n16515_));
  NOR2X1   g14079(.A(new_n16515_), .B(new_n2959_), .Y(new_n16516_));
  AND2X1   g14080(.A(new_n16516_), .B(new_n16513_), .Y(new_n16517_));
  AOI21X1  g14081(.A0(new_n13995_), .A1(pi0175), .B0(pi0766), .Y(new_n16518_));
  OAI21X1  g14082(.A0(new_n13996_), .A1(pi0175), .B0(new_n16518_), .Y(new_n16519_));
  AOI21X1  g14083(.A0(new_n12453_), .A1(new_n12104_), .B0(pi0175), .Y(new_n16520_));
  INVX1    g14084(.A(new_n16520_), .Y(new_n16521_));
  AOI21X1  g14085(.A0(new_n12929_), .A1(pi0175), .B0(new_n14977_), .Y(new_n16522_));
  AOI21X1  g14086(.A0(new_n16522_), .A1(new_n16521_), .B0(pi0039), .Y(new_n16523_));
  AOI21X1  g14087(.A0(new_n16523_), .A1(new_n16519_), .B0(pi0038), .Y(new_n16524_));
  INVX1    g14088(.A(new_n16524_), .Y(new_n16525_));
  NOR4X1   g14089(.A(new_n12211_), .B(new_n3003_), .C(new_n2740_), .D(new_n2555_), .Y(new_n16526_));
  AOI21X1  g14090(.A0(new_n16526_), .A1(new_n14977_), .B0(new_n12478_), .Y(new_n16527_));
  OAI21X1  g14091(.A0(new_n16527_), .A1(pi0039), .B0(new_n11203_), .Y(new_n16528_));
  OAI21X1  g14092(.A0(new_n16311_), .A1(new_n13576_), .B0(pi0175), .Y(new_n16529_));
  OAI21X1  g14093(.A0(new_n16529_), .A1(new_n14411_), .B0(pi0038), .Y(new_n16530_));
  INVX1    g14094(.A(new_n16530_), .Y(new_n16531_));
  AOI21X1  g14095(.A0(new_n16531_), .A1(new_n16528_), .B0(new_n15022_), .Y(new_n16532_));
  OAI21X1  g14096(.A0(new_n16525_), .A1(new_n16517_), .B0(new_n16532_), .Y(new_n16533_));
  AND2X1   g14097(.A(new_n16533_), .B(new_n3129_), .Y(new_n16534_));
  AOI22X1  g14098(.A0(new_n16534_), .A1(new_n16511_), .B0(new_n3810_), .B1(pi0175), .Y(new_n16535_));
  INVX1    g14099(.A(new_n16535_), .Y(new_n16536_));
  AOI21X1  g14100(.A0(new_n16475_), .A1(pi0625), .B0(pi1153), .Y(new_n16537_));
  OAI21X1  g14101(.A0(new_n16536_), .A1(pi0625), .B0(new_n16537_), .Y(new_n16538_));
  AND2X1   g14102(.A(new_n16446_), .B(new_n12584_), .Y(new_n16539_));
  AOI21X1  g14103(.A0(new_n16475_), .A1(new_n12493_), .B0(new_n12494_), .Y(new_n16540_));
  OAI21X1  g14104(.A0(new_n16536_), .A1(new_n12493_), .B0(new_n16540_), .Y(new_n16541_));
  AND2X1   g14105(.A(new_n16448_), .B(pi0608), .Y(new_n16542_));
  AOI22X1  g14106(.A0(new_n16542_), .A1(new_n16541_), .B0(new_n16539_), .B1(new_n16538_), .Y(new_n16543_));
  MX2X1    g14107(.A(new_n16543_), .B(new_n16536_), .S0(new_n11889_), .Y(new_n16544_));
  AOI21X1  g14108(.A0(new_n16450_), .A1(pi0609), .B0(pi1155), .Y(new_n16545_));
  OAI21X1  g14109(.A0(new_n16544_), .A1(pi0609), .B0(new_n16545_), .Y(new_n16546_));
  OAI21X1  g14110(.A0(new_n16478_), .A1(new_n12591_), .B0(new_n12596_), .Y(new_n16547_));
  INVX1    g14111(.A(new_n16547_), .Y(new_n16548_));
  AOI21X1  g14112(.A0(new_n16450_), .A1(new_n12590_), .B0(new_n12591_), .Y(new_n16549_));
  OAI21X1  g14113(.A0(new_n16544_), .A1(new_n12590_), .B0(new_n16549_), .Y(new_n16550_));
  OAI21X1  g14114(.A0(new_n16479_), .A1(pi1155), .B0(pi0660), .Y(new_n16551_));
  INVX1    g14115(.A(new_n16551_), .Y(new_n16552_));
  AOI22X1  g14116(.A0(new_n16552_), .A1(new_n16550_), .B0(new_n16548_), .B1(new_n16546_), .Y(new_n16553_));
  MX2X1    g14117(.A(new_n16553_), .B(new_n16544_), .S0(new_n11888_), .Y(new_n16554_));
  AOI21X1  g14118(.A0(new_n16451_), .A1(pi0618), .B0(pi1154), .Y(new_n16555_));
  OAI21X1  g14119(.A0(new_n16554_), .A1(pi0618), .B0(new_n16555_), .Y(new_n16556_));
  NOR2X1   g14120(.A(new_n16483_), .B(pi0627), .Y(new_n16557_));
  AOI21X1  g14121(.A0(new_n16451_), .A1(new_n12614_), .B0(new_n12615_), .Y(new_n16558_));
  OAI21X1  g14122(.A0(new_n16554_), .A1(new_n12614_), .B0(new_n16558_), .Y(new_n16559_));
  NOR2X1   g14123(.A(new_n16485_), .B(new_n12622_), .Y(new_n16560_));
  AOI22X1  g14124(.A0(new_n16560_), .A1(new_n16559_), .B0(new_n16557_), .B1(new_n16556_), .Y(new_n16561_));
  MX2X1    g14125(.A(new_n16561_), .B(new_n16554_), .S0(new_n11887_), .Y(new_n16562_));
  INVX1    g14126(.A(new_n16562_), .Y(new_n16563_));
  OAI21X1  g14127(.A0(new_n16453_), .A1(new_n12637_), .B0(new_n12638_), .Y(new_n16564_));
  AOI21X1  g14128(.A0(new_n16563_), .A1(new_n12637_), .B0(new_n16564_), .Y(new_n16565_));
  NOR3X1   g14129(.A(new_n16565_), .B(new_n16489_), .C(pi0648), .Y(new_n16566_));
  OAI21X1  g14130(.A0(new_n16453_), .A1(pi0619), .B0(pi1159), .Y(new_n16567_));
  AOI21X1  g14131(.A0(new_n16563_), .A1(pi0619), .B0(new_n16567_), .Y(new_n16568_));
  OR2X1    g14132(.A(new_n16491_), .B(new_n12645_), .Y(new_n16569_));
  OAI21X1  g14133(.A0(new_n16569_), .A1(new_n16568_), .B0(pi0789), .Y(new_n16570_));
  AOI21X1  g14134(.A0(new_n16562_), .A1(new_n11886_), .B0(new_n14264_), .Y(new_n16571_));
  OAI21X1  g14135(.A0(new_n16570_), .A1(new_n16566_), .B0(new_n16571_), .Y(new_n16572_));
  AOI21X1  g14136(.A0(new_n16434_), .A1(pi0626), .B0(new_n16352_), .Y(new_n16573_));
  OAI21X1  g14137(.A0(new_n16493_), .A1(pi0626), .B0(new_n16573_), .Y(new_n16574_));
  AOI21X1  g14138(.A0(new_n16434_), .A1(new_n12664_), .B0(new_n16356_), .Y(new_n16575_));
  OAI21X1  g14139(.A0(new_n16493_), .A1(new_n12664_), .B0(new_n16575_), .Y(new_n16576_));
  OR2X1    g14140(.A(new_n16454_), .B(new_n12770_), .Y(new_n16577_));
  NAND3X1  g14141(.A(new_n16577_), .B(new_n16576_), .C(new_n16574_), .Y(new_n16578_));
  AOI21X1  g14142(.A0(new_n16578_), .A1(pi0788), .B0(new_n14273_), .Y(new_n16579_));
  AOI22X1  g14143(.A0(new_n16579_), .A1(new_n16572_), .B0(new_n16509_), .B1(pi0792), .Y(new_n16580_));
  NOR2X1   g14144(.A(new_n16495_), .B(new_n14384_), .Y(new_n16581_));
  AND2X1   g14145(.A(new_n16461_), .B(new_n14386_), .Y(new_n16582_));
  AND2X1   g14146(.A(new_n16460_), .B(new_n14388_), .Y(new_n16583_));
  OR2X1    g14147(.A(new_n16583_), .B(new_n16582_), .Y(new_n16584_));
  OAI21X1  g14148(.A0(new_n16584_), .A1(new_n16581_), .B0(pi0787), .Y(new_n16585_));
  OAI21X1  g14149(.A0(new_n16580_), .A1(new_n14269_), .B0(new_n16585_), .Y(new_n16586_));
  OAI22X1  g14150(.A0(new_n16586_), .A1(new_n16507_), .B0(new_n16504_), .B1(new_n12897_), .Y(new_n16587_));
  OAI21X1  g14151(.A0(new_n6520_), .A1(pi0175), .B0(new_n12898_), .Y(new_n16588_));
  AOI21X1  g14152(.A0(new_n16587_), .A1(new_n6520_), .B0(new_n16588_), .Y(new_n16589_));
  AOI21X1  g14153(.A0(new_n16432_), .A1(new_n16431_), .B0(new_n16589_), .Y(po0332));
  AOI21X1  g14154(.A0(pi1093), .A1(pi1092), .B0(pi0176), .Y(new_n16591_));
  INVX1    g14155(.A(new_n16591_), .Y(new_n16592_));
  AOI21X1  g14156(.A0(new_n12178_), .A1(new_n15046_), .B0(new_n16591_), .Y(new_n16593_));
  AOI21X1  g14157(.A0(new_n12601_), .A1(new_n2739_), .B0(new_n16593_), .Y(new_n16594_));
  INVX1    g14158(.A(new_n16593_), .Y(new_n16595_));
  AOI21X1  g14159(.A0(new_n16595_), .A1(new_n12776_), .B0(new_n12591_), .Y(new_n16596_));
  AOI21X1  g14160(.A0(new_n16594_), .A1(new_n12779_), .B0(pi1155), .Y(new_n16597_));
  OAI21X1  g14161(.A0(new_n16597_), .A1(new_n16596_), .B0(pi0785), .Y(new_n16598_));
  OAI21X1  g14162(.A0(new_n16594_), .A1(pi0785), .B0(new_n16598_), .Y(new_n16599_));
  INVX1    g14163(.A(new_n16599_), .Y(new_n16600_));
  AOI21X1  g14164(.A0(new_n16600_), .A1(new_n12785_), .B0(new_n12615_), .Y(new_n16601_));
  AOI21X1  g14165(.A0(new_n16600_), .A1(new_n12788_), .B0(pi1154), .Y(new_n16602_));
  OR2X1    g14166(.A(new_n16602_), .B(new_n16601_), .Y(new_n16603_));
  MX2X1    g14167(.A(new_n16603_), .B(new_n16599_), .S0(new_n11887_), .Y(new_n16604_));
  AND2X1   g14168(.A(new_n16604_), .B(new_n11886_), .Y(new_n16605_));
  AOI21X1  g14169(.A0(new_n16591_), .A1(new_n12637_), .B0(new_n12638_), .Y(new_n16606_));
  OAI21X1  g14170(.A0(new_n16604_), .A1(new_n12637_), .B0(new_n16606_), .Y(new_n16607_));
  AOI21X1  g14171(.A0(new_n16591_), .A1(pi0619), .B0(pi1159), .Y(new_n16608_));
  OAI21X1  g14172(.A0(new_n16604_), .A1(pi0619), .B0(new_n16608_), .Y(new_n16609_));
  AOI21X1  g14173(.A0(new_n16609_), .A1(new_n16607_), .B0(new_n11886_), .Y(new_n16610_));
  NOR2X1   g14174(.A(new_n16610_), .B(new_n16605_), .Y(new_n16611_));
  INVX1    g14175(.A(new_n16611_), .Y(new_n16612_));
  MX2X1    g14176(.A(new_n16612_), .B(new_n16592_), .S0(new_n12841_), .Y(new_n16613_));
  MX2X1    g14177(.A(new_n16613_), .B(new_n16592_), .S0(new_n12711_), .Y(new_n16614_));
  INVX1    g14178(.A(pi0704), .Y(new_n16615_));
  AOI21X1  g14179(.A0(new_n12566_), .A1(new_n16615_), .B0(new_n16591_), .Y(new_n16616_));
  AND2X1   g14180(.A(new_n12566_), .B(new_n16615_), .Y(new_n16617_));
  AND2X1   g14181(.A(new_n16617_), .B(new_n12493_), .Y(new_n16618_));
  MX2X1    g14182(.A(new_n16591_), .B(pi0625), .S0(new_n16617_), .Y(new_n16619_));
  NOR2X1   g14183(.A(new_n16591_), .B(pi1153), .Y(new_n16620_));
  INVX1    g14184(.A(new_n16620_), .Y(new_n16621_));
  OAI22X1  g14185(.A0(new_n16621_), .A1(new_n16618_), .B0(new_n16619_), .B1(new_n12494_), .Y(new_n16622_));
  MX2X1    g14186(.A(new_n16622_), .B(new_n16616_), .S0(new_n11889_), .Y(new_n16623_));
  NOR4X1   g14187(.A(new_n16623_), .B(new_n12765_), .C(new_n12764_), .D(new_n12762_), .Y(new_n16624_));
  INVX1    g14188(.A(new_n16624_), .Y(new_n16625_));
  OR4X1    g14189(.A(new_n16625_), .B(new_n12870_), .C(new_n12851_), .D(pi0647), .Y(new_n16626_));
  NAND2X1  g14190(.A(new_n16591_), .B(pi0647), .Y(new_n16627_));
  NAND3X1  g14191(.A(new_n16627_), .B(new_n16626_), .C(new_n12706_), .Y(new_n16628_));
  INVX1    g14192(.A(new_n16628_), .Y(new_n16629_));
  NOR3X1   g14193(.A(new_n16625_), .B(new_n12870_), .C(new_n12851_), .Y(new_n16630_));
  MX2X1    g14194(.A(new_n16630_), .B(new_n16591_), .S0(new_n12705_), .Y(new_n16631_));
  INVX1    g14195(.A(new_n16631_), .Y(new_n16632_));
  AOI22X1  g14196(.A0(new_n16632_), .A1(new_n14386_), .B0(new_n16629_), .B1(pi0630), .Y(new_n16633_));
  INVX1    g14197(.A(new_n16633_), .Y(new_n16634_));
  AOI21X1  g14198(.A0(new_n16614_), .A1(new_n14385_), .B0(new_n16634_), .Y(new_n16635_));
  AOI21X1  g14199(.A0(new_n16592_), .A1(pi0626), .B0(new_n16352_), .Y(new_n16636_));
  OAI21X1  g14200(.A0(new_n16611_), .A1(pi0626), .B0(new_n16636_), .Y(new_n16637_));
  AOI21X1  g14201(.A0(new_n16592_), .A1(new_n12664_), .B0(new_n16356_), .Y(new_n16638_));
  OAI21X1  g14202(.A0(new_n16611_), .A1(new_n12664_), .B0(new_n16638_), .Y(new_n16639_));
  NAND2X1  g14203(.A(new_n16624_), .B(new_n12769_), .Y(new_n16640_));
  NAND3X1  g14204(.A(new_n16640_), .B(new_n16639_), .C(new_n16637_), .Y(new_n16641_));
  AND2X1   g14205(.A(new_n16641_), .B(pi0788), .Y(new_n16642_));
  INVX1    g14206(.A(new_n16642_), .Y(new_n16643_));
  NOR2X1   g14207(.A(new_n16616_), .B(new_n12120_), .Y(new_n16644_));
  MX2X1    g14208(.A(new_n16593_), .B(pi0625), .S0(new_n16644_), .Y(new_n16645_));
  OAI21X1  g14209(.A0(new_n16619_), .A1(new_n12494_), .B0(new_n12584_), .Y(new_n16646_));
  AOI21X1  g14210(.A0(new_n16645_), .A1(new_n16620_), .B0(new_n16646_), .Y(new_n16647_));
  AOI21X1  g14211(.A0(new_n16617_), .A1(new_n12493_), .B0(new_n16621_), .Y(new_n16648_));
  NOR3X1   g14212(.A(new_n16616_), .B(new_n12120_), .C(new_n12493_), .Y(new_n16649_));
  NOR3X1   g14213(.A(new_n16649_), .B(new_n16595_), .C(new_n12494_), .Y(new_n16650_));
  NOR3X1   g14214(.A(new_n16650_), .B(new_n16648_), .C(new_n12584_), .Y(new_n16651_));
  OAI21X1  g14215(.A0(new_n16651_), .A1(new_n16647_), .B0(pi0778), .Y(new_n16652_));
  OAI21X1  g14216(.A0(new_n16644_), .A1(new_n16595_), .B0(new_n11889_), .Y(new_n16653_));
  NAND2X1  g14217(.A(new_n16653_), .B(new_n16652_), .Y(new_n16654_));
  OAI21X1  g14218(.A0(new_n16623_), .A1(new_n12590_), .B0(new_n12591_), .Y(new_n16655_));
  AOI21X1  g14219(.A0(new_n16654_), .A1(new_n12590_), .B0(new_n16655_), .Y(new_n16656_));
  NOR3X1   g14220(.A(new_n16656_), .B(new_n16596_), .C(pi0660), .Y(new_n16657_));
  OAI21X1  g14221(.A0(new_n16623_), .A1(pi0609), .B0(pi1155), .Y(new_n16658_));
  AOI21X1  g14222(.A0(new_n16654_), .A1(pi0609), .B0(new_n16658_), .Y(new_n16659_));
  NOR3X1   g14223(.A(new_n16659_), .B(new_n16597_), .C(new_n12596_), .Y(new_n16660_));
  OAI21X1  g14224(.A0(new_n16660_), .A1(new_n16657_), .B0(pi0785), .Y(new_n16661_));
  NAND2X1  g14225(.A(new_n16654_), .B(new_n11888_), .Y(new_n16662_));
  AND2X1   g14226(.A(new_n16662_), .B(new_n16661_), .Y(new_n16663_));
  NOR3X1   g14227(.A(new_n16623_), .B(new_n12762_), .C(new_n12614_), .Y(new_n16664_));
  NOR2X1   g14228(.A(new_n16664_), .B(pi1154), .Y(new_n16665_));
  OAI21X1  g14229(.A0(new_n16663_), .A1(pi0618), .B0(new_n16665_), .Y(new_n16666_));
  NOR2X1   g14230(.A(new_n16601_), .B(pi0627), .Y(new_n16667_));
  NOR3X1   g14231(.A(new_n16623_), .B(new_n12762_), .C(pi0618), .Y(new_n16668_));
  NOR2X1   g14232(.A(new_n16668_), .B(new_n12615_), .Y(new_n16669_));
  OAI21X1  g14233(.A0(new_n16663_), .A1(new_n12614_), .B0(new_n16669_), .Y(new_n16670_));
  NOR2X1   g14234(.A(new_n16602_), .B(new_n12622_), .Y(new_n16671_));
  AOI22X1  g14235(.A0(new_n16671_), .A1(new_n16670_), .B0(new_n16667_), .B1(new_n16666_), .Y(new_n16672_));
  MX2X1    g14236(.A(new_n16672_), .B(new_n16663_), .S0(new_n11887_), .Y(new_n16673_));
  OR4X1    g14237(.A(new_n16623_), .B(new_n12764_), .C(new_n12762_), .D(new_n12637_), .Y(new_n16674_));
  AND2X1   g14238(.A(new_n16674_), .B(new_n12638_), .Y(new_n16675_));
  OAI21X1  g14239(.A0(new_n16673_), .A1(pi0619), .B0(new_n16675_), .Y(new_n16676_));
  AND2X1   g14240(.A(new_n16607_), .B(new_n12645_), .Y(new_n16677_));
  AND2X1   g14241(.A(new_n16677_), .B(new_n16676_), .Y(new_n16678_));
  NOR4X1   g14242(.A(new_n16623_), .B(new_n12764_), .C(new_n12762_), .D(pi0619), .Y(new_n16679_));
  NOR2X1   g14243(.A(new_n16679_), .B(new_n12638_), .Y(new_n16680_));
  OAI21X1  g14244(.A0(new_n16673_), .A1(new_n12637_), .B0(new_n16680_), .Y(new_n16681_));
  AND2X1   g14245(.A(new_n16609_), .B(pi0648), .Y(new_n16682_));
  AOI21X1  g14246(.A0(new_n16682_), .A1(new_n16681_), .B0(new_n11886_), .Y(new_n16683_));
  INVX1    g14247(.A(new_n16683_), .Y(new_n16684_));
  AOI21X1  g14248(.A0(new_n16673_), .A1(new_n11886_), .B0(new_n14264_), .Y(new_n16685_));
  OAI21X1  g14249(.A0(new_n16684_), .A1(new_n16678_), .B0(new_n16685_), .Y(new_n16686_));
  AOI21X1  g14250(.A0(new_n16686_), .A1(new_n16643_), .B0(new_n14273_), .Y(new_n16687_));
  INVX1    g14251(.A(new_n16613_), .Y(new_n16688_));
  AND2X1   g14252(.A(new_n16624_), .B(new_n12852_), .Y(new_n16689_));
  AOI22X1  g14253(.A0(new_n16689_), .A1(new_n14564_), .B0(new_n16688_), .B1(new_n12867_), .Y(new_n16690_));
  AOI22X1  g14254(.A0(new_n16689_), .A1(new_n14566_), .B0(new_n16688_), .B1(new_n12865_), .Y(new_n16691_));
  MX2X1    g14255(.A(new_n16691_), .B(new_n16690_), .S0(new_n12689_), .Y(new_n16692_));
  OAI21X1  g14256(.A0(new_n16692_), .A1(new_n11884_), .B0(new_n14562_), .Y(new_n16693_));
  OAI22X1  g14257(.A0(new_n16693_), .A1(new_n16687_), .B0(new_n16635_), .B1(new_n11883_), .Y(new_n16694_));
  AOI21X1  g14258(.A0(new_n16632_), .A1(pi1157), .B0(new_n16629_), .Y(new_n16695_));
  MX2X1    g14259(.A(new_n16695_), .B(new_n16630_), .S0(new_n11883_), .Y(new_n16696_));
  AOI21X1  g14260(.A0(new_n16696_), .A1(new_n12743_), .B0(new_n12739_), .Y(new_n16697_));
  OAI21X1  g14261(.A0(new_n16694_), .A1(new_n12743_), .B0(new_n16697_), .Y(new_n16698_));
  MX2X1    g14262(.A(new_n16614_), .B(new_n16592_), .S0(new_n12735_), .Y(new_n16699_));
  AOI21X1  g14263(.A0(new_n16591_), .A1(new_n12743_), .B0(pi0715), .Y(new_n16700_));
  OAI21X1  g14264(.A0(new_n16699_), .A1(new_n12743_), .B0(new_n16700_), .Y(new_n16701_));
  AND2X1   g14265(.A(new_n16701_), .B(pi1160), .Y(new_n16702_));
  AOI21X1  g14266(.A0(new_n16696_), .A1(pi0644), .B0(pi0715), .Y(new_n16703_));
  OAI21X1  g14267(.A0(new_n16694_), .A1(pi0644), .B0(new_n16703_), .Y(new_n16704_));
  AOI21X1  g14268(.A0(new_n16591_), .A1(pi0644), .B0(new_n12739_), .Y(new_n16705_));
  OAI21X1  g14269(.A0(new_n16699_), .A1(pi0644), .B0(new_n16705_), .Y(new_n16706_));
  AND2X1   g14270(.A(new_n16706_), .B(new_n11882_), .Y(new_n16707_));
  AOI22X1  g14271(.A0(new_n16707_), .A1(new_n16704_), .B0(new_n16702_), .B1(new_n16698_), .Y(new_n16708_));
  OR2X1    g14272(.A(new_n16694_), .B(pi0790), .Y(new_n16709_));
  AND2X1   g14273(.A(new_n16709_), .B(pi0832), .Y(new_n16710_));
  OAI21X1  g14274(.A0(new_n16708_), .A1(new_n12897_), .B0(new_n16710_), .Y(new_n16711_));
  AOI21X1  g14275(.A0(new_n13699_), .A1(new_n3129_), .B0(pi0176), .Y(new_n16712_));
  INVX1    g14276(.A(new_n16712_), .Y(new_n16713_));
  AND2X1   g14277(.A(new_n16436_), .B(new_n2996_), .Y(new_n16714_));
  OR4X1    g14278(.A(new_n16714_), .B(new_n12567_), .C(new_n3125_), .D(new_n3124_), .Y(new_n16715_));
  OAI21X1  g14279(.A0(new_n12953_), .A1(pi0038), .B0(new_n14017_), .Y(new_n16716_));
  OR2X1    g14280(.A(new_n16716_), .B(pi0176), .Y(new_n16717_));
  AND2X1   g14281(.A(new_n16717_), .B(new_n16615_), .Y(new_n16718_));
  INVX1    g14282(.A(new_n16718_), .Y(new_n16719_));
  AND2X1   g14283(.A(new_n12574_), .B(new_n6866_), .Y(new_n16720_));
  AOI21X1  g14284(.A0(new_n16720_), .A1(pi0704), .B0(new_n3810_), .Y(new_n16721_));
  AOI22X1  g14285(.A0(new_n16721_), .A1(new_n16719_), .B0(new_n16715_), .B1(pi0176), .Y(new_n16722_));
  OAI21X1  g14286(.A0(new_n16713_), .A1(pi0625), .B0(pi1153), .Y(new_n16723_));
  AOI21X1  g14287(.A0(new_n16722_), .A1(pi0625), .B0(new_n16723_), .Y(new_n16724_));
  OAI21X1  g14288(.A0(new_n16713_), .A1(new_n12493_), .B0(new_n12494_), .Y(new_n16725_));
  AOI21X1  g14289(.A0(new_n16722_), .A1(new_n12493_), .B0(new_n16725_), .Y(new_n16726_));
  NOR2X1   g14290(.A(new_n16726_), .B(new_n16724_), .Y(new_n16727_));
  MX2X1    g14291(.A(new_n16727_), .B(new_n16722_), .S0(new_n11889_), .Y(new_n16728_));
  MX2X1    g14292(.A(new_n16728_), .B(new_n16712_), .S0(new_n12618_), .Y(new_n16729_));
  AND2X1   g14293(.A(new_n16712_), .B(new_n12641_), .Y(new_n16730_));
  AOI21X1  g14294(.A0(new_n16729_), .A1(new_n14198_), .B0(new_n16730_), .Y(new_n16731_));
  MX2X1    g14295(.A(new_n16731_), .B(new_n16713_), .S0(new_n12659_), .Y(new_n16732_));
  MX2X1    g14296(.A(new_n16732_), .B(new_n16713_), .S0(new_n12691_), .Y(new_n16733_));
  MX2X1    g14297(.A(new_n16733_), .B(new_n16713_), .S0(pi0628), .Y(new_n16734_));
  MX2X1    g14298(.A(new_n16733_), .B(new_n16713_), .S0(new_n12683_), .Y(new_n16735_));
  MX2X1    g14299(.A(new_n16735_), .B(new_n16734_), .S0(new_n12684_), .Y(new_n16736_));
  MX2X1    g14300(.A(new_n16736_), .B(new_n16733_), .S0(new_n11884_), .Y(new_n16737_));
  MX2X1    g14301(.A(new_n16737_), .B(new_n16713_), .S0(pi0647), .Y(new_n16738_));
  MX2X1    g14302(.A(new_n16737_), .B(new_n16713_), .S0(new_n12705_), .Y(new_n16739_));
  MX2X1    g14303(.A(new_n16739_), .B(new_n16738_), .S0(new_n12706_), .Y(new_n16740_));
  OR2X1    g14304(.A(new_n16737_), .B(pi0787), .Y(new_n16741_));
  OAI21X1  g14305(.A0(new_n16740_), .A1(new_n11883_), .B0(new_n16741_), .Y(new_n16742_));
  AOI21X1  g14306(.A0(new_n16742_), .A1(new_n12743_), .B0(new_n12739_), .Y(new_n16743_));
  INVX1    g14307(.A(new_n13704_), .Y(new_n16744_));
  INVX1    g14308(.A(new_n13701_), .Y(new_n16745_));
  OAI21X1  g14309(.A0(new_n13977_), .A1(pi0038), .B0(new_n16745_), .Y(new_n16746_));
  MX2X1    g14310(.A(new_n16746_), .B(new_n16744_), .S0(new_n6866_), .Y(new_n16747_));
  MX2X1    g14311(.A(new_n16747_), .B(new_n16720_), .S0(pi0742), .Y(new_n16748_));
  MX2X1    g14312(.A(new_n16748_), .B(new_n6866_), .S0(new_n3810_), .Y(new_n16749_));
  MX2X1    g14313(.A(new_n16749_), .B(new_n16712_), .S0(new_n12601_), .Y(new_n16750_));
  NOR2X1   g14314(.A(new_n16749_), .B(new_n12601_), .Y(new_n16751_));
  AOI22X1  g14315(.A0(new_n16751_), .A1(pi0609), .B0(new_n16713_), .B1(new_n13430_), .Y(new_n16752_));
  AOI22X1  g14316(.A0(new_n16751_), .A1(new_n12590_), .B0(new_n16713_), .B1(new_n13436_), .Y(new_n16753_));
  MX2X1    g14317(.A(new_n16753_), .B(new_n16752_), .S0(pi1155), .Y(new_n16754_));
  MX2X1    g14318(.A(new_n16754_), .B(new_n16750_), .S0(new_n11888_), .Y(new_n16755_));
  OAI21X1  g14319(.A0(new_n16713_), .A1(pi0618), .B0(pi1154), .Y(new_n16756_));
  AOI21X1  g14320(.A0(new_n16755_), .A1(pi0618), .B0(new_n16756_), .Y(new_n16757_));
  OAI21X1  g14321(.A0(new_n16713_), .A1(new_n12614_), .B0(new_n12615_), .Y(new_n16758_));
  AOI21X1  g14322(.A0(new_n16755_), .A1(new_n12614_), .B0(new_n16758_), .Y(new_n16759_));
  NOR2X1   g14323(.A(new_n16759_), .B(new_n16757_), .Y(new_n16760_));
  MX2X1    g14324(.A(new_n16760_), .B(new_n16755_), .S0(new_n11887_), .Y(new_n16761_));
  OR2X1    g14325(.A(new_n16761_), .B(pi0789), .Y(new_n16762_));
  OAI21X1  g14326(.A0(new_n16713_), .A1(pi0619), .B0(pi1159), .Y(new_n16763_));
  AOI21X1  g14327(.A0(new_n16761_), .A1(pi0619), .B0(new_n16763_), .Y(new_n16764_));
  OAI21X1  g14328(.A0(new_n16713_), .A1(new_n12637_), .B0(new_n12638_), .Y(new_n16765_));
  AOI21X1  g14329(.A0(new_n16761_), .A1(new_n12637_), .B0(new_n16765_), .Y(new_n16766_));
  OAI21X1  g14330(.A0(new_n16766_), .A1(new_n16764_), .B0(pi0789), .Y(new_n16767_));
  AND2X1   g14331(.A(new_n16767_), .B(new_n16762_), .Y(new_n16768_));
  INVX1    g14332(.A(new_n16768_), .Y(new_n16769_));
  MX2X1    g14333(.A(new_n16769_), .B(new_n16713_), .S0(new_n12841_), .Y(new_n16770_));
  MX2X1    g14334(.A(new_n16770_), .B(new_n16713_), .S0(new_n12711_), .Y(new_n16771_));
  MX2X1    g14335(.A(new_n16771_), .B(new_n16713_), .S0(new_n12735_), .Y(new_n16772_));
  AOI21X1  g14336(.A0(new_n16712_), .A1(new_n12743_), .B0(pi0715), .Y(new_n16773_));
  OAI21X1  g14337(.A0(new_n16772_), .A1(new_n12743_), .B0(new_n16773_), .Y(new_n16774_));
  AND2X1   g14338(.A(new_n16774_), .B(pi1160), .Y(new_n16775_));
  INVX1    g14339(.A(new_n16775_), .Y(new_n16776_));
  AOI21X1  g14340(.A0(new_n16742_), .A1(pi0644), .B0(pi0715), .Y(new_n16777_));
  AOI21X1  g14341(.A0(new_n16712_), .A1(pi0644), .B0(new_n12739_), .Y(new_n16778_));
  OAI21X1  g14342(.A0(new_n16772_), .A1(pi0644), .B0(new_n16778_), .Y(new_n16779_));
  NAND2X1  g14343(.A(new_n16779_), .B(new_n11882_), .Y(new_n16780_));
  OAI22X1  g14344(.A0(new_n16780_), .A1(new_n16777_), .B0(new_n16776_), .B1(new_n16743_), .Y(new_n16781_));
  NAND2X1  g14345(.A(new_n16770_), .B(new_n14394_), .Y(new_n16782_));
  AOI22X1  g14346(.A0(new_n16735_), .A1(new_n12707_), .B0(new_n16734_), .B1(new_n12709_), .Y(new_n16783_));
  NAND2X1  g14347(.A(new_n16783_), .B(new_n16782_), .Y(new_n16784_));
  OAI21X1  g14348(.A0(new_n16712_), .A1(new_n12664_), .B0(new_n16351_), .Y(new_n16785_));
  AOI21X1  g14349(.A0(new_n16769_), .A1(new_n12664_), .B0(new_n16785_), .Y(new_n16786_));
  AOI21X1  g14350(.A0(new_n16767_), .A1(new_n16762_), .B0(new_n12664_), .Y(new_n16787_));
  OAI21X1  g14351(.A0(new_n16712_), .A1(pi0626), .B0(new_n16355_), .Y(new_n16788_));
  OAI22X1  g14352(.A0(new_n16788_), .A1(new_n16787_), .B0(new_n16732_), .B1(new_n12770_), .Y(new_n16789_));
  OAI21X1  g14353(.A0(new_n16789_), .A1(new_n16786_), .B0(pi0788), .Y(new_n16790_));
  NAND2X1  g14354(.A(new_n13672_), .B(new_n6866_), .Y(new_n16791_));
  NOR2X1   g14355(.A(new_n13673_), .B(pi0038), .Y(new_n16792_));
  OR2X1    g14356(.A(new_n13676_), .B(new_n16792_), .Y(new_n16793_));
  AOI21X1  g14357(.A0(new_n16793_), .A1(pi0176), .B0(new_n15046_), .Y(new_n16794_));
  NAND2X1  g14358(.A(new_n16794_), .B(new_n16791_), .Y(new_n16795_));
  MX2X1    g14359(.A(new_n13687_), .B(new_n13681_), .S0(pi0038), .Y(new_n16796_));
  OAI21X1  g14360(.A0(new_n13693_), .A1(new_n13690_), .B0(new_n6866_), .Y(new_n16797_));
  AND2X1   g14361(.A(new_n16797_), .B(new_n15046_), .Y(new_n16798_));
  OAI21X1  g14362(.A0(new_n16796_), .A1(new_n6866_), .B0(new_n16798_), .Y(new_n16799_));
  NAND3X1  g14363(.A(new_n16799_), .B(new_n16795_), .C(new_n16615_), .Y(new_n16800_));
  AOI21X1  g14364(.A0(new_n16748_), .A1(pi0704), .B0(new_n3810_), .Y(new_n16801_));
  AOI22X1  g14365(.A0(new_n16801_), .A1(new_n16800_), .B0(new_n3810_), .B1(pi0176), .Y(new_n16802_));
  INVX1    g14366(.A(new_n16802_), .Y(new_n16803_));
  AOI21X1  g14367(.A0(new_n16749_), .A1(pi0625), .B0(pi1153), .Y(new_n16804_));
  OAI21X1  g14368(.A0(new_n16803_), .A1(pi0625), .B0(new_n16804_), .Y(new_n16805_));
  NOR2X1   g14369(.A(new_n16724_), .B(pi0608), .Y(new_n16806_));
  AOI21X1  g14370(.A0(new_n16749_), .A1(new_n12493_), .B0(new_n12494_), .Y(new_n16807_));
  OAI21X1  g14371(.A0(new_n16803_), .A1(new_n12493_), .B0(new_n16807_), .Y(new_n16808_));
  NOR2X1   g14372(.A(new_n16726_), .B(new_n12584_), .Y(new_n16809_));
  AOI22X1  g14373(.A0(new_n16809_), .A1(new_n16808_), .B0(new_n16806_), .B1(new_n16805_), .Y(new_n16810_));
  MX2X1    g14374(.A(new_n16810_), .B(new_n16803_), .S0(new_n11889_), .Y(new_n16811_));
  AOI21X1  g14375(.A0(new_n16728_), .A1(pi0609), .B0(pi1155), .Y(new_n16812_));
  OAI21X1  g14376(.A0(new_n16811_), .A1(pi0609), .B0(new_n16812_), .Y(new_n16813_));
  OAI21X1  g14377(.A0(new_n16752_), .A1(new_n12591_), .B0(new_n12596_), .Y(new_n16814_));
  INVX1    g14378(.A(new_n16814_), .Y(new_n16815_));
  AOI21X1  g14379(.A0(new_n16728_), .A1(new_n12590_), .B0(new_n12591_), .Y(new_n16816_));
  OAI21X1  g14380(.A0(new_n16811_), .A1(new_n12590_), .B0(new_n16816_), .Y(new_n16817_));
  OAI21X1  g14381(.A0(new_n16753_), .A1(pi1155), .B0(pi0660), .Y(new_n16818_));
  INVX1    g14382(.A(new_n16818_), .Y(new_n16819_));
  AOI22X1  g14383(.A0(new_n16819_), .A1(new_n16817_), .B0(new_n16815_), .B1(new_n16813_), .Y(new_n16820_));
  MX2X1    g14384(.A(new_n16820_), .B(new_n16811_), .S0(new_n11888_), .Y(new_n16821_));
  AOI21X1  g14385(.A0(new_n16729_), .A1(pi0618), .B0(pi1154), .Y(new_n16822_));
  OAI21X1  g14386(.A0(new_n16821_), .A1(pi0618), .B0(new_n16822_), .Y(new_n16823_));
  NOR2X1   g14387(.A(new_n16757_), .B(pi0627), .Y(new_n16824_));
  AOI21X1  g14388(.A0(new_n16729_), .A1(new_n12614_), .B0(new_n12615_), .Y(new_n16825_));
  OAI21X1  g14389(.A0(new_n16821_), .A1(new_n12614_), .B0(new_n16825_), .Y(new_n16826_));
  NOR2X1   g14390(.A(new_n16759_), .B(new_n12622_), .Y(new_n16827_));
  AOI22X1  g14391(.A0(new_n16827_), .A1(new_n16826_), .B0(new_n16824_), .B1(new_n16823_), .Y(new_n16828_));
  MX2X1    g14392(.A(new_n16828_), .B(new_n16821_), .S0(new_n11887_), .Y(new_n16829_));
  INVX1    g14393(.A(new_n16829_), .Y(new_n16830_));
  OAI21X1  g14394(.A0(new_n16731_), .A1(new_n12637_), .B0(new_n12638_), .Y(new_n16831_));
  AOI21X1  g14395(.A0(new_n16830_), .A1(new_n12637_), .B0(new_n16831_), .Y(new_n16832_));
  NOR3X1   g14396(.A(new_n16832_), .B(new_n16764_), .C(pi0648), .Y(new_n16833_));
  OAI21X1  g14397(.A0(new_n16731_), .A1(pi0619), .B0(pi1159), .Y(new_n16834_));
  AOI21X1  g14398(.A0(new_n16830_), .A1(pi0619), .B0(new_n16834_), .Y(new_n16835_));
  OR2X1    g14399(.A(new_n16766_), .B(new_n12645_), .Y(new_n16836_));
  OAI21X1  g14400(.A0(new_n16836_), .A1(new_n16835_), .B0(pi0789), .Y(new_n16837_));
  AOI21X1  g14401(.A0(new_n16829_), .A1(new_n11886_), .B0(new_n14264_), .Y(new_n16838_));
  OAI21X1  g14402(.A0(new_n16837_), .A1(new_n16833_), .B0(new_n16838_), .Y(new_n16839_));
  AOI22X1  g14403(.A0(new_n16839_), .A1(new_n16790_), .B0(new_n16784_), .B1(pi0792), .Y(new_n16840_));
  OAI21X1  g14404(.A0(new_n16784_), .A1(new_n16350_), .B0(new_n14562_), .Y(new_n16841_));
  OR2X1    g14405(.A(new_n16841_), .B(new_n16840_), .Y(new_n16842_));
  NAND3X1  g14406(.A(new_n16779_), .B(new_n11882_), .C(new_n12743_), .Y(new_n16843_));
  AOI21X1  g14407(.A0(new_n16775_), .A1(pi0644), .B0(new_n12897_), .Y(new_n16844_));
  NAND2X1  g14408(.A(new_n16771_), .B(new_n14385_), .Y(new_n16845_));
  AOI22X1  g14409(.A0(new_n16739_), .A1(new_n14386_), .B0(new_n16738_), .B1(new_n14388_), .Y(new_n16846_));
  AOI21X1  g14410(.A0(new_n16846_), .A1(new_n16845_), .B0(new_n11883_), .Y(new_n16847_));
  AOI21X1  g14411(.A0(new_n16844_), .A1(new_n16843_), .B0(new_n16847_), .Y(new_n16848_));
  AOI22X1  g14412(.A0(new_n16848_), .A1(new_n16842_), .B0(new_n16781_), .B1(pi0790), .Y(new_n16849_));
  AOI21X1  g14413(.A0(po1038), .A1(new_n6866_), .B0(pi0832), .Y(new_n16850_));
  OAI21X1  g14414(.A0(new_n16849_), .A1(po1038), .B0(new_n16850_), .Y(new_n16851_));
  AND2X1   g14415(.A(new_n16851_), .B(new_n16711_), .Y(po0333));
  NOR2X1   g14416(.A(new_n3129_), .B(new_n7469_), .Y(new_n16853_));
  INVX1    g14417(.A(new_n16853_), .Y(new_n16854_));
  INVX1    g14418(.A(pi0686), .Y(new_n16855_));
  MX2X1    g14419(.A(new_n16744_), .B(new_n12574_), .S0(pi0757), .Y(new_n16856_));
  AOI21X1  g14420(.A0(new_n16745_), .A1(new_n7469_), .B0(pi0757), .Y(new_n16857_));
  AOI22X1  g14421(.A0(new_n16857_), .A1(new_n16746_), .B0(new_n16856_), .B1(new_n7469_), .Y(new_n16858_));
  OAI21X1  g14422(.A0(new_n13673_), .A1(new_n7469_), .B0(new_n2996_), .Y(new_n16859_));
  AOI21X1  g14423(.A0(new_n13671_), .A1(new_n7469_), .B0(new_n16859_), .Y(new_n16860_));
  OAI21X1  g14424(.A0(new_n12202_), .A1(pi0177), .B0(new_n12935_), .Y(new_n16861_));
  NAND2X1  g14425(.A(new_n16861_), .B(pi0757), .Y(new_n16862_));
  NOR2X1   g14426(.A(new_n13687_), .B(new_n7469_), .Y(new_n16863_));
  NOR2X1   g14427(.A(new_n13691_), .B(new_n13690_), .Y(new_n16864_));
  OAI21X1  g14428(.A0(new_n16864_), .A1(pi0177), .B0(new_n2996_), .Y(new_n16865_));
  NOR2X1   g14429(.A(new_n16865_), .B(new_n16863_), .Y(new_n16866_));
  OAI21X1  g14430(.A0(new_n13681_), .A1(new_n7469_), .B0(pi0038), .Y(new_n16867_));
  AOI21X1  g14431(.A0(new_n13692_), .A1(new_n7469_), .B0(new_n16867_), .Y(new_n16868_));
  OR2X1    g14432(.A(new_n16868_), .B(pi0757), .Y(new_n16869_));
  OAI22X1  g14433(.A0(new_n16869_), .A1(new_n16866_), .B0(new_n16862_), .B1(new_n16860_), .Y(new_n16870_));
  AOI21X1  g14434(.A0(new_n16870_), .A1(new_n16855_), .B0(new_n3810_), .Y(new_n16871_));
  OAI21X1  g14435(.A0(new_n16858_), .A1(new_n16855_), .B0(new_n16871_), .Y(new_n16872_));
  NAND3X1  g14436(.A(new_n16872_), .B(new_n16854_), .C(new_n12493_), .Y(new_n16873_));
  AOI21X1  g14437(.A0(new_n16858_), .A1(new_n3129_), .B0(new_n16853_), .Y(new_n16874_));
  AOI21X1  g14438(.A0(new_n16874_), .A1(pi0625), .B0(pi1153), .Y(new_n16875_));
  AOI21X1  g14439(.A0(new_n12955_), .A1(pi0177), .B0(pi0038), .Y(new_n16876_));
  OAI21X1  g14440(.A0(new_n12953_), .A1(pi0177), .B0(new_n16876_), .Y(new_n16877_));
  OAI21X1  g14441(.A0(new_n12202_), .A1(pi0177), .B0(new_n12567_), .Y(new_n16878_));
  NAND3X1  g14442(.A(new_n16878_), .B(new_n16877_), .C(new_n16855_), .Y(new_n16879_));
  AND2X1   g14443(.A(pi0686), .B(new_n7469_), .Y(new_n16880_));
  AOI21X1  g14444(.A0(new_n16880_), .A1(new_n12574_), .B0(new_n3810_), .Y(new_n16881_));
  AOI21X1  g14445(.A0(new_n16881_), .A1(new_n16879_), .B0(new_n16853_), .Y(new_n16882_));
  OAI21X1  g14446(.A0(new_n12574_), .A1(new_n3810_), .B0(new_n7469_), .Y(new_n16883_));
  OAI21X1  g14447(.A0(new_n16883_), .A1(pi0625), .B0(pi1153), .Y(new_n16884_));
  AOI21X1  g14448(.A0(new_n16882_), .A1(pi0625), .B0(new_n16884_), .Y(new_n16885_));
  OR2X1    g14449(.A(new_n16885_), .B(pi0608), .Y(new_n16886_));
  AOI21X1  g14450(.A0(new_n16875_), .A1(new_n16873_), .B0(new_n16886_), .Y(new_n16887_));
  NAND3X1  g14451(.A(new_n16872_), .B(new_n16854_), .C(pi0625), .Y(new_n16888_));
  AOI21X1  g14452(.A0(new_n16874_), .A1(new_n12493_), .B0(new_n12494_), .Y(new_n16889_));
  OAI21X1  g14453(.A0(new_n16883_), .A1(new_n12493_), .B0(new_n12494_), .Y(new_n16890_));
  AOI21X1  g14454(.A0(new_n16882_), .A1(new_n12493_), .B0(new_n16890_), .Y(new_n16891_));
  OR2X1    g14455(.A(new_n16891_), .B(new_n12584_), .Y(new_n16892_));
  AOI21X1  g14456(.A0(new_n16889_), .A1(new_n16888_), .B0(new_n16892_), .Y(new_n16893_));
  OAI21X1  g14457(.A0(new_n16893_), .A1(new_n16887_), .B0(pi0778), .Y(new_n16894_));
  NAND3X1  g14458(.A(new_n16872_), .B(new_n16854_), .C(new_n11889_), .Y(new_n16895_));
  NAND2X1  g14459(.A(new_n16895_), .B(new_n16894_), .Y(new_n16896_));
  OAI21X1  g14460(.A0(new_n16891_), .A1(new_n16885_), .B0(pi0778), .Y(new_n16897_));
  OAI21X1  g14461(.A0(new_n16882_), .A1(pi0778), .B0(new_n16897_), .Y(new_n16898_));
  OAI21X1  g14462(.A0(new_n16898_), .A1(new_n12590_), .B0(new_n12591_), .Y(new_n16899_));
  AOI21X1  g14463(.A0(new_n16896_), .A1(new_n12590_), .B0(new_n16899_), .Y(new_n16900_));
  NOR2X1   g14464(.A(new_n16874_), .B(new_n12601_), .Y(new_n16901_));
  AOI22X1  g14465(.A0(new_n16901_), .A1(pi0609), .B0(new_n16883_), .B1(new_n13430_), .Y(new_n16902_));
  OAI21X1  g14466(.A0(new_n16902_), .A1(new_n12591_), .B0(new_n12596_), .Y(new_n16903_));
  OAI21X1  g14467(.A0(new_n16898_), .A1(pi0609), .B0(pi1155), .Y(new_n16904_));
  AOI21X1  g14468(.A0(new_n16896_), .A1(pi0609), .B0(new_n16904_), .Y(new_n16905_));
  AOI22X1  g14469(.A0(new_n16901_), .A1(new_n12590_), .B0(new_n16883_), .B1(new_n13436_), .Y(new_n16906_));
  OAI21X1  g14470(.A0(new_n16906_), .A1(pi1155), .B0(pi0660), .Y(new_n16907_));
  OAI22X1  g14471(.A0(new_n16907_), .A1(new_n16905_), .B0(new_n16903_), .B1(new_n16900_), .Y(new_n16908_));
  MX2X1    g14472(.A(new_n16908_), .B(new_n16896_), .S0(new_n11888_), .Y(new_n16909_));
  MX2X1    g14473(.A(new_n16898_), .B(new_n16883_), .S0(new_n12618_), .Y(new_n16910_));
  OAI21X1  g14474(.A0(new_n16910_), .A1(new_n12614_), .B0(new_n12615_), .Y(new_n16911_));
  AOI21X1  g14475(.A0(new_n16909_), .A1(new_n12614_), .B0(new_n16911_), .Y(new_n16912_));
  INVX1    g14476(.A(new_n16883_), .Y(new_n16913_));
  MX2X1    g14477(.A(new_n16913_), .B(new_n16874_), .S0(new_n12623_), .Y(new_n16914_));
  MX2X1    g14478(.A(new_n16906_), .B(new_n16902_), .S0(pi1155), .Y(new_n16915_));
  MX2X1    g14479(.A(new_n16915_), .B(new_n16914_), .S0(new_n11888_), .Y(new_n16916_));
  OAI21X1  g14480(.A0(new_n16883_), .A1(pi0618), .B0(pi1154), .Y(new_n16917_));
  AOI21X1  g14481(.A0(new_n16916_), .A1(pi0618), .B0(new_n16917_), .Y(new_n16918_));
  OR2X1    g14482(.A(new_n16918_), .B(pi0627), .Y(new_n16919_));
  OAI21X1  g14483(.A0(new_n16910_), .A1(pi0618), .B0(pi1154), .Y(new_n16920_));
  AOI21X1  g14484(.A0(new_n16909_), .A1(pi0618), .B0(new_n16920_), .Y(new_n16921_));
  OAI21X1  g14485(.A0(new_n16883_), .A1(new_n12614_), .B0(new_n12615_), .Y(new_n16922_));
  AOI21X1  g14486(.A0(new_n16916_), .A1(new_n12614_), .B0(new_n16922_), .Y(new_n16923_));
  OR2X1    g14487(.A(new_n16923_), .B(new_n12622_), .Y(new_n16924_));
  OAI22X1  g14488(.A0(new_n16924_), .A1(new_n16921_), .B0(new_n16919_), .B1(new_n16912_), .Y(new_n16925_));
  MX2X1    g14489(.A(new_n16925_), .B(new_n16909_), .S0(new_n11887_), .Y(new_n16926_));
  MX2X1    g14490(.A(new_n16910_), .B(new_n16883_), .S0(new_n12641_), .Y(new_n16927_));
  OAI21X1  g14491(.A0(new_n16927_), .A1(new_n12637_), .B0(new_n12638_), .Y(new_n16928_));
  AOI21X1  g14492(.A0(new_n16926_), .A1(new_n12637_), .B0(new_n16928_), .Y(new_n16929_));
  OR2X1    g14493(.A(new_n16916_), .B(pi0781), .Y(new_n16930_));
  OAI21X1  g14494(.A0(new_n16923_), .A1(new_n16918_), .B0(pi0781), .Y(new_n16931_));
  NAND2X1  g14495(.A(new_n16931_), .B(new_n16930_), .Y(new_n16932_));
  AOI21X1  g14496(.A0(new_n16913_), .A1(new_n12637_), .B0(new_n12638_), .Y(new_n16933_));
  OAI21X1  g14497(.A0(new_n16932_), .A1(new_n12637_), .B0(new_n16933_), .Y(new_n16934_));
  NAND2X1  g14498(.A(new_n16934_), .B(new_n12645_), .Y(new_n16935_));
  OAI21X1  g14499(.A0(new_n16927_), .A1(pi0619), .B0(pi1159), .Y(new_n16936_));
  AOI21X1  g14500(.A0(new_n16926_), .A1(pi0619), .B0(new_n16936_), .Y(new_n16937_));
  AOI21X1  g14501(.A0(new_n16913_), .A1(pi0619), .B0(pi1159), .Y(new_n16938_));
  OAI21X1  g14502(.A0(new_n16932_), .A1(pi0619), .B0(new_n16938_), .Y(new_n16939_));
  NAND2X1  g14503(.A(new_n16939_), .B(pi0648), .Y(new_n16940_));
  OAI22X1  g14504(.A0(new_n16940_), .A1(new_n16937_), .B0(new_n16935_), .B1(new_n16929_), .Y(new_n16941_));
  MX2X1    g14505(.A(new_n16941_), .B(new_n16926_), .S0(new_n11886_), .Y(new_n16942_));
  MX2X1    g14506(.A(new_n16927_), .B(new_n16883_), .S0(new_n12659_), .Y(new_n16943_));
  AOI21X1  g14507(.A0(new_n16943_), .A1(pi0626), .B0(pi0641), .Y(new_n16944_));
  OAI21X1  g14508(.A0(new_n16942_), .A1(pi0626), .B0(new_n16944_), .Y(new_n16945_));
  NAND2X1  g14509(.A(new_n16939_), .B(new_n16934_), .Y(new_n16946_));
  MX2X1    g14510(.A(new_n16946_), .B(new_n16932_), .S0(new_n11886_), .Y(new_n16947_));
  OAI21X1  g14511(.A0(new_n16913_), .A1(new_n12664_), .B0(pi0641), .Y(new_n16948_));
  AOI21X1  g14512(.A0(new_n16947_), .A1(new_n12664_), .B0(new_n16948_), .Y(new_n16949_));
  NOR2X1   g14513(.A(new_n16949_), .B(pi1158), .Y(new_n16950_));
  AOI21X1  g14514(.A0(new_n16943_), .A1(new_n12664_), .B0(new_n12672_), .Y(new_n16951_));
  OAI21X1  g14515(.A0(new_n16942_), .A1(new_n12664_), .B0(new_n16951_), .Y(new_n16952_));
  OAI21X1  g14516(.A0(new_n16913_), .A1(pi0626), .B0(new_n12672_), .Y(new_n16953_));
  AOI21X1  g14517(.A0(new_n16947_), .A1(pi0626), .B0(new_n16953_), .Y(new_n16954_));
  NOR2X1   g14518(.A(new_n16954_), .B(new_n12676_), .Y(new_n16955_));
  AOI22X1  g14519(.A0(new_n16955_), .A1(new_n16952_), .B0(new_n16950_), .B1(new_n16945_), .Y(new_n16956_));
  MX2X1    g14520(.A(new_n16956_), .B(new_n16942_), .S0(new_n11885_), .Y(new_n16957_));
  MX2X1    g14521(.A(new_n16947_), .B(new_n16883_), .S0(new_n12841_), .Y(new_n16958_));
  OAI21X1  g14522(.A0(new_n16958_), .A1(new_n12683_), .B0(new_n12684_), .Y(new_n16959_));
  AOI21X1  g14523(.A0(new_n16957_), .A1(new_n12683_), .B0(new_n16959_), .Y(new_n16960_));
  MX2X1    g14524(.A(new_n16943_), .B(new_n16883_), .S0(new_n12691_), .Y(new_n16961_));
  AOI21X1  g14525(.A0(new_n16913_), .A1(new_n12683_), .B0(new_n12684_), .Y(new_n16962_));
  OAI21X1  g14526(.A0(new_n16961_), .A1(new_n12683_), .B0(new_n16962_), .Y(new_n16963_));
  NAND2X1  g14527(.A(new_n16963_), .B(new_n12689_), .Y(new_n16964_));
  OAI21X1  g14528(.A0(new_n16958_), .A1(pi0628), .B0(pi1156), .Y(new_n16965_));
  AOI21X1  g14529(.A0(new_n16957_), .A1(pi0628), .B0(new_n16965_), .Y(new_n16966_));
  AOI21X1  g14530(.A0(new_n16913_), .A1(pi0628), .B0(pi1156), .Y(new_n16967_));
  OAI21X1  g14531(.A0(new_n16961_), .A1(pi0628), .B0(new_n16967_), .Y(new_n16968_));
  NAND2X1  g14532(.A(new_n16968_), .B(pi0629), .Y(new_n16969_));
  OAI22X1  g14533(.A0(new_n16969_), .A1(new_n16966_), .B0(new_n16964_), .B1(new_n16960_), .Y(new_n16970_));
  AND2X1   g14534(.A(new_n16957_), .B(new_n11884_), .Y(new_n16971_));
  AOI21X1  g14535(.A0(new_n16970_), .A1(pi0792), .B0(new_n16971_), .Y(new_n16972_));
  MX2X1    g14536(.A(new_n16958_), .B(new_n16883_), .S0(new_n12711_), .Y(new_n16973_));
  INVX1    g14537(.A(new_n16973_), .Y(new_n16974_));
  AOI21X1  g14538(.A0(new_n16974_), .A1(pi0647), .B0(pi1157), .Y(new_n16975_));
  OAI21X1  g14539(.A0(new_n16972_), .A1(pi0647), .B0(new_n16975_), .Y(new_n16976_));
  INVX1    g14540(.A(new_n16961_), .Y(new_n16977_));
  AND2X1   g14541(.A(new_n16968_), .B(new_n16963_), .Y(new_n16978_));
  MX2X1    g14542(.A(new_n16978_), .B(new_n16977_), .S0(new_n11884_), .Y(new_n16979_));
  INVX1    g14543(.A(new_n16979_), .Y(new_n16980_));
  AOI21X1  g14544(.A0(new_n16913_), .A1(new_n12705_), .B0(new_n12706_), .Y(new_n16981_));
  OAI21X1  g14545(.A0(new_n16980_), .A1(new_n12705_), .B0(new_n16981_), .Y(new_n16982_));
  AND2X1   g14546(.A(new_n16982_), .B(new_n12723_), .Y(new_n16983_));
  AOI21X1  g14547(.A0(new_n16974_), .A1(new_n12705_), .B0(new_n12706_), .Y(new_n16984_));
  OAI21X1  g14548(.A0(new_n16972_), .A1(new_n12705_), .B0(new_n16984_), .Y(new_n16985_));
  AOI21X1  g14549(.A0(new_n16913_), .A1(pi0647), .B0(pi1157), .Y(new_n16986_));
  OAI21X1  g14550(.A0(new_n16980_), .A1(pi0647), .B0(new_n16986_), .Y(new_n16987_));
  AND2X1   g14551(.A(new_n16987_), .B(pi0630), .Y(new_n16988_));
  AOI22X1  g14552(.A0(new_n16988_), .A1(new_n16985_), .B0(new_n16983_), .B1(new_n16976_), .Y(new_n16989_));
  MX2X1    g14553(.A(new_n16989_), .B(new_n16972_), .S0(new_n11883_), .Y(new_n16990_));
  AND2X1   g14554(.A(new_n16987_), .B(new_n16982_), .Y(new_n16991_));
  MX2X1    g14555(.A(new_n16991_), .B(new_n16979_), .S0(new_n11883_), .Y(new_n16992_));
  AOI21X1  g14556(.A0(new_n16992_), .A1(new_n12743_), .B0(new_n12739_), .Y(new_n16993_));
  OAI21X1  g14557(.A0(new_n16990_), .A1(new_n12743_), .B0(new_n16993_), .Y(new_n16994_));
  MX2X1    g14558(.A(new_n16974_), .B(new_n16913_), .S0(new_n12735_), .Y(new_n16995_));
  OAI21X1  g14559(.A0(new_n16883_), .A1(pi0644), .B0(new_n12739_), .Y(new_n16996_));
  AOI21X1  g14560(.A0(new_n16995_), .A1(pi0644), .B0(new_n16996_), .Y(new_n16997_));
  NOR2X1   g14561(.A(new_n16997_), .B(new_n11882_), .Y(new_n16998_));
  AND2X1   g14562(.A(new_n16998_), .B(new_n16994_), .Y(new_n16999_));
  OR2X1    g14563(.A(new_n16972_), .B(pi0787), .Y(new_n17000_));
  OAI21X1  g14564(.A0(new_n16989_), .A1(new_n11883_), .B0(new_n17000_), .Y(new_n17001_));
  AND2X1   g14565(.A(new_n16992_), .B(pi0644), .Y(new_n17002_));
  OR2X1    g14566(.A(new_n17002_), .B(pi0715), .Y(new_n17003_));
  AOI21X1  g14567(.A0(new_n17001_), .A1(new_n12743_), .B0(new_n17003_), .Y(new_n17004_));
  OAI21X1  g14568(.A0(new_n16883_), .A1(new_n12743_), .B0(pi0715), .Y(new_n17005_));
  AOI21X1  g14569(.A0(new_n16995_), .A1(new_n12743_), .B0(new_n17005_), .Y(new_n17006_));
  OR2X1    g14570(.A(new_n17006_), .B(pi1160), .Y(new_n17007_));
  OAI21X1  g14571(.A0(new_n17007_), .A1(new_n17004_), .B0(pi0790), .Y(new_n17008_));
  AOI21X1  g14572(.A0(new_n16990_), .A1(new_n12897_), .B0(po1038), .Y(new_n17009_));
  OAI21X1  g14573(.A0(new_n17008_), .A1(new_n16999_), .B0(new_n17009_), .Y(new_n17010_));
  AOI21X1  g14574(.A0(po1038), .A1(new_n7469_), .B0(pi0832), .Y(new_n17011_));
  AOI21X1  g14575(.A0(pi1093), .A1(pi1092), .B0(pi0177), .Y(new_n17012_));
  INVX1    g14576(.A(new_n17012_), .Y(new_n17013_));
  AOI21X1  g14577(.A0(new_n12178_), .A1(new_n15065_), .B0(new_n17012_), .Y(new_n17014_));
  AOI21X1  g14578(.A0(new_n12601_), .A1(new_n2739_), .B0(new_n17014_), .Y(new_n17015_));
  INVX1    g14579(.A(new_n17014_), .Y(new_n17016_));
  AOI21X1  g14580(.A0(new_n17016_), .A1(new_n12776_), .B0(new_n12591_), .Y(new_n17017_));
  AOI21X1  g14581(.A0(new_n17015_), .A1(new_n12779_), .B0(pi1155), .Y(new_n17018_));
  OAI21X1  g14582(.A0(new_n17018_), .A1(new_n17017_), .B0(pi0785), .Y(new_n17019_));
  OAI21X1  g14583(.A0(new_n17015_), .A1(pi0785), .B0(new_n17019_), .Y(new_n17020_));
  INVX1    g14584(.A(new_n17020_), .Y(new_n17021_));
  AOI21X1  g14585(.A0(new_n17021_), .A1(new_n12785_), .B0(new_n12615_), .Y(new_n17022_));
  AOI21X1  g14586(.A0(new_n17021_), .A1(new_n12788_), .B0(pi1154), .Y(new_n17023_));
  OR2X1    g14587(.A(new_n17023_), .B(new_n17022_), .Y(new_n17024_));
  MX2X1    g14588(.A(new_n17024_), .B(new_n17020_), .S0(new_n11887_), .Y(new_n17025_));
  AND2X1   g14589(.A(new_n17025_), .B(new_n11886_), .Y(new_n17026_));
  AOI21X1  g14590(.A0(new_n17012_), .A1(new_n12637_), .B0(new_n12638_), .Y(new_n17027_));
  OAI21X1  g14591(.A0(new_n17025_), .A1(new_n12637_), .B0(new_n17027_), .Y(new_n17028_));
  AOI21X1  g14592(.A0(new_n17012_), .A1(pi0619), .B0(pi1159), .Y(new_n17029_));
  OAI21X1  g14593(.A0(new_n17025_), .A1(pi0619), .B0(new_n17029_), .Y(new_n17030_));
  AOI21X1  g14594(.A0(new_n17030_), .A1(new_n17028_), .B0(new_n11886_), .Y(new_n17031_));
  NOR2X1   g14595(.A(new_n17031_), .B(new_n17026_), .Y(new_n17032_));
  INVX1    g14596(.A(new_n17032_), .Y(new_n17033_));
  MX2X1    g14597(.A(new_n17033_), .B(new_n17013_), .S0(new_n12841_), .Y(new_n17034_));
  MX2X1    g14598(.A(new_n17034_), .B(new_n17013_), .S0(new_n12711_), .Y(new_n17035_));
  AOI21X1  g14599(.A0(new_n12566_), .A1(new_n16855_), .B0(new_n17012_), .Y(new_n17036_));
  AND2X1   g14600(.A(new_n12566_), .B(new_n16855_), .Y(new_n17037_));
  AND2X1   g14601(.A(new_n17037_), .B(new_n12493_), .Y(new_n17038_));
  MX2X1    g14602(.A(new_n17012_), .B(pi0625), .S0(new_n17037_), .Y(new_n17039_));
  NOR2X1   g14603(.A(new_n17012_), .B(pi1153), .Y(new_n17040_));
  INVX1    g14604(.A(new_n17040_), .Y(new_n17041_));
  OAI22X1  g14605(.A0(new_n17041_), .A1(new_n17038_), .B0(new_n17039_), .B1(new_n12494_), .Y(new_n17042_));
  MX2X1    g14606(.A(new_n17042_), .B(new_n17036_), .S0(new_n11889_), .Y(new_n17043_));
  NOR4X1   g14607(.A(new_n17043_), .B(new_n12765_), .C(new_n12764_), .D(new_n12762_), .Y(new_n17044_));
  INVX1    g14608(.A(new_n17044_), .Y(new_n17045_));
  NOR3X1   g14609(.A(new_n17045_), .B(new_n12870_), .C(new_n12851_), .Y(new_n17046_));
  INVX1    g14610(.A(new_n17046_), .Y(new_n17047_));
  AOI21X1  g14611(.A0(new_n17012_), .A1(pi0647), .B0(pi1157), .Y(new_n17048_));
  OAI21X1  g14612(.A0(new_n17047_), .A1(pi0647), .B0(new_n17048_), .Y(new_n17049_));
  MX2X1    g14613(.A(new_n17046_), .B(new_n17012_), .S0(new_n12705_), .Y(new_n17050_));
  OAI22X1  g14614(.A0(new_n17050_), .A1(new_n14387_), .B0(new_n17049_), .B1(new_n12723_), .Y(new_n17051_));
  AOI21X1  g14615(.A0(new_n17035_), .A1(new_n14385_), .B0(new_n17051_), .Y(new_n17052_));
  AOI21X1  g14616(.A0(new_n17013_), .A1(pi0626), .B0(new_n16352_), .Y(new_n17053_));
  OAI21X1  g14617(.A0(new_n17032_), .A1(pi0626), .B0(new_n17053_), .Y(new_n17054_));
  AOI21X1  g14618(.A0(new_n17013_), .A1(new_n12664_), .B0(new_n16356_), .Y(new_n17055_));
  OAI21X1  g14619(.A0(new_n17032_), .A1(new_n12664_), .B0(new_n17055_), .Y(new_n17056_));
  NAND2X1  g14620(.A(new_n17044_), .B(new_n12769_), .Y(new_n17057_));
  NAND3X1  g14621(.A(new_n17057_), .B(new_n17056_), .C(new_n17054_), .Y(new_n17058_));
  AND2X1   g14622(.A(new_n17058_), .B(pi0788), .Y(new_n17059_));
  INVX1    g14623(.A(new_n17059_), .Y(new_n17060_));
  NOR2X1   g14624(.A(new_n17036_), .B(new_n12120_), .Y(new_n17061_));
  NOR2X1   g14625(.A(new_n17061_), .B(new_n17016_), .Y(new_n17062_));
  INVX1    g14626(.A(new_n17062_), .Y(new_n17063_));
  MX2X1    g14627(.A(new_n17016_), .B(new_n12493_), .S0(new_n17061_), .Y(new_n17064_));
  NOR2X1   g14628(.A(new_n17064_), .B(new_n17041_), .Y(new_n17065_));
  OAI21X1  g14629(.A0(new_n17039_), .A1(new_n12494_), .B0(new_n12584_), .Y(new_n17066_));
  NOR3X1   g14630(.A(new_n17036_), .B(new_n12120_), .C(new_n12493_), .Y(new_n17067_));
  NOR3X1   g14631(.A(new_n17067_), .B(new_n17016_), .C(new_n12494_), .Y(new_n17068_));
  OAI21X1  g14632(.A0(new_n17041_), .A1(new_n17038_), .B0(pi0608), .Y(new_n17069_));
  OAI22X1  g14633(.A0(new_n17069_), .A1(new_n17068_), .B0(new_n17066_), .B1(new_n17065_), .Y(new_n17070_));
  MX2X1    g14634(.A(new_n17070_), .B(new_n17063_), .S0(new_n11889_), .Y(new_n17071_));
  OAI21X1  g14635(.A0(new_n17043_), .A1(new_n12590_), .B0(new_n12591_), .Y(new_n17072_));
  AOI21X1  g14636(.A0(new_n17071_), .A1(new_n12590_), .B0(new_n17072_), .Y(new_n17073_));
  NOR3X1   g14637(.A(new_n17073_), .B(new_n17017_), .C(pi0660), .Y(new_n17074_));
  OAI21X1  g14638(.A0(new_n17043_), .A1(pi0609), .B0(pi1155), .Y(new_n17075_));
  AOI21X1  g14639(.A0(new_n17071_), .A1(pi0609), .B0(new_n17075_), .Y(new_n17076_));
  NOR3X1   g14640(.A(new_n17076_), .B(new_n17018_), .C(new_n12596_), .Y(new_n17077_));
  OAI21X1  g14641(.A0(new_n17077_), .A1(new_n17074_), .B0(pi0785), .Y(new_n17078_));
  NAND2X1  g14642(.A(new_n17071_), .B(new_n11888_), .Y(new_n17079_));
  AND2X1   g14643(.A(new_n17079_), .B(new_n17078_), .Y(new_n17080_));
  NOR3X1   g14644(.A(new_n17043_), .B(new_n12762_), .C(new_n12614_), .Y(new_n17081_));
  NOR2X1   g14645(.A(new_n17081_), .B(pi1154), .Y(new_n17082_));
  OAI21X1  g14646(.A0(new_n17080_), .A1(pi0618), .B0(new_n17082_), .Y(new_n17083_));
  NOR2X1   g14647(.A(new_n17022_), .B(pi0627), .Y(new_n17084_));
  NOR3X1   g14648(.A(new_n17043_), .B(new_n12762_), .C(pi0618), .Y(new_n17085_));
  NOR2X1   g14649(.A(new_n17085_), .B(new_n12615_), .Y(new_n17086_));
  OAI21X1  g14650(.A0(new_n17080_), .A1(new_n12614_), .B0(new_n17086_), .Y(new_n17087_));
  NOR2X1   g14651(.A(new_n17023_), .B(new_n12622_), .Y(new_n17088_));
  AOI22X1  g14652(.A0(new_n17088_), .A1(new_n17087_), .B0(new_n17084_), .B1(new_n17083_), .Y(new_n17089_));
  MX2X1    g14653(.A(new_n17089_), .B(new_n17080_), .S0(new_n11887_), .Y(new_n17090_));
  OR4X1    g14654(.A(new_n17043_), .B(new_n12764_), .C(new_n12762_), .D(new_n12637_), .Y(new_n17091_));
  AND2X1   g14655(.A(new_n17091_), .B(new_n12638_), .Y(new_n17092_));
  OAI21X1  g14656(.A0(new_n17090_), .A1(pi0619), .B0(new_n17092_), .Y(new_n17093_));
  AND2X1   g14657(.A(new_n17028_), .B(new_n12645_), .Y(new_n17094_));
  AND2X1   g14658(.A(new_n17094_), .B(new_n17093_), .Y(new_n17095_));
  NOR4X1   g14659(.A(new_n17043_), .B(new_n12764_), .C(new_n12762_), .D(pi0619), .Y(new_n17096_));
  NOR2X1   g14660(.A(new_n17096_), .B(new_n12638_), .Y(new_n17097_));
  OAI21X1  g14661(.A0(new_n17090_), .A1(new_n12637_), .B0(new_n17097_), .Y(new_n17098_));
  AND2X1   g14662(.A(new_n17030_), .B(pi0648), .Y(new_n17099_));
  AOI21X1  g14663(.A0(new_n17099_), .A1(new_n17098_), .B0(new_n11886_), .Y(new_n17100_));
  INVX1    g14664(.A(new_n17100_), .Y(new_n17101_));
  AOI21X1  g14665(.A0(new_n17090_), .A1(new_n11886_), .B0(new_n14264_), .Y(new_n17102_));
  OAI21X1  g14666(.A0(new_n17101_), .A1(new_n17095_), .B0(new_n17102_), .Y(new_n17103_));
  AOI21X1  g14667(.A0(new_n17103_), .A1(new_n17060_), .B0(new_n14273_), .Y(new_n17104_));
  INVX1    g14668(.A(new_n17034_), .Y(new_n17105_));
  AND2X1   g14669(.A(new_n17044_), .B(new_n12852_), .Y(new_n17106_));
  AOI22X1  g14670(.A0(new_n17106_), .A1(new_n14564_), .B0(new_n17105_), .B1(new_n12867_), .Y(new_n17107_));
  AOI22X1  g14671(.A0(new_n17106_), .A1(new_n14566_), .B0(new_n17105_), .B1(new_n12865_), .Y(new_n17108_));
  MX2X1    g14672(.A(new_n17108_), .B(new_n17107_), .S0(new_n12689_), .Y(new_n17109_));
  OAI21X1  g14673(.A0(new_n17109_), .A1(new_n11884_), .B0(new_n14562_), .Y(new_n17110_));
  OAI22X1  g14674(.A0(new_n17110_), .A1(new_n17104_), .B0(new_n17052_), .B1(new_n11883_), .Y(new_n17111_));
  INVX1    g14675(.A(new_n17111_), .Y(new_n17112_));
  OAI21X1  g14676(.A0(new_n17050_), .A1(new_n12706_), .B0(new_n17049_), .Y(new_n17113_));
  MX2X1    g14677(.A(new_n17113_), .B(new_n17047_), .S0(new_n11883_), .Y(new_n17114_));
  OAI21X1  g14678(.A0(new_n17114_), .A1(pi0644), .B0(pi0715), .Y(new_n17115_));
  AOI21X1  g14679(.A0(new_n17112_), .A1(pi0644), .B0(new_n17115_), .Y(new_n17116_));
  OR4X1    g14680(.A(new_n12734_), .B(new_n2739_), .C(new_n11883_), .D(pi0177), .Y(new_n17117_));
  OAI21X1  g14681(.A0(new_n17035_), .A1(new_n12735_), .B0(new_n17117_), .Y(new_n17118_));
  OAI21X1  g14682(.A0(new_n17013_), .A1(pi0644), .B0(new_n12739_), .Y(new_n17119_));
  AOI21X1  g14683(.A0(new_n17118_), .A1(pi0644), .B0(new_n17119_), .Y(new_n17120_));
  OR2X1    g14684(.A(new_n17120_), .B(new_n11882_), .Y(new_n17121_));
  OAI21X1  g14685(.A0(new_n17114_), .A1(new_n12743_), .B0(new_n12739_), .Y(new_n17122_));
  AOI21X1  g14686(.A0(new_n17112_), .A1(new_n12743_), .B0(new_n17122_), .Y(new_n17123_));
  OAI21X1  g14687(.A0(new_n17013_), .A1(new_n12743_), .B0(pi0715), .Y(new_n17124_));
  AOI21X1  g14688(.A0(new_n17118_), .A1(new_n12743_), .B0(new_n17124_), .Y(new_n17125_));
  OR2X1    g14689(.A(new_n17125_), .B(pi1160), .Y(new_n17126_));
  OAI22X1  g14690(.A0(new_n17126_), .A1(new_n17123_), .B0(new_n17121_), .B1(new_n17116_), .Y(new_n17127_));
  OAI21X1  g14691(.A0(new_n17111_), .A1(pi0790), .B0(pi0832), .Y(new_n17128_));
  AOI21X1  g14692(.A0(new_n17127_), .A1(pi0790), .B0(new_n17128_), .Y(new_n17129_));
  AOI21X1  g14693(.A0(new_n17011_), .A1(new_n17010_), .B0(new_n17129_), .Y(po0334));
  AOI21X1  g14694(.A0(pi1093), .A1(pi1092), .B0(pi0178), .Y(new_n17131_));
  INVX1    g14695(.A(new_n17131_), .Y(new_n17132_));
  AOI21X1  g14696(.A0(new_n12178_), .A1(new_n15106_), .B0(new_n17131_), .Y(new_n17133_));
  AOI21X1  g14697(.A0(new_n12601_), .A1(new_n2739_), .B0(new_n17133_), .Y(new_n17134_));
  NAND2X1  g14698(.A(new_n12178_), .B(new_n15106_), .Y(new_n17135_));
  OAI21X1  g14699(.A0(new_n17135_), .A1(new_n13436_), .B0(new_n17134_), .Y(new_n17136_));
  AND2X1   g14700(.A(new_n17136_), .B(pi1155), .Y(new_n17137_));
  NOR2X1   g14701(.A(new_n17135_), .B(new_n13436_), .Y(new_n17138_));
  NOR3X1   g14702(.A(new_n17138_), .B(new_n17131_), .C(pi1155), .Y(new_n17139_));
  OAI21X1  g14703(.A0(new_n17139_), .A1(new_n17137_), .B0(pi0785), .Y(new_n17140_));
  OAI21X1  g14704(.A0(new_n17134_), .A1(pi0785), .B0(new_n17140_), .Y(new_n17141_));
  INVX1    g14705(.A(new_n17141_), .Y(new_n17142_));
  AOI21X1  g14706(.A0(new_n17142_), .A1(new_n12785_), .B0(new_n12615_), .Y(new_n17143_));
  AOI21X1  g14707(.A0(new_n17142_), .A1(new_n12788_), .B0(pi1154), .Y(new_n17144_));
  NOR2X1   g14708(.A(new_n17144_), .B(new_n17143_), .Y(new_n17145_));
  MX2X1    g14709(.A(new_n17145_), .B(new_n17142_), .S0(new_n11887_), .Y(new_n17146_));
  OR2X1    g14710(.A(new_n17146_), .B(pi0789), .Y(new_n17147_));
  AOI21X1  g14711(.A0(new_n17146_), .A1(new_n15910_), .B0(new_n12638_), .Y(new_n17148_));
  AOI21X1  g14712(.A0(new_n17146_), .A1(new_n15912_), .B0(pi1159), .Y(new_n17149_));
  OAI21X1  g14713(.A0(new_n17149_), .A1(new_n17148_), .B0(pi0789), .Y(new_n17150_));
  AND2X1   g14714(.A(new_n17150_), .B(new_n17147_), .Y(new_n17151_));
  INVX1    g14715(.A(new_n17151_), .Y(new_n17152_));
  MX2X1    g14716(.A(new_n17152_), .B(new_n17132_), .S0(new_n12841_), .Y(new_n17153_));
  MX2X1    g14717(.A(new_n17153_), .B(new_n17132_), .S0(new_n12711_), .Y(new_n17154_));
  AOI21X1  g14718(.A0(new_n12566_), .A1(new_n15112_), .B0(new_n17131_), .Y(new_n17155_));
  INVX1    g14719(.A(new_n17155_), .Y(new_n17156_));
  NOR3X1   g14720(.A(new_n13585_), .B(pi0688), .C(pi0625), .Y(new_n17157_));
  OR2X1    g14721(.A(new_n17157_), .B(new_n17155_), .Y(new_n17158_));
  NOR2X1   g14722(.A(new_n17131_), .B(pi1153), .Y(new_n17159_));
  INVX1    g14723(.A(new_n17159_), .Y(new_n17160_));
  OAI21X1  g14724(.A0(new_n17160_), .A1(new_n17157_), .B0(pi0778), .Y(new_n17161_));
  AOI21X1  g14725(.A0(new_n17158_), .A1(pi1153), .B0(new_n17161_), .Y(new_n17162_));
  AOI21X1  g14726(.A0(new_n17156_), .A1(new_n11889_), .B0(new_n17162_), .Y(new_n17163_));
  NOR4X1   g14727(.A(new_n17163_), .B(new_n12765_), .C(new_n12764_), .D(new_n12762_), .Y(new_n17164_));
  INVX1    g14728(.A(new_n17164_), .Y(new_n17165_));
  NOR3X1   g14729(.A(new_n17165_), .B(new_n12870_), .C(new_n12851_), .Y(new_n17166_));
  INVX1    g14730(.A(new_n17166_), .Y(new_n17167_));
  AOI21X1  g14731(.A0(new_n17131_), .A1(pi0647), .B0(pi1157), .Y(new_n17168_));
  OAI21X1  g14732(.A0(new_n17167_), .A1(pi0647), .B0(new_n17168_), .Y(new_n17169_));
  MX2X1    g14733(.A(new_n17166_), .B(new_n17131_), .S0(new_n12705_), .Y(new_n17170_));
  OAI22X1  g14734(.A0(new_n17170_), .A1(new_n14387_), .B0(new_n17169_), .B1(new_n12723_), .Y(new_n17171_));
  AOI21X1  g14735(.A0(new_n17154_), .A1(new_n14385_), .B0(new_n17171_), .Y(new_n17172_));
  NOR2X1   g14736(.A(new_n17172_), .B(new_n11883_), .Y(new_n17173_));
  AOI21X1  g14737(.A0(new_n17132_), .A1(pi0626), .B0(new_n16352_), .Y(new_n17174_));
  OAI21X1  g14738(.A0(new_n17151_), .A1(pi0626), .B0(new_n17174_), .Y(new_n17175_));
  AOI21X1  g14739(.A0(new_n17150_), .A1(new_n17147_), .B0(new_n12664_), .Y(new_n17176_));
  NOR2X1   g14740(.A(new_n17131_), .B(pi0626), .Y(new_n17177_));
  NOR3X1   g14741(.A(new_n17177_), .B(new_n17176_), .C(new_n16356_), .Y(new_n17178_));
  AOI21X1  g14742(.A0(new_n17164_), .A1(new_n12769_), .B0(new_n17178_), .Y(new_n17179_));
  AOI21X1  g14743(.A0(new_n17179_), .A1(new_n17175_), .B0(new_n11885_), .Y(new_n17180_));
  INVX1    g14744(.A(new_n17133_), .Y(new_n17181_));
  AOI21X1  g14745(.A0(new_n17156_), .A1(new_n12171_), .B0(new_n17181_), .Y(new_n17182_));
  NOR3X1   g14746(.A(new_n17155_), .B(new_n12120_), .C(new_n12493_), .Y(new_n17183_));
  OR2X1    g14747(.A(new_n17182_), .B(new_n17183_), .Y(new_n17184_));
  NOR2X1   g14748(.A(new_n17157_), .B(new_n17155_), .Y(new_n17185_));
  OAI21X1  g14749(.A0(new_n17185_), .A1(new_n12494_), .B0(new_n12584_), .Y(new_n17186_));
  AOI21X1  g14750(.A0(new_n17184_), .A1(new_n17159_), .B0(new_n17186_), .Y(new_n17187_));
  NOR3X1   g14751(.A(new_n17183_), .B(new_n17181_), .C(new_n12494_), .Y(new_n17188_));
  OAI21X1  g14752(.A0(new_n17160_), .A1(new_n17157_), .B0(pi0608), .Y(new_n17189_));
  NOR2X1   g14753(.A(new_n17189_), .B(new_n17188_), .Y(new_n17190_));
  OAI21X1  g14754(.A0(new_n17190_), .A1(new_n17187_), .B0(pi0778), .Y(new_n17191_));
  OAI21X1  g14755(.A0(new_n17182_), .A1(pi0778), .B0(new_n17191_), .Y(new_n17192_));
  OAI21X1  g14756(.A0(new_n17163_), .A1(new_n12590_), .B0(new_n12591_), .Y(new_n17193_));
  AOI21X1  g14757(.A0(new_n17192_), .A1(new_n12590_), .B0(new_n17193_), .Y(new_n17194_));
  NOR3X1   g14758(.A(new_n17194_), .B(new_n17137_), .C(pi0660), .Y(new_n17195_));
  OAI21X1  g14759(.A0(new_n17163_), .A1(pi0609), .B0(pi1155), .Y(new_n17196_));
  AOI21X1  g14760(.A0(new_n17192_), .A1(pi0609), .B0(new_n17196_), .Y(new_n17197_));
  NOR3X1   g14761(.A(new_n17197_), .B(new_n17139_), .C(new_n12596_), .Y(new_n17198_));
  OAI21X1  g14762(.A0(new_n17198_), .A1(new_n17195_), .B0(pi0785), .Y(new_n17199_));
  NAND2X1  g14763(.A(new_n17192_), .B(new_n11888_), .Y(new_n17200_));
  AND2X1   g14764(.A(new_n17200_), .B(new_n17199_), .Y(new_n17201_));
  NOR3X1   g14765(.A(new_n17163_), .B(new_n12762_), .C(new_n12614_), .Y(new_n17202_));
  NOR2X1   g14766(.A(new_n17202_), .B(pi1154), .Y(new_n17203_));
  OAI21X1  g14767(.A0(new_n17201_), .A1(pi0618), .B0(new_n17203_), .Y(new_n17204_));
  NOR2X1   g14768(.A(new_n17143_), .B(pi0627), .Y(new_n17205_));
  NOR3X1   g14769(.A(new_n17163_), .B(new_n12762_), .C(pi0618), .Y(new_n17206_));
  NOR2X1   g14770(.A(new_n17206_), .B(new_n12615_), .Y(new_n17207_));
  OAI21X1  g14771(.A0(new_n17201_), .A1(new_n12614_), .B0(new_n17207_), .Y(new_n17208_));
  NOR2X1   g14772(.A(new_n17144_), .B(new_n12622_), .Y(new_n17209_));
  AOI22X1  g14773(.A0(new_n17209_), .A1(new_n17208_), .B0(new_n17205_), .B1(new_n17204_), .Y(new_n17210_));
  MX2X1    g14774(.A(new_n17210_), .B(new_n17201_), .S0(new_n11887_), .Y(new_n17211_));
  OR4X1    g14775(.A(new_n17163_), .B(new_n12764_), .C(new_n12762_), .D(new_n12637_), .Y(new_n17212_));
  AND2X1   g14776(.A(new_n17212_), .B(new_n12638_), .Y(new_n17213_));
  OAI21X1  g14777(.A0(new_n17211_), .A1(pi0619), .B0(new_n17213_), .Y(new_n17214_));
  NOR2X1   g14778(.A(new_n17148_), .B(pi0648), .Y(new_n17215_));
  AND2X1   g14779(.A(new_n17215_), .B(new_n17214_), .Y(new_n17216_));
  INVX1    g14780(.A(new_n17216_), .Y(new_n17217_));
  NOR4X1   g14781(.A(new_n17163_), .B(new_n12764_), .C(new_n12762_), .D(pi0619), .Y(new_n17218_));
  NOR2X1   g14782(.A(new_n17218_), .B(new_n12638_), .Y(new_n17219_));
  OAI21X1  g14783(.A0(new_n17211_), .A1(new_n12637_), .B0(new_n17219_), .Y(new_n17220_));
  NOR2X1   g14784(.A(new_n17149_), .B(new_n12645_), .Y(new_n17221_));
  AOI21X1  g14785(.A0(new_n17221_), .A1(new_n17220_), .B0(new_n11886_), .Y(new_n17222_));
  AOI21X1  g14786(.A0(new_n17211_), .A1(new_n11886_), .B0(new_n14264_), .Y(new_n17223_));
  INVX1    g14787(.A(new_n17223_), .Y(new_n17224_));
  AOI21X1  g14788(.A0(new_n17222_), .A1(new_n17217_), .B0(new_n17224_), .Y(new_n17225_));
  OAI21X1  g14789(.A0(new_n17225_), .A1(new_n17180_), .B0(new_n16350_), .Y(new_n17226_));
  INVX1    g14790(.A(new_n17153_), .Y(new_n17227_));
  AND2X1   g14791(.A(new_n17164_), .B(new_n12852_), .Y(new_n17228_));
  AOI22X1  g14792(.A0(new_n17228_), .A1(new_n14564_), .B0(new_n17227_), .B1(new_n12867_), .Y(new_n17229_));
  AOI22X1  g14793(.A0(new_n17228_), .A1(new_n14566_), .B0(new_n17227_), .B1(new_n12865_), .Y(new_n17230_));
  MX2X1    g14794(.A(new_n17230_), .B(new_n17229_), .S0(new_n12689_), .Y(new_n17231_));
  OAI21X1  g14795(.A0(new_n17231_), .A1(new_n11884_), .B0(new_n14562_), .Y(new_n17232_));
  INVX1    g14796(.A(new_n17232_), .Y(new_n17233_));
  AOI21X1  g14797(.A0(new_n17233_), .A1(new_n17226_), .B0(new_n17173_), .Y(new_n17234_));
  OAI21X1  g14798(.A0(new_n17170_), .A1(new_n12706_), .B0(new_n17169_), .Y(new_n17235_));
  MX2X1    g14799(.A(new_n17235_), .B(new_n17167_), .S0(new_n11883_), .Y(new_n17236_));
  OAI21X1  g14800(.A0(new_n17236_), .A1(pi0644), .B0(pi0715), .Y(new_n17237_));
  AOI21X1  g14801(.A0(new_n17234_), .A1(pi0644), .B0(new_n17237_), .Y(new_n17238_));
  OR4X1    g14802(.A(new_n12734_), .B(new_n2739_), .C(new_n11883_), .D(pi0178), .Y(new_n17239_));
  OAI21X1  g14803(.A0(new_n17154_), .A1(new_n12735_), .B0(new_n17239_), .Y(new_n17240_));
  OAI21X1  g14804(.A0(new_n17132_), .A1(pi0644), .B0(new_n12739_), .Y(new_n17241_));
  AOI21X1  g14805(.A0(new_n17240_), .A1(pi0644), .B0(new_n17241_), .Y(new_n17242_));
  OR2X1    g14806(.A(new_n17242_), .B(new_n11882_), .Y(new_n17243_));
  OAI21X1  g14807(.A0(new_n17236_), .A1(new_n12743_), .B0(new_n12739_), .Y(new_n17244_));
  AOI21X1  g14808(.A0(new_n17234_), .A1(new_n12743_), .B0(new_n17244_), .Y(new_n17245_));
  OAI21X1  g14809(.A0(new_n17132_), .A1(new_n12743_), .B0(pi0715), .Y(new_n17246_));
  AOI21X1  g14810(.A0(new_n17240_), .A1(new_n12743_), .B0(new_n17246_), .Y(new_n17247_));
  OR2X1    g14811(.A(new_n17247_), .B(pi1160), .Y(new_n17248_));
  OAI22X1  g14812(.A0(new_n17248_), .A1(new_n17245_), .B0(new_n17243_), .B1(new_n17238_), .Y(new_n17249_));
  NAND2X1  g14813(.A(new_n17249_), .B(pi0790), .Y(new_n17250_));
  AOI21X1  g14814(.A0(new_n17234_), .A1(new_n12897_), .B0(new_n12898_), .Y(new_n17251_));
  INVX1    g14815(.A(new_n12691_), .Y(new_n17252_));
  AOI21X1  g14816(.A0(new_n13699_), .A1(new_n3129_), .B0(pi0178), .Y(new_n17253_));
  INVX1    g14817(.A(new_n17253_), .Y(new_n17254_));
  OAI21X1  g14818(.A0(new_n3810_), .A1(pi0688), .B0(new_n17253_), .Y(new_n17255_));
  AOI21X1  g14819(.A0(new_n12955_), .A1(pi0178), .B0(pi0038), .Y(new_n17256_));
  OAI22X1  g14820(.A0(new_n17256_), .A1(new_n3810_), .B0(new_n12953_), .B1(pi0178), .Y(new_n17257_));
  OAI21X1  g14821(.A0(new_n12202_), .A1(pi0178), .B0(new_n12567_), .Y(new_n17258_));
  NAND3X1  g14822(.A(new_n17258_), .B(new_n17257_), .C(new_n15112_), .Y(new_n17259_));
  AND2X1   g14823(.A(new_n17259_), .B(new_n17255_), .Y(new_n17260_));
  INVX1    g14824(.A(new_n17260_), .Y(new_n17261_));
  AOI21X1  g14825(.A0(new_n17253_), .A1(new_n12493_), .B0(new_n12494_), .Y(new_n17262_));
  OAI21X1  g14826(.A0(new_n17260_), .A1(new_n12493_), .B0(new_n17262_), .Y(new_n17263_));
  AOI21X1  g14827(.A0(new_n17253_), .A1(pi0625), .B0(pi1153), .Y(new_n17264_));
  OAI21X1  g14828(.A0(new_n17260_), .A1(pi0625), .B0(new_n17264_), .Y(new_n17265_));
  AND2X1   g14829(.A(new_n17265_), .B(new_n17263_), .Y(new_n17266_));
  MX2X1    g14830(.A(new_n17266_), .B(new_n17261_), .S0(new_n11889_), .Y(new_n17267_));
  MX2X1    g14831(.A(new_n17267_), .B(new_n17253_), .S0(new_n12618_), .Y(new_n17268_));
  INVX1    g14832(.A(new_n17268_), .Y(new_n17269_));
  MX2X1    g14833(.A(new_n17269_), .B(new_n17254_), .S0(new_n12641_), .Y(new_n17270_));
  INVX1    g14834(.A(new_n17270_), .Y(new_n17271_));
  MX2X1    g14835(.A(new_n17271_), .B(new_n17253_), .S0(new_n12659_), .Y(new_n17272_));
  AND2X1   g14836(.A(new_n17253_), .B(new_n12691_), .Y(new_n17273_));
  AOI21X1  g14837(.A0(new_n17272_), .A1(new_n17252_), .B0(new_n17273_), .Y(new_n17274_));
  AOI21X1  g14838(.A0(new_n17253_), .A1(new_n12683_), .B0(new_n12684_), .Y(new_n17275_));
  OAI21X1  g14839(.A0(new_n17274_), .A1(new_n12683_), .B0(new_n17275_), .Y(new_n17276_));
  AOI21X1  g14840(.A0(new_n17253_), .A1(pi0628), .B0(pi1156), .Y(new_n17277_));
  OAI21X1  g14841(.A0(new_n17274_), .A1(pi0628), .B0(new_n17277_), .Y(new_n17278_));
  AOI21X1  g14842(.A0(new_n17278_), .A1(new_n17276_), .B0(new_n11884_), .Y(new_n17279_));
  AOI21X1  g14843(.A0(new_n17274_), .A1(new_n11884_), .B0(new_n17279_), .Y(new_n17280_));
  MX2X1    g14844(.A(new_n17280_), .B(new_n17253_), .S0(pi0647), .Y(new_n17281_));
  MX2X1    g14845(.A(new_n17280_), .B(new_n17253_), .S0(new_n12705_), .Y(new_n17282_));
  MX2X1    g14846(.A(new_n17282_), .B(new_n17281_), .S0(new_n12706_), .Y(new_n17283_));
  MX2X1    g14847(.A(new_n17283_), .B(new_n17280_), .S0(new_n11883_), .Y(new_n17284_));
  AOI21X1  g14848(.A0(new_n17284_), .A1(new_n12743_), .B0(new_n12739_), .Y(new_n17285_));
  OAI22X1  g14849(.A0(new_n14342_), .A1(pi0760), .B0(new_n12202_), .B1(pi0178), .Y(new_n17286_));
  AOI21X1  g14850(.A0(new_n13977_), .A1(pi0178), .B0(pi0760), .Y(new_n17287_));
  OAI21X1  g14851(.A0(new_n12910_), .A1(pi0178), .B0(new_n17287_), .Y(new_n17288_));
  NAND3X1  g14852(.A(new_n12090_), .B(pi0760), .C(new_n10020_), .Y(new_n17289_));
  AOI21X1  g14853(.A0(new_n17289_), .A1(new_n17288_), .B0(pi0038), .Y(new_n17290_));
  AOI21X1  g14854(.A0(new_n17286_), .A1(pi0038), .B0(new_n17290_), .Y(new_n17291_));
  MX2X1    g14855(.A(new_n17291_), .B(pi0178), .S0(new_n3810_), .Y(new_n17292_));
  AND2X1   g14856(.A(new_n17292_), .B(new_n12623_), .Y(new_n17293_));
  AOI21X1  g14857(.A0(new_n17254_), .A1(new_n12601_), .B0(new_n17293_), .Y(new_n17294_));
  AOI22X1  g14858(.A0(new_n17293_), .A1(pi0609), .B0(new_n17254_), .B1(new_n13430_), .Y(new_n17295_));
  AOI22X1  g14859(.A0(new_n17293_), .A1(new_n12590_), .B0(new_n17254_), .B1(new_n13436_), .Y(new_n17296_));
  MX2X1    g14860(.A(new_n17296_), .B(new_n17295_), .S0(pi1155), .Y(new_n17297_));
  MX2X1    g14861(.A(new_n17297_), .B(new_n17294_), .S0(new_n11888_), .Y(new_n17298_));
  OAI21X1  g14862(.A0(new_n17254_), .A1(pi0618), .B0(pi1154), .Y(new_n17299_));
  AOI21X1  g14863(.A0(new_n17298_), .A1(pi0618), .B0(new_n17299_), .Y(new_n17300_));
  OAI21X1  g14864(.A0(new_n17254_), .A1(new_n12614_), .B0(new_n12615_), .Y(new_n17301_));
  AOI21X1  g14865(.A0(new_n17298_), .A1(new_n12614_), .B0(new_n17301_), .Y(new_n17302_));
  NOR2X1   g14866(.A(new_n17302_), .B(new_n17300_), .Y(new_n17303_));
  MX2X1    g14867(.A(new_n17303_), .B(new_n17298_), .S0(new_n11887_), .Y(new_n17304_));
  OAI21X1  g14868(.A0(new_n17254_), .A1(pi0619), .B0(pi1159), .Y(new_n17305_));
  AOI21X1  g14869(.A0(new_n17304_), .A1(pi0619), .B0(new_n17305_), .Y(new_n17306_));
  OAI21X1  g14870(.A0(new_n17254_), .A1(new_n12637_), .B0(new_n12638_), .Y(new_n17307_));
  AOI21X1  g14871(.A0(new_n17304_), .A1(new_n12637_), .B0(new_n17307_), .Y(new_n17308_));
  NOR2X1   g14872(.A(new_n17308_), .B(new_n17306_), .Y(new_n17309_));
  MX2X1    g14873(.A(new_n17309_), .B(new_n17304_), .S0(new_n11886_), .Y(new_n17310_));
  MX2X1    g14874(.A(new_n17310_), .B(new_n17253_), .S0(new_n12841_), .Y(new_n17311_));
  MX2X1    g14875(.A(new_n17311_), .B(new_n17253_), .S0(new_n12711_), .Y(new_n17312_));
  MX2X1    g14876(.A(new_n17312_), .B(new_n17253_), .S0(new_n12735_), .Y(new_n17313_));
  OAI21X1  g14877(.A0(new_n17254_), .A1(pi0644), .B0(new_n12739_), .Y(new_n17314_));
  AOI21X1  g14878(.A0(new_n17313_), .A1(pi0644), .B0(new_n17314_), .Y(new_n17315_));
  OR2X1    g14879(.A(new_n17315_), .B(new_n11882_), .Y(new_n17316_));
  AOI21X1  g14880(.A0(new_n17284_), .A1(pi0644), .B0(pi0715), .Y(new_n17317_));
  OAI21X1  g14881(.A0(new_n17254_), .A1(new_n12743_), .B0(pi0715), .Y(new_n17318_));
  AOI21X1  g14882(.A0(new_n17313_), .A1(new_n12743_), .B0(new_n17318_), .Y(new_n17319_));
  OR2X1    g14883(.A(new_n17319_), .B(pi1160), .Y(new_n17320_));
  OAI22X1  g14884(.A0(new_n17320_), .A1(new_n17317_), .B0(new_n17316_), .B1(new_n17285_), .Y(new_n17321_));
  NOR3X1   g14885(.A(new_n17319_), .B(pi1160), .C(pi0644), .Y(new_n17322_));
  NOR3X1   g14886(.A(new_n17315_), .B(new_n11882_), .C(new_n12743_), .Y(new_n17323_));
  NOR3X1   g14887(.A(new_n17323_), .B(new_n17322_), .C(new_n12897_), .Y(new_n17324_));
  MX2X1    g14888(.A(new_n17278_), .B(new_n17276_), .S0(new_n12689_), .Y(new_n17325_));
  OAI21X1  g14889(.A0(new_n17311_), .A1(new_n14395_), .B0(new_n17325_), .Y(new_n17326_));
  NAND2X1  g14890(.A(new_n17326_), .B(pi0792), .Y(new_n17327_));
  OR2X1    g14891(.A(new_n17291_), .B(new_n15112_), .Y(new_n17328_));
  OAI21X1  g14892(.A0(new_n12349_), .A1(new_n10020_), .B0(pi0760), .Y(new_n17329_));
  AOI21X1  g14893(.A0(new_n12289_), .A1(new_n10020_), .B0(new_n17329_), .Y(new_n17330_));
  OAI21X1  g14894(.A0(new_n12440_), .A1(pi0178), .B0(new_n15106_), .Y(new_n17331_));
  AOI21X1  g14895(.A0(new_n12401_), .A1(pi0178), .B0(new_n17331_), .Y(new_n17332_));
  OR2X1    g14896(.A(new_n17332_), .B(new_n2959_), .Y(new_n17333_));
  AND2X1   g14897(.A(new_n12467_), .B(pi0178), .Y(new_n17334_));
  OAI21X1  g14898(.A0(new_n12454_), .A1(pi0178), .B0(pi0760), .Y(new_n17335_));
  NOR4X1   g14899(.A(new_n13391_), .B(new_n12908_), .C(new_n12907_), .D(pi0178), .Y(new_n17336_));
  OAI21X1  g14900(.A0(new_n12929_), .A1(new_n10020_), .B0(new_n15106_), .Y(new_n17337_));
  OAI22X1  g14901(.A0(new_n17337_), .A1(new_n17336_), .B0(new_n17335_), .B1(new_n17334_), .Y(new_n17338_));
  AOI21X1  g14902(.A0(new_n17338_), .A1(new_n2959_), .B0(pi0038), .Y(new_n17339_));
  OAI21X1  g14903(.A0(new_n17333_), .A1(new_n17330_), .B0(new_n17339_), .Y(new_n17340_));
  OAI21X1  g14904(.A0(new_n12478_), .A1(pi0760), .B0(new_n13669_), .Y(new_n17341_));
  NAND2X1  g14905(.A(new_n17341_), .B(new_n10020_), .Y(new_n17342_));
  AOI21X1  g14906(.A0(new_n17135_), .A1(new_n14209_), .B0(new_n10020_), .Y(new_n17343_));
  AOI21X1  g14907(.A0(new_n17343_), .A1(new_n6857_), .B0(new_n2996_), .Y(new_n17344_));
  AOI21X1  g14908(.A0(new_n17344_), .A1(new_n17342_), .B0(pi0688), .Y(new_n17345_));
  AOI21X1  g14909(.A0(new_n17345_), .A1(new_n17340_), .B0(new_n3810_), .Y(new_n17346_));
  AOI22X1  g14910(.A0(new_n17346_), .A1(new_n17328_), .B0(new_n3810_), .B1(pi0178), .Y(new_n17347_));
  OAI21X1  g14911(.A0(new_n17292_), .A1(new_n12493_), .B0(new_n12494_), .Y(new_n17348_));
  AOI21X1  g14912(.A0(new_n17347_), .A1(new_n12493_), .B0(new_n17348_), .Y(new_n17349_));
  NAND2X1  g14913(.A(new_n17263_), .B(new_n12584_), .Y(new_n17350_));
  OAI21X1  g14914(.A0(new_n17292_), .A1(pi0625), .B0(pi1153), .Y(new_n17351_));
  AOI21X1  g14915(.A0(new_n17347_), .A1(pi0625), .B0(new_n17351_), .Y(new_n17352_));
  NAND2X1  g14916(.A(new_n17265_), .B(pi0608), .Y(new_n17353_));
  OAI22X1  g14917(.A0(new_n17353_), .A1(new_n17352_), .B0(new_n17350_), .B1(new_n17349_), .Y(new_n17354_));
  MX2X1    g14918(.A(new_n17354_), .B(new_n17347_), .S0(new_n11889_), .Y(new_n17355_));
  INVX1    g14919(.A(new_n17267_), .Y(new_n17356_));
  OAI21X1  g14920(.A0(new_n17356_), .A1(new_n12590_), .B0(new_n12591_), .Y(new_n17357_));
  AOI21X1  g14921(.A0(new_n17355_), .A1(new_n12590_), .B0(new_n17357_), .Y(new_n17358_));
  OAI21X1  g14922(.A0(new_n17295_), .A1(new_n12591_), .B0(new_n12596_), .Y(new_n17359_));
  OAI21X1  g14923(.A0(new_n17356_), .A1(pi0609), .B0(pi1155), .Y(new_n17360_));
  AOI21X1  g14924(.A0(new_n17355_), .A1(pi0609), .B0(new_n17360_), .Y(new_n17361_));
  OAI21X1  g14925(.A0(new_n17296_), .A1(pi1155), .B0(pi0660), .Y(new_n17362_));
  OAI22X1  g14926(.A0(new_n17362_), .A1(new_n17361_), .B0(new_n17359_), .B1(new_n17358_), .Y(new_n17363_));
  MX2X1    g14927(.A(new_n17363_), .B(new_n17355_), .S0(new_n11888_), .Y(new_n17364_));
  OAI21X1  g14928(.A0(new_n17269_), .A1(new_n12614_), .B0(new_n12615_), .Y(new_n17365_));
  AOI21X1  g14929(.A0(new_n17364_), .A1(new_n12614_), .B0(new_n17365_), .Y(new_n17366_));
  OR2X1    g14930(.A(new_n17300_), .B(pi0627), .Y(new_n17367_));
  OAI21X1  g14931(.A0(new_n17269_), .A1(pi0618), .B0(pi1154), .Y(new_n17368_));
  AOI21X1  g14932(.A0(new_n17364_), .A1(pi0618), .B0(new_n17368_), .Y(new_n17369_));
  OR2X1    g14933(.A(new_n17302_), .B(new_n12622_), .Y(new_n17370_));
  OAI22X1  g14934(.A0(new_n17370_), .A1(new_n17369_), .B0(new_n17367_), .B1(new_n17366_), .Y(new_n17371_));
  MX2X1    g14935(.A(new_n17371_), .B(new_n17364_), .S0(new_n11887_), .Y(new_n17372_));
  NAND2X1  g14936(.A(new_n17372_), .B(new_n12637_), .Y(new_n17373_));
  AOI21X1  g14937(.A0(new_n17271_), .A1(pi0619), .B0(pi1159), .Y(new_n17374_));
  OR2X1    g14938(.A(new_n17306_), .B(pi0648), .Y(new_n17375_));
  AOI21X1  g14939(.A0(new_n17374_), .A1(new_n17373_), .B0(new_n17375_), .Y(new_n17376_));
  NAND2X1  g14940(.A(new_n17372_), .B(pi0619), .Y(new_n17377_));
  AOI21X1  g14941(.A0(new_n17271_), .A1(new_n12637_), .B0(new_n12638_), .Y(new_n17378_));
  OR2X1    g14942(.A(new_n17308_), .B(new_n12645_), .Y(new_n17379_));
  AOI21X1  g14943(.A0(new_n17378_), .A1(new_n17377_), .B0(new_n17379_), .Y(new_n17380_));
  NOR3X1   g14944(.A(new_n17380_), .B(new_n17376_), .C(new_n11886_), .Y(new_n17381_));
  OAI21X1  g14945(.A0(new_n17372_), .A1(pi0789), .B0(new_n12842_), .Y(new_n17382_));
  AOI21X1  g14946(.A0(new_n17254_), .A1(pi0626), .B0(new_n16352_), .Y(new_n17383_));
  OAI21X1  g14947(.A0(new_n17310_), .A1(pi0626), .B0(new_n17383_), .Y(new_n17384_));
  AOI21X1  g14948(.A0(new_n17254_), .A1(new_n12664_), .B0(new_n16356_), .Y(new_n17385_));
  OAI21X1  g14949(.A0(new_n17310_), .A1(new_n12664_), .B0(new_n17385_), .Y(new_n17386_));
  NAND2X1  g14950(.A(new_n17272_), .B(new_n12769_), .Y(new_n17387_));
  NAND3X1  g14951(.A(new_n17387_), .B(new_n17386_), .C(new_n17384_), .Y(new_n17388_));
  AOI21X1  g14952(.A0(new_n17388_), .A1(pi0788), .B0(new_n14273_), .Y(new_n17389_));
  OAI21X1  g14953(.A0(new_n17382_), .A1(new_n17381_), .B0(new_n17389_), .Y(new_n17390_));
  AOI21X1  g14954(.A0(new_n17390_), .A1(new_n17327_), .B0(new_n14269_), .Y(new_n17391_));
  OR2X1    g14955(.A(new_n17312_), .B(new_n14384_), .Y(new_n17392_));
  OR2X1    g14956(.A(new_n17281_), .B(new_n14389_), .Y(new_n17393_));
  OR2X1    g14957(.A(new_n17282_), .B(new_n14387_), .Y(new_n17394_));
  NAND3X1  g14958(.A(new_n17394_), .B(new_n17393_), .C(new_n17392_), .Y(new_n17395_));
  AND2X1   g14959(.A(new_n17395_), .B(pi0787), .Y(new_n17396_));
  NOR3X1   g14960(.A(new_n17396_), .B(new_n17391_), .C(new_n17324_), .Y(new_n17397_));
  AOI21X1  g14961(.A0(new_n17321_), .A1(pi0790), .B0(new_n17397_), .Y(new_n17398_));
  OR2X1    g14962(.A(new_n17398_), .B(po1038), .Y(new_n17399_));
  AOI21X1  g14963(.A0(po1038), .A1(new_n10020_), .B0(pi0832), .Y(new_n17400_));
  AOI22X1  g14964(.A0(new_n17400_), .A1(new_n17399_), .B0(new_n17251_), .B1(new_n17250_), .Y(po0335));
  OAI21X1  g14965(.A0(new_n12202_), .A1(pi0179), .B0(new_n12935_), .Y(new_n17402_));
  OAI21X1  g14966(.A0(new_n12349_), .A1(new_n10461_), .B0(pi0039), .Y(new_n17403_));
  AOI21X1  g14967(.A0(new_n12289_), .A1(new_n10461_), .B0(new_n17403_), .Y(new_n17404_));
  OAI21X1  g14968(.A0(new_n12467_), .A1(new_n10461_), .B0(new_n2959_), .Y(new_n17405_));
  AOI21X1  g14969(.A0(new_n12454_), .A1(new_n10461_), .B0(new_n17405_), .Y(new_n17406_));
  OAI21X1  g14970(.A0(new_n17406_), .A1(new_n17404_), .B0(new_n2996_), .Y(new_n17407_));
  AOI21X1  g14971(.A0(new_n17407_), .A1(new_n17402_), .B0(new_n15091_), .Y(new_n17408_));
  OAI21X1  g14972(.A0(new_n13694_), .A1(pi0179), .B0(new_n15091_), .Y(new_n17409_));
  AOI21X1  g14973(.A0(new_n13688_), .A1(pi0179), .B0(new_n17409_), .Y(new_n17410_));
  NOR3X1   g14974(.A(new_n17410_), .B(new_n17408_), .C(pi0724), .Y(new_n17411_));
  AOI21X1  g14975(.A0(new_n16746_), .A1(new_n15091_), .B0(new_n10461_), .Y(new_n17412_));
  NOR3X1   g14976(.A(new_n13701_), .B(pi0741), .C(pi0179), .Y(new_n17413_));
  AOI21X1  g14977(.A0(new_n17413_), .A1(new_n13704_), .B0(new_n17412_), .Y(new_n17414_));
  OAI21X1  g14978(.A0(new_n12574_), .A1(new_n15091_), .B0(new_n17414_), .Y(new_n17415_));
  OAI21X1  g14979(.A0(new_n17415_), .A1(new_n15092_), .B0(new_n3129_), .Y(new_n17416_));
  OAI22X1  g14980(.A0(new_n17416_), .A1(new_n17411_), .B0(new_n3129_), .B1(new_n10461_), .Y(new_n17417_));
  NOR2X1   g14981(.A(new_n3129_), .B(new_n10461_), .Y(new_n17418_));
  AOI21X1  g14982(.A0(new_n17415_), .A1(new_n3129_), .B0(new_n17418_), .Y(new_n17419_));
  AOI21X1  g14983(.A0(new_n17419_), .A1(pi0625), .B0(pi1153), .Y(new_n17420_));
  OAI21X1  g14984(.A0(new_n17417_), .A1(pi0625), .B0(new_n17420_), .Y(new_n17421_));
  AOI21X1  g14985(.A0(new_n13699_), .A1(new_n3129_), .B0(pi0179), .Y(new_n17422_));
  OAI21X1  g14986(.A0(new_n3810_), .A1(pi0724), .B0(new_n17422_), .Y(new_n17423_));
  AOI21X1  g14987(.A0(new_n12955_), .A1(pi0179), .B0(pi0038), .Y(new_n17424_));
  OAI22X1  g14988(.A0(new_n17424_), .A1(new_n3810_), .B0(new_n12953_), .B1(pi0179), .Y(new_n17425_));
  OAI21X1  g14989(.A0(new_n12202_), .A1(pi0179), .B0(new_n12567_), .Y(new_n17426_));
  NAND3X1  g14990(.A(new_n17426_), .B(new_n17425_), .C(new_n15092_), .Y(new_n17427_));
  AOI21X1  g14991(.A0(new_n17427_), .A1(new_n17423_), .B0(new_n12493_), .Y(new_n17428_));
  OAI21X1  g14992(.A0(new_n12574_), .A1(new_n3810_), .B0(new_n10461_), .Y(new_n17429_));
  OAI21X1  g14993(.A0(new_n17429_), .A1(pi0625), .B0(pi1153), .Y(new_n17430_));
  OR2X1    g14994(.A(new_n17430_), .B(new_n17428_), .Y(new_n17431_));
  NAND3X1  g14995(.A(new_n17431_), .B(new_n17421_), .C(new_n12584_), .Y(new_n17432_));
  AOI21X1  g14996(.A0(new_n17419_), .A1(new_n12493_), .B0(new_n12494_), .Y(new_n17433_));
  OAI21X1  g14997(.A0(new_n17417_), .A1(new_n12493_), .B0(new_n17433_), .Y(new_n17434_));
  AOI21X1  g14998(.A0(new_n17427_), .A1(new_n17423_), .B0(pi0625), .Y(new_n17435_));
  OAI21X1  g14999(.A0(new_n17429_), .A1(new_n12493_), .B0(new_n12494_), .Y(new_n17436_));
  OR2X1    g15000(.A(new_n17436_), .B(new_n17435_), .Y(new_n17437_));
  NAND3X1  g15001(.A(new_n17437_), .B(new_n17434_), .C(pi0608), .Y(new_n17438_));
  AOI21X1  g15002(.A0(new_n17438_), .A1(new_n17432_), .B0(new_n11889_), .Y(new_n17439_));
  NOR2X1   g15003(.A(new_n17417_), .B(pi0778), .Y(new_n17440_));
  OR2X1    g15004(.A(new_n17440_), .B(new_n17439_), .Y(new_n17441_));
  AND2X1   g15005(.A(new_n17427_), .B(new_n17423_), .Y(new_n17442_));
  OAI22X1  g15006(.A0(new_n17436_), .A1(new_n17435_), .B0(new_n17430_), .B1(new_n17428_), .Y(new_n17443_));
  MX2X1    g15007(.A(new_n17443_), .B(new_n17442_), .S0(new_n11889_), .Y(new_n17444_));
  OAI21X1  g15008(.A0(new_n17444_), .A1(new_n12590_), .B0(new_n12591_), .Y(new_n17445_));
  AOI21X1  g15009(.A0(new_n17441_), .A1(new_n12590_), .B0(new_n17445_), .Y(new_n17446_));
  NOR2X1   g15010(.A(new_n17419_), .B(new_n12601_), .Y(new_n17447_));
  AOI22X1  g15011(.A0(new_n17447_), .A1(pi0609), .B0(new_n17429_), .B1(new_n13430_), .Y(new_n17448_));
  OAI21X1  g15012(.A0(new_n17448_), .A1(new_n12591_), .B0(new_n12596_), .Y(new_n17449_));
  OAI21X1  g15013(.A0(new_n17444_), .A1(pi0609), .B0(pi1155), .Y(new_n17450_));
  AOI21X1  g15014(.A0(new_n17441_), .A1(pi0609), .B0(new_n17450_), .Y(new_n17451_));
  AOI22X1  g15015(.A0(new_n17447_), .A1(new_n12590_), .B0(new_n17429_), .B1(new_n13436_), .Y(new_n17452_));
  OAI21X1  g15016(.A0(new_n17452_), .A1(pi1155), .B0(pi0660), .Y(new_n17453_));
  OAI22X1  g15017(.A0(new_n17453_), .A1(new_n17451_), .B0(new_n17449_), .B1(new_n17446_), .Y(new_n17454_));
  MX2X1    g15018(.A(new_n17454_), .B(new_n17441_), .S0(new_n11888_), .Y(new_n17455_));
  MX2X1    g15019(.A(new_n17444_), .B(new_n17429_), .S0(new_n12618_), .Y(new_n17456_));
  OAI21X1  g15020(.A0(new_n17456_), .A1(new_n12614_), .B0(new_n12615_), .Y(new_n17457_));
  AOI21X1  g15021(.A0(new_n17455_), .A1(new_n12614_), .B0(new_n17457_), .Y(new_n17458_));
  MX2X1    g15022(.A(new_n17422_), .B(new_n17419_), .S0(new_n12623_), .Y(new_n17459_));
  MX2X1    g15023(.A(new_n17452_), .B(new_n17448_), .S0(pi1155), .Y(new_n17460_));
  MX2X1    g15024(.A(new_n17460_), .B(new_n17459_), .S0(new_n11888_), .Y(new_n17461_));
  OAI21X1  g15025(.A0(new_n17429_), .A1(pi0618), .B0(pi1154), .Y(new_n17462_));
  AOI21X1  g15026(.A0(new_n17461_), .A1(pi0618), .B0(new_n17462_), .Y(new_n17463_));
  OR2X1    g15027(.A(new_n17463_), .B(pi0627), .Y(new_n17464_));
  OAI21X1  g15028(.A0(new_n17456_), .A1(pi0618), .B0(pi1154), .Y(new_n17465_));
  AOI21X1  g15029(.A0(new_n17455_), .A1(pi0618), .B0(new_n17465_), .Y(new_n17466_));
  OAI21X1  g15030(.A0(new_n17429_), .A1(new_n12614_), .B0(new_n12615_), .Y(new_n17467_));
  AOI21X1  g15031(.A0(new_n17461_), .A1(new_n12614_), .B0(new_n17467_), .Y(new_n17468_));
  OR2X1    g15032(.A(new_n17468_), .B(new_n12622_), .Y(new_n17469_));
  OAI22X1  g15033(.A0(new_n17469_), .A1(new_n17466_), .B0(new_n17464_), .B1(new_n17458_), .Y(new_n17470_));
  MX2X1    g15034(.A(new_n17470_), .B(new_n17455_), .S0(new_n11887_), .Y(new_n17471_));
  MX2X1    g15035(.A(new_n17456_), .B(new_n17429_), .S0(new_n12641_), .Y(new_n17472_));
  OAI21X1  g15036(.A0(new_n17472_), .A1(new_n12637_), .B0(new_n12638_), .Y(new_n17473_));
  AOI21X1  g15037(.A0(new_n17471_), .A1(new_n12637_), .B0(new_n17473_), .Y(new_n17474_));
  OR2X1    g15038(.A(new_n17461_), .B(pi0781), .Y(new_n17475_));
  OAI21X1  g15039(.A0(new_n17468_), .A1(new_n17463_), .B0(pi0781), .Y(new_n17476_));
  NAND2X1  g15040(.A(new_n17476_), .B(new_n17475_), .Y(new_n17477_));
  AOI21X1  g15041(.A0(new_n17422_), .A1(new_n12637_), .B0(new_n12638_), .Y(new_n17478_));
  OAI21X1  g15042(.A0(new_n17477_), .A1(new_n12637_), .B0(new_n17478_), .Y(new_n17479_));
  NAND2X1  g15043(.A(new_n17479_), .B(new_n12645_), .Y(new_n17480_));
  OAI21X1  g15044(.A0(new_n17472_), .A1(pi0619), .B0(pi1159), .Y(new_n17481_));
  AOI21X1  g15045(.A0(new_n17471_), .A1(pi0619), .B0(new_n17481_), .Y(new_n17482_));
  AOI21X1  g15046(.A0(new_n17422_), .A1(pi0619), .B0(pi1159), .Y(new_n17483_));
  OAI21X1  g15047(.A0(new_n17477_), .A1(pi0619), .B0(new_n17483_), .Y(new_n17484_));
  NAND2X1  g15048(.A(new_n17484_), .B(pi0648), .Y(new_n17485_));
  OAI22X1  g15049(.A0(new_n17485_), .A1(new_n17482_), .B0(new_n17480_), .B1(new_n17474_), .Y(new_n17486_));
  MX2X1    g15050(.A(new_n17486_), .B(new_n17471_), .S0(new_n11886_), .Y(new_n17487_));
  OR2X1    g15051(.A(new_n17487_), .B(pi0788), .Y(new_n17488_));
  MX2X1    g15052(.A(new_n17472_), .B(new_n17429_), .S0(new_n12659_), .Y(new_n17489_));
  AOI21X1  g15053(.A0(new_n17489_), .A1(pi0626), .B0(pi0641), .Y(new_n17490_));
  OAI21X1  g15054(.A0(new_n17487_), .A1(pi0626), .B0(new_n17490_), .Y(new_n17491_));
  AOI21X1  g15055(.A0(new_n17484_), .A1(new_n17479_), .B0(new_n11886_), .Y(new_n17492_));
  AOI21X1  g15056(.A0(new_n17477_), .A1(new_n11886_), .B0(new_n17492_), .Y(new_n17493_));
  AOI21X1  g15057(.A0(new_n17429_), .A1(pi0626), .B0(new_n12672_), .Y(new_n17494_));
  OAI21X1  g15058(.A0(new_n17493_), .A1(pi0626), .B0(new_n17494_), .Y(new_n17495_));
  AND2X1   g15059(.A(new_n17495_), .B(new_n12676_), .Y(new_n17496_));
  AOI21X1  g15060(.A0(new_n17489_), .A1(new_n12664_), .B0(new_n12672_), .Y(new_n17497_));
  OAI21X1  g15061(.A0(new_n17487_), .A1(new_n12664_), .B0(new_n17497_), .Y(new_n17498_));
  AOI21X1  g15062(.A0(new_n17429_), .A1(new_n12664_), .B0(pi0641), .Y(new_n17499_));
  OAI21X1  g15063(.A0(new_n17493_), .A1(new_n12664_), .B0(new_n17499_), .Y(new_n17500_));
  AND2X1   g15064(.A(new_n17500_), .B(pi1158), .Y(new_n17501_));
  AOI22X1  g15065(.A0(new_n17501_), .A1(new_n17498_), .B0(new_n17496_), .B1(new_n17491_), .Y(new_n17502_));
  OAI21X1  g15066(.A0(new_n17502_), .A1(new_n11885_), .B0(new_n17488_), .Y(new_n17503_));
  MX2X1    g15067(.A(new_n17493_), .B(new_n17422_), .S0(new_n12841_), .Y(new_n17504_));
  AOI21X1  g15068(.A0(new_n17504_), .A1(pi0628), .B0(pi1156), .Y(new_n17505_));
  OAI21X1  g15069(.A0(new_n17503_), .A1(pi0628), .B0(new_n17505_), .Y(new_n17506_));
  MX2X1    g15070(.A(new_n17489_), .B(new_n17429_), .S0(new_n12691_), .Y(new_n17507_));
  AOI21X1  g15071(.A0(new_n17422_), .A1(new_n12683_), .B0(new_n12684_), .Y(new_n17508_));
  OAI21X1  g15072(.A0(new_n17507_), .A1(new_n12683_), .B0(new_n17508_), .Y(new_n17509_));
  AND2X1   g15073(.A(new_n17509_), .B(new_n12689_), .Y(new_n17510_));
  AOI21X1  g15074(.A0(new_n17504_), .A1(new_n12683_), .B0(new_n12684_), .Y(new_n17511_));
  OAI21X1  g15075(.A0(new_n17503_), .A1(new_n12683_), .B0(new_n17511_), .Y(new_n17512_));
  AOI21X1  g15076(.A0(new_n17422_), .A1(pi0628), .B0(pi1156), .Y(new_n17513_));
  OAI21X1  g15077(.A0(new_n17507_), .A1(pi0628), .B0(new_n17513_), .Y(new_n17514_));
  AND2X1   g15078(.A(new_n17514_), .B(pi0629), .Y(new_n17515_));
  AOI22X1  g15079(.A0(new_n17515_), .A1(new_n17512_), .B0(new_n17510_), .B1(new_n17506_), .Y(new_n17516_));
  MX2X1    g15080(.A(new_n17516_), .B(new_n17503_), .S0(new_n11884_), .Y(new_n17517_));
  MX2X1    g15081(.A(new_n17504_), .B(new_n17422_), .S0(new_n12711_), .Y(new_n17518_));
  AOI21X1  g15082(.A0(new_n17518_), .A1(pi0647), .B0(pi1157), .Y(new_n17519_));
  OAI21X1  g15083(.A0(new_n17517_), .A1(pi0647), .B0(new_n17519_), .Y(new_n17520_));
  AOI21X1  g15084(.A0(new_n17514_), .A1(new_n17509_), .B0(new_n11884_), .Y(new_n17521_));
  AOI21X1  g15085(.A0(new_n17507_), .A1(new_n11884_), .B0(new_n17521_), .Y(new_n17522_));
  INVX1    g15086(.A(new_n17522_), .Y(new_n17523_));
  AOI21X1  g15087(.A0(new_n17422_), .A1(new_n12705_), .B0(new_n12706_), .Y(new_n17524_));
  OAI21X1  g15088(.A0(new_n17523_), .A1(new_n12705_), .B0(new_n17524_), .Y(new_n17525_));
  AND2X1   g15089(.A(new_n17525_), .B(new_n12723_), .Y(new_n17526_));
  AOI21X1  g15090(.A0(new_n17518_), .A1(new_n12705_), .B0(new_n12706_), .Y(new_n17527_));
  OAI21X1  g15091(.A0(new_n17517_), .A1(new_n12705_), .B0(new_n17527_), .Y(new_n17528_));
  AOI21X1  g15092(.A0(new_n17422_), .A1(pi0647), .B0(pi1157), .Y(new_n17529_));
  OAI21X1  g15093(.A0(new_n17523_), .A1(pi0647), .B0(new_n17529_), .Y(new_n17530_));
  AND2X1   g15094(.A(new_n17530_), .B(pi0630), .Y(new_n17531_));
  AOI22X1  g15095(.A0(new_n17531_), .A1(new_n17528_), .B0(new_n17526_), .B1(new_n17520_), .Y(new_n17532_));
  OR2X1    g15096(.A(new_n17517_), .B(pi0787), .Y(new_n17533_));
  OAI21X1  g15097(.A0(new_n17532_), .A1(new_n11883_), .B0(new_n17533_), .Y(new_n17534_));
  NAND2X1  g15098(.A(new_n17530_), .B(new_n17525_), .Y(new_n17535_));
  MX2X1    g15099(.A(new_n17535_), .B(new_n17523_), .S0(new_n11883_), .Y(new_n17536_));
  OAI21X1  g15100(.A0(new_n17536_), .A1(pi0644), .B0(pi0715), .Y(new_n17537_));
  AOI21X1  g15101(.A0(new_n17534_), .A1(pi0644), .B0(new_n17537_), .Y(new_n17538_));
  MX2X1    g15102(.A(new_n17518_), .B(new_n17422_), .S0(new_n12735_), .Y(new_n17539_));
  OAI21X1  g15103(.A0(new_n17429_), .A1(pi0644), .B0(new_n12739_), .Y(new_n17540_));
  AOI21X1  g15104(.A0(new_n17539_), .A1(pi0644), .B0(new_n17540_), .Y(new_n17541_));
  NOR3X1   g15105(.A(new_n17541_), .B(new_n17538_), .C(new_n11882_), .Y(new_n17542_));
  OAI21X1  g15106(.A0(new_n17536_), .A1(new_n12743_), .B0(new_n12739_), .Y(new_n17543_));
  AOI21X1  g15107(.A0(new_n17534_), .A1(new_n12743_), .B0(new_n17543_), .Y(new_n17544_));
  OAI21X1  g15108(.A0(new_n17429_), .A1(new_n12743_), .B0(pi0715), .Y(new_n17545_));
  AOI21X1  g15109(.A0(new_n17539_), .A1(new_n12743_), .B0(new_n17545_), .Y(new_n17546_));
  OR2X1    g15110(.A(new_n17546_), .B(pi1160), .Y(new_n17547_));
  OAI21X1  g15111(.A0(new_n17547_), .A1(new_n17544_), .B0(pi0790), .Y(new_n17548_));
  MX2X1    g15112(.A(new_n17532_), .B(new_n17517_), .S0(new_n11883_), .Y(new_n17549_));
  AOI21X1  g15113(.A0(new_n17549_), .A1(new_n12897_), .B0(po1038), .Y(new_n17550_));
  OAI21X1  g15114(.A0(new_n17548_), .A1(new_n17542_), .B0(new_n17550_), .Y(new_n17551_));
  AOI21X1  g15115(.A0(po1038), .A1(new_n10461_), .B0(pi0832), .Y(new_n17552_));
  AOI21X1  g15116(.A0(pi1093), .A1(pi1092), .B0(pi0179), .Y(new_n17553_));
  INVX1    g15117(.A(new_n17553_), .Y(new_n17554_));
  AOI21X1  g15118(.A0(new_n12178_), .A1(new_n15091_), .B0(new_n17553_), .Y(new_n17555_));
  AOI21X1  g15119(.A0(new_n12601_), .A1(new_n2739_), .B0(new_n17555_), .Y(new_n17556_));
  INVX1    g15120(.A(new_n17555_), .Y(new_n17557_));
  AOI21X1  g15121(.A0(new_n17557_), .A1(new_n12776_), .B0(new_n12591_), .Y(new_n17558_));
  AOI21X1  g15122(.A0(new_n17556_), .A1(new_n12779_), .B0(pi1155), .Y(new_n17559_));
  OAI21X1  g15123(.A0(new_n17559_), .A1(new_n17558_), .B0(pi0785), .Y(new_n17560_));
  OAI21X1  g15124(.A0(new_n17556_), .A1(pi0785), .B0(new_n17560_), .Y(new_n17561_));
  INVX1    g15125(.A(new_n17561_), .Y(new_n17562_));
  AOI21X1  g15126(.A0(new_n17562_), .A1(new_n12785_), .B0(new_n12615_), .Y(new_n17563_));
  AOI21X1  g15127(.A0(new_n17562_), .A1(new_n12788_), .B0(pi1154), .Y(new_n17564_));
  OR2X1    g15128(.A(new_n17564_), .B(new_n17563_), .Y(new_n17565_));
  MX2X1    g15129(.A(new_n17565_), .B(new_n17561_), .S0(new_n11887_), .Y(new_n17566_));
  AND2X1   g15130(.A(new_n17566_), .B(new_n11886_), .Y(new_n17567_));
  AOI21X1  g15131(.A0(new_n17553_), .A1(new_n12637_), .B0(new_n12638_), .Y(new_n17568_));
  OAI21X1  g15132(.A0(new_n17566_), .A1(new_n12637_), .B0(new_n17568_), .Y(new_n17569_));
  AOI21X1  g15133(.A0(new_n17553_), .A1(pi0619), .B0(pi1159), .Y(new_n17570_));
  OAI21X1  g15134(.A0(new_n17566_), .A1(pi0619), .B0(new_n17570_), .Y(new_n17571_));
  AOI21X1  g15135(.A0(new_n17571_), .A1(new_n17569_), .B0(new_n11886_), .Y(new_n17572_));
  NOR2X1   g15136(.A(new_n17572_), .B(new_n17567_), .Y(new_n17573_));
  INVX1    g15137(.A(new_n17573_), .Y(new_n17574_));
  MX2X1    g15138(.A(new_n17574_), .B(new_n17554_), .S0(new_n12841_), .Y(new_n17575_));
  MX2X1    g15139(.A(new_n17575_), .B(new_n17554_), .S0(new_n12711_), .Y(new_n17576_));
  AOI21X1  g15140(.A0(new_n12566_), .A1(new_n15092_), .B0(new_n17553_), .Y(new_n17577_));
  AND2X1   g15141(.A(new_n12566_), .B(new_n15092_), .Y(new_n17578_));
  AND2X1   g15142(.A(new_n17578_), .B(new_n12493_), .Y(new_n17579_));
  MX2X1    g15143(.A(new_n17553_), .B(pi0625), .S0(new_n17578_), .Y(new_n17580_));
  NOR2X1   g15144(.A(new_n17553_), .B(pi1153), .Y(new_n17581_));
  INVX1    g15145(.A(new_n17581_), .Y(new_n17582_));
  OAI22X1  g15146(.A0(new_n17582_), .A1(new_n17579_), .B0(new_n17580_), .B1(new_n12494_), .Y(new_n17583_));
  MX2X1    g15147(.A(new_n17583_), .B(new_n17577_), .S0(new_n11889_), .Y(new_n17584_));
  NOR4X1   g15148(.A(new_n17584_), .B(new_n12765_), .C(new_n12764_), .D(new_n12762_), .Y(new_n17585_));
  INVX1    g15149(.A(new_n17585_), .Y(new_n17586_));
  NOR3X1   g15150(.A(new_n17586_), .B(new_n12870_), .C(new_n12851_), .Y(new_n17587_));
  INVX1    g15151(.A(new_n17587_), .Y(new_n17588_));
  AOI21X1  g15152(.A0(new_n17553_), .A1(pi0647), .B0(pi1157), .Y(new_n17589_));
  OAI21X1  g15153(.A0(new_n17588_), .A1(pi0647), .B0(new_n17589_), .Y(new_n17590_));
  MX2X1    g15154(.A(new_n17587_), .B(new_n17553_), .S0(new_n12705_), .Y(new_n17591_));
  OAI22X1  g15155(.A0(new_n17591_), .A1(new_n14387_), .B0(new_n17590_), .B1(new_n12723_), .Y(new_n17592_));
  AOI21X1  g15156(.A0(new_n17576_), .A1(new_n14385_), .B0(new_n17592_), .Y(new_n17593_));
  AOI21X1  g15157(.A0(new_n17554_), .A1(pi0626), .B0(new_n16352_), .Y(new_n17594_));
  OAI21X1  g15158(.A0(new_n17573_), .A1(pi0626), .B0(new_n17594_), .Y(new_n17595_));
  AOI21X1  g15159(.A0(new_n17554_), .A1(new_n12664_), .B0(new_n16356_), .Y(new_n17596_));
  OAI21X1  g15160(.A0(new_n17573_), .A1(new_n12664_), .B0(new_n17596_), .Y(new_n17597_));
  NAND2X1  g15161(.A(new_n17585_), .B(new_n12769_), .Y(new_n17598_));
  NAND3X1  g15162(.A(new_n17598_), .B(new_n17597_), .C(new_n17595_), .Y(new_n17599_));
  AND2X1   g15163(.A(new_n17599_), .B(pi0788), .Y(new_n17600_));
  INVX1    g15164(.A(new_n17600_), .Y(new_n17601_));
  NOR2X1   g15165(.A(new_n17577_), .B(new_n12120_), .Y(new_n17602_));
  NOR2X1   g15166(.A(new_n17602_), .B(new_n17557_), .Y(new_n17603_));
  INVX1    g15167(.A(new_n17603_), .Y(new_n17604_));
  MX2X1    g15168(.A(new_n17557_), .B(new_n12493_), .S0(new_n17602_), .Y(new_n17605_));
  NOR2X1   g15169(.A(new_n17605_), .B(new_n17582_), .Y(new_n17606_));
  OAI21X1  g15170(.A0(new_n17580_), .A1(new_n12494_), .B0(new_n12584_), .Y(new_n17607_));
  NOR3X1   g15171(.A(new_n17577_), .B(new_n12120_), .C(new_n12493_), .Y(new_n17608_));
  NOR3X1   g15172(.A(new_n17608_), .B(new_n17557_), .C(new_n12494_), .Y(new_n17609_));
  OAI21X1  g15173(.A0(new_n17582_), .A1(new_n17579_), .B0(pi0608), .Y(new_n17610_));
  OAI22X1  g15174(.A0(new_n17610_), .A1(new_n17609_), .B0(new_n17607_), .B1(new_n17606_), .Y(new_n17611_));
  MX2X1    g15175(.A(new_n17611_), .B(new_n17604_), .S0(new_n11889_), .Y(new_n17612_));
  OAI21X1  g15176(.A0(new_n17584_), .A1(new_n12590_), .B0(new_n12591_), .Y(new_n17613_));
  AOI21X1  g15177(.A0(new_n17612_), .A1(new_n12590_), .B0(new_n17613_), .Y(new_n17614_));
  NOR3X1   g15178(.A(new_n17614_), .B(new_n17558_), .C(pi0660), .Y(new_n17615_));
  OAI21X1  g15179(.A0(new_n17584_), .A1(pi0609), .B0(pi1155), .Y(new_n17616_));
  AOI21X1  g15180(.A0(new_n17612_), .A1(pi0609), .B0(new_n17616_), .Y(new_n17617_));
  NOR3X1   g15181(.A(new_n17617_), .B(new_n17559_), .C(new_n12596_), .Y(new_n17618_));
  OAI21X1  g15182(.A0(new_n17618_), .A1(new_n17615_), .B0(pi0785), .Y(new_n17619_));
  NAND2X1  g15183(.A(new_n17612_), .B(new_n11888_), .Y(new_n17620_));
  AND2X1   g15184(.A(new_n17620_), .B(new_n17619_), .Y(new_n17621_));
  NOR3X1   g15185(.A(new_n17584_), .B(new_n12762_), .C(new_n12614_), .Y(new_n17622_));
  NOR2X1   g15186(.A(new_n17622_), .B(pi1154), .Y(new_n17623_));
  OAI21X1  g15187(.A0(new_n17621_), .A1(pi0618), .B0(new_n17623_), .Y(new_n17624_));
  NOR2X1   g15188(.A(new_n17563_), .B(pi0627), .Y(new_n17625_));
  NOR3X1   g15189(.A(new_n17584_), .B(new_n12762_), .C(pi0618), .Y(new_n17626_));
  NOR2X1   g15190(.A(new_n17626_), .B(new_n12615_), .Y(new_n17627_));
  OAI21X1  g15191(.A0(new_n17621_), .A1(new_n12614_), .B0(new_n17627_), .Y(new_n17628_));
  NOR2X1   g15192(.A(new_n17564_), .B(new_n12622_), .Y(new_n17629_));
  AOI22X1  g15193(.A0(new_n17629_), .A1(new_n17628_), .B0(new_n17625_), .B1(new_n17624_), .Y(new_n17630_));
  MX2X1    g15194(.A(new_n17630_), .B(new_n17621_), .S0(new_n11887_), .Y(new_n17631_));
  OR4X1    g15195(.A(new_n17584_), .B(new_n12764_), .C(new_n12762_), .D(new_n12637_), .Y(new_n17632_));
  AND2X1   g15196(.A(new_n17632_), .B(new_n12638_), .Y(new_n17633_));
  OAI21X1  g15197(.A0(new_n17631_), .A1(pi0619), .B0(new_n17633_), .Y(new_n17634_));
  AND2X1   g15198(.A(new_n17569_), .B(new_n12645_), .Y(new_n17635_));
  AND2X1   g15199(.A(new_n17635_), .B(new_n17634_), .Y(new_n17636_));
  NOR4X1   g15200(.A(new_n17584_), .B(new_n12764_), .C(new_n12762_), .D(pi0619), .Y(new_n17637_));
  NOR2X1   g15201(.A(new_n17637_), .B(new_n12638_), .Y(new_n17638_));
  OAI21X1  g15202(.A0(new_n17631_), .A1(new_n12637_), .B0(new_n17638_), .Y(new_n17639_));
  AND2X1   g15203(.A(new_n17571_), .B(pi0648), .Y(new_n17640_));
  AOI21X1  g15204(.A0(new_n17640_), .A1(new_n17639_), .B0(new_n11886_), .Y(new_n17641_));
  INVX1    g15205(.A(new_n17641_), .Y(new_n17642_));
  AOI21X1  g15206(.A0(new_n17631_), .A1(new_n11886_), .B0(new_n14264_), .Y(new_n17643_));
  OAI21X1  g15207(.A0(new_n17642_), .A1(new_n17636_), .B0(new_n17643_), .Y(new_n17644_));
  AOI21X1  g15208(.A0(new_n17644_), .A1(new_n17601_), .B0(new_n14273_), .Y(new_n17645_));
  INVX1    g15209(.A(new_n17575_), .Y(new_n17646_));
  AND2X1   g15210(.A(new_n17585_), .B(new_n12852_), .Y(new_n17647_));
  AOI22X1  g15211(.A0(new_n17647_), .A1(new_n14564_), .B0(new_n17646_), .B1(new_n12867_), .Y(new_n17648_));
  AOI22X1  g15212(.A0(new_n17647_), .A1(new_n14566_), .B0(new_n17646_), .B1(new_n12865_), .Y(new_n17649_));
  MX2X1    g15213(.A(new_n17649_), .B(new_n17648_), .S0(new_n12689_), .Y(new_n17650_));
  OAI21X1  g15214(.A0(new_n17650_), .A1(new_n11884_), .B0(new_n14562_), .Y(new_n17651_));
  OAI22X1  g15215(.A0(new_n17651_), .A1(new_n17645_), .B0(new_n17593_), .B1(new_n11883_), .Y(new_n17652_));
  INVX1    g15216(.A(new_n17652_), .Y(new_n17653_));
  OAI21X1  g15217(.A0(new_n17591_), .A1(new_n12706_), .B0(new_n17590_), .Y(new_n17654_));
  MX2X1    g15218(.A(new_n17654_), .B(new_n17588_), .S0(new_n11883_), .Y(new_n17655_));
  OAI21X1  g15219(.A0(new_n17655_), .A1(pi0644), .B0(pi0715), .Y(new_n17656_));
  AOI21X1  g15220(.A0(new_n17653_), .A1(pi0644), .B0(new_n17656_), .Y(new_n17657_));
  OR4X1    g15221(.A(new_n12734_), .B(new_n2739_), .C(new_n11883_), .D(pi0179), .Y(new_n17658_));
  OAI21X1  g15222(.A0(new_n17576_), .A1(new_n12735_), .B0(new_n17658_), .Y(new_n17659_));
  OAI21X1  g15223(.A0(new_n17554_), .A1(pi0644), .B0(new_n12739_), .Y(new_n17660_));
  AOI21X1  g15224(.A0(new_n17659_), .A1(pi0644), .B0(new_n17660_), .Y(new_n17661_));
  OR2X1    g15225(.A(new_n17661_), .B(new_n11882_), .Y(new_n17662_));
  OAI21X1  g15226(.A0(new_n17655_), .A1(new_n12743_), .B0(new_n12739_), .Y(new_n17663_));
  AOI21X1  g15227(.A0(new_n17653_), .A1(new_n12743_), .B0(new_n17663_), .Y(new_n17664_));
  OAI21X1  g15228(.A0(new_n17554_), .A1(new_n12743_), .B0(pi0715), .Y(new_n17665_));
  AOI21X1  g15229(.A0(new_n17659_), .A1(new_n12743_), .B0(new_n17665_), .Y(new_n17666_));
  OR2X1    g15230(.A(new_n17666_), .B(pi1160), .Y(new_n17667_));
  OAI22X1  g15231(.A0(new_n17667_), .A1(new_n17664_), .B0(new_n17662_), .B1(new_n17657_), .Y(new_n17668_));
  OAI21X1  g15232(.A0(new_n17652_), .A1(pi0790), .B0(pi0832), .Y(new_n17669_));
  AOI21X1  g15233(.A0(new_n17668_), .A1(pi0790), .B0(new_n17669_), .Y(new_n17670_));
  AOI21X1  g15234(.A0(new_n17552_), .A1(new_n17551_), .B0(new_n17670_), .Y(po0336));
  AOI21X1  g15235(.A0(pi1093), .A1(pi1092), .B0(pi0180), .Y(new_n17672_));
  INVX1    g15236(.A(new_n17672_), .Y(new_n17673_));
  AOI21X1  g15237(.A0(new_n12178_), .A1(new_n15141_), .B0(new_n17672_), .Y(new_n17674_));
  AOI21X1  g15238(.A0(new_n12601_), .A1(new_n2739_), .B0(new_n17674_), .Y(new_n17675_));
  NAND2X1  g15239(.A(new_n12178_), .B(new_n15141_), .Y(new_n17676_));
  OAI21X1  g15240(.A0(new_n17676_), .A1(new_n13436_), .B0(new_n17675_), .Y(new_n17677_));
  AND2X1   g15241(.A(new_n17677_), .B(pi1155), .Y(new_n17678_));
  NOR2X1   g15242(.A(new_n17676_), .B(new_n13436_), .Y(new_n17679_));
  NOR3X1   g15243(.A(new_n17679_), .B(new_n17672_), .C(pi1155), .Y(new_n17680_));
  OAI21X1  g15244(.A0(new_n17680_), .A1(new_n17678_), .B0(pi0785), .Y(new_n17681_));
  OAI21X1  g15245(.A0(new_n17675_), .A1(pi0785), .B0(new_n17681_), .Y(new_n17682_));
  INVX1    g15246(.A(new_n17682_), .Y(new_n17683_));
  AOI21X1  g15247(.A0(new_n17683_), .A1(new_n12785_), .B0(new_n12615_), .Y(new_n17684_));
  AOI21X1  g15248(.A0(new_n17683_), .A1(new_n12788_), .B0(pi1154), .Y(new_n17685_));
  NOR2X1   g15249(.A(new_n17685_), .B(new_n17684_), .Y(new_n17686_));
  MX2X1    g15250(.A(new_n17686_), .B(new_n17683_), .S0(new_n11887_), .Y(new_n17687_));
  OR2X1    g15251(.A(new_n17687_), .B(pi0789), .Y(new_n17688_));
  AOI21X1  g15252(.A0(new_n17687_), .A1(new_n15910_), .B0(new_n12638_), .Y(new_n17689_));
  AOI21X1  g15253(.A0(new_n17687_), .A1(new_n15912_), .B0(pi1159), .Y(new_n17690_));
  OAI21X1  g15254(.A0(new_n17690_), .A1(new_n17689_), .B0(pi0789), .Y(new_n17691_));
  AND2X1   g15255(.A(new_n17691_), .B(new_n17688_), .Y(new_n17692_));
  INVX1    g15256(.A(new_n17692_), .Y(new_n17693_));
  MX2X1    g15257(.A(new_n17693_), .B(new_n17673_), .S0(new_n12841_), .Y(new_n17694_));
  MX2X1    g15258(.A(new_n17694_), .B(new_n17673_), .S0(new_n12711_), .Y(new_n17695_));
  AOI21X1  g15259(.A0(new_n12566_), .A1(new_n15160_), .B0(new_n17672_), .Y(new_n17696_));
  INVX1    g15260(.A(new_n17696_), .Y(new_n17697_));
  NOR3X1   g15261(.A(new_n13585_), .B(pi0702), .C(pi0625), .Y(new_n17698_));
  OR2X1    g15262(.A(new_n17698_), .B(new_n17696_), .Y(new_n17699_));
  NOR2X1   g15263(.A(new_n17672_), .B(pi1153), .Y(new_n17700_));
  INVX1    g15264(.A(new_n17700_), .Y(new_n17701_));
  OAI21X1  g15265(.A0(new_n17701_), .A1(new_n17698_), .B0(pi0778), .Y(new_n17702_));
  AOI21X1  g15266(.A0(new_n17699_), .A1(pi1153), .B0(new_n17702_), .Y(new_n17703_));
  AOI21X1  g15267(.A0(new_n17697_), .A1(new_n11889_), .B0(new_n17703_), .Y(new_n17704_));
  NOR4X1   g15268(.A(new_n17704_), .B(new_n12765_), .C(new_n12764_), .D(new_n12762_), .Y(new_n17705_));
  INVX1    g15269(.A(new_n17705_), .Y(new_n17706_));
  NOR3X1   g15270(.A(new_n17706_), .B(new_n12870_), .C(new_n12851_), .Y(new_n17707_));
  INVX1    g15271(.A(new_n17707_), .Y(new_n17708_));
  AOI21X1  g15272(.A0(new_n17672_), .A1(pi0647), .B0(pi1157), .Y(new_n17709_));
  OAI21X1  g15273(.A0(new_n17708_), .A1(pi0647), .B0(new_n17709_), .Y(new_n17710_));
  MX2X1    g15274(.A(new_n17707_), .B(new_n17672_), .S0(new_n12705_), .Y(new_n17711_));
  OAI22X1  g15275(.A0(new_n17711_), .A1(new_n14387_), .B0(new_n17710_), .B1(new_n12723_), .Y(new_n17712_));
  AOI21X1  g15276(.A0(new_n17695_), .A1(new_n14385_), .B0(new_n17712_), .Y(new_n17713_));
  NOR2X1   g15277(.A(new_n17713_), .B(new_n11883_), .Y(new_n17714_));
  AOI21X1  g15278(.A0(new_n17673_), .A1(pi0626), .B0(new_n16352_), .Y(new_n17715_));
  OAI21X1  g15279(.A0(new_n17692_), .A1(pi0626), .B0(new_n17715_), .Y(new_n17716_));
  AOI21X1  g15280(.A0(new_n17691_), .A1(new_n17688_), .B0(new_n12664_), .Y(new_n17717_));
  NOR2X1   g15281(.A(new_n17672_), .B(pi0626), .Y(new_n17718_));
  NOR3X1   g15282(.A(new_n17718_), .B(new_n17717_), .C(new_n16356_), .Y(new_n17719_));
  AOI21X1  g15283(.A0(new_n17705_), .A1(new_n12769_), .B0(new_n17719_), .Y(new_n17720_));
  AOI21X1  g15284(.A0(new_n17720_), .A1(new_n17716_), .B0(new_n11885_), .Y(new_n17721_));
  INVX1    g15285(.A(new_n17674_), .Y(new_n17722_));
  AOI21X1  g15286(.A0(new_n17697_), .A1(new_n12171_), .B0(new_n17722_), .Y(new_n17723_));
  NOR3X1   g15287(.A(new_n17696_), .B(new_n12120_), .C(new_n12493_), .Y(new_n17724_));
  OR2X1    g15288(.A(new_n17723_), .B(new_n17724_), .Y(new_n17725_));
  NOR2X1   g15289(.A(new_n17698_), .B(new_n17696_), .Y(new_n17726_));
  OAI21X1  g15290(.A0(new_n17726_), .A1(new_n12494_), .B0(new_n12584_), .Y(new_n17727_));
  AOI21X1  g15291(.A0(new_n17725_), .A1(new_n17700_), .B0(new_n17727_), .Y(new_n17728_));
  NOR3X1   g15292(.A(new_n17724_), .B(new_n17722_), .C(new_n12494_), .Y(new_n17729_));
  OAI21X1  g15293(.A0(new_n17701_), .A1(new_n17698_), .B0(pi0608), .Y(new_n17730_));
  NOR2X1   g15294(.A(new_n17730_), .B(new_n17729_), .Y(new_n17731_));
  OAI21X1  g15295(.A0(new_n17731_), .A1(new_n17728_), .B0(pi0778), .Y(new_n17732_));
  OAI21X1  g15296(.A0(new_n17723_), .A1(pi0778), .B0(new_n17732_), .Y(new_n17733_));
  OAI21X1  g15297(.A0(new_n17704_), .A1(new_n12590_), .B0(new_n12591_), .Y(new_n17734_));
  AOI21X1  g15298(.A0(new_n17733_), .A1(new_n12590_), .B0(new_n17734_), .Y(new_n17735_));
  NOR3X1   g15299(.A(new_n17735_), .B(new_n17678_), .C(pi0660), .Y(new_n17736_));
  OAI21X1  g15300(.A0(new_n17704_), .A1(pi0609), .B0(pi1155), .Y(new_n17737_));
  AOI21X1  g15301(.A0(new_n17733_), .A1(pi0609), .B0(new_n17737_), .Y(new_n17738_));
  NOR3X1   g15302(.A(new_n17738_), .B(new_n17680_), .C(new_n12596_), .Y(new_n17739_));
  OAI21X1  g15303(.A0(new_n17739_), .A1(new_n17736_), .B0(pi0785), .Y(new_n17740_));
  NAND2X1  g15304(.A(new_n17733_), .B(new_n11888_), .Y(new_n17741_));
  AND2X1   g15305(.A(new_n17741_), .B(new_n17740_), .Y(new_n17742_));
  NOR3X1   g15306(.A(new_n17704_), .B(new_n12762_), .C(new_n12614_), .Y(new_n17743_));
  NOR2X1   g15307(.A(new_n17743_), .B(pi1154), .Y(new_n17744_));
  OAI21X1  g15308(.A0(new_n17742_), .A1(pi0618), .B0(new_n17744_), .Y(new_n17745_));
  NOR2X1   g15309(.A(new_n17684_), .B(pi0627), .Y(new_n17746_));
  NOR3X1   g15310(.A(new_n17704_), .B(new_n12762_), .C(pi0618), .Y(new_n17747_));
  NOR2X1   g15311(.A(new_n17747_), .B(new_n12615_), .Y(new_n17748_));
  OAI21X1  g15312(.A0(new_n17742_), .A1(new_n12614_), .B0(new_n17748_), .Y(new_n17749_));
  NOR2X1   g15313(.A(new_n17685_), .B(new_n12622_), .Y(new_n17750_));
  AOI22X1  g15314(.A0(new_n17750_), .A1(new_n17749_), .B0(new_n17746_), .B1(new_n17745_), .Y(new_n17751_));
  MX2X1    g15315(.A(new_n17751_), .B(new_n17742_), .S0(new_n11887_), .Y(new_n17752_));
  OR4X1    g15316(.A(new_n17704_), .B(new_n12764_), .C(new_n12762_), .D(new_n12637_), .Y(new_n17753_));
  AND2X1   g15317(.A(new_n17753_), .B(new_n12638_), .Y(new_n17754_));
  OAI21X1  g15318(.A0(new_n17752_), .A1(pi0619), .B0(new_n17754_), .Y(new_n17755_));
  NOR2X1   g15319(.A(new_n17689_), .B(pi0648), .Y(new_n17756_));
  AND2X1   g15320(.A(new_n17756_), .B(new_n17755_), .Y(new_n17757_));
  INVX1    g15321(.A(new_n17757_), .Y(new_n17758_));
  NOR4X1   g15322(.A(new_n17704_), .B(new_n12764_), .C(new_n12762_), .D(pi0619), .Y(new_n17759_));
  NOR2X1   g15323(.A(new_n17759_), .B(new_n12638_), .Y(new_n17760_));
  OAI21X1  g15324(.A0(new_n17752_), .A1(new_n12637_), .B0(new_n17760_), .Y(new_n17761_));
  NOR2X1   g15325(.A(new_n17690_), .B(new_n12645_), .Y(new_n17762_));
  AOI21X1  g15326(.A0(new_n17762_), .A1(new_n17761_), .B0(new_n11886_), .Y(new_n17763_));
  AOI21X1  g15327(.A0(new_n17752_), .A1(new_n11886_), .B0(new_n14264_), .Y(new_n17764_));
  INVX1    g15328(.A(new_n17764_), .Y(new_n17765_));
  AOI21X1  g15329(.A0(new_n17763_), .A1(new_n17758_), .B0(new_n17765_), .Y(new_n17766_));
  OAI21X1  g15330(.A0(new_n17766_), .A1(new_n17721_), .B0(new_n16350_), .Y(new_n17767_));
  INVX1    g15331(.A(new_n17694_), .Y(new_n17768_));
  AND2X1   g15332(.A(new_n17705_), .B(new_n12852_), .Y(new_n17769_));
  AOI22X1  g15333(.A0(new_n17769_), .A1(new_n14564_), .B0(new_n17768_), .B1(new_n12867_), .Y(new_n17770_));
  AOI22X1  g15334(.A0(new_n17769_), .A1(new_n14566_), .B0(new_n17768_), .B1(new_n12865_), .Y(new_n17771_));
  MX2X1    g15335(.A(new_n17771_), .B(new_n17770_), .S0(new_n12689_), .Y(new_n17772_));
  OAI21X1  g15336(.A0(new_n17772_), .A1(new_n11884_), .B0(new_n14562_), .Y(new_n17773_));
  INVX1    g15337(.A(new_n17773_), .Y(new_n17774_));
  AOI21X1  g15338(.A0(new_n17774_), .A1(new_n17767_), .B0(new_n17714_), .Y(new_n17775_));
  OAI21X1  g15339(.A0(new_n17711_), .A1(new_n12706_), .B0(new_n17710_), .Y(new_n17776_));
  MX2X1    g15340(.A(new_n17776_), .B(new_n17708_), .S0(new_n11883_), .Y(new_n17777_));
  OAI21X1  g15341(.A0(new_n17777_), .A1(pi0644), .B0(pi0715), .Y(new_n17778_));
  AOI21X1  g15342(.A0(new_n17775_), .A1(pi0644), .B0(new_n17778_), .Y(new_n17779_));
  OR4X1    g15343(.A(new_n12734_), .B(new_n2739_), .C(new_n11883_), .D(pi0180), .Y(new_n17780_));
  OAI21X1  g15344(.A0(new_n17695_), .A1(new_n12735_), .B0(new_n17780_), .Y(new_n17781_));
  OAI21X1  g15345(.A0(new_n17673_), .A1(pi0644), .B0(new_n12739_), .Y(new_n17782_));
  AOI21X1  g15346(.A0(new_n17781_), .A1(pi0644), .B0(new_n17782_), .Y(new_n17783_));
  OR2X1    g15347(.A(new_n17783_), .B(new_n11882_), .Y(new_n17784_));
  OAI21X1  g15348(.A0(new_n17777_), .A1(new_n12743_), .B0(new_n12739_), .Y(new_n17785_));
  AOI21X1  g15349(.A0(new_n17775_), .A1(new_n12743_), .B0(new_n17785_), .Y(new_n17786_));
  OAI21X1  g15350(.A0(new_n17673_), .A1(new_n12743_), .B0(pi0715), .Y(new_n17787_));
  AOI21X1  g15351(.A0(new_n17781_), .A1(new_n12743_), .B0(new_n17787_), .Y(new_n17788_));
  OR2X1    g15352(.A(new_n17788_), .B(pi1160), .Y(new_n17789_));
  OAI22X1  g15353(.A0(new_n17789_), .A1(new_n17786_), .B0(new_n17784_), .B1(new_n17779_), .Y(new_n17790_));
  NAND2X1  g15354(.A(new_n17790_), .B(pi0790), .Y(new_n17791_));
  AOI21X1  g15355(.A0(new_n17775_), .A1(new_n12897_), .B0(new_n12898_), .Y(new_n17792_));
  AOI21X1  g15356(.A0(new_n13699_), .A1(new_n3129_), .B0(pi0180), .Y(new_n17793_));
  INVX1    g15357(.A(new_n17793_), .Y(new_n17794_));
  OAI21X1  g15358(.A0(new_n3810_), .A1(pi0702), .B0(new_n17793_), .Y(new_n17795_));
  AOI21X1  g15359(.A0(new_n12955_), .A1(pi0180), .B0(pi0038), .Y(new_n17796_));
  OAI22X1  g15360(.A0(new_n17796_), .A1(new_n3810_), .B0(new_n12953_), .B1(pi0180), .Y(new_n17797_));
  OAI21X1  g15361(.A0(new_n12202_), .A1(pi0180), .B0(new_n12567_), .Y(new_n17798_));
  NAND3X1  g15362(.A(new_n17798_), .B(new_n17797_), .C(new_n15160_), .Y(new_n17799_));
  AND2X1   g15363(.A(new_n17799_), .B(new_n17795_), .Y(new_n17800_));
  INVX1    g15364(.A(new_n17800_), .Y(new_n17801_));
  AOI21X1  g15365(.A0(new_n17793_), .A1(new_n12493_), .B0(new_n12494_), .Y(new_n17802_));
  OAI21X1  g15366(.A0(new_n17800_), .A1(new_n12493_), .B0(new_n17802_), .Y(new_n17803_));
  AOI21X1  g15367(.A0(new_n17793_), .A1(pi0625), .B0(pi1153), .Y(new_n17804_));
  OAI21X1  g15368(.A0(new_n17800_), .A1(pi0625), .B0(new_n17804_), .Y(new_n17805_));
  AND2X1   g15369(.A(new_n17805_), .B(new_n17803_), .Y(new_n17806_));
  MX2X1    g15370(.A(new_n17806_), .B(new_n17801_), .S0(new_n11889_), .Y(new_n17807_));
  MX2X1    g15371(.A(new_n17807_), .B(new_n17793_), .S0(new_n12618_), .Y(new_n17808_));
  INVX1    g15372(.A(new_n17808_), .Y(new_n17809_));
  MX2X1    g15373(.A(new_n17809_), .B(new_n17794_), .S0(new_n12641_), .Y(new_n17810_));
  INVX1    g15374(.A(new_n17810_), .Y(new_n17811_));
  MX2X1    g15375(.A(new_n17811_), .B(new_n17793_), .S0(new_n12659_), .Y(new_n17812_));
  AND2X1   g15376(.A(new_n17793_), .B(new_n12691_), .Y(new_n17813_));
  AOI21X1  g15377(.A0(new_n17812_), .A1(new_n17252_), .B0(new_n17813_), .Y(new_n17814_));
  AOI21X1  g15378(.A0(new_n17793_), .A1(new_n12683_), .B0(new_n12684_), .Y(new_n17815_));
  OAI21X1  g15379(.A0(new_n17814_), .A1(new_n12683_), .B0(new_n17815_), .Y(new_n17816_));
  AOI21X1  g15380(.A0(new_n17793_), .A1(pi0628), .B0(pi1156), .Y(new_n17817_));
  OAI21X1  g15381(.A0(new_n17814_), .A1(pi0628), .B0(new_n17817_), .Y(new_n17818_));
  AOI21X1  g15382(.A0(new_n17818_), .A1(new_n17816_), .B0(new_n11884_), .Y(new_n17819_));
  AOI21X1  g15383(.A0(new_n17814_), .A1(new_n11884_), .B0(new_n17819_), .Y(new_n17820_));
  MX2X1    g15384(.A(new_n17820_), .B(new_n17793_), .S0(pi0647), .Y(new_n17821_));
  MX2X1    g15385(.A(new_n17820_), .B(new_n17793_), .S0(new_n12705_), .Y(new_n17822_));
  MX2X1    g15386(.A(new_n17822_), .B(new_n17821_), .S0(new_n12706_), .Y(new_n17823_));
  MX2X1    g15387(.A(new_n17823_), .B(new_n17820_), .S0(new_n11883_), .Y(new_n17824_));
  AOI21X1  g15388(.A0(new_n17824_), .A1(new_n12743_), .B0(new_n12739_), .Y(new_n17825_));
  OAI22X1  g15389(.A0(new_n12904_), .A1(new_n5225_), .B0(new_n12089_), .B1(new_n15141_), .Y(new_n17826_));
  OR2X1    g15390(.A(pi0753), .B(pi0180), .Y(new_n17827_));
  OAI22X1  g15391(.A0(new_n12168_), .A1(new_n5225_), .B0(new_n11948_), .B1(new_n15141_), .Y(new_n17828_));
  AOI22X1  g15392(.A0(new_n17828_), .A1(new_n2959_), .B0(pi0753), .B1(pi0180), .Y(new_n17829_));
  OAI21X1  g15393(.A0(new_n17827_), .A1(new_n12910_), .B0(new_n17829_), .Y(new_n17830_));
  AOI21X1  g15394(.A0(new_n17826_), .A1(pi0039), .B0(new_n17830_), .Y(new_n17831_));
  AOI21X1  g15395(.A0(new_n12901_), .A1(new_n5225_), .B0(new_n2996_), .Y(new_n17832_));
  OAI21X1  g15396(.A0(new_n14342_), .A1(pi0753), .B0(new_n17832_), .Y(new_n17833_));
  OAI21X1  g15397(.A0(new_n17831_), .A1(pi0038), .B0(new_n17833_), .Y(new_n17834_));
  MX2X1    g15398(.A(new_n17834_), .B(pi0180), .S0(new_n3810_), .Y(new_n17835_));
  AND2X1   g15399(.A(new_n17835_), .B(new_n12623_), .Y(new_n17836_));
  AOI21X1  g15400(.A0(new_n17794_), .A1(new_n12601_), .B0(new_n17836_), .Y(new_n17837_));
  AOI22X1  g15401(.A0(new_n17836_), .A1(pi0609), .B0(new_n17794_), .B1(new_n13430_), .Y(new_n17838_));
  AOI22X1  g15402(.A0(new_n17836_), .A1(new_n12590_), .B0(new_n17794_), .B1(new_n13436_), .Y(new_n17839_));
  MX2X1    g15403(.A(new_n17839_), .B(new_n17838_), .S0(pi1155), .Y(new_n17840_));
  MX2X1    g15404(.A(new_n17840_), .B(new_n17837_), .S0(new_n11888_), .Y(new_n17841_));
  OAI21X1  g15405(.A0(new_n17794_), .A1(pi0618), .B0(pi1154), .Y(new_n17842_));
  AOI21X1  g15406(.A0(new_n17841_), .A1(pi0618), .B0(new_n17842_), .Y(new_n17843_));
  OAI21X1  g15407(.A0(new_n17794_), .A1(new_n12614_), .B0(new_n12615_), .Y(new_n17844_));
  AOI21X1  g15408(.A0(new_n17841_), .A1(new_n12614_), .B0(new_n17844_), .Y(new_n17845_));
  NOR2X1   g15409(.A(new_n17845_), .B(new_n17843_), .Y(new_n17846_));
  MX2X1    g15410(.A(new_n17846_), .B(new_n17841_), .S0(new_n11887_), .Y(new_n17847_));
  OAI21X1  g15411(.A0(new_n17794_), .A1(pi0619), .B0(pi1159), .Y(new_n17848_));
  AOI21X1  g15412(.A0(new_n17847_), .A1(pi0619), .B0(new_n17848_), .Y(new_n17849_));
  OAI21X1  g15413(.A0(new_n17794_), .A1(new_n12637_), .B0(new_n12638_), .Y(new_n17850_));
  AOI21X1  g15414(.A0(new_n17847_), .A1(new_n12637_), .B0(new_n17850_), .Y(new_n17851_));
  NOR2X1   g15415(.A(new_n17851_), .B(new_n17849_), .Y(new_n17852_));
  MX2X1    g15416(.A(new_n17852_), .B(new_n17847_), .S0(new_n11886_), .Y(new_n17853_));
  MX2X1    g15417(.A(new_n17853_), .B(new_n17793_), .S0(new_n12841_), .Y(new_n17854_));
  MX2X1    g15418(.A(new_n17854_), .B(new_n17793_), .S0(new_n12711_), .Y(new_n17855_));
  MX2X1    g15419(.A(new_n17855_), .B(new_n17793_), .S0(new_n12735_), .Y(new_n17856_));
  OAI21X1  g15420(.A0(new_n17794_), .A1(pi0644), .B0(new_n12739_), .Y(new_n17857_));
  AOI21X1  g15421(.A0(new_n17856_), .A1(pi0644), .B0(new_n17857_), .Y(new_n17858_));
  OR2X1    g15422(.A(new_n17858_), .B(new_n11882_), .Y(new_n17859_));
  AOI21X1  g15423(.A0(new_n17824_), .A1(pi0644), .B0(pi0715), .Y(new_n17860_));
  OAI21X1  g15424(.A0(new_n17794_), .A1(new_n12743_), .B0(pi0715), .Y(new_n17861_));
  AOI21X1  g15425(.A0(new_n17856_), .A1(new_n12743_), .B0(new_n17861_), .Y(new_n17862_));
  OR2X1    g15426(.A(new_n17862_), .B(pi1160), .Y(new_n17863_));
  OAI22X1  g15427(.A0(new_n17863_), .A1(new_n17860_), .B0(new_n17859_), .B1(new_n17825_), .Y(new_n17864_));
  NOR3X1   g15428(.A(new_n17862_), .B(pi1160), .C(pi0644), .Y(new_n17865_));
  NOR3X1   g15429(.A(new_n17858_), .B(new_n11882_), .C(new_n12743_), .Y(new_n17866_));
  NOR3X1   g15430(.A(new_n17866_), .B(new_n17865_), .C(new_n12897_), .Y(new_n17867_));
  MX2X1    g15431(.A(new_n17818_), .B(new_n17816_), .S0(new_n12689_), .Y(new_n17868_));
  OAI21X1  g15432(.A0(new_n17854_), .A1(new_n14395_), .B0(new_n17868_), .Y(new_n17869_));
  NAND2X1  g15433(.A(new_n17869_), .B(pi0792), .Y(new_n17870_));
  OR2X1    g15434(.A(new_n17834_), .B(new_n15160_), .Y(new_n17871_));
  OAI21X1  g15435(.A0(new_n12349_), .A1(new_n5225_), .B0(pi0753), .Y(new_n17872_));
  AOI21X1  g15436(.A0(new_n12289_), .A1(new_n5225_), .B0(new_n17872_), .Y(new_n17873_));
  OAI21X1  g15437(.A0(new_n12440_), .A1(pi0180), .B0(new_n15141_), .Y(new_n17874_));
  AOI21X1  g15438(.A0(new_n12401_), .A1(pi0180), .B0(new_n17874_), .Y(new_n17875_));
  OR2X1    g15439(.A(new_n17875_), .B(new_n2959_), .Y(new_n17876_));
  AND2X1   g15440(.A(new_n12467_), .B(pi0180), .Y(new_n17877_));
  OAI21X1  g15441(.A0(new_n12454_), .A1(pi0180), .B0(pi0753), .Y(new_n17878_));
  NOR4X1   g15442(.A(new_n13391_), .B(new_n12908_), .C(new_n12907_), .D(pi0180), .Y(new_n17879_));
  OAI21X1  g15443(.A0(new_n12929_), .A1(new_n5225_), .B0(new_n15141_), .Y(new_n17880_));
  OAI22X1  g15444(.A0(new_n17880_), .A1(new_n17879_), .B0(new_n17878_), .B1(new_n17877_), .Y(new_n17881_));
  AOI21X1  g15445(.A0(new_n17881_), .A1(new_n2959_), .B0(pi0038), .Y(new_n17882_));
  OAI21X1  g15446(.A0(new_n17876_), .A1(new_n17873_), .B0(new_n17882_), .Y(new_n17883_));
  OAI21X1  g15447(.A0(new_n12478_), .A1(pi0753), .B0(new_n13669_), .Y(new_n17884_));
  NAND2X1  g15448(.A(new_n17884_), .B(new_n5225_), .Y(new_n17885_));
  AOI21X1  g15449(.A0(new_n17676_), .A1(new_n14209_), .B0(new_n5225_), .Y(new_n17886_));
  AOI21X1  g15450(.A0(new_n17886_), .A1(new_n6857_), .B0(new_n2996_), .Y(new_n17887_));
  AOI21X1  g15451(.A0(new_n17887_), .A1(new_n17885_), .B0(pi0702), .Y(new_n17888_));
  AOI21X1  g15452(.A0(new_n17888_), .A1(new_n17883_), .B0(new_n3810_), .Y(new_n17889_));
  AOI22X1  g15453(.A0(new_n17889_), .A1(new_n17871_), .B0(new_n3810_), .B1(pi0180), .Y(new_n17890_));
  OAI21X1  g15454(.A0(new_n17835_), .A1(new_n12493_), .B0(new_n12494_), .Y(new_n17891_));
  AOI21X1  g15455(.A0(new_n17890_), .A1(new_n12493_), .B0(new_n17891_), .Y(new_n17892_));
  NAND2X1  g15456(.A(new_n17803_), .B(new_n12584_), .Y(new_n17893_));
  OAI21X1  g15457(.A0(new_n17835_), .A1(pi0625), .B0(pi1153), .Y(new_n17894_));
  AOI21X1  g15458(.A0(new_n17890_), .A1(pi0625), .B0(new_n17894_), .Y(new_n17895_));
  NAND2X1  g15459(.A(new_n17805_), .B(pi0608), .Y(new_n17896_));
  OAI22X1  g15460(.A0(new_n17896_), .A1(new_n17895_), .B0(new_n17893_), .B1(new_n17892_), .Y(new_n17897_));
  MX2X1    g15461(.A(new_n17897_), .B(new_n17890_), .S0(new_n11889_), .Y(new_n17898_));
  INVX1    g15462(.A(new_n17807_), .Y(new_n17899_));
  OAI21X1  g15463(.A0(new_n17899_), .A1(new_n12590_), .B0(new_n12591_), .Y(new_n17900_));
  AOI21X1  g15464(.A0(new_n17898_), .A1(new_n12590_), .B0(new_n17900_), .Y(new_n17901_));
  OAI21X1  g15465(.A0(new_n17838_), .A1(new_n12591_), .B0(new_n12596_), .Y(new_n17902_));
  OAI21X1  g15466(.A0(new_n17899_), .A1(pi0609), .B0(pi1155), .Y(new_n17903_));
  AOI21X1  g15467(.A0(new_n17898_), .A1(pi0609), .B0(new_n17903_), .Y(new_n17904_));
  OAI21X1  g15468(.A0(new_n17839_), .A1(pi1155), .B0(pi0660), .Y(new_n17905_));
  OAI22X1  g15469(.A0(new_n17905_), .A1(new_n17904_), .B0(new_n17902_), .B1(new_n17901_), .Y(new_n17906_));
  MX2X1    g15470(.A(new_n17906_), .B(new_n17898_), .S0(new_n11888_), .Y(new_n17907_));
  OAI21X1  g15471(.A0(new_n17809_), .A1(new_n12614_), .B0(new_n12615_), .Y(new_n17908_));
  AOI21X1  g15472(.A0(new_n17907_), .A1(new_n12614_), .B0(new_n17908_), .Y(new_n17909_));
  OR2X1    g15473(.A(new_n17843_), .B(pi0627), .Y(new_n17910_));
  OAI21X1  g15474(.A0(new_n17809_), .A1(pi0618), .B0(pi1154), .Y(new_n17911_));
  AOI21X1  g15475(.A0(new_n17907_), .A1(pi0618), .B0(new_n17911_), .Y(new_n17912_));
  OR2X1    g15476(.A(new_n17845_), .B(new_n12622_), .Y(new_n17913_));
  OAI22X1  g15477(.A0(new_n17913_), .A1(new_n17912_), .B0(new_n17910_), .B1(new_n17909_), .Y(new_n17914_));
  MX2X1    g15478(.A(new_n17914_), .B(new_n17907_), .S0(new_n11887_), .Y(new_n17915_));
  NAND2X1  g15479(.A(new_n17915_), .B(new_n12637_), .Y(new_n17916_));
  AOI21X1  g15480(.A0(new_n17811_), .A1(pi0619), .B0(pi1159), .Y(new_n17917_));
  OR2X1    g15481(.A(new_n17849_), .B(pi0648), .Y(new_n17918_));
  AOI21X1  g15482(.A0(new_n17917_), .A1(new_n17916_), .B0(new_n17918_), .Y(new_n17919_));
  NAND2X1  g15483(.A(new_n17915_), .B(pi0619), .Y(new_n17920_));
  AOI21X1  g15484(.A0(new_n17811_), .A1(new_n12637_), .B0(new_n12638_), .Y(new_n17921_));
  OR2X1    g15485(.A(new_n17851_), .B(new_n12645_), .Y(new_n17922_));
  AOI21X1  g15486(.A0(new_n17921_), .A1(new_n17920_), .B0(new_n17922_), .Y(new_n17923_));
  NOR3X1   g15487(.A(new_n17923_), .B(new_n17919_), .C(new_n11886_), .Y(new_n17924_));
  OAI21X1  g15488(.A0(new_n17915_), .A1(pi0789), .B0(new_n12842_), .Y(new_n17925_));
  AOI21X1  g15489(.A0(new_n17794_), .A1(pi0626), .B0(new_n16352_), .Y(new_n17926_));
  OAI21X1  g15490(.A0(new_n17853_), .A1(pi0626), .B0(new_n17926_), .Y(new_n17927_));
  AOI21X1  g15491(.A0(new_n17794_), .A1(new_n12664_), .B0(new_n16356_), .Y(new_n17928_));
  OAI21X1  g15492(.A0(new_n17853_), .A1(new_n12664_), .B0(new_n17928_), .Y(new_n17929_));
  NAND2X1  g15493(.A(new_n17812_), .B(new_n12769_), .Y(new_n17930_));
  NAND3X1  g15494(.A(new_n17930_), .B(new_n17929_), .C(new_n17927_), .Y(new_n17931_));
  AOI21X1  g15495(.A0(new_n17931_), .A1(pi0788), .B0(new_n14273_), .Y(new_n17932_));
  OAI21X1  g15496(.A0(new_n17925_), .A1(new_n17924_), .B0(new_n17932_), .Y(new_n17933_));
  AOI21X1  g15497(.A0(new_n17933_), .A1(new_n17870_), .B0(new_n14269_), .Y(new_n17934_));
  OR2X1    g15498(.A(new_n17855_), .B(new_n14384_), .Y(new_n17935_));
  OR2X1    g15499(.A(new_n17821_), .B(new_n14389_), .Y(new_n17936_));
  OR2X1    g15500(.A(new_n17822_), .B(new_n14387_), .Y(new_n17937_));
  NAND3X1  g15501(.A(new_n17937_), .B(new_n17936_), .C(new_n17935_), .Y(new_n17938_));
  AND2X1   g15502(.A(new_n17938_), .B(pi0787), .Y(new_n17939_));
  NOR3X1   g15503(.A(new_n17939_), .B(new_n17934_), .C(new_n17867_), .Y(new_n17940_));
  AOI21X1  g15504(.A0(new_n17864_), .A1(pi0790), .B0(new_n17940_), .Y(new_n17941_));
  OR2X1    g15505(.A(new_n17941_), .B(po1038), .Y(new_n17942_));
  AOI21X1  g15506(.A0(po1038), .A1(new_n5225_), .B0(pi0832), .Y(new_n17943_));
  AOI22X1  g15507(.A0(new_n17943_), .A1(new_n17942_), .B0(new_n17792_), .B1(new_n17791_), .Y(po0337));
  AOI21X1  g15508(.A0(pi1093), .A1(pi1092), .B0(pi0181), .Y(new_n17945_));
  INVX1    g15509(.A(new_n17945_), .Y(new_n17946_));
  AOI21X1  g15510(.A0(new_n12178_), .A1(new_n15172_), .B0(new_n17945_), .Y(new_n17947_));
  AOI21X1  g15511(.A0(new_n12601_), .A1(new_n2739_), .B0(new_n17947_), .Y(new_n17948_));
  NAND2X1  g15512(.A(new_n12178_), .B(new_n15172_), .Y(new_n17949_));
  OAI21X1  g15513(.A0(new_n17949_), .A1(new_n13436_), .B0(new_n17948_), .Y(new_n17950_));
  AND2X1   g15514(.A(new_n17950_), .B(pi1155), .Y(new_n17951_));
  NOR2X1   g15515(.A(new_n17949_), .B(new_n13436_), .Y(new_n17952_));
  NOR3X1   g15516(.A(new_n17952_), .B(new_n17945_), .C(pi1155), .Y(new_n17953_));
  OAI21X1  g15517(.A0(new_n17953_), .A1(new_n17951_), .B0(pi0785), .Y(new_n17954_));
  OAI21X1  g15518(.A0(new_n17948_), .A1(pi0785), .B0(new_n17954_), .Y(new_n17955_));
  INVX1    g15519(.A(new_n17955_), .Y(new_n17956_));
  AOI21X1  g15520(.A0(new_n17956_), .A1(new_n12785_), .B0(new_n12615_), .Y(new_n17957_));
  AOI21X1  g15521(.A0(new_n17956_), .A1(new_n12788_), .B0(pi1154), .Y(new_n17958_));
  NOR2X1   g15522(.A(new_n17958_), .B(new_n17957_), .Y(new_n17959_));
  MX2X1    g15523(.A(new_n17959_), .B(new_n17956_), .S0(new_n11887_), .Y(new_n17960_));
  OR2X1    g15524(.A(new_n17960_), .B(pi0789), .Y(new_n17961_));
  AOI21X1  g15525(.A0(new_n17960_), .A1(new_n15910_), .B0(new_n12638_), .Y(new_n17962_));
  AOI21X1  g15526(.A0(new_n17960_), .A1(new_n15912_), .B0(pi1159), .Y(new_n17963_));
  OAI21X1  g15527(.A0(new_n17963_), .A1(new_n17962_), .B0(pi0789), .Y(new_n17964_));
  AND2X1   g15528(.A(new_n17964_), .B(new_n17961_), .Y(new_n17965_));
  INVX1    g15529(.A(new_n17965_), .Y(new_n17966_));
  MX2X1    g15530(.A(new_n17966_), .B(new_n17946_), .S0(new_n12841_), .Y(new_n17967_));
  MX2X1    g15531(.A(new_n17967_), .B(new_n17946_), .S0(new_n12711_), .Y(new_n17968_));
  AOI21X1  g15532(.A0(new_n12566_), .A1(new_n15191_), .B0(new_n17945_), .Y(new_n17969_));
  INVX1    g15533(.A(new_n17969_), .Y(new_n17970_));
  NOR3X1   g15534(.A(new_n13585_), .B(pi0709), .C(pi0625), .Y(new_n17971_));
  OR2X1    g15535(.A(new_n17971_), .B(new_n17969_), .Y(new_n17972_));
  NOR2X1   g15536(.A(new_n17945_), .B(pi1153), .Y(new_n17973_));
  INVX1    g15537(.A(new_n17973_), .Y(new_n17974_));
  OAI21X1  g15538(.A0(new_n17974_), .A1(new_n17971_), .B0(pi0778), .Y(new_n17975_));
  AOI21X1  g15539(.A0(new_n17972_), .A1(pi1153), .B0(new_n17975_), .Y(new_n17976_));
  AOI21X1  g15540(.A0(new_n17970_), .A1(new_n11889_), .B0(new_n17976_), .Y(new_n17977_));
  NOR4X1   g15541(.A(new_n17977_), .B(new_n12765_), .C(new_n12764_), .D(new_n12762_), .Y(new_n17978_));
  INVX1    g15542(.A(new_n17978_), .Y(new_n17979_));
  NOR3X1   g15543(.A(new_n17979_), .B(new_n12870_), .C(new_n12851_), .Y(new_n17980_));
  INVX1    g15544(.A(new_n17980_), .Y(new_n17981_));
  AOI21X1  g15545(.A0(new_n17945_), .A1(pi0647), .B0(pi1157), .Y(new_n17982_));
  OAI21X1  g15546(.A0(new_n17981_), .A1(pi0647), .B0(new_n17982_), .Y(new_n17983_));
  MX2X1    g15547(.A(new_n17980_), .B(new_n17945_), .S0(new_n12705_), .Y(new_n17984_));
  OAI22X1  g15548(.A0(new_n17984_), .A1(new_n14387_), .B0(new_n17983_), .B1(new_n12723_), .Y(new_n17985_));
  AOI21X1  g15549(.A0(new_n17968_), .A1(new_n14385_), .B0(new_n17985_), .Y(new_n17986_));
  NOR2X1   g15550(.A(new_n17986_), .B(new_n11883_), .Y(new_n17987_));
  AOI21X1  g15551(.A0(new_n17946_), .A1(pi0626), .B0(new_n16352_), .Y(new_n17988_));
  OAI21X1  g15552(.A0(new_n17965_), .A1(pi0626), .B0(new_n17988_), .Y(new_n17989_));
  AOI21X1  g15553(.A0(new_n17964_), .A1(new_n17961_), .B0(new_n12664_), .Y(new_n17990_));
  NOR2X1   g15554(.A(new_n17945_), .B(pi0626), .Y(new_n17991_));
  NOR3X1   g15555(.A(new_n17991_), .B(new_n17990_), .C(new_n16356_), .Y(new_n17992_));
  AOI21X1  g15556(.A0(new_n17978_), .A1(new_n12769_), .B0(new_n17992_), .Y(new_n17993_));
  AOI21X1  g15557(.A0(new_n17993_), .A1(new_n17989_), .B0(new_n11885_), .Y(new_n17994_));
  INVX1    g15558(.A(new_n17947_), .Y(new_n17995_));
  AOI21X1  g15559(.A0(new_n17970_), .A1(new_n12171_), .B0(new_n17995_), .Y(new_n17996_));
  NOR3X1   g15560(.A(new_n17969_), .B(new_n12120_), .C(new_n12493_), .Y(new_n17997_));
  OR2X1    g15561(.A(new_n17996_), .B(new_n17997_), .Y(new_n17998_));
  NOR2X1   g15562(.A(new_n17971_), .B(new_n17969_), .Y(new_n17999_));
  OAI21X1  g15563(.A0(new_n17999_), .A1(new_n12494_), .B0(new_n12584_), .Y(new_n18000_));
  AOI21X1  g15564(.A0(new_n17998_), .A1(new_n17973_), .B0(new_n18000_), .Y(new_n18001_));
  NOR3X1   g15565(.A(new_n17997_), .B(new_n17995_), .C(new_n12494_), .Y(new_n18002_));
  OAI21X1  g15566(.A0(new_n17974_), .A1(new_n17971_), .B0(pi0608), .Y(new_n18003_));
  NOR2X1   g15567(.A(new_n18003_), .B(new_n18002_), .Y(new_n18004_));
  OAI21X1  g15568(.A0(new_n18004_), .A1(new_n18001_), .B0(pi0778), .Y(new_n18005_));
  OAI21X1  g15569(.A0(new_n17996_), .A1(pi0778), .B0(new_n18005_), .Y(new_n18006_));
  OAI21X1  g15570(.A0(new_n17977_), .A1(new_n12590_), .B0(new_n12591_), .Y(new_n18007_));
  AOI21X1  g15571(.A0(new_n18006_), .A1(new_n12590_), .B0(new_n18007_), .Y(new_n18008_));
  NOR3X1   g15572(.A(new_n18008_), .B(new_n17951_), .C(pi0660), .Y(new_n18009_));
  OAI21X1  g15573(.A0(new_n17977_), .A1(pi0609), .B0(pi1155), .Y(new_n18010_));
  AOI21X1  g15574(.A0(new_n18006_), .A1(pi0609), .B0(new_n18010_), .Y(new_n18011_));
  NOR3X1   g15575(.A(new_n18011_), .B(new_n17953_), .C(new_n12596_), .Y(new_n18012_));
  OAI21X1  g15576(.A0(new_n18012_), .A1(new_n18009_), .B0(pi0785), .Y(new_n18013_));
  NAND2X1  g15577(.A(new_n18006_), .B(new_n11888_), .Y(new_n18014_));
  AND2X1   g15578(.A(new_n18014_), .B(new_n18013_), .Y(new_n18015_));
  NOR3X1   g15579(.A(new_n17977_), .B(new_n12762_), .C(new_n12614_), .Y(new_n18016_));
  NOR2X1   g15580(.A(new_n18016_), .B(pi1154), .Y(new_n18017_));
  OAI21X1  g15581(.A0(new_n18015_), .A1(pi0618), .B0(new_n18017_), .Y(new_n18018_));
  NOR2X1   g15582(.A(new_n17957_), .B(pi0627), .Y(new_n18019_));
  NOR3X1   g15583(.A(new_n17977_), .B(new_n12762_), .C(pi0618), .Y(new_n18020_));
  NOR2X1   g15584(.A(new_n18020_), .B(new_n12615_), .Y(new_n18021_));
  OAI21X1  g15585(.A0(new_n18015_), .A1(new_n12614_), .B0(new_n18021_), .Y(new_n18022_));
  NOR2X1   g15586(.A(new_n17958_), .B(new_n12622_), .Y(new_n18023_));
  AOI22X1  g15587(.A0(new_n18023_), .A1(new_n18022_), .B0(new_n18019_), .B1(new_n18018_), .Y(new_n18024_));
  MX2X1    g15588(.A(new_n18024_), .B(new_n18015_), .S0(new_n11887_), .Y(new_n18025_));
  OR4X1    g15589(.A(new_n17977_), .B(new_n12764_), .C(new_n12762_), .D(new_n12637_), .Y(new_n18026_));
  AND2X1   g15590(.A(new_n18026_), .B(new_n12638_), .Y(new_n18027_));
  OAI21X1  g15591(.A0(new_n18025_), .A1(pi0619), .B0(new_n18027_), .Y(new_n18028_));
  NOR2X1   g15592(.A(new_n17962_), .B(pi0648), .Y(new_n18029_));
  AND2X1   g15593(.A(new_n18029_), .B(new_n18028_), .Y(new_n18030_));
  INVX1    g15594(.A(new_n18030_), .Y(new_n18031_));
  NOR4X1   g15595(.A(new_n17977_), .B(new_n12764_), .C(new_n12762_), .D(pi0619), .Y(new_n18032_));
  NOR2X1   g15596(.A(new_n18032_), .B(new_n12638_), .Y(new_n18033_));
  OAI21X1  g15597(.A0(new_n18025_), .A1(new_n12637_), .B0(new_n18033_), .Y(new_n18034_));
  NOR2X1   g15598(.A(new_n17963_), .B(new_n12645_), .Y(new_n18035_));
  AOI21X1  g15599(.A0(new_n18035_), .A1(new_n18034_), .B0(new_n11886_), .Y(new_n18036_));
  AOI21X1  g15600(.A0(new_n18025_), .A1(new_n11886_), .B0(new_n14264_), .Y(new_n18037_));
  INVX1    g15601(.A(new_n18037_), .Y(new_n18038_));
  AOI21X1  g15602(.A0(new_n18036_), .A1(new_n18031_), .B0(new_n18038_), .Y(new_n18039_));
  OAI21X1  g15603(.A0(new_n18039_), .A1(new_n17994_), .B0(new_n16350_), .Y(new_n18040_));
  INVX1    g15604(.A(new_n17967_), .Y(new_n18041_));
  AND2X1   g15605(.A(new_n17978_), .B(new_n12852_), .Y(new_n18042_));
  AOI22X1  g15606(.A0(new_n18042_), .A1(new_n14564_), .B0(new_n18041_), .B1(new_n12867_), .Y(new_n18043_));
  AOI22X1  g15607(.A0(new_n18042_), .A1(new_n14566_), .B0(new_n18041_), .B1(new_n12865_), .Y(new_n18044_));
  MX2X1    g15608(.A(new_n18044_), .B(new_n18043_), .S0(new_n12689_), .Y(new_n18045_));
  OAI21X1  g15609(.A0(new_n18045_), .A1(new_n11884_), .B0(new_n14562_), .Y(new_n18046_));
  INVX1    g15610(.A(new_n18046_), .Y(new_n18047_));
  AOI21X1  g15611(.A0(new_n18047_), .A1(new_n18040_), .B0(new_n17987_), .Y(new_n18048_));
  OAI21X1  g15612(.A0(new_n17984_), .A1(new_n12706_), .B0(new_n17983_), .Y(new_n18049_));
  MX2X1    g15613(.A(new_n18049_), .B(new_n17981_), .S0(new_n11883_), .Y(new_n18050_));
  OAI21X1  g15614(.A0(new_n18050_), .A1(pi0644), .B0(pi0715), .Y(new_n18051_));
  AOI21X1  g15615(.A0(new_n18048_), .A1(pi0644), .B0(new_n18051_), .Y(new_n18052_));
  OR4X1    g15616(.A(new_n12734_), .B(new_n2739_), .C(new_n11883_), .D(pi0181), .Y(new_n18053_));
  OAI21X1  g15617(.A0(new_n17968_), .A1(new_n12735_), .B0(new_n18053_), .Y(new_n18054_));
  OAI21X1  g15618(.A0(new_n17946_), .A1(pi0644), .B0(new_n12739_), .Y(new_n18055_));
  AOI21X1  g15619(.A0(new_n18054_), .A1(pi0644), .B0(new_n18055_), .Y(new_n18056_));
  OR2X1    g15620(.A(new_n18056_), .B(new_n11882_), .Y(new_n18057_));
  OAI21X1  g15621(.A0(new_n18050_), .A1(new_n12743_), .B0(new_n12739_), .Y(new_n18058_));
  AOI21X1  g15622(.A0(new_n18048_), .A1(new_n12743_), .B0(new_n18058_), .Y(new_n18059_));
  OAI21X1  g15623(.A0(new_n17946_), .A1(new_n12743_), .B0(pi0715), .Y(new_n18060_));
  AOI21X1  g15624(.A0(new_n18054_), .A1(new_n12743_), .B0(new_n18060_), .Y(new_n18061_));
  OR2X1    g15625(.A(new_n18061_), .B(pi1160), .Y(new_n18062_));
  OAI22X1  g15626(.A0(new_n18062_), .A1(new_n18059_), .B0(new_n18057_), .B1(new_n18052_), .Y(new_n18063_));
  NAND2X1  g15627(.A(new_n18063_), .B(pi0790), .Y(new_n18064_));
  AOI21X1  g15628(.A0(new_n18048_), .A1(new_n12897_), .B0(new_n12898_), .Y(new_n18065_));
  AOI21X1  g15629(.A0(new_n13699_), .A1(new_n3129_), .B0(pi0181), .Y(new_n18066_));
  INVX1    g15630(.A(new_n18066_), .Y(new_n18067_));
  OAI21X1  g15631(.A0(new_n3810_), .A1(pi0709), .B0(new_n18066_), .Y(new_n18068_));
  AOI21X1  g15632(.A0(new_n12955_), .A1(pi0181), .B0(pi0038), .Y(new_n18069_));
  OAI22X1  g15633(.A0(new_n18069_), .A1(new_n3810_), .B0(new_n12953_), .B1(pi0181), .Y(new_n18070_));
  OAI21X1  g15634(.A0(new_n12202_), .A1(pi0181), .B0(new_n12567_), .Y(new_n18071_));
  NAND3X1  g15635(.A(new_n18071_), .B(new_n18070_), .C(new_n15191_), .Y(new_n18072_));
  AND2X1   g15636(.A(new_n18072_), .B(new_n18068_), .Y(new_n18073_));
  INVX1    g15637(.A(new_n18073_), .Y(new_n18074_));
  AOI21X1  g15638(.A0(new_n18066_), .A1(new_n12493_), .B0(new_n12494_), .Y(new_n18075_));
  OAI21X1  g15639(.A0(new_n18073_), .A1(new_n12493_), .B0(new_n18075_), .Y(new_n18076_));
  AOI21X1  g15640(.A0(new_n18066_), .A1(pi0625), .B0(pi1153), .Y(new_n18077_));
  OAI21X1  g15641(.A0(new_n18073_), .A1(pi0625), .B0(new_n18077_), .Y(new_n18078_));
  AND2X1   g15642(.A(new_n18078_), .B(new_n18076_), .Y(new_n18079_));
  MX2X1    g15643(.A(new_n18079_), .B(new_n18074_), .S0(new_n11889_), .Y(new_n18080_));
  MX2X1    g15644(.A(new_n18080_), .B(new_n18066_), .S0(new_n12618_), .Y(new_n18081_));
  INVX1    g15645(.A(new_n18081_), .Y(new_n18082_));
  MX2X1    g15646(.A(new_n18082_), .B(new_n18067_), .S0(new_n12641_), .Y(new_n18083_));
  INVX1    g15647(.A(new_n18083_), .Y(new_n18084_));
  MX2X1    g15648(.A(new_n18084_), .B(new_n18066_), .S0(new_n12659_), .Y(new_n18085_));
  AND2X1   g15649(.A(new_n18066_), .B(new_n12691_), .Y(new_n18086_));
  AOI21X1  g15650(.A0(new_n18085_), .A1(new_n17252_), .B0(new_n18086_), .Y(new_n18087_));
  AOI21X1  g15651(.A0(new_n18066_), .A1(new_n12683_), .B0(new_n12684_), .Y(new_n18088_));
  OAI21X1  g15652(.A0(new_n18087_), .A1(new_n12683_), .B0(new_n18088_), .Y(new_n18089_));
  AOI21X1  g15653(.A0(new_n18066_), .A1(pi0628), .B0(pi1156), .Y(new_n18090_));
  OAI21X1  g15654(.A0(new_n18087_), .A1(pi0628), .B0(new_n18090_), .Y(new_n18091_));
  AOI21X1  g15655(.A0(new_n18091_), .A1(new_n18089_), .B0(new_n11884_), .Y(new_n18092_));
  AOI21X1  g15656(.A0(new_n18087_), .A1(new_n11884_), .B0(new_n18092_), .Y(new_n18093_));
  MX2X1    g15657(.A(new_n18093_), .B(new_n18066_), .S0(pi0647), .Y(new_n18094_));
  MX2X1    g15658(.A(new_n18093_), .B(new_n18066_), .S0(new_n12705_), .Y(new_n18095_));
  MX2X1    g15659(.A(new_n18095_), .B(new_n18094_), .S0(new_n12706_), .Y(new_n18096_));
  MX2X1    g15660(.A(new_n18096_), .B(new_n18093_), .S0(new_n11883_), .Y(new_n18097_));
  AOI21X1  g15661(.A0(new_n18097_), .A1(new_n12743_), .B0(new_n12739_), .Y(new_n18098_));
  OAI22X1  g15662(.A0(new_n12904_), .A1(new_n5226_), .B0(new_n12089_), .B1(new_n15172_), .Y(new_n18099_));
  OR2X1    g15663(.A(pi0754), .B(pi0181), .Y(new_n18100_));
  OAI22X1  g15664(.A0(new_n12168_), .A1(new_n5226_), .B0(new_n11948_), .B1(new_n15172_), .Y(new_n18101_));
  AOI22X1  g15665(.A0(new_n18101_), .A1(new_n2959_), .B0(pi0754), .B1(pi0181), .Y(new_n18102_));
  OAI21X1  g15666(.A0(new_n18100_), .A1(new_n12910_), .B0(new_n18102_), .Y(new_n18103_));
  AOI21X1  g15667(.A0(new_n18099_), .A1(pi0039), .B0(new_n18103_), .Y(new_n18104_));
  AOI21X1  g15668(.A0(new_n12901_), .A1(new_n5226_), .B0(new_n2996_), .Y(new_n18105_));
  OAI21X1  g15669(.A0(new_n14342_), .A1(pi0754), .B0(new_n18105_), .Y(new_n18106_));
  OAI21X1  g15670(.A0(new_n18104_), .A1(pi0038), .B0(new_n18106_), .Y(new_n18107_));
  MX2X1    g15671(.A(new_n18107_), .B(pi0181), .S0(new_n3810_), .Y(new_n18108_));
  AND2X1   g15672(.A(new_n18108_), .B(new_n12623_), .Y(new_n18109_));
  AOI21X1  g15673(.A0(new_n18067_), .A1(new_n12601_), .B0(new_n18109_), .Y(new_n18110_));
  AOI22X1  g15674(.A0(new_n18109_), .A1(pi0609), .B0(new_n18067_), .B1(new_n13430_), .Y(new_n18111_));
  AOI22X1  g15675(.A0(new_n18109_), .A1(new_n12590_), .B0(new_n18067_), .B1(new_n13436_), .Y(new_n18112_));
  MX2X1    g15676(.A(new_n18112_), .B(new_n18111_), .S0(pi1155), .Y(new_n18113_));
  MX2X1    g15677(.A(new_n18113_), .B(new_n18110_), .S0(new_n11888_), .Y(new_n18114_));
  OAI21X1  g15678(.A0(new_n18067_), .A1(pi0618), .B0(pi1154), .Y(new_n18115_));
  AOI21X1  g15679(.A0(new_n18114_), .A1(pi0618), .B0(new_n18115_), .Y(new_n18116_));
  OAI21X1  g15680(.A0(new_n18067_), .A1(new_n12614_), .B0(new_n12615_), .Y(new_n18117_));
  AOI21X1  g15681(.A0(new_n18114_), .A1(new_n12614_), .B0(new_n18117_), .Y(new_n18118_));
  NOR2X1   g15682(.A(new_n18118_), .B(new_n18116_), .Y(new_n18119_));
  MX2X1    g15683(.A(new_n18119_), .B(new_n18114_), .S0(new_n11887_), .Y(new_n18120_));
  OAI21X1  g15684(.A0(new_n18067_), .A1(pi0619), .B0(pi1159), .Y(new_n18121_));
  AOI21X1  g15685(.A0(new_n18120_), .A1(pi0619), .B0(new_n18121_), .Y(new_n18122_));
  OAI21X1  g15686(.A0(new_n18067_), .A1(new_n12637_), .B0(new_n12638_), .Y(new_n18123_));
  AOI21X1  g15687(.A0(new_n18120_), .A1(new_n12637_), .B0(new_n18123_), .Y(new_n18124_));
  NOR2X1   g15688(.A(new_n18124_), .B(new_n18122_), .Y(new_n18125_));
  MX2X1    g15689(.A(new_n18125_), .B(new_n18120_), .S0(new_n11886_), .Y(new_n18126_));
  MX2X1    g15690(.A(new_n18126_), .B(new_n18066_), .S0(new_n12841_), .Y(new_n18127_));
  MX2X1    g15691(.A(new_n18127_), .B(new_n18066_), .S0(new_n12711_), .Y(new_n18128_));
  MX2X1    g15692(.A(new_n18128_), .B(new_n18066_), .S0(new_n12735_), .Y(new_n18129_));
  OAI21X1  g15693(.A0(new_n18067_), .A1(pi0644), .B0(new_n12739_), .Y(new_n18130_));
  AOI21X1  g15694(.A0(new_n18129_), .A1(pi0644), .B0(new_n18130_), .Y(new_n18131_));
  OR2X1    g15695(.A(new_n18131_), .B(new_n11882_), .Y(new_n18132_));
  AOI21X1  g15696(.A0(new_n18097_), .A1(pi0644), .B0(pi0715), .Y(new_n18133_));
  OAI21X1  g15697(.A0(new_n18067_), .A1(new_n12743_), .B0(pi0715), .Y(new_n18134_));
  AOI21X1  g15698(.A0(new_n18129_), .A1(new_n12743_), .B0(new_n18134_), .Y(new_n18135_));
  OR2X1    g15699(.A(new_n18135_), .B(pi1160), .Y(new_n18136_));
  OAI22X1  g15700(.A0(new_n18136_), .A1(new_n18133_), .B0(new_n18132_), .B1(new_n18098_), .Y(new_n18137_));
  NOR3X1   g15701(.A(new_n18135_), .B(pi1160), .C(pi0644), .Y(new_n18138_));
  NOR3X1   g15702(.A(new_n18131_), .B(new_n11882_), .C(new_n12743_), .Y(new_n18139_));
  NOR3X1   g15703(.A(new_n18139_), .B(new_n18138_), .C(new_n12897_), .Y(new_n18140_));
  MX2X1    g15704(.A(new_n18091_), .B(new_n18089_), .S0(new_n12689_), .Y(new_n18141_));
  OAI21X1  g15705(.A0(new_n18127_), .A1(new_n14395_), .B0(new_n18141_), .Y(new_n18142_));
  NAND2X1  g15706(.A(new_n18142_), .B(pi0792), .Y(new_n18143_));
  OR2X1    g15707(.A(new_n18107_), .B(new_n15191_), .Y(new_n18144_));
  OAI21X1  g15708(.A0(new_n12349_), .A1(new_n5226_), .B0(pi0754), .Y(new_n18145_));
  AOI21X1  g15709(.A0(new_n12289_), .A1(new_n5226_), .B0(new_n18145_), .Y(new_n18146_));
  OAI21X1  g15710(.A0(new_n12440_), .A1(pi0181), .B0(new_n15172_), .Y(new_n18147_));
  AOI21X1  g15711(.A0(new_n12401_), .A1(pi0181), .B0(new_n18147_), .Y(new_n18148_));
  OR2X1    g15712(.A(new_n18148_), .B(new_n2959_), .Y(new_n18149_));
  AND2X1   g15713(.A(new_n12467_), .B(pi0181), .Y(new_n18150_));
  OAI21X1  g15714(.A0(new_n12454_), .A1(pi0181), .B0(pi0754), .Y(new_n18151_));
  NOR4X1   g15715(.A(new_n13391_), .B(new_n12908_), .C(new_n12907_), .D(pi0181), .Y(new_n18152_));
  OAI21X1  g15716(.A0(new_n12929_), .A1(new_n5226_), .B0(new_n15172_), .Y(new_n18153_));
  OAI22X1  g15717(.A0(new_n18153_), .A1(new_n18152_), .B0(new_n18151_), .B1(new_n18150_), .Y(new_n18154_));
  AOI21X1  g15718(.A0(new_n18154_), .A1(new_n2959_), .B0(pi0038), .Y(new_n18155_));
  OAI21X1  g15719(.A0(new_n18149_), .A1(new_n18146_), .B0(new_n18155_), .Y(new_n18156_));
  OAI21X1  g15720(.A0(new_n12478_), .A1(pi0754), .B0(new_n13669_), .Y(new_n18157_));
  NAND2X1  g15721(.A(new_n18157_), .B(new_n5226_), .Y(new_n18158_));
  AOI21X1  g15722(.A0(new_n17949_), .A1(new_n14209_), .B0(new_n5226_), .Y(new_n18159_));
  AOI21X1  g15723(.A0(new_n18159_), .A1(new_n6857_), .B0(new_n2996_), .Y(new_n18160_));
  AOI21X1  g15724(.A0(new_n18160_), .A1(new_n18158_), .B0(pi0709), .Y(new_n18161_));
  AOI21X1  g15725(.A0(new_n18161_), .A1(new_n18156_), .B0(new_n3810_), .Y(new_n18162_));
  AOI22X1  g15726(.A0(new_n18162_), .A1(new_n18144_), .B0(new_n3810_), .B1(pi0181), .Y(new_n18163_));
  OAI21X1  g15727(.A0(new_n18108_), .A1(new_n12493_), .B0(new_n12494_), .Y(new_n18164_));
  AOI21X1  g15728(.A0(new_n18163_), .A1(new_n12493_), .B0(new_n18164_), .Y(new_n18165_));
  NAND2X1  g15729(.A(new_n18076_), .B(new_n12584_), .Y(new_n18166_));
  OAI21X1  g15730(.A0(new_n18108_), .A1(pi0625), .B0(pi1153), .Y(new_n18167_));
  AOI21X1  g15731(.A0(new_n18163_), .A1(pi0625), .B0(new_n18167_), .Y(new_n18168_));
  NAND2X1  g15732(.A(new_n18078_), .B(pi0608), .Y(new_n18169_));
  OAI22X1  g15733(.A0(new_n18169_), .A1(new_n18168_), .B0(new_n18166_), .B1(new_n18165_), .Y(new_n18170_));
  MX2X1    g15734(.A(new_n18170_), .B(new_n18163_), .S0(new_n11889_), .Y(new_n18171_));
  INVX1    g15735(.A(new_n18080_), .Y(new_n18172_));
  OAI21X1  g15736(.A0(new_n18172_), .A1(new_n12590_), .B0(new_n12591_), .Y(new_n18173_));
  AOI21X1  g15737(.A0(new_n18171_), .A1(new_n12590_), .B0(new_n18173_), .Y(new_n18174_));
  OAI21X1  g15738(.A0(new_n18111_), .A1(new_n12591_), .B0(new_n12596_), .Y(new_n18175_));
  OAI21X1  g15739(.A0(new_n18172_), .A1(pi0609), .B0(pi1155), .Y(new_n18176_));
  AOI21X1  g15740(.A0(new_n18171_), .A1(pi0609), .B0(new_n18176_), .Y(new_n18177_));
  OAI21X1  g15741(.A0(new_n18112_), .A1(pi1155), .B0(pi0660), .Y(new_n18178_));
  OAI22X1  g15742(.A0(new_n18178_), .A1(new_n18177_), .B0(new_n18175_), .B1(new_n18174_), .Y(new_n18179_));
  MX2X1    g15743(.A(new_n18179_), .B(new_n18171_), .S0(new_n11888_), .Y(new_n18180_));
  OAI21X1  g15744(.A0(new_n18082_), .A1(new_n12614_), .B0(new_n12615_), .Y(new_n18181_));
  AOI21X1  g15745(.A0(new_n18180_), .A1(new_n12614_), .B0(new_n18181_), .Y(new_n18182_));
  OR2X1    g15746(.A(new_n18116_), .B(pi0627), .Y(new_n18183_));
  OAI21X1  g15747(.A0(new_n18082_), .A1(pi0618), .B0(pi1154), .Y(new_n18184_));
  AOI21X1  g15748(.A0(new_n18180_), .A1(pi0618), .B0(new_n18184_), .Y(new_n18185_));
  OR2X1    g15749(.A(new_n18118_), .B(new_n12622_), .Y(new_n18186_));
  OAI22X1  g15750(.A0(new_n18186_), .A1(new_n18185_), .B0(new_n18183_), .B1(new_n18182_), .Y(new_n18187_));
  MX2X1    g15751(.A(new_n18187_), .B(new_n18180_), .S0(new_n11887_), .Y(new_n18188_));
  NAND2X1  g15752(.A(new_n18188_), .B(new_n12637_), .Y(new_n18189_));
  AOI21X1  g15753(.A0(new_n18084_), .A1(pi0619), .B0(pi1159), .Y(new_n18190_));
  OR2X1    g15754(.A(new_n18122_), .B(pi0648), .Y(new_n18191_));
  AOI21X1  g15755(.A0(new_n18190_), .A1(new_n18189_), .B0(new_n18191_), .Y(new_n18192_));
  NAND2X1  g15756(.A(new_n18188_), .B(pi0619), .Y(new_n18193_));
  AOI21X1  g15757(.A0(new_n18084_), .A1(new_n12637_), .B0(new_n12638_), .Y(new_n18194_));
  OR2X1    g15758(.A(new_n18124_), .B(new_n12645_), .Y(new_n18195_));
  AOI21X1  g15759(.A0(new_n18194_), .A1(new_n18193_), .B0(new_n18195_), .Y(new_n18196_));
  NOR3X1   g15760(.A(new_n18196_), .B(new_n18192_), .C(new_n11886_), .Y(new_n18197_));
  OAI21X1  g15761(.A0(new_n18188_), .A1(pi0789), .B0(new_n12842_), .Y(new_n18198_));
  AOI21X1  g15762(.A0(new_n18067_), .A1(pi0626), .B0(new_n16352_), .Y(new_n18199_));
  OAI21X1  g15763(.A0(new_n18126_), .A1(pi0626), .B0(new_n18199_), .Y(new_n18200_));
  AOI21X1  g15764(.A0(new_n18067_), .A1(new_n12664_), .B0(new_n16356_), .Y(new_n18201_));
  OAI21X1  g15765(.A0(new_n18126_), .A1(new_n12664_), .B0(new_n18201_), .Y(new_n18202_));
  NAND2X1  g15766(.A(new_n18085_), .B(new_n12769_), .Y(new_n18203_));
  NAND3X1  g15767(.A(new_n18203_), .B(new_n18202_), .C(new_n18200_), .Y(new_n18204_));
  AOI21X1  g15768(.A0(new_n18204_), .A1(pi0788), .B0(new_n14273_), .Y(new_n18205_));
  OAI21X1  g15769(.A0(new_n18198_), .A1(new_n18197_), .B0(new_n18205_), .Y(new_n18206_));
  AOI21X1  g15770(.A0(new_n18206_), .A1(new_n18143_), .B0(new_n14269_), .Y(new_n18207_));
  OR2X1    g15771(.A(new_n18128_), .B(new_n14384_), .Y(new_n18208_));
  OR2X1    g15772(.A(new_n18094_), .B(new_n14389_), .Y(new_n18209_));
  OR2X1    g15773(.A(new_n18095_), .B(new_n14387_), .Y(new_n18210_));
  NAND3X1  g15774(.A(new_n18210_), .B(new_n18209_), .C(new_n18208_), .Y(new_n18211_));
  AND2X1   g15775(.A(new_n18211_), .B(pi0787), .Y(new_n18212_));
  NOR3X1   g15776(.A(new_n18212_), .B(new_n18207_), .C(new_n18140_), .Y(new_n18213_));
  AOI21X1  g15777(.A0(new_n18137_), .A1(pi0790), .B0(new_n18213_), .Y(new_n18214_));
  OR2X1    g15778(.A(new_n18214_), .B(po1038), .Y(new_n18215_));
  AOI21X1  g15779(.A0(po1038), .A1(new_n5226_), .B0(pi0832), .Y(new_n18216_));
  AOI22X1  g15780(.A0(new_n18216_), .A1(new_n18215_), .B0(new_n18065_), .B1(new_n18064_), .Y(po0338));
  AOI21X1  g15781(.A0(pi1093), .A1(pi1092), .B0(pi0182), .Y(new_n18218_));
  INVX1    g15782(.A(new_n18218_), .Y(new_n18219_));
  AOI21X1  g15783(.A0(new_n12178_), .A1(new_n15203_), .B0(new_n18218_), .Y(new_n18220_));
  AOI21X1  g15784(.A0(new_n12601_), .A1(new_n2739_), .B0(new_n18220_), .Y(new_n18221_));
  NAND2X1  g15785(.A(new_n12178_), .B(new_n15203_), .Y(new_n18222_));
  OAI21X1  g15786(.A0(new_n18222_), .A1(new_n13436_), .B0(new_n18221_), .Y(new_n18223_));
  AND2X1   g15787(.A(new_n18223_), .B(pi1155), .Y(new_n18224_));
  NOR2X1   g15788(.A(new_n18222_), .B(new_n13436_), .Y(new_n18225_));
  NOR3X1   g15789(.A(new_n18225_), .B(new_n18218_), .C(pi1155), .Y(new_n18226_));
  OAI21X1  g15790(.A0(new_n18226_), .A1(new_n18224_), .B0(pi0785), .Y(new_n18227_));
  OAI21X1  g15791(.A0(new_n18221_), .A1(pi0785), .B0(new_n18227_), .Y(new_n18228_));
  INVX1    g15792(.A(new_n18228_), .Y(new_n18229_));
  AOI21X1  g15793(.A0(new_n18229_), .A1(new_n12785_), .B0(new_n12615_), .Y(new_n18230_));
  AOI21X1  g15794(.A0(new_n18229_), .A1(new_n12788_), .B0(pi1154), .Y(new_n18231_));
  NOR2X1   g15795(.A(new_n18231_), .B(new_n18230_), .Y(new_n18232_));
  MX2X1    g15796(.A(new_n18232_), .B(new_n18229_), .S0(new_n11887_), .Y(new_n18233_));
  OR2X1    g15797(.A(new_n18233_), .B(pi0789), .Y(new_n18234_));
  AOI21X1  g15798(.A0(new_n18233_), .A1(new_n15910_), .B0(new_n12638_), .Y(new_n18235_));
  AOI21X1  g15799(.A0(new_n18233_), .A1(new_n15912_), .B0(pi1159), .Y(new_n18236_));
  OAI21X1  g15800(.A0(new_n18236_), .A1(new_n18235_), .B0(pi0789), .Y(new_n18237_));
  AND2X1   g15801(.A(new_n18237_), .B(new_n18234_), .Y(new_n18238_));
  INVX1    g15802(.A(new_n18238_), .Y(new_n18239_));
  MX2X1    g15803(.A(new_n18239_), .B(new_n18219_), .S0(new_n12841_), .Y(new_n18240_));
  MX2X1    g15804(.A(new_n18240_), .B(new_n18219_), .S0(new_n12711_), .Y(new_n18241_));
  AOI21X1  g15805(.A0(new_n12566_), .A1(new_n15209_), .B0(new_n18218_), .Y(new_n18242_));
  INVX1    g15806(.A(new_n18242_), .Y(new_n18243_));
  NOR3X1   g15807(.A(new_n13585_), .B(pi0734), .C(pi0625), .Y(new_n18244_));
  OR2X1    g15808(.A(new_n18244_), .B(new_n18242_), .Y(new_n18245_));
  NOR2X1   g15809(.A(new_n18218_), .B(pi1153), .Y(new_n18246_));
  INVX1    g15810(.A(new_n18246_), .Y(new_n18247_));
  OAI21X1  g15811(.A0(new_n18247_), .A1(new_n18244_), .B0(pi0778), .Y(new_n18248_));
  AOI21X1  g15812(.A0(new_n18245_), .A1(pi1153), .B0(new_n18248_), .Y(new_n18249_));
  AOI21X1  g15813(.A0(new_n18243_), .A1(new_n11889_), .B0(new_n18249_), .Y(new_n18250_));
  NOR4X1   g15814(.A(new_n18250_), .B(new_n12765_), .C(new_n12764_), .D(new_n12762_), .Y(new_n18251_));
  INVX1    g15815(.A(new_n18251_), .Y(new_n18252_));
  NOR3X1   g15816(.A(new_n18252_), .B(new_n12870_), .C(new_n12851_), .Y(new_n18253_));
  INVX1    g15817(.A(new_n18253_), .Y(new_n18254_));
  AOI21X1  g15818(.A0(new_n18218_), .A1(pi0647), .B0(pi1157), .Y(new_n18255_));
  OAI21X1  g15819(.A0(new_n18254_), .A1(pi0647), .B0(new_n18255_), .Y(new_n18256_));
  MX2X1    g15820(.A(new_n18253_), .B(new_n18218_), .S0(new_n12705_), .Y(new_n18257_));
  OAI22X1  g15821(.A0(new_n18257_), .A1(new_n14387_), .B0(new_n18256_), .B1(new_n12723_), .Y(new_n18258_));
  AOI21X1  g15822(.A0(new_n18241_), .A1(new_n14385_), .B0(new_n18258_), .Y(new_n18259_));
  NOR2X1   g15823(.A(new_n18259_), .B(new_n11883_), .Y(new_n18260_));
  AOI21X1  g15824(.A0(new_n18219_), .A1(pi0626), .B0(new_n16352_), .Y(new_n18261_));
  OAI21X1  g15825(.A0(new_n18238_), .A1(pi0626), .B0(new_n18261_), .Y(new_n18262_));
  AOI21X1  g15826(.A0(new_n18237_), .A1(new_n18234_), .B0(new_n12664_), .Y(new_n18263_));
  NOR2X1   g15827(.A(new_n18218_), .B(pi0626), .Y(new_n18264_));
  NOR3X1   g15828(.A(new_n18264_), .B(new_n18263_), .C(new_n16356_), .Y(new_n18265_));
  AOI21X1  g15829(.A0(new_n18251_), .A1(new_n12769_), .B0(new_n18265_), .Y(new_n18266_));
  AOI21X1  g15830(.A0(new_n18266_), .A1(new_n18262_), .B0(new_n11885_), .Y(new_n18267_));
  INVX1    g15831(.A(new_n18220_), .Y(new_n18268_));
  AOI21X1  g15832(.A0(new_n18243_), .A1(new_n12171_), .B0(new_n18268_), .Y(new_n18269_));
  NOR3X1   g15833(.A(new_n18242_), .B(new_n12120_), .C(new_n12493_), .Y(new_n18270_));
  OR2X1    g15834(.A(new_n18269_), .B(new_n18270_), .Y(new_n18271_));
  NOR2X1   g15835(.A(new_n18244_), .B(new_n18242_), .Y(new_n18272_));
  OAI21X1  g15836(.A0(new_n18272_), .A1(new_n12494_), .B0(new_n12584_), .Y(new_n18273_));
  AOI21X1  g15837(.A0(new_n18271_), .A1(new_n18246_), .B0(new_n18273_), .Y(new_n18274_));
  NOR3X1   g15838(.A(new_n18270_), .B(new_n18268_), .C(new_n12494_), .Y(new_n18275_));
  OAI21X1  g15839(.A0(new_n18247_), .A1(new_n18244_), .B0(pi0608), .Y(new_n18276_));
  NOR2X1   g15840(.A(new_n18276_), .B(new_n18275_), .Y(new_n18277_));
  OAI21X1  g15841(.A0(new_n18277_), .A1(new_n18274_), .B0(pi0778), .Y(new_n18278_));
  OAI21X1  g15842(.A0(new_n18269_), .A1(pi0778), .B0(new_n18278_), .Y(new_n18279_));
  OAI21X1  g15843(.A0(new_n18250_), .A1(new_n12590_), .B0(new_n12591_), .Y(new_n18280_));
  AOI21X1  g15844(.A0(new_n18279_), .A1(new_n12590_), .B0(new_n18280_), .Y(new_n18281_));
  NOR3X1   g15845(.A(new_n18281_), .B(new_n18224_), .C(pi0660), .Y(new_n18282_));
  OAI21X1  g15846(.A0(new_n18250_), .A1(pi0609), .B0(pi1155), .Y(new_n18283_));
  AOI21X1  g15847(.A0(new_n18279_), .A1(pi0609), .B0(new_n18283_), .Y(new_n18284_));
  NOR3X1   g15848(.A(new_n18284_), .B(new_n18226_), .C(new_n12596_), .Y(new_n18285_));
  OAI21X1  g15849(.A0(new_n18285_), .A1(new_n18282_), .B0(pi0785), .Y(new_n18286_));
  NAND2X1  g15850(.A(new_n18279_), .B(new_n11888_), .Y(new_n18287_));
  AND2X1   g15851(.A(new_n18287_), .B(new_n18286_), .Y(new_n18288_));
  NOR3X1   g15852(.A(new_n18250_), .B(new_n12762_), .C(new_n12614_), .Y(new_n18289_));
  NOR2X1   g15853(.A(new_n18289_), .B(pi1154), .Y(new_n18290_));
  OAI21X1  g15854(.A0(new_n18288_), .A1(pi0618), .B0(new_n18290_), .Y(new_n18291_));
  NOR2X1   g15855(.A(new_n18230_), .B(pi0627), .Y(new_n18292_));
  NOR3X1   g15856(.A(new_n18250_), .B(new_n12762_), .C(pi0618), .Y(new_n18293_));
  NOR2X1   g15857(.A(new_n18293_), .B(new_n12615_), .Y(new_n18294_));
  OAI21X1  g15858(.A0(new_n18288_), .A1(new_n12614_), .B0(new_n18294_), .Y(new_n18295_));
  NOR2X1   g15859(.A(new_n18231_), .B(new_n12622_), .Y(new_n18296_));
  AOI22X1  g15860(.A0(new_n18296_), .A1(new_n18295_), .B0(new_n18292_), .B1(new_n18291_), .Y(new_n18297_));
  MX2X1    g15861(.A(new_n18297_), .B(new_n18288_), .S0(new_n11887_), .Y(new_n18298_));
  OR4X1    g15862(.A(new_n18250_), .B(new_n12764_), .C(new_n12762_), .D(new_n12637_), .Y(new_n18299_));
  AND2X1   g15863(.A(new_n18299_), .B(new_n12638_), .Y(new_n18300_));
  OAI21X1  g15864(.A0(new_n18298_), .A1(pi0619), .B0(new_n18300_), .Y(new_n18301_));
  NOR2X1   g15865(.A(new_n18235_), .B(pi0648), .Y(new_n18302_));
  AND2X1   g15866(.A(new_n18302_), .B(new_n18301_), .Y(new_n18303_));
  INVX1    g15867(.A(new_n18303_), .Y(new_n18304_));
  NOR4X1   g15868(.A(new_n18250_), .B(new_n12764_), .C(new_n12762_), .D(pi0619), .Y(new_n18305_));
  NOR2X1   g15869(.A(new_n18305_), .B(new_n12638_), .Y(new_n18306_));
  OAI21X1  g15870(.A0(new_n18298_), .A1(new_n12637_), .B0(new_n18306_), .Y(new_n18307_));
  NOR2X1   g15871(.A(new_n18236_), .B(new_n12645_), .Y(new_n18308_));
  AOI21X1  g15872(.A0(new_n18308_), .A1(new_n18307_), .B0(new_n11886_), .Y(new_n18309_));
  AOI21X1  g15873(.A0(new_n18298_), .A1(new_n11886_), .B0(new_n14264_), .Y(new_n18310_));
  INVX1    g15874(.A(new_n18310_), .Y(new_n18311_));
  AOI21X1  g15875(.A0(new_n18309_), .A1(new_n18304_), .B0(new_n18311_), .Y(new_n18312_));
  OAI21X1  g15876(.A0(new_n18312_), .A1(new_n18267_), .B0(new_n16350_), .Y(new_n18313_));
  INVX1    g15877(.A(new_n18240_), .Y(new_n18314_));
  AND2X1   g15878(.A(new_n18251_), .B(new_n12852_), .Y(new_n18315_));
  AOI22X1  g15879(.A0(new_n18315_), .A1(new_n14564_), .B0(new_n18314_), .B1(new_n12867_), .Y(new_n18316_));
  AOI22X1  g15880(.A0(new_n18315_), .A1(new_n14566_), .B0(new_n18314_), .B1(new_n12865_), .Y(new_n18317_));
  MX2X1    g15881(.A(new_n18317_), .B(new_n18316_), .S0(new_n12689_), .Y(new_n18318_));
  OAI21X1  g15882(.A0(new_n18318_), .A1(new_n11884_), .B0(new_n14562_), .Y(new_n18319_));
  INVX1    g15883(.A(new_n18319_), .Y(new_n18320_));
  AOI21X1  g15884(.A0(new_n18320_), .A1(new_n18313_), .B0(new_n18260_), .Y(new_n18321_));
  OAI21X1  g15885(.A0(new_n18257_), .A1(new_n12706_), .B0(new_n18256_), .Y(new_n18322_));
  MX2X1    g15886(.A(new_n18322_), .B(new_n18254_), .S0(new_n11883_), .Y(new_n18323_));
  OAI21X1  g15887(.A0(new_n18323_), .A1(pi0644), .B0(pi0715), .Y(new_n18324_));
  AOI21X1  g15888(.A0(new_n18321_), .A1(pi0644), .B0(new_n18324_), .Y(new_n18325_));
  OR4X1    g15889(.A(new_n12734_), .B(new_n2739_), .C(new_n11883_), .D(pi0182), .Y(new_n18326_));
  OAI21X1  g15890(.A0(new_n18241_), .A1(new_n12735_), .B0(new_n18326_), .Y(new_n18327_));
  OAI21X1  g15891(.A0(new_n18219_), .A1(pi0644), .B0(new_n12739_), .Y(new_n18328_));
  AOI21X1  g15892(.A0(new_n18327_), .A1(pi0644), .B0(new_n18328_), .Y(new_n18329_));
  OR2X1    g15893(.A(new_n18329_), .B(new_n11882_), .Y(new_n18330_));
  OAI21X1  g15894(.A0(new_n18323_), .A1(new_n12743_), .B0(new_n12739_), .Y(new_n18331_));
  AOI21X1  g15895(.A0(new_n18321_), .A1(new_n12743_), .B0(new_n18331_), .Y(new_n18332_));
  OAI21X1  g15896(.A0(new_n18219_), .A1(new_n12743_), .B0(pi0715), .Y(new_n18333_));
  AOI21X1  g15897(.A0(new_n18327_), .A1(new_n12743_), .B0(new_n18333_), .Y(new_n18334_));
  OR2X1    g15898(.A(new_n18334_), .B(pi1160), .Y(new_n18335_));
  OAI22X1  g15899(.A0(new_n18335_), .A1(new_n18332_), .B0(new_n18330_), .B1(new_n18325_), .Y(new_n18336_));
  NAND2X1  g15900(.A(new_n18336_), .B(pi0790), .Y(new_n18337_));
  AOI21X1  g15901(.A0(new_n18321_), .A1(new_n12897_), .B0(new_n12898_), .Y(new_n18338_));
  AOI21X1  g15902(.A0(new_n13699_), .A1(new_n3129_), .B0(pi0182), .Y(new_n18339_));
  INVX1    g15903(.A(new_n18339_), .Y(new_n18340_));
  OAI21X1  g15904(.A0(new_n3810_), .A1(pi0734), .B0(new_n18339_), .Y(new_n18341_));
  AOI21X1  g15905(.A0(new_n12955_), .A1(pi0182), .B0(pi0038), .Y(new_n18342_));
  OAI22X1  g15906(.A0(new_n18342_), .A1(new_n3810_), .B0(new_n12953_), .B1(pi0182), .Y(new_n18343_));
  OAI21X1  g15907(.A0(new_n12202_), .A1(pi0182), .B0(new_n12567_), .Y(new_n18344_));
  NAND3X1  g15908(.A(new_n18344_), .B(new_n18343_), .C(new_n15209_), .Y(new_n18345_));
  AND2X1   g15909(.A(new_n18345_), .B(new_n18341_), .Y(new_n18346_));
  INVX1    g15910(.A(new_n18346_), .Y(new_n18347_));
  AOI21X1  g15911(.A0(new_n18339_), .A1(new_n12493_), .B0(new_n12494_), .Y(new_n18348_));
  OAI21X1  g15912(.A0(new_n18346_), .A1(new_n12493_), .B0(new_n18348_), .Y(new_n18349_));
  AOI21X1  g15913(.A0(new_n18339_), .A1(pi0625), .B0(pi1153), .Y(new_n18350_));
  OAI21X1  g15914(.A0(new_n18346_), .A1(pi0625), .B0(new_n18350_), .Y(new_n18351_));
  AND2X1   g15915(.A(new_n18351_), .B(new_n18349_), .Y(new_n18352_));
  MX2X1    g15916(.A(new_n18352_), .B(new_n18347_), .S0(new_n11889_), .Y(new_n18353_));
  MX2X1    g15917(.A(new_n18353_), .B(new_n18339_), .S0(new_n12618_), .Y(new_n18354_));
  INVX1    g15918(.A(new_n18354_), .Y(new_n18355_));
  MX2X1    g15919(.A(new_n18355_), .B(new_n18340_), .S0(new_n12641_), .Y(new_n18356_));
  INVX1    g15920(.A(new_n18356_), .Y(new_n18357_));
  MX2X1    g15921(.A(new_n18357_), .B(new_n18339_), .S0(new_n12659_), .Y(new_n18358_));
  AND2X1   g15922(.A(new_n18339_), .B(new_n12691_), .Y(new_n18359_));
  AOI21X1  g15923(.A0(new_n18358_), .A1(new_n17252_), .B0(new_n18359_), .Y(new_n18360_));
  AOI21X1  g15924(.A0(new_n18339_), .A1(new_n12683_), .B0(new_n12684_), .Y(new_n18361_));
  OAI21X1  g15925(.A0(new_n18360_), .A1(new_n12683_), .B0(new_n18361_), .Y(new_n18362_));
  AOI21X1  g15926(.A0(new_n18339_), .A1(pi0628), .B0(pi1156), .Y(new_n18363_));
  OAI21X1  g15927(.A0(new_n18360_), .A1(pi0628), .B0(new_n18363_), .Y(new_n18364_));
  AOI21X1  g15928(.A0(new_n18364_), .A1(new_n18362_), .B0(new_n11884_), .Y(new_n18365_));
  AOI21X1  g15929(.A0(new_n18360_), .A1(new_n11884_), .B0(new_n18365_), .Y(new_n18366_));
  MX2X1    g15930(.A(new_n18366_), .B(new_n18339_), .S0(pi0647), .Y(new_n18367_));
  MX2X1    g15931(.A(new_n18366_), .B(new_n18339_), .S0(new_n12705_), .Y(new_n18368_));
  MX2X1    g15932(.A(new_n18368_), .B(new_n18367_), .S0(new_n12706_), .Y(new_n18369_));
  MX2X1    g15933(.A(new_n18369_), .B(new_n18366_), .S0(new_n11883_), .Y(new_n18370_));
  AOI21X1  g15934(.A0(new_n18370_), .A1(new_n12743_), .B0(new_n12739_), .Y(new_n18371_));
  OAI22X1  g15935(.A0(new_n14342_), .A1(pi0756), .B0(new_n12202_), .B1(pi0182), .Y(new_n18372_));
  AOI21X1  g15936(.A0(new_n13977_), .A1(pi0182), .B0(pi0756), .Y(new_n18373_));
  OAI21X1  g15937(.A0(new_n12910_), .A1(pi0182), .B0(new_n18373_), .Y(new_n18374_));
  NAND3X1  g15938(.A(new_n12090_), .B(pi0756), .C(new_n5227_), .Y(new_n18375_));
  AOI21X1  g15939(.A0(new_n18375_), .A1(new_n18374_), .B0(pi0038), .Y(new_n18376_));
  AOI21X1  g15940(.A0(new_n18372_), .A1(pi0038), .B0(new_n18376_), .Y(new_n18377_));
  MX2X1    g15941(.A(new_n18377_), .B(pi0182), .S0(new_n3810_), .Y(new_n18378_));
  AND2X1   g15942(.A(new_n18378_), .B(new_n12623_), .Y(new_n18379_));
  AOI21X1  g15943(.A0(new_n18340_), .A1(new_n12601_), .B0(new_n18379_), .Y(new_n18380_));
  AOI22X1  g15944(.A0(new_n18379_), .A1(pi0609), .B0(new_n18340_), .B1(new_n13430_), .Y(new_n18381_));
  AOI22X1  g15945(.A0(new_n18379_), .A1(new_n12590_), .B0(new_n18340_), .B1(new_n13436_), .Y(new_n18382_));
  MX2X1    g15946(.A(new_n18382_), .B(new_n18381_), .S0(pi1155), .Y(new_n18383_));
  MX2X1    g15947(.A(new_n18383_), .B(new_n18380_), .S0(new_n11888_), .Y(new_n18384_));
  OAI21X1  g15948(.A0(new_n18340_), .A1(pi0618), .B0(pi1154), .Y(new_n18385_));
  AOI21X1  g15949(.A0(new_n18384_), .A1(pi0618), .B0(new_n18385_), .Y(new_n18386_));
  OAI21X1  g15950(.A0(new_n18340_), .A1(new_n12614_), .B0(new_n12615_), .Y(new_n18387_));
  AOI21X1  g15951(.A0(new_n18384_), .A1(new_n12614_), .B0(new_n18387_), .Y(new_n18388_));
  NOR2X1   g15952(.A(new_n18388_), .B(new_n18386_), .Y(new_n18389_));
  MX2X1    g15953(.A(new_n18389_), .B(new_n18384_), .S0(new_n11887_), .Y(new_n18390_));
  OAI21X1  g15954(.A0(new_n18340_), .A1(pi0619), .B0(pi1159), .Y(new_n18391_));
  AOI21X1  g15955(.A0(new_n18390_), .A1(pi0619), .B0(new_n18391_), .Y(new_n18392_));
  OAI21X1  g15956(.A0(new_n18340_), .A1(new_n12637_), .B0(new_n12638_), .Y(new_n18393_));
  AOI21X1  g15957(.A0(new_n18390_), .A1(new_n12637_), .B0(new_n18393_), .Y(new_n18394_));
  NOR2X1   g15958(.A(new_n18394_), .B(new_n18392_), .Y(new_n18395_));
  MX2X1    g15959(.A(new_n18395_), .B(new_n18390_), .S0(new_n11886_), .Y(new_n18396_));
  MX2X1    g15960(.A(new_n18396_), .B(new_n18339_), .S0(new_n12841_), .Y(new_n18397_));
  MX2X1    g15961(.A(new_n18397_), .B(new_n18339_), .S0(new_n12711_), .Y(new_n18398_));
  MX2X1    g15962(.A(new_n18398_), .B(new_n18339_), .S0(new_n12735_), .Y(new_n18399_));
  OAI21X1  g15963(.A0(new_n18340_), .A1(pi0644), .B0(new_n12739_), .Y(new_n18400_));
  AOI21X1  g15964(.A0(new_n18399_), .A1(pi0644), .B0(new_n18400_), .Y(new_n18401_));
  OR2X1    g15965(.A(new_n18401_), .B(new_n11882_), .Y(new_n18402_));
  AOI21X1  g15966(.A0(new_n18370_), .A1(pi0644), .B0(pi0715), .Y(new_n18403_));
  OAI21X1  g15967(.A0(new_n18340_), .A1(new_n12743_), .B0(pi0715), .Y(new_n18404_));
  AOI21X1  g15968(.A0(new_n18399_), .A1(new_n12743_), .B0(new_n18404_), .Y(new_n18405_));
  OR2X1    g15969(.A(new_n18405_), .B(pi1160), .Y(new_n18406_));
  OAI22X1  g15970(.A0(new_n18406_), .A1(new_n18403_), .B0(new_n18402_), .B1(new_n18371_), .Y(new_n18407_));
  NOR3X1   g15971(.A(new_n18405_), .B(pi1160), .C(pi0644), .Y(new_n18408_));
  NOR3X1   g15972(.A(new_n18401_), .B(new_n11882_), .C(new_n12743_), .Y(new_n18409_));
  NOR3X1   g15973(.A(new_n18409_), .B(new_n18408_), .C(new_n12897_), .Y(new_n18410_));
  MX2X1    g15974(.A(new_n18364_), .B(new_n18362_), .S0(new_n12689_), .Y(new_n18411_));
  OAI21X1  g15975(.A0(new_n18397_), .A1(new_n14395_), .B0(new_n18411_), .Y(new_n18412_));
  NAND2X1  g15976(.A(new_n18412_), .B(pi0792), .Y(new_n18413_));
  OR2X1    g15977(.A(new_n18377_), .B(new_n15209_), .Y(new_n18414_));
  OAI21X1  g15978(.A0(new_n12349_), .A1(new_n5227_), .B0(pi0756), .Y(new_n18415_));
  AOI21X1  g15979(.A0(new_n12289_), .A1(new_n5227_), .B0(new_n18415_), .Y(new_n18416_));
  OAI21X1  g15980(.A0(new_n12440_), .A1(pi0182), .B0(new_n15203_), .Y(new_n18417_));
  AOI21X1  g15981(.A0(new_n12401_), .A1(pi0182), .B0(new_n18417_), .Y(new_n18418_));
  OR2X1    g15982(.A(new_n18418_), .B(new_n2959_), .Y(new_n18419_));
  AND2X1   g15983(.A(new_n12467_), .B(pi0182), .Y(new_n18420_));
  OAI21X1  g15984(.A0(new_n12454_), .A1(pi0182), .B0(pi0756), .Y(new_n18421_));
  NOR4X1   g15985(.A(new_n13391_), .B(new_n12908_), .C(new_n12907_), .D(pi0182), .Y(new_n18422_));
  OAI21X1  g15986(.A0(new_n12929_), .A1(new_n5227_), .B0(new_n15203_), .Y(new_n18423_));
  OAI22X1  g15987(.A0(new_n18423_), .A1(new_n18422_), .B0(new_n18421_), .B1(new_n18420_), .Y(new_n18424_));
  AOI21X1  g15988(.A0(new_n18424_), .A1(new_n2959_), .B0(pi0038), .Y(new_n18425_));
  OAI21X1  g15989(.A0(new_n18419_), .A1(new_n18416_), .B0(new_n18425_), .Y(new_n18426_));
  OAI21X1  g15990(.A0(new_n12478_), .A1(pi0756), .B0(new_n13669_), .Y(new_n18427_));
  NAND2X1  g15991(.A(new_n18427_), .B(new_n5227_), .Y(new_n18428_));
  AOI21X1  g15992(.A0(new_n18222_), .A1(new_n14209_), .B0(new_n5227_), .Y(new_n18429_));
  AOI21X1  g15993(.A0(new_n18429_), .A1(new_n6857_), .B0(new_n2996_), .Y(new_n18430_));
  AOI21X1  g15994(.A0(new_n18430_), .A1(new_n18428_), .B0(pi0734), .Y(new_n18431_));
  AOI21X1  g15995(.A0(new_n18431_), .A1(new_n18426_), .B0(new_n3810_), .Y(new_n18432_));
  AOI22X1  g15996(.A0(new_n18432_), .A1(new_n18414_), .B0(new_n3810_), .B1(pi0182), .Y(new_n18433_));
  OAI21X1  g15997(.A0(new_n18378_), .A1(new_n12493_), .B0(new_n12494_), .Y(new_n18434_));
  AOI21X1  g15998(.A0(new_n18433_), .A1(new_n12493_), .B0(new_n18434_), .Y(new_n18435_));
  NAND2X1  g15999(.A(new_n18349_), .B(new_n12584_), .Y(new_n18436_));
  OAI21X1  g16000(.A0(new_n18378_), .A1(pi0625), .B0(pi1153), .Y(new_n18437_));
  AOI21X1  g16001(.A0(new_n18433_), .A1(pi0625), .B0(new_n18437_), .Y(new_n18438_));
  NAND2X1  g16002(.A(new_n18351_), .B(pi0608), .Y(new_n18439_));
  OAI22X1  g16003(.A0(new_n18439_), .A1(new_n18438_), .B0(new_n18436_), .B1(new_n18435_), .Y(new_n18440_));
  MX2X1    g16004(.A(new_n18440_), .B(new_n18433_), .S0(new_n11889_), .Y(new_n18441_));
  INVX1    g16005(.A(new_n18353_), .Y(new_n18442_));
  OAI21X1  g16006(.A0(new_n18442_), .A1(new_n12590_), .B0(new_n12591_), .Y(new_n18443_));
  AOI21X1  g16007(.A0(new_n18441_), .A1(new_n12590_), .B0(new_n18443_), .Y(new_n18444_));
  OAI21X1  g16008(.A0(new_n18381_), .A1(new_n12591_), .B0(new_n12596_), .Y(new_n18445_));
  OAI21X1  g16009(.A0(new_n18442_), .A1(pi0609), .B0(pi1155), .Y(new_n18446_));
  AOI21X1  g16010(.A0(new_n18441_), .A1(pi0609), .B0(new_n18446_), .Y(new_n18447_));
  OAI21X1  g16011(.A0(new_n18382_), .A1(pi1155), .B0(pi0660), .Y(new_n18448_));
  OAI22X1  g16012(.A0(new_n18448_), .A1(new_n18447_), .B0(new_n18445_), .B1(new_n18444_), .Y(new_n18449_));
  MX2X1    g16013(.A(new_n18449_), .B(new_n18441_), .S0(new_n11888_), .Y(new_n18450_));
  OAI21X1  g16014(.A0(new_n18355_), .A1(new_n12614_), .B0(new_n12615_), .Y(new_n18451_));
  AOI21X1  g16015(.A0(new_n18450_), .A1(new_n12614_), .B0(new_n18451_), .Y(new_n18452_));
  OR2X1    g16016(.A(new_n18386_), .B(pi0627), .Y(new_n18453_));
  OAI21X1  g16017(.A0(new_n18355_), .A1(pi0618), .B0(pi1154), .Y(new_n18454_));
  AOI21X1  g16018(.A0(new_n18450_), .A1(pi0618), .B0(new_n18454_), .Y(new_n18455_));
  OR2X1    g16019(.A(new_n18388_), .B(new_n12622_), .Y(new_n18456_));
  OAI22X1  g16020(.A0(new_n18456_), .A1(new_n18455_), .B0(new_n18453_), .B1(new_n18452_), .Y(new_n18457_));
  MX2X1    g16021(.A(new_n18457_), .B(new_n18450_), .S0(new_n11887_), .Y(new_n18458_));
  NAND2X1  g16022(.A(new_n18458_), .B(new_n12637_), .Y(new_n18459_));
  AOI21X1  g16023(.A0(new_n18357_), .A1(pi0619), .B0(pi1159), .Y(new_n18460_));
  OR2X1    g16024(.A(new_n18392_), .B(pi0648), .Y(new_n18461_));
  AOI21X1  g16025(.A0(new_n18460_), .A1(new_n18459_), .B0(new_n18461_), .Y(new_n18462_));
  NAND2X1  g16026(.A(new_n18458_), .B(pi0619), .Y(new_n18463_));
  AOI21X1  g16027(.A0(new_n18357_), .A1(new_n12637_), .B0(new_n12638_), .Y(new_n18464_));
  OR2X1    g16028(.A(new_n18394_), .B(new_n12645_), .Y(new_n18465_));
  AOI21X1  g16029(.A0(new_n18464_), .A1(new_n18463_), .B0(new_n18465_), .Y(new_n18466_));
  NOR3X1   g16030(.A(new_n18466_), .B(new_n18462_), .C(new_n11886_), .Y(new_n18467_));
  OAI21X1  g16031(.A0(new_n18458_), .A1(pi0789), .B0(new_n12842_), .Y(new_n18468_));
  AOI21X1  g16032(.A0(new_n18340_), .A1(pi0626), .B0(new_n16352_), .Y(new_n18469_));
  OAI21X1  g16033(.A0(new_n18396_), .A1(pi0626), .B0(new_n18469_), .Y(new_n18470_));
  AOI21X1  g16034(.A0(new_n18340_), .A1(new_n12664_), .B0(new_n16356_), .Y(new_n18471_));
  OAI21X1  g16035(.A0(new_n18396_), .A1(new_n12664_), .B0(new_n18471_), .Y(new_n18472_));
  NAND2X1  g16036(.A(new_n18358_), .B(new_n12769_), .Y(new_n18473_));
  NAND3X1  g16037(.A(new_n18473_), .B(new_n18472_), .C(new_n18470_), .Y(new_n18474_));
  AOI21X1  g16038(.A0(new_n18474_), .A1(pi0788), .B0(new_n14273_), .Y(new_n18475_));
  OAI21X1  g16039(.A0(new_n18468_), .A1(new_n18467_), .B0(new_n18475_), .Y(new_n18476_));
  AOI21X1  g16040(.A0(new_n18476_), .A1(new_n18413_), .B0(new_n14269_), .Y(new_n18477_));
  OR2X1    g16041(.A(new_n18398_), .B(new_n14384_), .Y(new_n18478_));
  OR2X1    g16042(.A(new_n18367_), .B(new_n14389_), .Y(new_n18479_));
  OR2X1    g16043(.A(new_n18368_), .B(new_n14387_), .Y(new_n18480_));
  NAND3X1  g16044(.A(new_n18480_), .B(new_n18479_), .C(new_n18478_), .Y(new_n18481_));
  AND2X1   g16045(.A(new_n18481_), .B(pi0787), .Y(new_n18482_));
  NOR3X1   g16046(.A(new_n18482_), .B(new_n18477_), .C(new_n18410_), .Y(new_n18483_));
  AOI21X1  g16047(.A0(new_n18407_), .A1(pi0790), .B0(new_n18483_), .Y(new_n18484_));
  OR2X1    g16048(.A(new_n18484_), .B(po1038), .Y(new_n18485_));
  AOI21X1  g16049(.A0(po1038), .A1(new_n5227_), .B0(pi0832), .Y(new_n18486_));
  AOI22X1  g16050(.A0(new_n18486_), .A1(new_n18485_), .B0(new_n18338_), .B1(new_n18337_), .Y(po0339));
  AOI21X1  g16051(.A0(pi1093), .A1(pi1092), .B0(pi0183), .Y(new_n18488_));
  INVX1    g16052(.A(new_n18488_), .Y(new_n18489_));
  AOI21X1  g16053(.A0(new_n12178_), .A1(new_n14782_), .B0(new_n18488_), .Y(new_n18490_));
  AOI21X1  g16054(.A0(new_n12601_), .A1(new_n2739_), .B0(new_n18490_), .Y(new_n18491_));
  NAND2X1  g16055(.A(new_n12178_), .B(new_n14782_), .Y(new_n18492_));
  OAI21X1  g16056(.A0(new_n18492_), .A1(new_n13436_), .B0(new_n18491_), .Y(new_n18493_));
  AND2X1   g16057(.A(new_n18493_), .B(pi1155), .Y(new_n18494_));
  NOR2X1   g16058(.A(new_n18492_), .B(new_n13436_), .Y(new_n18495_));
  NOR3X1   g16059(.A(new_n18495_), .B(new_n18488_), .C(pi1155), .Y(new_n18496_));
  OAI21X1  g16060(.A0(new_n18496_), .A1(new_n18494_), .B0(pi0785), .Y(new_n18497_));
  OAI21X1  g16061(.A0(new_n18491_), .A1(pi0785), .B0(new_n18497_), .Y(new_n18498_));
  INVX1    g16062(.A(new_n18498_), .Y(new_n18499_));
  AOI21X1  g16063(.A0(new_n18499_), .A1(new_n12785_), .B0(new_n12615_), .Y(new_n18500_));
  AOI21X1  g16064(.A0(new_n18499_), .A1(new_n12788_), .B0(pi1154), .Y(new_n18501_));
  NOR2X1   g16065(.A(new_n18501_), .B(new_n18500_), .Y(new_n18502_));
  MX2X1    g16066(.A(new_n18502_), .B(new_n18499_), .S0(new_n11887_), .Y(new_n18503_));
  OR2X1    g16067(.A(new_n18503_), .B(pi0789), .Y(new_n18504_));
  AOI21X1  g16068(.A0(new_n18503_), .A1(new_n15910_), .B0(new_n12638_), .Y(new_n18505_));
  AOI21X1  g16069(.A0(new_n18503_), .A1(new_n15912_), .B0(pi1159), .Y(new_n18506_));
  OAI21X1  g16070(.A0(new_n18506_), .A1(new_n18505_), .B0(pi0789), .Y(new_n18507_));
  AND2X1   g16071(.A(new_n18507_), .B(new_n18504_), .Y(new_n18508_));
  INVX1    g16072(.A(new_n18508_), .Y(new_n18509_));
  MX2X1    g16073(.A(new_n18509_), .B(new_n18489_), .S0(new_n12841_), .Y(new_n18510_));
  MX2X1    g16074(.A(new_n18510_), .B(new_n18489_), .S0(new_n12711_), .Y(new_n18511_));
  AOI21X1  g16075(.A0(new_n12566_), .A1(new_n14788_), .B0(new_n18488_), .Y(new_n18512_));
  INVX1    g16076(.A(new_n18512_), .Y(new_n18513_));
  NOR3X1   g16077(.A(new_n13585_), .B(pi0725), .C(pi0625), .Y(new_n18514_));
  OR2X1    g16078(.A(new_n18514_), .B(new_n18512_), .Y(new_n18515_));
  NOR2X1   g16079(.A(new_n18488_), .B(pi1153), .Y(new_n18516_));
  INVX1    g16080(.A(new_n18516_), .Y(new_n18517_));
  OAI21X1  g16081(.A0(new_n18517_), .A1(new_n18514_), .B0(pi0778), .Y(new_n18518_));
  AOI21X1  g16082(.A0(new_n18515_), .A1(pi1153), .B0(new_n18518_), .Y(new_n18519_));
  AOI21X1  g16083(.A0(new_n18513_), .A1(new_n11889_), .B0(new_n18519_), .Y(new_n18520_));
  NOR4X1   g16084(.A(new_n18520_), .B(new_n12765_), .C(new_n12764_), .D(new_n12762_), .Y(new_n18521_));
  INVX1    g16085(.A(new_n18521_), .Y(new_n18522_));
  NOR3X1   g16086(.A(new_n18522_), .B(new_n12870_), .C(new_n12851_), .Y(new_n18523_));
  INVX1    g16087(.A(new_n18523_), .Y(new_n18524_));
  AOI21X1  g16088(.A0(new_n18488_), .A1(pi0647), .B0(pi1157), .Y(new_n18525_));
  OAI21X1  g16089(.A0(new_n18524_), .A1(pi0647), .B0(new_n18525_), .Y(new_n18526_));
  MX2X1    g16090(.A(new_n18523_), .B(new_n18488_), .S0(new_n12705_), .Y(new_n18527_));
  OAI22X1  g16091(.A0(new_n18527_), .A1(new_n14387_), .B0(new_n18526_), .B1(new_n12723_), .Y(new_n18528_));
  AOI21X1  g16092(.A0(new_n18511_), .A1(new_n14385_), .B0(new_n18528_), .Y(new_n18529_));
  NOR2X1   g16093(.A(new_n18529_), .B(new_n11883_), .Y(new_n18530_));
  AOI21X1  g16094(.A0(new_n18489_), .A1(pi0626), .B0(new_n16352_), .Y(new_n18531_));
  OAI21X1  g16095(.A0(new_n18508_), .A1(pi0626), .B0(new_n18531_), .Y(new_n18532_));
  AOI21X1  g16096(.A0(new_n18507_), .A1(new_n18504_), .B0(new_n12664_), .Y(new_n18533_));
  NOR2X1   g16097(.A(new_n18488_), .B(pi0626), .Y(new_n18534_));
  NOR3X1   g16098(.A(new_n18534_), .B(new_n18533_), .C(new_n16356_), .Y(new_n18535_));
  AOI21X1  g16099(.A0(new_n18521_), .A1(new_n12769_), .B0(new_n18535_), .Y(new_n18536_));
  AOI21X1  g16100(.A0(new_n18536_), .A1(new_n18532_), .B0(new_n11885_), .Y(new_n18537_));
  INVX1    g16101(.A(new_n18490_), .Y(new_n18538_));
  AOI21X1  g16102(.A0(new_n18513_), .A1(new_n12171_), .B0(new_n18538_), .Y(new_n18539_));
  NOR3X1   g16103(.A(new_n18512_), .B(new_n12120_), .C(new_n12493_), .Y(new_n18540_));
  OR2X1    g16104(.A(new_n18539_), .B(new_n18540_), .Y(new_n18541_));
  NOR2X1   g16105(.A(new_n18514_), .B(new_n18512_), .Y(new_n18542_));
  OAI21X1  g16106(.A0(new_n18542_), .A1(new_n12494_), .B0(new_n12584_), .Y(new_n18543_));
  AOI21X1  g16107(.A0(new_n18541_), .A1(new_n18516_), .B0(new_n18543_), .Y(new_n18544_));
  NOR3X1   g16108(.A(new_n18540_), .B(new_n18538_), .C(new_n12494_), .Y(new_n18545_));
  OAI21X1  g16109(.A0(new_n18517_), .A1(new_n18514_), .B0(pi0608), .Y(new_n18546_));
  NOR2X1   g16110(.A(new_n18546_), .B(new_n18545_), .Y(new_n18547_));
  OAI21X1  g16111(.A0(new_n18547_), .A1(new_n18544_), .B0(pi0778), .Y(new_n18548_));
  OAI21X1  g16112(.A0(new_n18539_), .A1(pi0778), .B0(new_n18548_), .Y(new_n18549_));
  OAI21X1  g16113(.A0(new_n18520_), .A1(new_n12590_), .B0(new_n12591_), .Y(new_n18550_));
  AOI21X1  g16114(.A0(new_n18549_), .A1(new_n12590_), .B0(new_n18550_), .Y(new_n18551_));
  NOR3X1   g16115(.A(new_n18551_), .B(new_n18494_), .C(pi0660), .Y(new_n18552_));
  OAI21X1  g16116(.A0(new_n18520_), .A1(pi0609), .B0(pi1155), .Y(new_n18553_));
  AOI21X1  g16117(.A0(new_n18549_), .A1(pi0609), .B0(new_n18553_), .Y(new_n18554_));
  NOR3X1   g16118(.A(new_n18554_), .B(new_n18496_), .C(new_n12596_), .Y(new_n18555_));
  OAI21X1  g16119(.A0(new_n18555_), .A1(new_n18552_), .B0(pi0785), .Y(new_n18556_));
  NAND2X1  g16120(.A(new_n18549_), .B(new_n11888_), .Y(new_n18557_));
  AND2X1   g16121(.A(new_n18557_), .B(new_n18556_), .Y(new_n18558_));
  NOR3X1   g16122(.A(new_n18520_), .B(new_n12762_), .C(new_n12614_), .Y(new_n18559_));
  NOR2X1   g16123(.A(new_n18559_), .B(pi1154), .Y(new_n18560_));
  OAI21X1  g16124(.A0(new_n18558_), .A1(pi0618), .B0(new_n18560_), .Y(new_n18561_));
  NOR2X1   g16125(.A(new_n18500_), .B(pi0627), .Y(new_n18562_));
  NOR3X1   g16126(.A(new_n18520_), .B(new_n12762_), .C(pi0618), .Y(new_n18563_));
  NOR2X1   g16127(.A(new_n18563_), .B(new_n12615_), .Y(new_n18564_));
  OAI21X1  g16128(.A0(new_n18558_), .A1(new_n12614_), .B0(new_n18564_), .Y(new_n18565_));
  NOR2X1   g16129(.A(new_n18501_), .B(new_n12622_), .Y(new_n18566_));
  AOI22X1  g16130(.A0(new_n18566_), .A1(new_n18565_), .B0(new_n18562_), .B1(new_n18561_), .Y(new_n18567_));
  MX2X1    g16131(.A(new_n18567_), .B(new_n18558_), .S0(new_n11887_), .Y(new_n18568_));
  OR4X1    g16132(.A(new_n18520_), .B(new_n12764_), .C(new_n12762_), .D(new_n12637_), .Y(new_n18569_));
  AND2X1   g16133(.A(new_n18569_), .B(new_n12638_), .Y(new_n18570_));
  OAI21X1  g16134(.A0(new_n18568_), .A1(pi0619), .B0(new_n18570_), .Y(new_n18571_));
  NOR2X1   g16135(.A(new_n18505_), .B(pi0648), .Y(new_n18572_));
  AND2X1   g16136(.A(new_n18572_), .B(new_n18571_), .Y(new_n18573_));
  INVX1    g16137(.A(new_n18573_), .Y(new_n18574_));
  NOR4X1   g16138(.A(new_n18520_), .B(new_n12764_), .C(new_n12762_), .D(pi0619), .Y(new_n18575_));
  NOR2X1   g16139(.A(new_n18575_), .B(new_n12638_), .Y(new_n18576_));
  OAI21X1  g16140(.A0(new_n18568_), .A1(new_n12637_), .B0(new_n18576_), .Y(new_n18577_));
  NOR2X1   g16141(.A(new_n18506_), .B(new_n12645_), .Y(new_n18578_));
  AOI21X1  g16142(.A0(new_n18578_), .A1(new_n18577_), .B0(new_n11886_), .Y(new_n18579_));
  AOI21X1  g16143(.A0(new_n18568_), .A1(new_n11886_), .B0(new_n14264_), .Y(new_n18580_));
  INVX1    g16144(.A(new_n18580_), .Y(new_n18581_));
  AOI21X1  g16145(.A0(new_n18579_), .A1(new_n18574_), .B0(new_n18581_), .Y(new_n18582_));
  OAI21X1  g16146(.A0(new_n18582_), .A1(new_n18537_), .B0(new_n16350_), .Y(new_n18583_));
  INVX1    g16147(.A(new_n18510_), .Y(new_n18584_));
  AND2X1   g16148(.A(new_n18521_), .B(new_n12852_), .Y(new_n18585_));
  AOI22X1  g16149(.A0(new_n18585_), .A1(new_n14564_), .B0(new_n18584_), .B1(new_n12867_), .Y(new_n18586_));
  AOI22X1  g16150(.A0(new_n18585_), .A1(new_n14566_), .B0(new_n18584_), .B1(new_n12865_), .Y(new_n18587_));
  MX2X1    g16151(.A(new_n18587_), .B(new_n18586_), .S0(new_n12689_), .Y(new_n18588_));
  OAI21X1  g16152(.A0(new_n18588_), .A1(new_n11884_), .B0(new_n14562_), .Y(new_n18589_));
  INVX1    g16153(.A(new_n18589_), .Y(new_n18590_));
  AOI21X1  g16154(.A0(new_n18590_), .A1(new_n18583_), .B0(new_n18530_), .Y(new_n18591_));
  OAI21X1  g16155(.A0(new_n18527_), .A1(new_n12706_), .B0(new_n18526_), .Y(new_n18592_));
  MX2X1    g16156(.A(new_n18592_), .B(new_n18524_), .S0(new_n11883_), .Y(new_n18593_));
  OAI21X1  g16157(.A0(new_n18593_), .A1(pi0644), .B0(pi0715), .Y(new_n18594_));
  AOI21X1  g16158(.A0(new_n18591_), .A1(pi0644), .B0(new_n18594_), .Y(new_n18595_));
  OR4X1    g16159(.A(new_n12734_), .B(new_n2739_), .C(new_n11883_), .D(pi0183), .Y(new_n18596_));
  OAI21X1  g16160(.A0(new_n18511_), .A1(new_n12735_), .B0(new_n18596_), .Y(new_n18597_));
  OAI21X1  g16161(.A0(new_n18489_), .A1(pi0644), .B0(new_n12739_), .Y(new_n18598_));
  AOI21X1  g16162(.A0(new_n18597_), .A1(pi0644), .B0(new_n18598_), .Y(new_n18599_));
  OR2X1    g16163(.A(new_n18599_), .B(new_n11882_), .Y(new_n18600_));
  OAI21X1  g16164(.A0(new_n18593_), .A1(new_n12743_), .B0(new_n12739_), .Y(new_n18601_));
  AOI21X1  g16165(.A0(new_n18591_), .A1(new_n12743_), .B0(new_n18601_), .Y(new_n18602_));
  OAI21X1  g16166(.A0(new_n18489_), .A1(new_n12743_), .B0(pi0715), .Y(new_n18603_));
  AOI21X1  g16167(.A0(new_n18597_), .A1(new_n12743_), .B0(new_n18603_), .Y(new_n18604_));
  OR2X1    g16168(.A(new_n18604_), .B(pi1160), .Y(new_n18605_));
  OAI22X1  g16169(.A0(new_n18605_), .A1(new_n18602_), .B0(new_n18600_), .B1(new_n18595_), .Y(new_n18606_));
  NAND2X1  g16170(.A(new_n18606_), .B(pi0790), .Y(new_n18607_));
  AOI21X1  g16171(.A0(new_n18591_), .A1(new_n12897_), .B0(new_n12898_), .Y(new_n18608_));
  AOI21X1  g16172(.A0(new_n13699_), .A1(new_n3129_), .B0(pi0183), .Y(new_n18609_));
  INVX1    g16173(.A(new_n18609_), .Y(new_n18610_));
  OAI21X1  g16174(.A0(new_n3810_), .A1(pi0725), .B0(new_n18609_), .Y(new_n18611_));
  AOI21X1  g16175(.A0(new_n12955_), .A1(pi0183), .B0(pi0038), .Y(new_n18612_));
  OAI22X1  g16176(.A0(new_n18612_), .A1(new_n3810_), .B0(new_n12953_), .B1(pi0183), .Y(new_n18613_));
  OAI21X1  g16177(.A0(new_n12202_), .A1(pi0183), .B0(new_n12567_), .Y(new_n18614_));
  NAND3X1  g16178(.A(new_n18614_), .B(new_n18613_), .C(new_n14788_), .Y(new_n18615_));
  AND2X1   g16179(.A(new_n18615_), .B(new_n18611_), .Y(new_n18616_));
  INVX1    g16180(.A(new_n18616_), .Y(new_n18617_));
  AOI21X1  g16181(.A0(new_n18609_), .A1(new_n12493_), .B0(new_n12494_), .Y(new_n18618_));
  OAI21X1  g16182(.A0(new_n18616_), .A1(new_n12493_), .B0(new_n18618_), .Y(new_n18619_));
  AOI21X1  g16183(.A0(new_n18609_), .A1(pi0625), .B0(pi1153), .Y(new_n18620_));
  OAI21X1  g16184(.A0(new_n18616_), .A1(pi0625), .B0(new_n18620_), .Y(new_n18621_));
  AND2X1   g16185(.A(new_n18621_), .B(new_n18619_), .Y(new_n18622_));
  MX2X1    g16186(.A(new_n18622_), .B(new_n18617_), .S0(new_n11889_), .Y(new_n18623_));
  MX2X1    g16187(.A(new_n18623_), .B(new_n18609_), .S0(new_n12618_), .Y(new_n18624_));
  INVX1    g16188(.A(new_n18624_), .Y(new_n18625_));
  MX2X1    g16189(.A(new_n18625_), .B(new_n18610_), .S0(new_n12641_), .Y(new_n18626_));
  INVX1    g16190(.A(new_n18626_), .Y(new_n18627_));
  MX2X1    g16191(.A(new_n18627_), .B(new_n18609_), .S0(new_n12659_), .Y(new_n18628_));
  AND2X1   g16192(.A(new_n18609_), .B(new_n12691_), .Y(new_n18629_));
  AOI21X1  g16193(.A0(new_n18628_), .A1(new_n17252_), .B0(new_n18629_), .Y(new_n18630_));
  AOI21X1  g16194(.A0(new_n18609_), .A1(new_n12683_), .B0(new_n12684_), .Y(new_n18631_));
  OAI21X1  g16195(.A0(new_n18630_), .A1(new_n12683_), .B0(new_n18631_), .Y(new_n18632_));
  AOI21X1  g16196(.A0(new_n18609_), .A1(pi0628), .B0(pi1156), .Y(new_n18633_));
  OAI21X1  g16197(.A0(new_n18630_), .A1(pi0628), .B0(new_n18633_), .Y(new_n18634_));
  AOI21X1  g16198(.A0(new_n18634_), .A1(new_n18632_), .B0(new_n11884_), .Y(new_n18635_));
  AOI21X1  g16199(.A0(new_n18630_), .A1(new_n11884_), .B0(new_n18635_), .Y(new_n18636_));
  MX2X1    g16200(.A(new_n18636_), .B(new_n18609_), .S0(pi0647), .Y(new_n18637_));
  MX2X1    g16201(.A(new_n18636_), .B(new_n18609_), .S0(new_n12705_), .Y(new_n18638_));
  MX2X1    g16202(.A(new_n18638_), .B(new_n18637_), .S0(new_n12706_), .Y(new_n18639_));
  MX2X1    g16203(.A(new_n18639_), .B(new_n18636_), .S0(new_n11883_), .Y(new_n18640_));
  AOI21X1  g16204(.A0(new_n18640_), .A1(new_n12743_), .B0(new_n12739_), .Y(new_n18641_));
  OAI22X1  g16205(.A0(new_n14342_), .A1(pi0755), .B0(new_n12202_), .B1(pi0183), .Y(new_n18642_));
  AOI21X1  g16206(.A0(new_n13977_), .A1(pi0183), .B0(pi0755), .Y(new_n18643_));
  OAI21X1  g16207(.A0(new_n12910_), .A1(pi0183), .B0(new_n18643_), .Y(new_n18644_));
  NAND3X1  g16208(.A(new_n12090_), .B(pi0755), .C(new_n6928_), .Y(new_n18645_));
  AOI21X1  g16209(.A0(new_n18645_), .A1(new_n18644_), .B0(pi0038), .Y(new_n18646_));
  AOI21X1  g16210(.A0(new_n18642_), .A1(pi0038), .B0(new_n18646_), .Y(new_n18647_));
  MX2X1    g16211(.A(new_n18647_), .B(pi0183), .S0(new_n3810_), .Y(new_n18648_));
  AND2X1   g16212(.A(new_n18648_), .B(new_n12623_), .Y(new_n18649_));
  AOI21X1  g16213(.A0(new_n18610_), .A1(new_n12601_), .B0(new_n18649_), .Y(new_n18650_));
  AOI22X1  g16214(.A0(new_n18649_), .A1(pi0609), .B0(new_n18610_), .B1(new_n13430_), .Y(new_n18651_));
  AOI22X1  g16215(.A0(new_n18649_), .A1(new_n12590_), .B0(new_n18610_), .B1(new_n13436_), .Y(new_n18652_));
  MX2X1    g16216(.A(new_n18652_), .B(new_n18651_), .S0(pi1155), .Y(new_n18653_));
  MX2X1    g16217(.A(new_n18653_), .B(new_n18650_), .S0(new_n11888_), .Y(new_n18654_));
  OAI21X1  g16218(.A0(new_n18610_), .A1(pi0618), .B0(pi1154), .Y(new_n18655_));
  AOI21X1  g16219(.A0(new_n18654_), .A1(pi0618), .B0(new_n18655_), .Y(new_n18656_));
  OAI21X1  g16220(.A0(new_n18610_), .A1(new_n12614_), .B0(new_n12615_), .Y(new_n18657_));
  AOI21X1  g16221(.A0(new_n18654_), .A1(new_n12614_), .B0(new_n18657_), .Y(new_n18658_));
  NOR2X1   g16222(.A(new_n18658_), .B(new_n18656_), .Y(new_n18659_));
  MX2X1    g16223(.A(new_n18659_), .B(new_n18654_), .S0(new_n11887_), .Y(new_n18660_));
  OAI21X1  g16224(.A0(new_n18610_), .A1(pi0619), .B0(pi1159), .Y(new_n18661_));
  AOI21X1  g16225(.A0(new_n18660_), .A1(pi0619), .B0(new_n18661_), .Y(new_n18662_));
  OAI21X1  g16226(.A0(new_n18610_), .A1(new_n12637_), .B0(new_n12638_), .Y(new_n18663_));
  AOI21X1  g16227(.A0(new_n18660_), .A1(new_n12637_), .B0(new_n18663_), .Y(new_n18664_));
  NOR2X1   g16228(.A(new_n18664_), .B(new_n18662_), .Y(new_n18665_));
  MX2X1    g16229(.A(new_n18665_), .B(new_n18660_), .S0(new_n11886_), .Y(new_n18666_));
  MX2X1    g16230(.A(new_n18666_), .B(new_n18609_), .S0(new_n12841_), .Y(new_n18667_));
  MX2X1    g16231(.A(new_n18667_), .B(new_n18609_), .S0(new_n12711_), .Y(new_n18668_));
  MX2X1    g16232(.A(new_n18668_), .B(new_n18609_), .S0(new_n12735_), .Y(new_n18669_));
  OAI21X1  g16233(.A0(new_n18610_), .A1(pi0644), .B0(new_n12739_), .Y(new_n18670_));
  AOI21X1  g16234(.A0(new_n18669_), .A1(pi0644), .B0(new_n18670_), .Y(new_n18671_));
  OR2X1    g16235(.A(new_n18671_), .B(new_n11882_), .Y(new_n18672_));
  AOI21X1  g16236(.A0(new_n18640_), .A1(pi0644), .B0(pi0715), .Y(new_n18673_));
  OAI21X1  g16237(.A0(new_n18610_), .A1(new_n12743_), .B0(pi0715), .Y(new_n18674_));
  AOI21X1  g16238(.A0(new_n18669_), .A1(new_n12743_), .B0(new_n18674_), .Y(new_n18675_));
  OR2X1    g16239(.A(new_n18675_), .B(pi1160), .Y(new_n18676_));
  OAI22X1  g16240(.A0(new_n18676_), .A1(new_n18673_), .B0(new_n18672_), .B1(new_n18641_), .Y(new_n18677_));
  NOR3X1   g16241(.A(new_n18675_), .B(pi1160), .C(pi0644), .Y(new_n18678_));
  NOR3X1   g16242(.A(new_n18671_), .B(new_n11882_), .C(new_n12743_), .Y(new_n18679_));
  NOR3X1   g16243(.A(new_n18679_), .B(new_n18678_), .C(new_n12897_), .Y(new_n18680_));
  MX2X1    g16244(.A(new_n18634_), .B(new_n18632_), .S0(new_n12689_), .Y(new_n18681_));
  OAI21X1  g16245(.A0(new_n18667_), .A1(new_n14395_), .B0(new_n18681_), .Y(new_n18682_));
  NAND2X1  g16246(.A(new_n18682_), .B(pi0792), .Y(new_n18683_));
  OR2X1    g16247(.A(new_n18647_), .B(new_n14788_), .Y(new_n18684_));
  OAI21X1  g16248(.A0(new_n12349_), .A1(new_n6928_), .B0(pi0755), .Y(new_n18685_));
  AOI21X1  g16249(.A0(new_n12289_), .A1(new_n6928_), .B0(new_n18685_), .Y(new_n18686_));
  OAI21X1  g16250(.A0(new_n12440_), .A1(pi0183), .B0(new_n14782_), .Y(new_n18687_));
  AOI21X1  g16251(.A0(new_n12401_), .A1(pi0183), .B0(new_n18687_), .Y(new_n18688_));
  OR2X1    g16252(.A(new_n18688_), .B(new_n2959_), .Y(new_n18689_));
  AND2X1   g16253(.A(new_n12467_), .B(pi0183), .Y(new_n18690_));
  OAI21X1  g16254(.A0(new_n12454_), .A1(pi0183), .B0(pi0755), .Y(new_n18691_));
  NOR4X1   g16255(.A(new_n13391_), .B(new_n12908_), .C(new_n12907_), .D(pi0183), .Y(new_n18692_));
  OAI21X1  g16256(.A0(new_n12929_), .A1(new_n6928_), .B0(new_n14782_), .Y(new_n18693_));
  OAI22X1  g16257(.A0(new_n18693_), .A1(new_n18692_), .B0(new_n18691_), .B1(new_n18690_), .Y(new_n18694_));
  AOI21X1  g16258(.A0(new_n18694_), .A1(new_n2959_), .B0(pi0038), .Y(new_n18695_));
  OAI21X1  g16259(.A0(new_n18689_), .A1(new_n18686_), .B0(new_n18695_), .Y(new_n18696_));
  OAI21X1  g16260(.A0(new_n12478_), .A1(pi0755), .B0(new_n13669_), .Y(new_n18697_));
  NAND2X1  g16261(.A(new_n18697_), .B(new_n6928_), .Y(new_n18698_));
  AOI21X1  g16262(.A0(new_n18492_), .A1(new_n14209_), .B0(new_n6928_), .Y(new_n18699_));
  AOI21X1  g16263(.A0(new_n18699_), .A1(new_n6857_), .B0(new_n2996_), .Y(new_n18700_));
  AOI21X1  g16264(.A0(new_n18700_), .A1(new_n18698_), .B0(pi0725), .Y(new_n18701_));
  AOI21X1  g16265(.A0(new_n18701_), .A1(new_n18696_), .B0(new_n3810_), .Y(new_n18702_));
  AOI22X1  g16266(.A0(new_n18702_), .A1(new_n18684_), .B0(new_n3810_), .B1(pi0183), .Y(new_n18703_));
  OAI21X1  g16267(.A0(new_n18648_), .A1(new_n12493_), .B0(new_n12494_), .Y(new_n18704_));
  AOI21X1  g16268(.A0(new_n18703_), .A1(new_n12493_), .B0(new_n18704_), .Y(new_n18705_));
  NAND2X1  g16269(.A(new_n18619_), .B(new_n12584_), .Y(new_n18706_));
  OAI21X1  g16270(.A0(new_n18648_), .A1(pi0625), .B0(pi1153), .Y(new_n18707_));
  AOI21X1  g16271(.A0(new_n18703_), .A1(pi0625), .B0(new_n18707_), .Y(new_n18708_));
  NAND2X1  g16272(.A(new_n18621_), .B(pi0608), .Y(new_n18709_));
  OAI22X1  g16273(.A0(new_n18709_), .A1(new_n18708_), .B0(new_n18706_), .B1(new_n18705_), .Y(new_n18710_));
  MX2X1    g16274(.A(new_n18710_), .B(new_n18703_), .S0(new_n11889_), .Y(new_n18711_));
  INVX1    g16275(.A(new_n18623_), .Y(new_n18712_));
  OAI21X1  g16276(.A0(new_n18712_), .A1(new_n12590_), .B0(new_n12591_), .Y(new_n18713_));
  AOI21X1  g16277(.A0(new_n18711_), .A1(new_n12590_), .B0(new_n18713_), .Y(new_n18714_));
  OAI21X1  g16278(.A0(new_n18651_), .A1(new_n12591_), .B0(new_n12596_), .Y(new_n18715_));
  OAI21X1  g16279(.A0(new_n18712_), .A1(pi0609), .B0(pi1155), .Y(new_n18716_));
  AOI21X1  g16280(.A0(new_n18711_), .A1(pi0609), .B0(new_n18716_), .Y(new_n18717_));
  OAI21X1  g16281(.A0(new_n18652_), .A1(pi1155), .B0(pi0660), .Y(new_n18718_));
  OAI22X1  g16282(.A0(new_n18718_), .A1(new_n18717_), .B0(new_n18715_), .B1(new_n18714_), .Y(new_n18719_));
  MX2X1    g16283(.A(new_n18719_), .B(new_n18711_), .S0(new_n11888_), .Y(new_n18720_));
  OAI21X1  g16284(.A0(new_n18625_), .A1(new_n12614_), .B0(new_n12615_), .Y(new_n18721_));
  AOI21X1  g16285(.A0(new_n18720_), .A1(new_n12614_), .B0(new_n18721_), .Y(new_n18722_));
  OR2X1    g16286(.A(new_n18656_), .B(pi0627), .Y(new_n18723_));
  OAI21X1  g16287(.A0(new_n18625_), .A1(pi0618), .B0(pi1154), .Y(new_n18724_));
  AOI21X1  g16288(.A0(new_n18720_), .A1(pi0618), .B0(new_n18724_), .Y(new_n18725_));
  OR2X1    g16289(.A(new_n18658_), .B(new_n12622_), .Y(new_n18726_));
  OAI22X1  g16290(.A0(new_n18726_), .A1(new_n18725_), .B0(new_n18723_), .B1(new_n18722_), .Y(new_n18727_));
  MX2X1    g16291(.A(new_n18727_), .B(new_n18720_), .S0(new_n11887_), .Y(new_n18728_));
  NAND2X1  g16292(.A(new_n18728_), .B(new_n12637_), .Y(new_n18729_));
  AOI21X1  g16293(.A0(new_n18627_), .A1(pi0619), .B0(pi1159), .Y(new_n18730_));
  OR2X1    g16294(.A(new_n18662_), .B(pi0648), .Y(new_n18731_));
  AOI21X1  g16295(.A0(new_n18730_), .A1(new_n18729_), .B0(new_n18731_), .Y(new_n18732_));
  NAND2X1  g16296(.A(new_n18728_), .B(pi0619), .Y(new_n18733_));
  AOI21X1  g16297(.A0(new_n18627_), .A1(new_n12637_), .B0(new_n12638_), .Y(new_n18734_));
  OR2X1    g16298(.A(new_n18664_), .B(new_n12645_), .Y(new_n18735_));
  AOI21X1  g16299(.A0(new_n18734_), .A1(new_n18733_), .B0(new_n18735_), .Y(new_n18736_));
  NOR3X1   g16300(.A(new_n18736_), .B(new_n18732_), .C(new_n11886_), .Y(new_n18737_));
  OAI21X1  g16301(.A0(new_n18728_), .A1(pi0789), .B0(new_n12842_), .Y(new_n18738_));
  AOI21X1  g16302(.A0(new_n18610_), .A1(pi0626), .B0(new_n16352_), .Y(new_n18739_));
  OAI21X1  g16303(.A0(new_n18666_), .A1(pi0626), .B0(new_n18739_), .Y(new_n18740_));
  AOI21X1  g16304(.A0(new_n18610_), .A1(new_n12664_), .B0(new_n16356_), .Y(new_n18741_));
  OAI21X1  g16305(.A0(new_n18666_), .A1(new_n12664_), .B0(new_n18741_), .Y(new_n18742_));
  NAND2X1  g16306(.A(new_n18628_), .B(new_n12769_), .Y(new_n18743_));
  NAND3X1  g16307(.A(new_n18743_), .B(new_n18742_), .C(new_n18740_), .Y(new_n18744_));
  AOI21X1  g16308(.A0(new_n18744_), .A1(pi0788), .B0(new_n14273_), .Y(new_n18745_));
  OAI21X1  g16309(.A0(new_n18738_), .A1(new_n18737_), .B0(new_n18745_), .Y(new_n18746_));
  AOI21X1  g16310(.A0(new_n18746_), .A1(new_n18683_), .B0(new_n14269_), .Y(new_n18747_));
  OR2X1    g16311(.A(new_n18668_), .B(new_n14384_), .Y(new_n18748_));
  OR2X1    g16312(.A(new_n18637_), .B(new_n14389_), .Y(new_n18749_));
  OR2X1    g16313(.A(new_n18638_), .B(new_n14387_), .Y(new_n18750_));
  NAND3X1  g16314(.A(new_n18750_), .B(new_n18749_), .C(new_n18748_), .Y(new_n18751_));
  AND2X1   g16315(.A(new_n18751_), .B(pi0787), .Y(new_n18752_));
  NOR3X1   g16316(.A(new_n18752_), .B(new_n18747_), .C(new_n18680_), .Y(new_n18753_));
  AOI21X1  g16317(.A0(new_n18677_), .A1(pi0790), .B0(new_n18753_), .Y(new_n18754_));
  OR2X1    g16318(.A(new_n18754_), .B(po1038), .Y(new_n18755_));
  AOI21X1  g16319(.A0(po1038), .A1(new_n6928_), .B0(pi0832), .Y(new_n18756_));
  AOI22X1  g16320(.A0(new_n18756_), .A1(new_n18755_), .B0(new_n18608_), .B1(new_n18607_), .Y(po0340));
  AOI21X1  g16321(.A0(pi1093), .A1(pi1092), .B0(pi0184), .Y(new_n18758_));
  INVX1    g16322(.A(new_n18758_), .Y(new_n18759_));
  AOI21X1  g16323(.A0(new_n12178_), .A1(new_n15329_), .B0(new_n18758_), .Y(new_n18760_));
  AOI21X1  g16324(.A0(new_n12601_), .A1(new_n2739_), .B0(new_n18760_), .Y(new_n18761_));
  NAND2X1  g16325(.A(new_n12178_), .B(new_n15329_), .Y(new_n18762_));
  OAI21X1  g16326(.A0(new_n18762_), .A1(new_n13436_), .B0(new_n18761_), .Y(new_n18763_));
  AND2X1   g16327(.A(new_n18763_), .B(pi1155), .Y(new_n18764_));
  NOR2X1   g16328(.A(new_n18762_), .B(new_n13436_), .Y(new_n18765_));
  NOR3X1   g16329(.A(new_n18765_), .B(new_n18758_), .C(pi1155), .Y(new_n18766_));
  OAI21X1  g16330(.A0(new_n18766_), .A1(new_n18764_), .B0(pi0785), .Y(new_n18767_));
  OAI21X1  g16331(.A0(new_n18761_), .A1(pi0785), .B0(new_n18767_), .Y(new_n18768_));
  INVX1    g16332(.A(new_n18768_), .Y(new_n18769_));
  AOI21X1  g16333(.A0(new_n18769_), .A1(new_n12785_), .B0(new_n12615_), .Y(new_n18770_));
  AOI21X1  g16334(.A0(new_n18769_), .A1(new_n12788_), .B0(pi1154), .Y(new_n18771_));
  NOR2X1   g16335(.A(new_n18771_), .B(new_n18770_), .Y(new_n18772_));
  MX2X1    g16336(.A(new_n18772_), .B(new_n18769_), .S0(new_n11887_), .Y(new_n18773_));
  OR2X1    g16337(.A(new_n18773_), .B(pi0789), .Y(new_n18774_));
  AOI21X1  g16338(.A0(new_n18773_), .A1(new_n15910_), .B0(new_n12638_), .Y(new_n18775_));
  AOI21X1  g16339(.A0(new_n18773_), .A1(new_n15912_), .B0(pi1159), .Y(new_n18776_));
  OAI21X1  g16340(.A0(new_n18776_), .A1(new_n18775_), .B0(pi0789), .Y(new_n18777_));
  AND2X1   g16341(.A(new_n18777_), .B(new_n18774_), .Y(new_n18778_));
  INVX1    g16342(.A(new_n18778_), .Y(new_n18779_));
  MX2X1    g16343(.A(new_n18779_), .B(new_n18759_), .S0(new_n12841_), .Y(new_n18780_));
  MX2X1    g16344(.A(new_n18780_), .B(new_n18759_), .S0(new_n12711_), .Y(new_n18781_));
  AOI21X1  g16345(.A0(new_n12566_), .A1(new_n15335_), .B0(new_n18758_), .Y(new_n18782_));
  INVX1    g16346(.A(new_n18782_), .Y(new_n18783_));
  NOR3X1   g16347(.A(new_n13585_), .B(pi0737), .C(pi0625), .Y(new_n18784_));
  OR2X1    g16348(.A(new_n18784_), .B(new_n18782_), .Y(new_n18785_));
  NOR2X1   g16349(.A(new_n18758_), .B(pi1153), .Y(new_n18786_));
  INVX1    g16350(.A(new_n18786_), .Y(new_n18787_));
  OAI21X1  g16351(.A0(new_n18787_), .A1(new_n18784_), .B0(pi0778), .Y(new_n18788_));
  AOI21X1  g16352(.A0(new_n18785_), .A1(pi1153), .B0(new_n18788_), .Y(new_n18789_));
  AOI21X1  g16353(.A0(new_n18783_), .A1(new_n11889_), .B0(new_n18789_), .Y(new_n18790_));
  NOR4X1   g16354(.A(new_n18790_), .B(new_n12765_), .C(new_n12764_), .D(new_n12762_), .Y(new_n18791_));
  INVX1    g16355(.A(new_n18791_), .Y(new_n18792_));
  NOR3X1   g16356(.A(new_n18792_), .B(new_n12870_), .C(new_n12851_), .Y(new_n18793_));
  INVX1    g16357(.A(new_n18793_), .Y(new_n18794_));
  AOI21X1  g16358(.A0(new_n18758_), .A1(pi0647), .B0(pi1157), .Y(new_n18795_));
  OAI21X1  g16359(.A0(new_n18794_), .A1(pi0647), .B0(new_n18795_), .Y(new_n18796_));
  MX2X1    g16360(.A(new_n18793_), .B(new_n18758_), .S0(new_n12705_), .Y(new_n18797_));
  OAI22X1  g16361(.A0(new_n18797_), .A1(new_n14387_), .B0(new_n18796_), .B1(new_n12723_), .Y(new_n18798_));
  AOI21X1  g16362(.A0(new_n18781_), .A1(new_n14385_), .B0(new_n18798_), .Y(new_n18799_));
  NOR2X1   g16363(.A(new_n18799_), .B(new_n11883_), .Y(new_n18800_));
  AOI21X1  g16364(.A0(new_n18759_), .A1(pi0626), .B0(new_n16352_), .Y(new_n18801_));
  OAI21X1  g16365(.A0(new_n18778_), .A1(pi0626), .B0(new_n18801_), .Y(new_n18802_));
  AOI21X1  g16366(.A0(new_n18777_), .A1(new_n18774_), .B0(new_n12664_), .Y(new_n18803_));
  NOR2X1   g16367(.A(new_n18758_), .B(pi0626), .Y(new_n18804_));
  NOR3X1   g16368(.A(new_n18804_), .B(new_n18803_), .C(new_n16356_), .Y(new_n18805_));
  AOI21X1  g16369(.A0(new_n18791_), .A1(new_n12769_), .B0(new_n18805_), .Y(new_n18806_));
  AOI21X1  g16370(.A0(new_n18806_), .A1(new_n18802_), .B0(new_n11885_), .Y(new_n18807_));
  INVX1    g16371(.A(new_n18760_), .Y(new_n18808_));
  AOI21X1  g16372(.A0(new_n18783_), .A1(new_n12171_), .B0(new_n18808_), .Y(new_n18809_));
  NOR3X1   g16373(.A(new_n18782_), .B(new_n12120_), .C(new_n12493_), .Y(new_n18810_));
  OR2X1    g16374(.A(new_n18809_), .B(new_n18810_), .Y(new_n18811_));
  NOR2X1   g16375(.A(new_n18784_), .B(new_n18782_), .Y(new_n18812_));
  OAI21X1  g16376(.A0(new_n18812_), .A1(new_n12494_), .B0(new_n12584_), .Y(new_n18813_));
  AOI21X1  g16377(.A0(new_n18811_), .A1(new_n18786_), .B0(new_n18813_), .Y(new_n18814_));
  NOR3X1   g16378(.A(new_n18810_), .B(new_n18808_), .C(new_n12494_), .Y(new_n18815_));
  OAI21X1  g16379(.A0(new_n18787_), .A1(new_n18784_), .B0(pi0608), .Y(new_n18816_));
  NOR2X1   g16380(.A(new_n18816_), .B(new_n18815_), .Y(new_n18817_));
  OAI21X1  g16381(.A0(new_n18817_), .A1(new_n18814_), .B0(pi0778), .Y(new_n18818_));
  OAI21X1  g16382(.A0(new_n18809_), .A1(pi0778), .B0(new_n18818_), .Y(new_n18819_));
  OAI21X1  g16383(.A0(new_n18790_), .A1(new_n12590_), .B0(new_n12591_), .Y(new_n18820_));
  AOI21X1  g16384(.A0(new_n18819_), .A1(new_n12590_), .B0(new_n18820_), .Y(new_n18821_));
  NOR3X1   g16385(.A(new_n18821_), .B(new_n18764_), .C(pi0660), .Y(new_n18822_));
  OAI21X1  g16386(.A0(new_n18790_), .A1(pi0609), .B0(pi1155), .Y(new_n18823_));
  AOI21X1  g16387(.A0(new_n18819_), .A1(pi0609), .B0(new_n18823_), .Y(new_n18824_));
  NOR3X1   g16388(.A(new_n18824_), .B(new_n18766_), .C(new_n12596_), .Y(new_n18825_));
  OAI21X1  g16389(.A0(new_n18825_), .A1(new_n18822_), .B0(pi0785), .Y(new_n18826_));
  NAND2X1  g16390(.A(new_n18819_), .B(new_n11888_), .Y(new_n18827_));
  AND2X1   g16391(.A(new_n18827_), .B(new_n18826_), .Y(new_n18828_));
  NOR3X1   g16392(.A(new_n18790_), .B(new_n12762_), .C(new_n12614_), .Y(new_n18829_));
  NOR2X1   g16393(.A(new_n18829_), .B(pi1154), .Y(new_n18830_));
  OAI21X1  g16394(.A0(new_n18828_), .A1(pi0618), .B0(new_n18830_), .Y(new_n18831_));
  NOR2X1   g16395(.A(new_n18770_), .B(pi0627), .Y(new_n18832_));
  NOR3X1   g16396(.A(new_n18790_), .B(new_n12762_), .C(pi0618), .Y(new_n18833_));
  NOR2X1   g16397(.A(new_n18833_), .B(new_n12615_), .Y(new_n18834_));
  OAI21X1  g16398(.A0(new_n18828_), .A1(new_n12614_), .B0(new_n18834_), .Y(new_n18835_));
  NOR2X1   g16399(.A(new_n18771_), .B(new_n12622_), .Y(new_n18836_));
  AOI22X1  g16400(.A0(new_n18836_), .A1(new_n18835_), .B0(new_n18832_), .B1(new_n18831_), .Y(new_n18837_));
  MX2X1    g16401(.A(new_n18837_), .B(new_n18828_), .S0(new_n11887_), .Y(new_n18838_));
  OR4X1    g16402(.A(new_n18790_), .B(new_n12764_), .C(new_n12762_), .D(new_n12637_), .Y(new_n18839_));
  AND2X1   g16403(.A(new_n18839_), .B(new_n12638_), .Y(new_n18840_));
  OAI21X1  g16404(.A0(new_n18838_), .A1(pi0619), .B0(new_n18840_), .Y(new_n18841_));
  NOR2X1   g16405(.A(new_n18775_), .B(pi0648), .Y(new_n18842_));
  AND2X1   g16406(.A(new_n18842_), .B(new_n18841_), .Y(new_n18843_));
  INVX1    g16407(.A(new_n18843_), .Y(new_n18844_));
  NOR4X1   g16408(.A(new_n18790_), .B(new_n12764_), .C(new_n12762_), .D(pi0619), .Y(new_n18845_));
  NOR2X1   g16409(.A(new_n18845_), .B(new_n12638_), .Y(new_n18846_));
  OAI21X1  g16410(.A0(new_n18838_), .A1(new_n12637_), .B0(new_n18846_), .Y(new_n18847_));
  NOR2X1   g16411(.A(new_n18776_), .B(new_n12645_), .Y(new_n18848_));
  AOI21X1  g16412(.A0(new_n18848_), .A1(new_n18847_), .B0(new_n11886_), .Y(new_n18849_));
  AOI21X1  g16413(.A0(new_n18838_), .A1(new_n11886_), .B0(new_n14264_), .Y(new_n18850_));
  INVX1    g16414(.A(new_n18850_), .Y(new_n18851_));
  AOI21X1  g16415(.A0(new_n18849_), .A1(new_n18844_), .B0(new_n18851_), .Y(new_n18852_));
  OAI21X1  g16416(.A0(new_n18852_), .A1(new_n18807_), .B0(new_n16350_), .Y(new_n18853_));
  INVX1    g16417(.A(new_n18780_), .Y(new_n18854_));
  AND2X1   g16418(.A(new_n18791_), .B(new_n12852_), .Y(new_n18855_));
  AOI22X1  g16419(.A0(new_n18855_), .A1(new_n14564_), .B0(new_n18854_), .B1(new_n12867_), .Y(new_n18856_));
  AOI22X1  g16420(.A0(new_n18855_), .A1(new_n14566_), .B0(new_n18854_), .B1(new_n12865_), .Y(new_n18857_));
  MX2X1    g16421(.A(new_n18857_), .B(new_n18856_), .S0(new_n12689_), .Y(new_n18858_));
  OAI21X1  g16422(.A0(new_n18858_), .A1(new_n11884_), .B0(new_n14562_), .Y(new_n18859_));
  INVX1    g16423(.A(new_n18859_), .Y(new_n18860_));
  AOI21X1  g16424(.A0(new_n18860_), .A1(new_n18853_), .B0(new_n18800_), .Y(new_n18861_));
  OAI21X1  g16425(.A0(new_n18797_), .A1(new_n12706_), .B0(new_n18796_), .Y(new_n18862_));
  MX2X1    g16426(.A(new_n18862_), .B(new_n18794_), .S0(new_n11883_), .Y(new_n18863_));
  OAI21X1  g16427(.A0(new_n18863_), .A1(pi0644), .B0(pi0715), .Y(new_n18864_));
  AOI21X1  g16428(.A0(new_n18861_), .A1(pi0644), .B0(new_n18864_), .Y(new_n18865_));
  OR4X1    g16429(.A(new_n12734_), .B(new_n2739_), .C(new_n11883_), .D(pi0184), .Y(new_n18866_));
  OAI21X1  g16430(.A0(new_n18781_), .A1(new_n12735_), .B0(new_n18866_), .Y(new_n18867_));
  OAI21X1  g16431(.A0(new_n18759_), .A1(pi0644), .B0(new_n12739_), .Y(new_n18868_));
  AOI21X1  g16432(.A0(new_n18867_), .A1(pi0644), .B0(new_n18868_), .Y(new_n18869_));
  OR2X1    g16433(.A(new_n18869_), .B(new_n11882_), .Y(new_n18870_));
  OAI21X1  g16434(.A0(new_n18863_), .A1(new_n12743_), .B0(new_n12739_), .Y(new_n18871_));
  AOI21X1  g16435(.A0(new_n18861_), .A1(new_n12743_), .B0(new_n18871_), .Y(new_n18872_));
  OAI21X1  g16436(.A0(new_n18759_), .A1(new_n12743_), .B0(pi0715), .Y(new_n18873_));
  AOI21X1  g16437(.A0(new_n18867_), .A1(new_n12743_), .B0(new_n18873_), .Y(new_n18874_));
  OR2X1    g16438(.A(new_n18874_), .B(pi1160), .Y(new_n18875_));
  OAI22X1  g16439(.A0(new_n18875_), .A1(new_n18872_), .B0(new_n18870_), .B1(new_n18865_), .Y(new_n18876_));
  NAND2X1  g16440(.A(new_n18876_), .B(pi0790), .Y(new_n18877_));
  AOI21X1  g16441(.A0(new_n18861_), .A1(new_n12897_), .B0(new_n12898_), .Y(new_n18878_));
  AOI21X1  g16442(.A0(new_n13699_), .A1(new_n3129_), .B0(pi0184), .Y(new_n18879_));
  INVX1    g16443(.A(new_n18879_), .Y(new_n18880_));
  OAI21X1  g16444(.A0(new_n3810_), .A1(pi0737), .B0(new_n18879_), .Y(new_n18881_));
  AOI21X1  g16445(.A0(new_n12955_), .A1(pi0184), .B0(pi0038), .Y(new_n18882_));
  OAI22X1  g16446(.A0(new_n18882_), .A1(new_n3810_), .B0(new_n12953_), .B1(pi0184), .Y(new_n18883_));
  OAI21X1  g16447(.A0(new_n12202_), .A1(pi0184), .B0(new_n12567_), .Y(new_n18884_));
  NAND3X1  g16448(.A(new_n18884_), .B(new_n18883_), .C(new_n15335_), .Y(new_n18885_));
  AND2X1   g16449(.A(new_n18885_), .B(new_n18881_), .Y(new_n18886_));
  INVX1    g16450(.A(new_n18886_), .Y(new_n18887_));
  AOI21X1  g16451(.A0(new_n18879_), .A1(new_n12493_), .B0(new_n12494_), .Y(new_n18888_));
  OAI21X1  g16452(.A0(new_n18886_), .A1(new_n12493_), .B0(new_n18888_), .Y(new_n18889_));
  AOI21X1  g16453(.A0(new_n18879_), .A1(pi0625), .B0(pi1153), .Y(new_n18890_));
  OAI21X1  g16454(.A0(new_n18886_), .A1(pi0625), .B0(new_n18890_), .Y(new_n18891_));
  AND2X1   g16455(.A(new_n18891_), .B(new_n18889_), .Y(new_n18892_));
  MX2X1    g16456(.A(new_n18892_), .B(new_n18887_), .S0(new_n11889_), .Y(new_n18893_));
  MX2X1    g16457(.A(new_n18893_), .B(new_n18879_), .S0(new_n12618_), .Y(new_n18894_));
  INVX1    g16458(.A(new_n18894_), .Y(new_n18895_));
  MX2X1    g16459(.A(new_n18895_), .B(new_n18880_), .S0(new_n12641_), .Y(new_n18896_));
  INVX1    g16460(.A(new_n18896_), .Y(new_n18897_));
  MX2X1    g16461(.A(new_n18897_), .B(new_n18879_), .S0(new_n12659_), .Y(new_n18898_));
  AND2X1   g16462(.A(new_n18879_), .B(new_n12691_), .Y(new_n18899_));
  AOI21X1  g16463(.A0(new_n18898_), .A1(new_n17252_), .B0(new_n18899_), .Y(new_n18900_));
  AOI21X1  g16464(.A0(new_n18879_), .A1(new_n12683_), .B0(new_n12684_), .Y(new_n18901_));
  OAI21X1  g16465(.A0(new_n18900_), .A1(new_n12683_), .B0(new_n18901_), .Y(new_n18902_));
  AOI21X1  g16466(.A0(new_n18879_), .A1(pi0628), .B0(pi1156), .Y(new_n18903_));
  OAI21X1  g16467(.A0(new_n18900_), .A1(pi0628), .B0(new_n18903_), .Y(new_n18904_));
  AOI21X1  g16468(.A0(new_n18904_), .A1(new_n18902_), .B0(new_n11884_), .Y(new_n18905_));
  AOI21X1  g16469(.A0(new_n18900_), .A1(new_n11884_), .B0(new_n18905_), .Y(new_n18906_));
  MX2X1    g16470(.A(new_n18906_), .B(new_n18879_), .S0(pi0647), .Y(new_n18907_));
  MX2X1    g16471(.A(new_n18906_), .B(new_n18879_), .S0(new_n12705_), .Y(new_n18908_));
  MX2X1    g16472(.A(new_n18908_), .B(new_n18907_), .S0(new_n12706_), .Y(new_n18909_));
  MX2X1    g16473(.A(new_n18909_), .B(new_n18906_), .S0(new_n11883_), .Y(new_n18910_));
  AOI21X1  g16474(.A0(new_n18910_), .A1(new_n12743_), .B0(new_n12739_), .Y(new_n18911_));
  OAI22X1  g16475(.A0(new_n14342_), .A1(pi0777), .B0(new_n12202_), .B1(pi0184), .Y(new_n18912_));
  AOI21X1  g16476(.A0(new_n13977_), .A1(pi0184), .B0(pi0777), .Y(new_n18913_));
  OAI21X1  g16477(.A0(new_n12910_), .A1(pi0184), .B0(new_n18913_), .Y(new_n18914_));
  NAND3X1  g16478(.A(new_n12090_), .B(pi0777), .C(new_n8717_), .Y(new_n18915_));
  AOI21X1  g16479(.A0(new_n18915_), .A1(new_n18914_), .B0(pi0038), .Y(new_n18916_));
  AOI21X1  g16480(.A0(new_n18912_), .A1(pi0038), .B0(new_n18916_), .Y(new_n18917_));
  MX2X1    g16481(.A(new_n18917_), .B(pi0184), .S0(new_n3810_), .Y(new_n18918_));
  AND2X1   g16482(.A(new_n18918_), .B(new_n12623_), .Y(new_n18919_));
  AOI21X1  g16483(.A0(new_n18880_), .A1(new_n12601_), .B0(new_n18919_), .Y(new_n18920_));
  AOI22X1  g16484(.A0(new_n18919_), .A1(pi0609), .B0(new_n18880_), .B1(new_n13430_), .Y(new_n18921_));
  AOI22X1  g16485(.A0(new_n18919_), .A1(new_n12590_), .B0(new_n18880_), .B1(new_n13436_), .Y(new_n18922_));
  MX2X1    g16486(.A(new_n18922_), .B(new_n18921_), .S0(pi1155), .Y(new_n18923_));
  MX2X1    g16487(.A(new_n18923_), .B(new_n18920_), .S0(new_n11888_), .Y(new_n18924_));
  OAI21X1  g16488(.A0(new_n18880_), .A1(pi0618), .B0(pi1154), .Y(new_n18925_));
  AOI21X1  g16489(.A0(new_n18924_), .A1(pi0618), .B0(new_n18925_), .Y(new_n18926_));
  OAI21X1  g16490(.A0(new_n18880_), .A1(new_n12614_), .B0(new_n12615_), .Y(new_n18927_));
  AOI21X1  g16491(.A0(new_n18924_), .A1(new_n12614_), .B0(new_n18927_), .Y(new_n18928_));
  NOR2X1   g16492(.A(new_n18928_), .B(new_n18926_), .Y(new_n18929_));
  MX2X1    g16493(.A(new_n18929_), .B(new_n18924_), .S0(new_n11887_), .Y(new_n18930_));
  OAI21X1  g16494(.A0(new_n18880_), .A1(pi0619), .B0(pi1159), .Y(new_n18931_));
  AOI21X1  g16495(.A0(new_n18930_), .A1(pi0619), .B0(new_n18931_), .Y(new_n18932_));
  OAI21X1  g16496(.A0(new_n18880_), .A1(new_n12637_), .B0(new_n12638_), .Y(new_n18933_));
  AOI21X1  g16497(.A0(new_n18930_), .A1(new_n12637_), .B0(new_n18933_), .Y(new_n18934_));
  NOR2X1   g16498(.A(new_n18934_), .B(new_n18932_), .Y(new_n18935_));
  MX2X1    g16499(.A(new_n18935_), .B(new_n18930_), .S0(new_n11886_), .Y(new_n18936_));
  MX2X1    g16500(.A(new_n18936_), .B(new_n18879_), .S0(new_n12841_), .Y(new_n18937_));
  MX2X1    g16501(.A(new_n18937_), .B(new_n18879_), .S0(new_n12711_), .Y(new_n18938_));
  MX2X1    g16502(.A(new_n18938_), .B(new_n18879_), .S0(new_n12735_), .Y(new_n18939_));
  OAI21X1  g16503(.A0(new_n18880_), .A1(pi0644), .B0(new_n12739_), .Y(new_n18940_));
  AOI21X1  g16504(.A0(new_n18939_), .A1(pi0644), .B0(new_n18940_), .Y(new_n18941_));
  OR2X1    g16505(.A(new_n18941_), .B(new_n11882_), .Y(new_n18942_));
  AOI21X1  g16506(.A0(new_n18910_), .A1(pi0644), .B0(pi0715), .Y(new_n18943_));
  OAI21X1  g16507(.A0(new_n18880_), .A1(new_n12743_), .B0(pi0715), .Y(new_n18944_));
  AOI21X1  g16508(.A0(new_n18939_), .A1(new_n12743_), .B0(new_n18944_), .Y(new_n18945_));
  OR2X1    g16509(.A(new_n18945_), .B(pi1160), .Y(new_n18946_));
  OAI22X1  g16510(.A0(new_n18946_), .A1(new_n18943_), .B0(new_n18942_), .B1(new_n18911_), .Y(new_n18947_));
  NOR3X1   g16511(.A(new_n18945_), .B(pi1160), .C(pi0644), .Y(new_n18948_));
  NOR3X1   g16512(.A(new_n18941_), .B(new_n11882_), .C(new_n12743_), .Y(new_n18949_));
  NOR3X1   g16513(.A(new_n18949_), .B(new_n18948_), .C(new_n12897_), .Y(new_n18950_));
  MX2X1    g16514(.A(new_n18904_), .B(new_n18902_), .S0(new_n12689_), .Y(new_n18951_));
  OAI21X1  g16515(.A0(new_n18937_), .A1(new_n14395_), .B0(new_n18951_), .Y(new_n18952_));
  NAND2X1  g16516(.A(new_n18952_), .B(pi0792), .Y(new_n18953_));
  OR2X1    g16517(.A(new_n18917_), .B(new_n15335_), .Y(new_n18954_));
  OAI21X1  g16518(.A0(new_n12349_), .A1(new_n8717_), .B0(pi0777), .Y(new_n18955_));
  AOI21X1  g16519(.A0(new_n12289_), .A1(new_n8717_), .B0(new_n18955_), .Y(new_n18956_));
  OAI21X1  g16520(.A0(new_n12440_), .A1(pi0184), .B0(new_n15329_), .Y(new_n18957_));
  AOI21X1  g16521(.A0(new_n12401_), .A1(pi0184), .B0(new_n18957_), .Y(new_n18958_));
  OR2X1    g16522(.A(new_n18958_), .B(new_n2959_), .Y(new_n18959_));
  AND2X1   g16523(.A(new_n12467_), .B(pi0184), .Y(new_n18960_));
  OAI21X1  g16524(.A0(new_n12454_), .A1(pi0184), .B0(pi0777), .Y(new_n18961_));
  NOR4X1   g16525(.A(new_n13391_), .B(new_n12908_), .C(new_n12907_), .D(pi0184), .Y(new_n18962_));
  OAI21X1  g16526(.A0(new_n12929_), .A1(new_n8717_), .B0(new_n15329_), .Y(new_n18963_));
  OAI22X1  g16527(.A0(new_n18963_), .A1(new_n18962_), .B0(new_n18961_), .B1(new_n18960_), .Y(new_n18964_));
  AOI21X1  g16528(.A0(new_n18964_), .A1(new_n2959_), .B0(pi0038), .Y(new_n18965_));
  OAI21X1  g16529(.A0(new_n18959_), .A1(new_n18956_), .B0(new_n18965_), .Y(new_n18966_));
  OAI21X1  g16530(.A0(new_n12478_), .A1(pi0777), .B0(new_n13669_), .Y(new_n18967_));
  NAND2X1  g16531(.A(new_n18967_), .B(new_n8717_), .Y(new_n18968_));
  AOI21X1  g16532(.A0(new_n18762_), .A1(new_n14209_), .B0(new_n8717_), .Y(new_n18969_));
  AOI21X1  g16533(.A0(new_n18969_), .A1(new_n6857_), .B0(new_n2996_), .Y(new_n18970_));
  AOI21X1  g16534(.A0(new_n18970_), .A1(new_n18968_), .B0(pi0737), .Y(new_n18971_));
  AOI21X1  g16535(.A0(new_n18971_), .A1(new_n18966_), .B0(new_n3810_), .Y(new_n18972_));
  AOI22X1  g16536(.A0(new_n18972_), .A1(new_n18954_), .B0(new_n3810_), .B1(pi0184), .Y(new_n18973_));
  OAI21X1  g16537(.A0(new_n18918_), .A1(new_n12493_), .B0(new_n12494_), .Y(new_n18974_));
  AOI21X1  g16538(.A0(new_n18973_), .A1(new_n12493_), .B0(new_n18974_), .Y(new_n18975_));
  NAND2X1  g16539(.A(new_n18889_), .B(new_n12584_), .Y(new_n18976_));
  OAI21X1  g16540(.A0(new_n18918_), .A1(pi0625), .B0(pi1153), .Y(new_n18977_));
  AOI21X1  g16541(.A0(new_n18973_), .A1(pi0625), .B0(new_n18977_), .Y(new_n18978_));
  NAND2X1  g16542(.A(new_n18891_), .B(pi0608), .Y(new_n18979_));
  OAI22X1  g16543(.A0(new_n18979_), .A1(new_n18978_), .B0(new_n18976_), .B1(new_n18975_), .Y(new_n18980_));
  MX2X1    g16544(.A(new_n18980_), .B(new_n18973_), .S0(new_n11889_), .Y(new_n18981_));
  INVX1    g16545(.A(new_n18893_), .Y(new_n18982_));
  OAI21X1  g16546(.A0(new_n18982_), .A1(new_n12590_), .B0(new_n12591_), .Y(new_n18983_));
  AOI21X1  g16547(.A0(new_n18981_), .A1(new_n12590_), .B0(new_n18983_), .Y(new_n18984_));
  OAI21X1  g16548(.A0(new_n18921_), .A1(new_n12591_), .B0(new_n12596_), .Y(new_n18985_));
  OAI21X1  g16549(.A0(new_n18982_), .A1(pi0609), .B0(pi1155), .Y(new_n18986_));
  AOI21X1  g16550(.A0(new_n18981_), .A1(pi0609), .B0(new_n18986_), .Y(new_n18987_));
  OAI21X1  g16551(.A0(new_n18922_), .A1(pi1155), .B0(pi0660), .Y(new_n18988_));
  OAI22X1  g16552(.A0(new_n18988_), .A1(new_n18987_), .B0(new_n18985_), .B1(new_n18984_), .Y(new_n18989_));
  MX2X1    g16553(.A(new_n18989_), .B(new_n18981_), .S0(new_n11888_), .Y(new_n18990_));
  OAI21X1  g16554(.A0(new_n18895_), .A1(new_n12614_), .B0(new_n12615_), .Y(new_n18991_));
  AOI21X1  g16555(.A0(new_n18990_), .A1(new_n12614_), .B0(new_n18991_), .Y(new_n18992_));
  OR2X1    g16556(.A(new_n18926_), .B(pi0627), .Y(new_n18993_));
  OAI21X1  g16557(.A0(new_n18895_), .A1(pi0618), .B0(pi1154), .Y(new_n18994_));
  AOI21X1  g16558(.A0(new_n18990_), .A1(pi0618), .B0(new_n18994_), .Y(new_n18995_));
  OR2X1    g16559(.A(new_n18928_), .B(new_n12622_), .Y(new_n18996_));
  OAI22X1  g16560(.A0(new_n18996_), .A1(new_n18995_), .B0(new_n18993_), .B1(new_n18992_), .Y(new_n18997_));
  MX2X1    g16561(.A(new_n18997_), .B(new_n18990_), .S0(new_n11887_), .Y(new_n18998_));
  NAND2X1  g16562(.A(new_n18998_), .B(new_n12637_), .Y(new_n18999_));
  AOI21X1  g16563(.A0(new_n18897_), .A1(pi0619), .B0(pi1159), .Y(new_n19000_));
  OR2X1    g16564(.A(new_n18932_), .B(pi0648), .Y(new_n19001_));
  AOI21X1  g16565(.A0(new_n19000_), .A1(new_n18999_), .B0(new_n19001_), .Y(new_n19002_));
  NAND2X1  g16566(.A(new_n18998_), .B(pi0619), .Y(new_n19003_));
  AOI21X1  g16567(.A0(new_n18897_), .A1(new_n12637_), .B0(new_n12638_), .Y(new_n19004_));
  OR2X1    g16568(.A(new_n18934_), .B(new_n12645_), .Y(new_n19005_));
  AOI21X1  g16569(.A0(new_n19004_), .A1(new_n19003_), .B0(new_n19005_), .Y(new_n19006_));
  NOR3X1   g16570(.A(new_n19006_), .B(new_n19002_), .C(new_n11886_), .Y(new_n19007_));
  OAI21X1  g16571(.A0(new_n18998_), .A1(pi0789), .B0(new_n12842_), .Y(new_n19008_));
  AOI21X1  g16572(.A0(new_n18880_), .A1(pi0626), .B0(new_n16352_), .Y(new_n19009_));
  OAI21X1  g16573(.A0(new_n18936_), .A1(pi0626), .B0(new_n19009_), .Y(new_n19010_));
  AOI21X1  g16574(.A0(new_n18880_), .A1(new_n12664_), .B0(new_n16356_), .Y(new_n19011_));
  OAI21X1  g16575(.A0(new_n18936_), .A1(new_n12664_), .B0(new_n19011_), .Y(new_n19012_));
  NAND2X1  g16576(.A(new_n18898_), .B(new_n12769_), .Y(new_n19013_));
  NAND3X1  g16577(.A(new_n19013_), .B(new_n19012_), .C(new_n19010_), .Y(new_n19014_));
  AOI21X1  g16578(.A0(new_n19014_), .A1(pi0788), .B0(new_n14273_), .Y(new_n19015_));
  OAI21X1  g16579(.A0(new_n19008_), .A1(new_n19007_), .B0(new_n19015_), .Y(new_n19016_));
  AOI21X1  g16580(.A0(new_n19016_), .A1(new_n18953_), .B0(new_n14269_), .Y(new_n19017_));
  OR2X1    g16581(.A(new_n18938_), .B(new_n14384_), .Y(new_n19018_));
  OR2X1    g16582(.A(new_n18907_), .B(new_n14389_), .Y(new_n19019_));
  OR2X1    g16583(.A(new_n18908_), .B(new_n14387_), .Y(new_n19020_));
  NAND3X1  g16584(.A(new_n19020_), .B(new_n19019_), .C(new_n19018_), .Y(new_n19021_));
  AND2X1   g16585(.A(new_n19021_), .B(pi0787), .Y(new_n19022_));
  NOR3X1   g16586(.A(new_n19022_), .B(new_n19017_), .C(new_n18950_), .Y(new_n19023_));
  AOI21X1  g16587(.A0(new_n18947_), .A1(pi0790), .B0(new_n19023_), .Y(new_n19024_));
  OR2X1    g16588(.A(new_n19024_), .B(po1038), .Y(new_n19025_));
  AOI21X1  g16589(.A0(po1038), .A1(new_n8717_), .B0(pi0832), .Y(new_n19026_));
  AOI22X1  g16590(.A0(new_n19026_), .A1(new_n19025_), .B0(new_n18878_), .B1(new_n18877_), .Y(po0341));
  AOI21X1  g16591(.A0(pi1093), .A1(pi1092), .B0(pi0185), .Y(new_n19028_));
  INVX1    g16592(.A(new_n19028_), .Y(new_n19029_));
  AOI21X1  g16593(.A0(new_n12178_), .A1(new_n14820_), .B0(new_n19028_), .Y(new_n19030_));
  AOI21X1  g16594(.A0(new_n12601_), .A1(new_n2739_), .B0(new_n19030_), .Y(new_n19031_));
  NAND2X1  g16595(.A(new_n12178_), .B(new_n14820_), .Y(new_n19032_));
  OAI21X1  g16596(.A0(new_n19032_), .A1(new_n13436_), .B0(new_n19031_), .Y(new_n19033_));
  AND2X1   g16597(.A(new_n19033_), .B(pi1155), .Y(new_n19034_));
  NOR2X1   g16598(.A(new_n19032_), .B(new_n13436_), .Y(new_n19035_));
  NOR3X1   g16599(.A(new_n19035_), .B(new_n19028_), .C(pi1155), .Y(new_n19036_));
  OAI21X1  g16600(.A0(new_n19036_), .A1(new_n19034_), .B0(pi0785), .Y(new_n19037_));
  OAI21X1  g16601(.A0(new_n19031_), .A1(pi0785), .B0(new_n19037_), .Y(new_n19038_));
  INVX1    g16602(.A(new_n19038_), .Y(new_n19039_));
  AOI21X1  g16603(.A0(new_n19039_), .A1(new_n12785_), .B0(new_n12615_), .Y(new_n19040_));
  AOI21X1  g16604(.A0(new_n19039_), .A1(new_n12788_), .B0(pi1154), .Y(new_n19041_));
  NOR2X1   g16605(.A(new_n19041_), .B(new_n19040_), .Y(new_n19042_));
  MX2X1    g16606(.A(new_n19042_), .B(new_n19039_), .S0(new_n11887_), .Y(new_n19043_));
  OR2X1    g16607(.A(new_n19043_), .B(pi0789), .Y(new_n19044_));
  AOI21X1  g16608(.A0(new_n19043_), .A1(new_n15910_), .B0(new_n12638_), .Y(new_n19045_));
  AOI21X1  g16609(.A0(new_n19043_), .A1(new_n15912_), .B0(pi1159), .Y(new_n19046_));
  OAI21X1  g16610(.A0(new_n19046_), .A1(new_n19045_), .B0(pi0789), .Y(new_n19047_));
  AND2X1   g16611(.A(new_n19047_), .B(new_n19044_), .Y(new_n19048_));
  INVX1    g16612(.A(new_n19048_), .Y(new_n19049_));
  MX2X1    g16613(.A(new_n19049_), .B(new_n19029_), .S0(new_n12841_), .Y(new_n19050_));
  MX2X1    g16614(.A(new_n19050_), .B(new_n19029_), .S0(new_n12711_), .Y(new_n19051_));
  AOI21X1  g16615(.A0(new_n12566_), .A1(new_n14840_), .B0(new_n19028_), .Y(new_n19052_));
  INVX1    g16616(.A(new_n19052_), .Y(new_n19053_));
  NOR3X1   g16617(.A(new_n13585_), .B(pi0701), .C(pi0625), .Y(new_n19054_));
  OR2X1    g16618(.A(new_n19054_), .B(new_n19052_), .Y(new_n19055_));
  NOR2X1   g16619(.A(new_n19028_), .B(pi1153), .Y(new_n19056_));
  INVX1    g16620(.A(new_n19056_), .Y(new_n19057_));
  OAI21X1  g16621(.A0(new_n19057_), .A1(new_n19054_), .B0(pi0778), .Y(new_n19058_));
  AOI21X1  g16622(.A0(new_n19055_), .A1(pi1153), .B0(new_n19058_), .Y(new_n19059_));
  AOI21X1  g16623(.A0(new_n19053_), .A1(new_n11889_), .B0(new_n19059_), .Y(new_n19060_));
  NOR4X1   g16624(.A(new_n19060_), .B(new_n12765_), .C(new_n12764_), .D(new_n12762_), .Y(new_n19061_));
  INVX1    g16625(.A(new_n19061_), .Y(new_n19062_));
  NOR3X1   g16626(.A(new_n19062_), .B(new_n12870_), .C(new_n12851_), .Y(new_n19063_));
  INVX1    g16627(.A(new_n19063_), .Y(new_n19064_));
  AOI21X1  g16628(.A0(new_n19028_), .A1(pi0647), .B0(pi1157), .Y(new_n19065_));
  OAI21X1  g16629(.A0(new_n19064_), .A1(pi0647), .B0(new_n19065_), .Y(new_n19066_));
  MX2X1    g16630(.A(new_n19063_), .B(new_n19028_), .S0(new_n12705_), .Y(new_n19067_));
  OAI22X1  g16631(.A0(new_n19067_), .A1(new_n14387_), .B0(new_n19066_), .B1(new_n12723_), .Y(new_n19068_));
  AOI21X1  g16632(.A0(new_n19051_), .A1(new_n14385_), .B0(new_n19068_), .Y(new_n19069_));
  NOR2X1   g16633(.A(new_n19069_), .B(new_n11883_), .Y(new_n19070_));
  AOI21X1  g16634(.A0(new_n19029_), .A1(pi0626), .B0(new_n16352_), .Y(new_n19071_));
  OAI21X1  g16635(.A0(new_n19048_), .A1(pi0626), .B0(new_n19071_), .Y(new_n19072_));
  AOI21X1  g16636(.A0(new_n19047_), .A1(new_n19044_), .B0(new_n12664_), .Y(new_n19073_));
  NOR2X1   g16637(.A(new_n19028_), .B(pi0626), .Y(new_n19074_));
  NOR3X1   g16638(.A(new_n19074_), .B(new_n19073_), .C(new_n16356_), .Y(new_n19075_));
  AOI21X1  g16639(.A0(new_n19061_), .A1(new_n12769_), .B0(new_n19075_), .Y(new_n19076_));
  AOI21X1  g16640(.A0(new_n19076_), .A1(new_n19072_), .B0(new_n11885_), .Y(new_n19077_));
  INVX1    g16641(.A(new_n19030_), .Y(new_n19078_));
  AOI21X1  g16642(.A0(new_n19053_), .A1(new_n12171_), .B0(new_n19078_), .Y(new_n19079_));
  NOR3X1   g16643(.A(new_n19052_), .B(new_n12120_), .C(new_n12493_), .Y(new_n19080_));
  OR2X1    g16644(.A(new_n19079_), .B(new_n19080_), .Y(new_n19081_));
  NOR2X1   g16645(.A(new_n19054_), .B(new_n19052_), .Y(new_n19082_));
  OAI21X1  g16646(.A0(new_n19082_), .A1(new_n12494_), .B0(new_n12584_), .Y(new_n19083_));
  AOI21X1  g16647(.A0(new_n19081_), .A1(new_n19056_), .B0(new_n19083_), .Y(new_n19084_));
  NOR3X1   g16648(.A(new_n19080_), .B(new_n19078_), .C(new_n12494_), .Y(new_n19085_));
  OAI21X1  g16649(.A0(new_n19057_), .A1(new_n19054_), .B0(pi0608), .Y(new_n19086_));
  NOR2X1   g16650(.A(new_n19086_), .B(new_n19085_), .Y(new_n19087_));
  OAI21X1  g16651(.A0(new_n19087_), .A1(new_n19084_), .B0(pi0778), .Y(new_n19088_));
  OAI21X1  g16652(.A0(new_n19079_), .A1(pi0778), .B0(new_n19088_), .Y(new_n19089_));
  OAI21X1  g16653(.A0(new_n19060_), .A1(new_n12590_), .B0(new_n12591_), .Y(new_n19090_));
  AOI21X1  g16654(.A0(new_n19089_), .A1(new_n12590_), .B0(new_n19090_), .Y(new_n19091_));
  NOR3X1   g16655(.A(new_n19091_), .B(new_n19034_), .C(pi0660), .Y(new_n19092_));
  OAI21X1  g16656(.A0(new_n19060_), .A1(pi0609), .B0(pi1155), .Y(new_n19093_));
  AOI21X1  g16657(.A0(new_n19089_), .A1(pi0609), .B0(new_n19093_), .Y(new_n19094_));
  NOR3X1   g16658(.A(new_n19094_), .B(new_n19036_), .C(new_n12596_), .Y(new_n19095_));
  OAI21X1  g16659(.A0(new_n19095_), .A1(new_n19092_), .B0(pi0785), .Y(new_n19096_));
  NAND2X1  g16660(.A(new_n19089_), .B(new_n11888_), .Y(new_n19097_));
  AND2X1   g16661(.A(new_n19097_), .B(new_n19096_), .Y(new_n19098_));
  NOR3X1   g16662(.A(new_n19060_), .B(new_n12762_), .C(new_n12614_), .Y(new_n19099_));
  NOR2X1   g16663(.A(new_n19099_), .B(pi1154), .Y(new_n19100_));
  OAI21X1  g16664(.A0(new_n19098_), .A1(pi0618), .B0(new_n19100_), .Y(new_n19101_));
  NOR2X1   g16665(.A(new_n19040_), .B(pi0627), .Y(new_n19102_));
  NOR3X1   g16666(.A(new_n19060_), .B(new_n12762_), .C(pi0618), .Y(new_n19103_));
  NOR2X1   g16667(.A(new_n19103_), .B(new_n12615_), .Y(new_n19104_));
  OAI21X1  g16668(.A0(new_n19098_), .A1(new_n12614_), .B0(new_n19104_), .Y(new_n19105_));
  NOR2X1   g16669(.A(new_n19041_), .B(new_n12622_), .Y(new_n19106_));
  AOI22X1  g16670(.A0(new_n19106_), .A1(new_n19105_), .B0(new_n19102_), .B1(new_n19101_), .Y(new_n19107_));
  MX2X1    g16671(.A(new_n19107_), .B(new_n19098_), .S0(new_n11887_), .Y(new_n19108_));
  OR4X1    g16672(.A(new_n19060_), .B(new_n12764_), .C(new_n12762_), .D(new_n12637_), .Y(new_n19109_));
  AND2X1   g16673(.A(new_n19109_), .B(new_n12638_), .Y(new_n19110_));
  OAI21X1  g16674(.A0(new_n19108_), .A1(pi0619), .B0(new_n19110_), .Y(new_n19111_));
  NOR2X1   g16675(.A(new_n19045_), .B(pi0648), .Y(new_n19112_));
  AND2X1   g16676(.A(new_n19112_), .B(new_n19111_), .Y(new_n19113_));
  INVX1    g16677(.A(new_n19113_), .Y(new_n19114_));
  NOR4X1   g16678(.A(new_n19060_), .B(new_n12764_), .C(new_n12762_), .D(pi0619), .Y(new_n19115_));
  NOR2X1   g16679(.A(new_n19115_), .B(new_n12638_), .Y(new_n19116_));
  OAI21X1  g16680(.A0(new_n19108_), .A1(new_n12637_), .B0(new_n19116_), .Y(new_n19117_));
  NOR2X1   g16681(.A(new_n19046_), .B(new_n12645_), .Y(new_n19118_));
  AOI21X1  g16682(.A0(new_n19118_), .A1(new_n19117_), .B0(new_n11886_), .Y(new_n19119_));
  AOI21X1  g16683(.A0(new_n19108_), .A1(new_n11886_), .B0(new_n14264_), .Y(new_n19120_));
  INVX1    g16684(.A(new_n19120_), .Y(new_n19121_));
  AOI21X1  g16685(.A0(new_n19119_), .A1(new_n19114_), .B0(new_n19121_), .Y(new_n19122_));
  OAI21X1  g16686(.A0(new_n19122_), .A1(new_n19077_), .B0(new_n16350_), .Y(new_n19123_));
  INVX1    g16687(.A(new_n19050_), .Y(new_n19124_));
  AND2X1   g16688(.A(new_n19061_), .B(new_n12852_), .Y(new_n19125_));
  AOI22X1  g16689(.A0(new_n19125_), .A1(new_n14564_), .B0(new_n19124_), .B1(new_n12867_), .Y(new_n19126_));
  AOI22X1  g16690(.A0(new_n19125_), .A1(new_n14566_), .B0(new_n19124_), .B1(new_n12865_), .Y(new_n19127_));
  MX2X1    g16691(.A(new_n19127_), .B(new_n19126_), .S0(new_n12689_), .Y(new_n19128_));
  OAI21X1  g16692(.A0(new_n19128_), .A1(new_n11884_), .B0(new_n14562_), .Y(new_n19129_));
  INVX1    g16693(.A(new_n19129_), .Y(new_n19130_));
  AOI21X1  g16694(.A0(new_n19130_), .A1(new_n19123_), .B0(new_n19070_), .Y(new_n19131_));
  OAI21X1  g16695(.A0(new_n19067_), .A1(new_n12706_), .B0(new_n19066_), .Y(new_n19132_));
  MX2X1    g16696(.A(new_n19132_), .B(new_n19064_), .S0(new_n11883_), .Y(new_n19133_));
  OAI21X1  g16697(.A0(new_n19133_), .A1(pi0644), .B0(pi0715), .Y(new_n19134_));
  AOI21X1  g16698(.A0(new_n19131_), .A1(pi0644), .B0(new_n19134_), .Y(new_n19135_));
  OR4X1    g16699(.A(new_n12734_), .B(new_n2739_), .C(new_n11883_), .D(pi0185), .Y(new_n19136_));
  OAI21X1  g16700(.A0(new_n19051_), .A1(new_n12735_), .B0(new_n19136_), .Y(new_n19137_));
  OAI21X1  g16701(.A0(new_n19029_), .A1(pi0644), .B0(new_n12739_), .Y(new_n19138_));
  AOI21X1  g16702(.A0(new_n19137_), .A1(pi0644), .B0(new_n19138_), .Y(new_n19139_));
  OR2X1    g16703(.A(new_n19139_), .B(new_n11882_), .Y(new_n19140_));
  OAI21X1  g16704(.A0(new_n19133_), .A1(new_n12743_), .B0(new_n12739_), .Y(new_n19141_));
  AOI21X1  g16705(.A0(new_n19131_), .A1(new_n12743_), .B0(new_n19141_), .Y(new_n19142_));
  OAI21X1  g16706(.A0(new_n19029_), .A1(new_n12743_), .B0(pi0715), .Y(new_n19143_));
  AOI21X1  g16707(.A0(new_n19137_), .A1(new_n12743_), .B0(new_n19143_), .Y(new_n19144_));
  OR2X1    g16708(.A(new_n19144_), .B(pi1160), .Y(new_n19145_));
  OAI22X1  g16709(.A0(new_n19145_), .A1(new_n19142_), .B0(new_n19140_), .B1(new_n19135_), .Y(new_n19146_));
  NAND2X1  g16710(.A(new_n19146_), .B(pi0790), .Y(new_n19147_));
  AOI21X1  g16711(.A0(new_n19131_), .A1(new_n12897_), .B0(new_n12898_), .Y(new_n19148_));
  AOI21X1  g16712(.A0(new_n13699_), .A1(new_n3129_), .B0(pi0185), .Y(new_n19149_));
  INVX1    g16713(.A(new_n19149_), .Y(new_n19150_));
  OAI21X1  g16714(.A0(new_n3810_), .A1(pi0701), .B0(new_n19149_), .Y(new_n19151_));
  AOI21X1  g16715(.A0(new_n12955_), .A1(pi0185), .B0(pi0038), .Y(new_n19152_));
  OAI22X1  g16716(.A0(new_n19152_), .A1(new_n3810_), .B0(new_n12953_), .B1(pi0185), .Y(new_n19153_));
  OAI21X1  g16717(.A0(new_n12202_), .A1(pi0185), .B0(new_n12567_), .Y(new_n19154_));
  NAND3X1  g16718(.A(new_n19154_), .B(new_n19153_), .C(new_n14840_), .Y(new_n19155_));
  AND2X1   g16719(.A(new_n19155_), .B(new_n19151_), .Y(new_n19156_));
  INVX1    g16720(.A(new_n19156_), .Y(new_n19157_));
  AOI21X1  g16721(.A0(new_n19149_), .A1(new_n12493_), .B0(new_n12494_), .Y(new_n19158_));
  OAI21X1  g16722(.A0(new_n19156_), .A1(new_n12493_), .B0(new_n19158_), .Y(new_n19159_));
  AOI21X1  g16723(.A0(new_n19149_), .A1(pi0625), .B0(pi1153), .Y(new_n19160_));
  OAI21X1  g16724(.A0(new_n19156_), .A1(pi0625), .B0(new_n19160_), .Y(new_n19161_));
  AND2X1   g16725(.A(new_n19161_), .B(new_n19159_), .Y(new_n19162_));
  MX2X1    g16726(.A(new_n19162_), .B(new_n19157_), .S0(new_n11889_), .Y(new_n19163_));
  MX2X1    g16727(.A(new_n19163_), .B(new_n19149_), .S0(new_n12618_), .Y(new_n19164_));
  INVX1    g16728(.A(new_n19164_), .Y(new_n19165_));
  MX2X1    g16729(.A(new_n19165_), .B(new_n19150_), .S0(new_n12641_), .Y(new_n19166_));
  INVX1    g16730(.A(new_n19166_), .Y(new_n19167_));
  MX2X1    g16731(.A(new_n19167_), .B(new_n19149_), .S0(new_n12659_), .Y(new_n19168_));
  AND2X1   g16732(.A(new_n19149_), .B(new_n12691_), .Y(new_n19169_));
  AOI21X1  g16733(.A0(new_n19168_), .A1(new_n17252_), .B0(new_n19169_), .Y(new_n19170_));
  AOI21X1  g16734(.A0(new_n19149_), .A1(new_n12683_), .B0(new_n12684_), .Y(new_n19171_));
  OAI21X1  g16735(.A0(new_n19170_), .A1(new_n12683_), .B0(new_n19171_), .Y(new_n19172_));
  AOI21X1  g16736(.A0(new_n19149_), .A1(pi0628), .B0(pi1156), .Y(new_n19173_));
  OAI21X1  g16737(.A0(new_n19170_), .A1(pi0628), .B0(new_n19173_), .Y(new_n19174_));
  AOI21X1  g16738(.A0(new_n19174_), .A1(new_n19172_), .B0(new_n11884_), .Y(new_n19175_));
  AOI21X1  g16739(.A0(new_n19170_), .A1(new_n11884_), .B0(new_n19175_), .Y(new_n19176_));
  MX2X1    g16740(.A(new_n19176_), .B(new_n19149_), .S0(pi0647), .Y(new_n19177_));
  MX2X1    g16741(.A(new_n19176_), .B(new_n19149_), .S0(new_n12705_), .Y(new_n19178_));
  MX2X1    g16742(.A(new_n19178_), .B(new_n19177_), .S0(new_n12706_), .Y(new_n19179_));
  MX2X1    g16743(.A(new_n19179_), .B(new_n19176_), .S0(new_n11883_), .Y(new_n19180_));
  AOI21X1  g16744(.A0(new_n19180_), .A1(new_n12743_), .B0(new_n12739_), .Y(new_n19181_));
  OAI22X1  g16745(.A0(new_n12904_), .A1(new_n9996_), .B0(new_n12089_), .B1(new_n14820_), .Y(new_n19182_));
  OR2X1    g16746(.A(pi0751), .B(pi0185), .Y(new_n19183_));
  OAI22X1  g16747(.A0(new_n12168_), .A1(new_n9996_), .B0(new_n11948_), .B1(new_n14820_), .Y(new_n19184_));
  AOI22X1  g16748(.A0(new_n19184_), .A1(new_n2959_), .B0(pi0751), .B1(pi0185), .Y(new_n19185_));
  OAI21X1  g16749(.A0(new_n19183_), .A1(new_n12910_), .B0(new_n19185_), .Y(new_n19186_));
  AOI21X1  g16750(.A0(new_n19182_), .A1(pi0039), .B0(new_n19186_), .Y(new_n19187_));
  AOI21X1  g16751(.A0(new_n12901_), .A1(new_n9996_), .B0(new_n2996_), .Y(new_n19188_));
  OAI21X1  g16752(.A0(new_n14342_), .A1(pi0751), .B0(new_n19188_), .Y(new_n19189_));
  OAI21X1  g16753(.A0(new_n19187_), .A1(pi0038), .B0(new_n19189_), .Y(new_n19190_));
  MX2X1    g16754(.A(new_n19190_), .B(pi0185), .S0(new_n3810_), .Y(new_n19191_));
  AND2X1   g16755(.A(new_n19191_), .B(new_n12623_), .Y(new_n19192_));
  AOI21X1  g16756(.A0(new_n19150_), .A1(new_n12601_), .B0(new_n19192_), .Y(new_n19193_));
  AOI22X1  g16757(.A0(new_n19192_), .A1(pi0609), .B0(new_n19150_), .B1(new_n13430_), .Y(new_n19194_));
  AOI22X1  g16758(.A0(new_n19192_), .A1(new_n12590_), .B0(new_n19150_), .B1(new_n13436_), .Y(new_n19195_));
  MX2X1    g16759(.A(new_n19195_), .B(new_n19194_), .S0(pi1155), .Y(new_n19196_));
  MX2X1    g16760(.A(new_n19196_), .B(new_n19193_), .S0(new_n11888_), .Y(new_n19197_));
  OAI21X1  g16761(.A0(new_n19150_), .A1(pi0618), .B0(pi1154), .Y(new_n19198_));
  AOI21X1  g16762(.A0(new_n19197_), .A1(pi0618), .B0(new_n19198_), .Y(new_n19199_));
  OAI21X1  g16763(.A0(new_n19150_), .A1(new_n12614_), .B0(new_n12615_), .Y(new_n19200_));
  AOI21X1  g16764(.A0(new_n19197_), .A1(new_n12614_), .B0(new_n19200_), .Y(new_n19201_));
  NOR2X1   g16765(.A(new_n19201_), .B(new_n19199_), .Y(new_n19202_));
  MX2X1    g16766(.A(new_n19202_), .B(new_n19197_), .S0(new_n11887_), .Y(new_n19203_));
  OAI21X1  g16767(.A0(new_n19150_), .A1(pi0619), .B0(pi1159), .Y(new_n19204_));
  AOI21X1  g16768(.A0(new_n19203_), .A1(pi0619), .B0(new_n19204_), .Y(new_n19205_));
  OAI21X1  g16769(.A0(new_n19150_), .A1(new_n12637_), .B0(new_n12638_), .Y(new_n19206_));
  AOI21X1  g16770(.A0(new_n19203_), .A1(new_n12637_), .B0(new_n19206_), .Y(new_n19207_));
  NOR2X1   g16771(.A(new_n19207_), .B(new_n19205_), .Y(new_n19208_));
  MX2X1    g16772(.A(new_n19208_), .B(new_n19203_), .S0(new_n11886_), .Y(new_n19209_));
  MX2X1    g16773(.A(new_n19209_), .B(new_n19149_), .S0(new_n12841_), .Y(new_n19210_));
  MX2X1    g16774(.A(new_n19210_), .B(new_n19149_), .S0(new_n12711_), .Y(new_n19211_));
  MX2X1    g16775(.A(new_n19211_), .B(new_n19149_), .S0(new_n12735_), .Y(new_n19212_));
  OAI21X1  g16776(.A0(new_n19150_), .A1(pi0644), .B0(new_n12739_), .Y(new_n19213_));
  AOI21X1  g16777(.A0(new_n19212_), .A1(pi0644), .B0(new_n19213_), .Y(new_n19214_));
  OR2X1    g16778(.A(new_n19214_), .B(new_n11882_), .Y(new_n19215_));
  AOI21X1  g16779(.A0(new_n19180_), .A1(pi0644), .B0(pi0715), .Y(new_n19216_));
  OAI21X1  g16780(.A0(new_n19150_), .A1(new_n12743_), .B0(pi0715), .Y(new_n19217_));
  AOI21X1  g16781(.A0(new_n19212_), .A1(new_n12743_), .B0(new_n19217_), .Y(new_n19218_));
  OR2X1    g16782(.A(new_n19218_), .B(pi1160), .Y(new_n19219_));
  OAI22X1  g16783(.A0(new_n19219_), .A1(new_n19216_), .B0(new_n19215_), .B1(new_n19181_), .Y(new_n19220_));
  NOR3X1   g16784(.A(new_n19218_), .B(pi1160), .C(pi0644), .Y(new_n19221_));
  NOR3X1   g16785(.A(new_n19214_), .B(new_n11882_), .C(new_n12743_), .Y(new_n19222_));
  NOR3X1   g16786(.A(new_n19222_), .B(new_n19221_), .C(new_n12897_), .Y(new_n19223_));
  MX2X1    g16787(.A(new_n19174_), .B(new_n19172_), .S0(new_n12689_), .Y(new_n19224_));
  OAI21X1  g16788(.A0(new_n19210_), .A1(new_n14395_), .B0(new_n19224_), .Y(new_n19225_));
  NAND2X1  g16789(.A(new_n19225_), .B(pi0792), .Y(new_n19226_));
  OR2X1    g16790(.A(new_n19190_), .B(new_n14840_), .Y(new_n19227_));
  OAI21X1  g16791(.A0(new_n12349_), .A1(new_n9996_), .B0(pi0751), .Y(new_n19228_));
  AOI21X1  g16792(.A0(new_n12289_), .A1(new_n9996_), .B0(new_n19228_), .Y(new_n19229_));
  OAI21X1  g16793(.A0(new_n12440_), .A1(pi0185), .B0(new_n14820_), .Y(new_n19230_));
  AOI21X1  g16794(.A0(new_n12401_), .A1(pi0185), .B0(new_n19230_), .Y(new_n19231_));
  OR2X1    g16795(.A(new_n19231_), .B(new_n2959_), .Y(new_n19232_));
  AND2X1   g16796(.A(new_n12467_), .B(pi0185), .Y(new_n19233_));
  OAI21X1  g16797(.A0(new_n12454_), .A1(pi0185), .B0(pi0751), .Y(new_n19234_));
  NOR4X1   g16798(.A(new_n13391_), .B(new_n12908_), .C(new_n12907_), .D(pi0185), .Y(new_n19235_));
  OAI21X1  g16799(.A0(new_n12929_), .A1(new_n9996_), .B0(new_n14820_), .Y(new_n19236_));
  OAI22X1  g16800(.A0(new_n19236_), .A1(new_n19235_), .B0(new_n19234_), .B1(new_n19233_), .Y(new_n19237_));
  AOI21X1  g16801(.A0(new_n19237_), .A1(new_n2959_), .B0(pi0038), .Y(new_n19238_));
  OAI21X1  g16802(.A0(new_n19232_), .A1(new_n19229_), .B0(new_n19238_), .Y(new_n19239_));
  OAI21X1  g16803(.A0(new_n12478_), .A1(pi0751), .B0(new_n13669_), .Y(new_n19240_));
  NAND2X1  g16804(.A(new_n19240_), .B(new_n9996_), .Y(new_n19241_));
  AOI21X1  g16805(.A0(new_n19032_), .A1(new_n14209_), .B0(new_n9996_), .Y(new_n19242_));
  AOI21X1  g16806(.A0(new_n19242_), .A1(new_n6857_), .B0(new_n2996_), .Y(new_n19243_));
  AOI21X1  g16807(.A0(new_n19243_), .A1(new_n19241_), .B0(pi0701), .Y(new_n19244_));
  AOI21X1  g16808(.A0(new_n19244_), .A1(new_n19239_), .B0(new_n3810_), .Y(new_n19245_));
  AOI22X1  g16809(.A0(new_n19245_), .A1(new_n19227_), .B0(new_n3810_), .B1(pi0185), .Y(new_n19246_));
  OAI21X1  g16810(.A0(new_n19191_), .A1(new_n12493_), .B0(new_n12494_), .Y(new_n19247_));
  AOI21X1  g16811(.A0(new_n19246_), .A1(new_n12493_), .B0(new_n19247_), .Y(new_n19248_));
  NAND2X1  g16812(.A(new_n19159_), .B(new_n12584_), .Y(new_n19249_));
  OAI21X1  g16813(.A0(new_n19191_), .A1(pi0625), .B0(pi1153), .Y(new_n19250_));
  AOI21X1  g16814(.A0(new_n19246_), .A1(pi0625), .B0(new_n19250_), .Y(new_n19251_));
  NAND2X1  g16815(.A(new_n19161_), .B(pi0608), .Y(new_n19252_));
  OAI22X1  g16816(.A0(new_n19252_), .A1(new_n19251_), .B0(new_n19249_), .B1(new_n19248_), .Y(new_n19253_));
  MX2X1    g16817(.A(new_n19253_), .B(new_n19246_), .S0(new_n11889_), .Y(new_n19254_));
  INVX1    g16818(.A(new_n19163_), .Y(new_n19255_));
  OAI21X1  g16819(.A0(new_n19255_), .A1(new_n12590_), .B0(new_n12591_), .Y(new_n19256_));
  AOI21X1  g16820(.A0(new_n19254_), .A1(new_n12590_), .B0(new_n19256_), .Y(new_n19257_));
  OAI21X1  g16821(.A0(new_n19194_), .A1(new_n12591_), .B0(new_n12596_), .Y(new_n19258_));
  OAI21X1  g16822(.A0(new_n19255_), .A1(pi0609), .B0(pi1155), .Y(new_n19259_));
  AOI21X1  g16823(.A0(new_n19254_), .A1(pi0609), .B0(new_n19259_), .Y(new_n19260_));
  OAI21X1  g16824(.A0(new_n19195_), .A1(pi1155), .B0(pi0660), .Y(new_n19261_));
  OAI22X1  g16825(.A0(new_n19261_), .A1(new_n19260_), .B0(new_n19258_), .B1(new_n19257_), .Y(new_n19262_));
  MX2X1    g16826(.A(new_n19262_), .B(new_n19254_), .S0(new_n11888_), .Y(new_n19263_));
  OAI21X1  g16827(.A0(new_n19165_), .A1(new_n12614_), .B0(new_n12615_), .Y(new_n19264_));
  AOI21X1  g16828(.A0(new_n19263_), .A1(new_n12614_), .B0(new_n19264_), .Y(new_n19265_));
  OR2X1    g16829(.A(new_n19199_), .B(pi0627), .Y(new_n19266_));
  OAI21X1  g16830(.A0(new_n19165_), .A1(pi0618), .B0(pi1154), .Y(new_n19267_));
  AOI21X1  g16831(.A0(new_n19263_), .A1(pi0618), .B0(new_n19267_), .Y(new_n19268_));
  OR2X1    g16832(.A(new_n19201_), .B(new_n12622_), .Y(new_n19269_));
  OAI22X1  g16833(.A0(new_n19269_), .A1(new_n19268_), .B0(new_n19266_), .B1(new_n19265_), .Y(new_n19270_));
  MX2X1    g16834(.A(new_n19270_), .B(new_n19263_), .S0(new_n11887_), .Y(new_n19271_));
  NAND2X1  g16835(.A(new_n19271_), .B(new_n12637_), .Y(new_n19272_));
  AOI21X1  g16836(.A0(new_n19167_), .A1(pi0619), .B0(pi1159), .Y(new_n19273_));
  OR2X1    g16837(.A(new_n19205_), .B(pi0648), .Y(new_n19274_));
  AOI21X1  g16838(.A0(new_n19273_), .A1(new_n19272_), .B0(new_n19274_), .Y(new_n19275_));
  NAND2X1  g16839(.A(new_n19271_), .B(pi0619), .Y(new_n19276_));
  AOI21X1  g16840(.A0(new_n19167_), .A1(new_n12637_), .B0(new_n12638_), .Y(new_n19277_));
  OR2X1    g16841(.A(new_n19207_), .B(new_n12645_), .Y(new_n19278_));
  AOI21X1  g16842(.A0(new_n19277_), .A1(new_n19276_), .B0(new_n19278_), .Y(new_n19279_));
  NOR3X1   g16843(.A(new_n19279_), .B(new_n19275_), .C(new_n11886_), .Y(new_n19280_));
  OAI21X1  g16844(.A0(new_n19271_), .A1(pi0789), .B0(new_n12842_), .Y(new_n19281_));
  AOI21X1  g16845(.A0(new_n19150_), .A1(pi0626), .B0(new_n16352_), .Y(new_n19282_));
  OAI21X1  g16846(.A0(new_n19209_), .A1(pi0626), .B0(new_n19282_), .Y(new_n19283_));
  AOI21X1  g16847(.A0(new_n19150_), .A1(new_n12664_), .B0(new_n16356_), .Y(new_n19284_));
  OAI21X1  g16848(.A0(new_n19209_), .A1(new_n12664_), .B0(new_n19284_), .Y(new_n19285_));
  NAND2X1  g16849(.A(new_n19168_), .B(new_n12769_), .Y(new_n19286_));
  NAND3X1  g16850(.A(new_n19286_), .B(new_n19285_), .C(new_n19283_), .Y(new_n19287_));
  AOI21X1  g16851(.A0(new_n19287_), .A1(pi0788), .B0(new_n14273_), .Y(new_n19288_));
  OAI21X1  g16852(.A0(new_n19281_), .A1(new_n19280_), .B0(new_n19288_), .Y(new_n19289_));
  AOI21X1  g16853(.A0(new_n19289_), .A1(new_n19226_), .B0(new_n14269_), .Y(new_n19290_));
  OR2X1    g16854(.A(new_n19211_), .B(new_n14384_), .Y(new_n19291_));
  OR2X1    g16855(.A(new_n19177_), .B(new_n14389_), .Y(new_n19292_));
  OR2X1    g16856(.A(new_n19178_), .B(new_n14387_), .Y(new_n19293_));
  NAND3X1  g16857(.A(new_n19293_), .B(new_n19292_), .C(new_n19291_), .Y(new_n19294_));
  AND2X1   g16858(.A(new_n19294_), .B(pi0787), .Y(new_n19295_));
  NOR3X1   g16859(.A(new_n19295_), .B(new_n19290_), .C(new_n19223_), .Y(new_n19296_));
  AOI21X1  g16860(.A0(new_n19220_), .A1(pi0790), .B0(new_n19296_), .Y(new_n19297_));
  OR2X1    g16861(.A(new_n19297_), .B(po1038), .Y(new_n19298_));
  AOI21X1  g16862(.A0(po1038), .A1(new_n9996_), .B0(pi0832), .Y(new_n19299_));
  AOI22X1  g16863(.A0(new_n19299_), .A1(new_n19298_), .B0(new_n19148_), .B1(new_n19147_), .Y(po0342));
  NOR2X1   g16864(.A(new_n13676_), .B(new_n15370_), .Y(new_n19301_));
  OAI21X1  g16865(.A0(new_n13674_), .A1(new_n6861_), .B0(new_n19301_), .Y(new_n19302_));
  AOI21X1  g16866(.A0(new_n13672_), .A1(new_n6861_), .B0(new_n19302_), .Y(new_n19303_));
  OAI21X1  g16867(.A0(new_n13694_), .A1(pi0186), .B0(new_n15370_), .Y(new_n19304_));
  AOI21X1  g16868(.A0(new_n13688_), .A1(pi0186), .B0(new_n19304_), .Y(new_n19305_));
  OR2X1    g16869(.A(new_n19305_), .B(new_n15364_), .Y(new_n19306_));
  OR2X1    g16870(.A(new_n19306_), .B(new_n19303_), .Y(new_n19307_));
  OAI21X1  g16871(.A0(new_n13699_), .A1(pi0186), .B0(pi0752), .Y(new_n19308_));
  AOI21X1  g16872(.A0(new_n12199_), .A1(new_n2996_), .B0(new_n6861_), .Y(new_n19309_));
  NOR2X1   g16873(.A(pi0752), .B(pi0186), .Y(new_n19310_));
  AOI21X1  g16874(.A0(new_n19310_), .A1(new_n13704_), .B0(new_n19309_), .Y(new_n19311_));
  OR2X1    g16875(.A(new_n19311_), .B(new_n13701_), .Y(new_n19312_));
  AND2X1   g16876(.A(new_n19312_), .B(new_n19308_), .Y(new_n19313_));
  AOI21X1  g16877(.A0(new_n19313_), .A1(new_n15364_), .B0(new_n3810_), .Y(new_n19314_));
  AOI22X1  g16878(.A0(new_n19314_), .A1(new_n19307_), .B0(new_n3810_), .B1(pi0186), .Y(new_n19315_));
  NAND2X1  g16879(.A(new_n19312_), .B(new_n19308_), .Y(new_n19316_));
  MX2X1    g16880(.A(new_n19316_), .B(pi0186), .S0(new_n3810_), .Y(new_n19317_));
  OAI21X1  g16881(.A0(new_n19317_), .A1(new_n12493_), .B0(new_n12494_), .Y(new_n19318_));
  AOI21X1  g16882(.A0(new_n19315_), .A1(new_n12493_), .B0(new_n19318_), .Y(new_n19319_));
  NAND3X1  g16883(.A(new_n12574_), .B(new_n15364_), .C(new_n6861_), .Y(new_n19320_));
  AOI21X1  g16884(.A0(new_n12955_), .A1(pi0186), .B0(pi0038), .Y(new_n19321_));
  OAI21X1  g16885(.A0(new_n12953_), .A1(pi0186), .B0(new_n19321_), .Y(new_n19322_));
  OR2X1    g16886(.A(new_n12202_), .B(pi0186), .Y(new_n19323_));
  AOI21X1  g16887(.A0(new_n19323_), .A1(new_n12567_), .B0(new_n15364_), .Y(new_n19324_));
  AOI21X1  g16888(.A0(new_n19324_), .A1(new_n19322_), .B0(new_n3810_), .Y(new_n19325_));
  AOI22X1  g16889(.A0(new_n19325_), .A1(new_n19320_), .B0(new_n3810_), .B1(pi0186), .Y(new_n19326_));
  OAI21X1  g16890(.A0(new_n12574_), .A1(new_n3810_), .B0(new_n6861_), .Y(new_n19327_));
  OAI21X1  g16891(.A0(new_n19327_), .A1(pi0625), .B0(pi1153), .Y(new_n19328_));
  AOI21X1  g16892(.A0(new_n19326_), .A1(pi0625), .B0(new_n19328_), .Y(new_n19329_));
  OR2X1    g16893(.A(new_n19329_), .B(pi0608), .Y(new_n19330_));
  OAI21X1  g16894(.A0(new_n19317_), .A1(pi0625), .B0(pi1153), .Y(new_n19331_));
  AOI21X1  g16895(.A0(new_n19315_), .A1(pi0625), .B0(new_n19331_), .Y(new_n19332_));
  OAI21X1  g16896(.A0(new_n19327_), .A1(new_n12493_), .B0(new_n12494_), .Y(new_n19333_));
  AOI21X1  g16897(.A0(new_n19326_), .A1(new_n12493_), .B0(new_n19333_), .Y(new_n19334_));
  OR2X1    g16898(.A(new_n19334_), .B(new_n12584_), .Y(new_n19335_));
  OAI22X1  g16899(.A0(new_n19335_), .A1(new_n19332_), .B0(new_n19330_), .B1(new_n19319_), .Y(new_n19336_));
  MX2X1    g16900(.A(new_n19336_), .B(new_n19315_), .S0(new_n11889_), .Y(new_n19337_));
  OAI21X1  g16901(.A0(new_n19334_), .A1(new_n19329_), .B0(pi0778), .Y(new_n19338_));
  OAI21X1  g16902(.A0(new_n19326_), .A1(pi0778), .B0(new_n19338_), .Y(new_n19339_));
  OAI21X1  g16903(.A0(new_n19339_), .A1(new_n12590_), .B0(new_n12591_), .Y(new_n19340_));
  AOI21X1  g16904(.A0(new_n19337_), .A1(new_n12590_), .B0(new_n19340_), .Y(new_n19341_));
  INVX1    g16905(.A(new_n19327_), .Y(new_n19342_));
  NAND2X1  g16906(.A(new_n19317_), .B(new_n12623_), .Y(new_n19343_));
  OAI22X1  g16907(.A0(new_n19343_), .A1(new_n12590_), .B0(new_n19342_), .B1(new_n12599_), .Y(new_n19344_));
  NAND2X1  g16908(.A(new_n19344_), .B(pi1155), .Y(new_n19345_));
  NAND2X1  g16909(.A(new_n19345_), .B(new_n12596_), .Y(new_n19346_));
  OAI21X1  g16910(.A0(new_n19339_), .A1(pi0609), .B0(pi1155), .Y(new_n19347_));
  AOI21X1  g16911(.A0(new_n19337_), .A1(pi0609), .B0(new_n19347_), .Y(new_n19348_));
  OAI22X1  g16912(.A0(new_n19343_), .A1(pi0609), .B0(new_n19342_), .B1(new_n12608_), .Y(new_n19349_));
  NAND2X1  g16913(.A(new_n19349_), .B(new_n12591_), .Y(new_n19350_));
  NAND2X1  g16914(.A(new_n19350_), .B(pi0660), .Y(new_n19351_));
  OAI22X1  g16915(.A0(new_n19351_), .A1(new_n19348_), .B0(new_n19346_), .B1(new_n19341_), .Y(new_n19352_));
  MX2X1    g16916(.A(new_n19352_), .B(new_n19337_), .S0(new_n11888_), .Y(new_n19353_));
  MX2X1    g16917(.A(new_n19339_), .B(new_n19327_), .S0(new_n12618_), .Y(new_n19354_));
  OAI21X1  g16918(.A0(new_n19354_), .A1(new_n12614_), .B0(new_n12615_), .Y(new_n19355_));
  AOI21X1  g16919(.A0(new_n19353_), .A1(new_n12614_), .B0(new_n19355_), .Y(new_n19356_));
  MX2X1    g16920(.A(new_n19327_), .B(new_n19317_), .S0(new_n12623_), .Y(new_n19357_));
  AOI21X1  g16921(.A0(new_n19350_), .A1(new_n19345_), .B0(new_n11888_), .Y(new_n19358_));
  AOI21X1  g16922(.A0(new_n19357_), .A1(new_n11888_), .B0(new_n19358_), .Y(new_n19359_));
  OAI21X1  g16923(.A0(new_n19327_), .A1(pi0618), .B0(pi1154), .Y(new_n19360_));
  AOI21X1  g16924(.A0(new_n19359_), .A1(pi0618), .B0(new_n19360_), .Y(new_n19361_));
  OR2X1    g16925(.A(new_n19361_), .B(pi0627), .Y(new_n19362_));
  OAI21X1  g16926(.A0(new_n19354_), .A1(pi0618), .B0(pi1154), .Y(new_n19363_));
  AOI21X1  g16927(.A0(new_n19353_), .A1(pi0618), .B0(new_n19363_), .Y(new_n19364_));
  OAI21X1  g16928(.A0(new_n19327_), .A1(new_n12614_), .B0(new_n12615_), .Y(new_n19365_));
  AOI21X1  g16929(.A0(new_n19359_), .A1(new_n12614_), .B0(new_n19365_), .Y(new_n19366_));
  OR2X1    g16930(.A(new_n19366_), .B(new_n12622_), .Y(new_n19367_));
  OAI22X1  g16931(.A0(new_n19367_), .A1(new_n19364_), .B0(new_n19362_), .B1(new_n19356_), .Y(new_n19368_));
  MX2X1    g16932(.A(new_n19368_), .B(new_n19353_), .S0(new_n11887_), .Y(new_n19369_));
  MX2X1    g16933(.A(new_n19354_), .B(new_n19327_), .S0(new_n12641_), .Y(new_n19370_));
  OAI21X1  g16934(.A0(new_n19370_), .A1(new_n12637_), .B0(new_n12638_), .Y(new_n19371_));
  AOI21X1  g16935(.A0(new_n19369_), .A1(new_n12637_), .B0(new_n19371_), .Y(new_n19372_));
  NOR2X1   g16936(.A(new_n19366_), .B(new_n19361_), .Y(new_n19373_));
  MX2X1    g16937(.A(new_n19373_), .B(new_n19359_), .S0(new_n11887_), .Y(new_n19374_));
  OAI21X1  g16938(.A0(new_n19327_), .A1(pi0619), .B0(pi1159), .Y(new_n19375_));
  AOI21X1  g16939(.A0(new_n19374_), .A1(pi0619), .B0(new_n19375_), .Y(new_n19376_));
  OR2X1    g16940(.A(new_n19376_), .B(pi0648), .Y(new_n19377_));
  OAI21X1  g16941(.A0(new_n19370_), .A1(pi0619), .B0(pi1159), .Y(new_n19378_));
  AOI21X1  g16942(.A0(new_n19369_), .A1(pi0619), .B0(new_n19378_), .Y(new_n19379_));
  OAI21X1  g16943(.A0(new_n19327_), .A1(new_n12637_), .B0(new_n12638_), .Y(new_n19380_));
  AOI21X1  g16944(.A0(new_n19374_), .A1(new_n12637_), .B0(new_n19380_), .Y(new_n19381_));
  OR2X1    g16945(.A(new_n19381_), .B(new_n12645_), .Y(new_n19382_));
  OAI22X1  g16946(.A0(new_n19382_), .A1(new_n19379_), .B0(new_n19377_), .B1(new_n19372_), .Y(new_n19383_));
  MX2X1    g16947(.A(new_n19383_), .B(new_n19369_), .S0(new_n11886_), .Y(new_n19384_));
  MX2X1    g16948(.A(new_n19370_), .B(new_n19327_), .S0(new_n12659_), .Y(new_n19385_));
  AOI21X1  g16949(.A0(new_n19385_), .A1(pi0626), .B0(pi0641), .Y(new_n19386_));
  OAI21X1  g16950(.A0(new_n19384_), .A1(pi0626), .B0(new_n19386_), .Y(new_n19387_));
  OR2X1    g16951(.A(new_n19374_), .B(pi0789), .Y(new_n19388_));
  OAI21X1  g16952(.A0(new_n19381_), .A1(new_n19376_), .B0(pi0789), .Y(new_n19389_));
  NAND2X1  g16953(.A(new_n19389_), .B(new_n19388_), .Y(new_n19390_));
  NAND2X1  g16954(.A(new_n19390_), .B(new_n12664_), .Y(new_n19391_));
  AOI21X1  g16955(.A0(new_n19327_), .A1(pi0626), .B0(new_n12672_), .Y(new_n19392_));
  AOI21X1  g16956(.A0(new_n19392_), .A1(new_n19391_), .B0(pi1158), .Y(new_n19393_));
  AOI21X1  g16957(.A0(new_n19385_), .A1(new_n12664_), .B0(new_n12672_), .Y(new_n19394_));
  OAI21X1  g16958(.A0(new_n19384_), .A1(new_n12664_), .B0(new_n19394_), .Y(new_n19395_));
  NAND2X1  g16959(.A(new_n19390_), .B(pi0626), .Y(new_n19396_));
  AOI21X1  g16960(.A0(new_n19327_), .A1(new_n12664_), .B0(pi0641), .Y(new_n19397_));
  AOI21X1  g16961(.A0(new_n19397_), .A1(new_n19396_), .B0(new_n12676_), .Y(new_n19398_));
  AOI22X1  g16962(.A0(new_n19398_), .A1(new_n19395_), .B0(new_n19393_), .B1(new_n19387_), .Y(new_n19399_));
  MX2X1    g16963(.A(new_n19399_), .B(new_n19384_), .S0(new_n11885_), .Y(new_n19400_));
  MX2X1    g16964(.A(new_n19390_), .B(new_n19327_), .S0(new_n12841_), .Y(new_n19401_));
  OAI21X1  g16965(.A0(new_n19401_), .A1(new_n12683_), .B0(new_n12684_), .Y(new_n19402_));
  AOI21X1  g16966(.A0(new_n19400_), .A1(new_n12683_), .B0(new_n19402_), .Y(new_n19403_));
  MX2X1    g16967(.A(new_n19385_), .B(new_n19327_), .S0(new_n12691_), .Y(new_n19404_));
  AOI21X1  g16968(.A0(new_n19342_), .A1(new_n12683_), .B0(new_n12684_), .Y(new_n19405_));
  OAI21X1  g16969(.A0(new_n19404_), .A1(new_n12683_), .B0(new_n19405_), .Y(new_n19406_));
  AND2X1   g16970(.A(new_n19406_), .B(new_n12689_), .Y(new_n19407_));
  INVX1    g16971(.A(new_n19407_), .Y(new_n19408_));
  OAI21X1  g16972(.A0(new_n19401_), .A1(pi0628), .B0(pi1156), .Y(new_n19409_));
  AOI21X1  g16973(.A0(new_n19400_), .A1(pi0628), .B0(new_n19409_), .Y(new_n19410_));
  AOI21X1  g16974(.A0(new_n19342_), .A1(pi0628), .B0(pi1156), .Y(new_n19411_));
  OAI21X1  g16975(.A0(new_n19404_), .A1(pi0628), .B0(new_n19411_), .Y(new_n19412_));
  AND2X1   g16976(.A(new_n19412_), .B(pi0629), .Y(new_n19413_));
  INVX1    g16977(.A(new_n19413_), .Y(new_n19414_));
  OAI22X1  g16978(.A0(new_n19414_), .A1(new_n19410_), .B0(new_n19408_), .B1(new_n19403_), .Y(new_n19415_));
  MX2X1    g16979(.A(new_n19415_), .B(new_n19400_), .S0(new_n11884_), .Y(new_n19416_));
  MX2X1    g16980(.A(new_n19401_), .B(new_n19327_), .S0(new_n12711_), .Y(new_n19417_));
  OAI21X1  g16981(.A0(new_n19417_), .A1(new_n12705_), .B0(new_n12706_), .Y(new_n19418_));
  AOI21X1  g16982(.A0(new_n19416_), .A1(new_n12705_), .B0(new_n19418_), .Y(new_n19419_));
  AOI21X1  g16983(.A0(new_n19412_), .A1(new_n19406_), .B0(new_n11884_), .Y(new_n19420_));
  AOI21X1  g16984(.A0(new_n19404_), .A1(new_n11884_), .B0(new_n19420_), .Y(new_n19421_));
  OAI21X1  g16985(.A0(new_n19327_), .A1(pi0647), .B0(pi1157), .Y(new_n19422_));
  AOI21X1  g16986(.A0(new_n19421_), .A1(pi0647), .B0(new_n19422_), .Y(new_n19423_));
  NOR2X1   g16987(.A(new_n19423_), .B(pi0630), .Y(new_n19424_));
  INVX1    g16988(.A(new_n19424_), .Y(new_n19425_));
  OAI21X1  g16989(.A0(new_n19417_), .A1(pi0647), .B0(pi1157), .Y(new_n19426_));
  AOI21X1  g16990(.A0(new_n19416_), .A1(pi0647), .B0(new_n19426_), .Y(new_n19427_));
  OAI21X1  g16991(.A0(new_n19327_), .A1(new_n12705_), .B0(new_n12706_), .Y(new_n19428_));
  AOI21X1  g16992(.A0(new_n19421_), .A1(new_n12705_), .B0(new_n19428_), .Y(new_n19429_));
  NOR2X1   g16993(.A(new_n19429_), .B(new_n12723_), .Y(new_n19430_));
  INVX1    g16994(.A(new_n19430_), .Y(new_n19431_));
  OAI22X1  g16995(.A0(new_n19431_), .A1(new_n19427_), .B0(new_n19425_), .B1(new_n19419_), .Y(new_n19432_));
  MX2X1    g16996(.A(new_n19432_), .B(new_n19416_), .S0(new_n11883_), .Y(new_n19433_));
  OAI21X1  g16997(.A0(new_n19429_), .A1(new_n19423_), .B0(pi0787), .Y(new_n19434_));
  OAI21X1  g16998(.A0(new_n19421_), .A1(pi0787), .B0(new_n19434_), .Y(new_n19435_));
  OAI21X1  g16999(.A0(new_n19435_), .A1(pi0644), .B0(pi0715), .Y(new_n19436_));
  AOI21X1  g17000(.A0(new_n19433_), .A1(pi0644), .B0(new_n19436_), .Y(new_n19437_));
  AND2X1   g17001(.A(new_n19327_), .B(new_n12735_), .Y(new_n19438_));
  AOI21X1  g17002(.A0(new_n19417_), .A1(new_n12736_), .B0(new_n19438_), .Y(new_n19439_));
  OAI21X1  g17003(.A0(new_n19327_), .A1(pi0644), .B0(new_n12739_), .Y(new_n19440_));
  AOI21X1  g17004(.A0(new_n19439_), .A1(pi0644), .B0(new_n19440_), .Y(new_n19441_));
  NOR3X1   g17005(.A(new_n19441_), .B(new_n19437_), .C(new_n11882_), .Y(new_n19442_));
  OAI21X1  g17006(.A0(new_n19435_), .A1(new_n12743_), .B0(new_n12739_), .Y(new_n19443_));
  AOI21X1  g17007(.A0(new_n19433_), .A1(new_n12743_), .B0(new_n19443_), .Y(new_n19444_));
  OAI21X1  g17008(.A0(new_n19327_), .A1(new_n12743_), .B0(pi0715), .Y(new_n19445_));
  AOI21X1  g17009(.A0(new_n19439_), .A1(new_n12743_), .B0(new_n19445_), .Y(new_n19446_));
  OR2X1    g17010(.A(new_n19446_), .B(pi1160), .Y(new_n19447_));
  OAI21X1  g17011(.A0(new_n19447_), .A1(new_n19444_), .B0(pi0790), .Y(new_n19448_));
  OR2X1    g17012(.A(new_n19433_), .B(pi0790), .Y(new_n19449_));
  AND2X1   g17013(.A(new_n19449_), .B(new_n6520_), .Y(new_n19450_));
  OAI21X1  g17014(.A0(new_n19448_), .A1(new_n19442_), .B0(new_n19450_), .Y(new_n19451_));
  AOI21X1  g17015(.A0(po1038), .A1(new_n6861_), .B0(pi0832), .Y(new_n19452_));
  AOI21X1  g17016(.A0(pi1093), .A1(pi1092), .B0(pi0186), .Y(new_n19453_));
  INVX1    g17017(.A(new_n19453_), .Y(new_n19454_));
  AOI21X1  g17018(.A0(new_n12178_), .A1(new_n15370_), .B0(new_n19453_), .Y(new_n19455_));
  AOI21X1  g17019(.A0(new_n12601_), .A1(new_n2739_), .B0(new_n19455_), .Y(new_n19456_));
  INVX1    g17020(.A(new_n19455_), .Y(new_n19457_));
  AOI21X1  g17021(.A0(new_n19457_), .A1(new_n12776_), .B0(new_n12591_), .Y(new_n19458_));
  AOI21X1  g17022(.A0(new_n19456_), .A1(new_n12779_), .B0(pi1155), .Y(new_n19459_));
  OAI21X1  g17023(.A0(new_n19459_), .A1(new_n19458_), .B0(pi0785), .Y(new_n19460_));
  OAI21X1  g17024(.A0(new_n19456_), .A1(pi0785), .B0(new_n19460_), .Y(new_n19461_));
  INVX1    g17025(.A(new_n19461_), .Y(new_n19462_));
  AOI21X1  g17026(.A0(new_n19462_), .A1(new_n12785_), .B0(new_n12615_), .Y(new_n19463_));
  AOI21X1  g17027(.A0(new_n19462_), .A1(new_n12788_), .B0(pi1154), .Y(new_n19464_));
  OR2X1    g17028(.A(new_n19464_), .B(new_n19463_), .Y(new_n19465_));
  MX2X1    g17029(.A(new_n19465_), .B(new_n19461_), .S0(new_n11887_), .Y(new_n19466_));
  AND2X1   g17030(.A(new_n19466_), .B(new_n11886_), .Y(new_n19467_));
  AOI21X1  g17031(.A0(new_n19453_), .A1(new_n12637_), .B0(new_n12638_), .Y(new_n19468_));
  OAI21X1  g17032(.A0(new_n19466_), .A1(new_n12637_), .B0(new_n19468_), .Y(new_n19469_));
  AOI21X1  g17033(.A0(new_n19453_), .A1(pi0619), .B0(pi1159), .Y(new_n19470_));
  OAI21X1  g17034(.A0(new_n19466_), .A1(pi0619), .B0(new_n19470_), .Y(new_n19471_));
  AOI21X1  g17035(.A0(new_n19471_), .A1(new_n19469_), .B0(new_n11886_), .Y(new_n19472_));
  NOR2X1   g17036(.A(new_n19472_), .B(new_n19467_), .Y(new_n19473_));
  INVX1    g17037(.A(new_n19473_), .Y(new_n19474_));
  MX2X1    g17038(.A(new_n19474_), .B(new_n19454_), .S0(new_n12841_), .Y(new_n19475_));
  MX2X1    g17039(.A(new_n19475_), .B(new_n19454_), .S0(new_n12711_), .Y(new_n19476_));
  AOI21X1  g17040(.A0(new_n12566_), .A1(pi0703), .B0(new_n19453_), .Y(new_n19477_));
  AND2X1   g17041(.A(new_n12566_), .B(pi0703), .Y(new_n19478_));
  AND2X1   g17042(.A(new_n19478_), .B(new_n12493_), .Y(new_n19479_));
  MX2X1    g17043(.A(new_n19453_), .B(pi0625), .S0(new_n19478_), .Y(new_n19480_));
  NOR2X1   g17044(.A(new_n19453_), .B(pi1153), .Y(new_n19481_));
  INVX1    g17045(.A(new_n19481_), .Y(new_n19482_));
  OAI22X1  g17046(.A0(new_n19482_), .A1(new_n19479_), .B0(new_n19480_), .B1(new_n12494_), .Y(new_n19483_));
  MX2X1    g17047(.A(new_n19483_), .B(new_n19477_), .S0(new_n11889_), .Y(new_n19484_));
  NOR4X1   g17048(.A(new_n19484_), .B(new_n12765_), .C(new_n12764_), .D(new_n12762_), .Y(new_n19485_));
  INVX1    g17049(.A(new_n19485_), .Y(new_n19486_));
  NOR3X1   g17050(.A(new_n19486_), .B(new_n12870_), .C(new_n12851_), .Y(new_n19487_));
  INVX1    g17051(.A(new_n19487_), .Y(new_n19488_));
  AOI21X1  g17052(.A0(new_n19453_), .A1(pi0647), .B0(pi1157), .Y(new_n19489_));
  OAI21X1  g17053(.A0(new_n19488_), .A1(pi0647), .B0(new_n19489_), .Y(new_n19490_));
  MX2X1    g17054(.A(new_n19487_), .B(new_n19453_), .S0(new_n12705_), .Y(new_n19491_));
  OAI22X1  g17055(.A0(new_n19491_), .A1(new_n14387_), .B0(new_n19490_), .B1(new_n12723_), .Y(new_n19492_));
  AOI21X1  g17056(.A0(new_n19476_), .A1(new_n14385_), .B0(new_n19492_), .Y(new_n19493_));
  AOI21X1  g17057(.A0(new_n19454_), .A1(pi0626), .B0(new_n16352_), .Y(new_n19494_));
  OAI21X1  g17058(.A0(new_n19473_), .A1(pi0626), .B0(new_n19494_), .Y(new_n19495_));
  AOI21X1  g17059(.A0(new_n19454_), .A1(new_n12664_), .B0(new_n16356_), .Y(new_n19496_));
  OAI21X1  g17060(.A0(new_n19473_), .A1(new_n12664_), .B0(new_n19496_), .Y(new_n19497_));
  NAND2X1  g17061(.A(new_n19485_), .B(new_n12769_), .Y(new_n19498_));
  NAND3X1  g17062(.A(new_n19498_), .B(new_n19497_), .C(new_n19495_), .Y(new_n19499_));
  AND2X1   g17063(.A(new_n19499_), .B(pi0788), .Y(new_n19500_));
  INVX1    g17064(.A(new_n19500_), .Y(new_n19501_));
  NOR2X1   g17065(.A(new_n19477_), .B(new_n12120_), .Y(new_n19502_));
  NOR2X1   g17066(.A(new_n19502_), .B(new_n19457_), .Y(new_n19503_));
  INVX1    g17067(.A(new_n19503_), .Y(new_n19504_));
  MX2X1    g17068(.A(new_n19457_), .B(new_n12493_), .S0(new_n19502_), .Y(new_n19505_));
  NOR2X1   g17069(.A(new_n19505_), .B(new_n19482_), .Y(new_n19506_));
  OAI21X1  g17070(.A0(new_n19480_), .A1(new_n12494_), .B0(new_n12584_), .Y(new_n19507_));
  NOR3X1   g17071(.A(new_n19477_), .B(new_n12120_), .C(new_n12493_), .Y(new_n19508_));
  NOR3X1   g17072(.A(new_n19508_), .B(new_n19457_), .C(new_n12494_), .Y(new_n19509_));
  OAI21X1  g17073(.A0(new_n19482_), .A1(new_n19479_), .B0(pi0608), .Y(new_n19510_));
  OAI22X1  g17074(.A0(new_n19510_), .A1(new_n19509_), .B0(new_n19507_), .B1(new_n19506_), .Y(new_n19511_));
  MX2X1    g17075(.A(new_n19511_), .B(new_n19504_), .S0(new_n11889_), .Y(new_n19512_));
  OAI21X1  g17076(.A0(new_n19484_), .A1(new_n12590_), .B0(new_n12591_), .Y(new_n19513_));
  AOI21X1  g17077(.A0(new_n19512_), .A1(new_n12590_), .B0(new_n19513_), .Y(new_n19514_));
  NOR3X1   g17078(.A(new_n19514_), .B(new_n19458_), .C(pi0660), .Y(new_n19515_));
  OAI21X1  g17079(.A0(new_n19484_), .A1(pi0609), .B0(pi1155), .Y(new_n19516_));
  AOI21X1  g17080(.A0(new_n19512_), .A1(pi0609), .B0(new_n19516_), .Y(new_n19517_));
  NOR3X1   g17081(.A(new_n19517_), .B(new_n19459_), .C(new_n12596_), .Y(new_n19518_));
  OAI21X1  g17082(.A0(new_n19518_), .A1(new_n19515_), .B0(pi0785), .Y(new_n19519_));
  NAND2X1  g17083(.A(new_n19512_), .B(new_n11888_), .Y(new_n19520_));
  AND2X1   g17084(.A(new_n19520_), .B(new_n19519_), .Y(new_n19521_));
  NOR3X1   g17085(.A(new_n19484_), .B(new_n12762_), .C(new_n12614_), .Y(new_n19522_));
  NOR2X1   g17086(.A(new_n19522_), .B(pi1154), .Y(new_n19523_));
  OAI21X1  g17087(.A0(new_n19521_), .A1(pi0618), .B0(new_n19523_), .Y(new_n19524_));
  NOR2X1   g17088(.A(new_n19463_), .B(pi0627), .Y(new_n19525_));
  NOR3X1   g17089(.A(new_n19484_), .B(new_n12762_), .C(pi0618), .Y(new_n19526_));
  NOR2X1   g17090(.A(new_n19526_), .B(new_n12615_), .Y(new_n19527_));
  OAI21X1  g17091(.A0(new_n19521_), .A1(new_n12614_), .B0(new_n19527_), .Y(new_n19528_));
  NOR2X1   g17092(.A(new_n19464_), .B(new_n12622_), .Y(new_n19529_));
  AOI22X1  g17093(.A0(new_n19529_), .A1(new_n19528_), .B0(new_n19525_), .B1(new_n19524_), .Y(new_n19530_));
  MX2X1    g17094(.A(new_n19530_), .B(new_n19521_), .S0(new_n11887_), .Y(new_n19531_));
  OR4X1    g17095(.A(new_n19484_), .B(new_n12764_), .C(new_n12762_), .D(new_n12637_), .Y(new_n19532_));
  AND2X1   g17096(.A(new_n19532_), .B(new_n12638_), .Y(new_n19533_));
  OAI21X1  g17097(.A0(new_n19531_), .A1(pi0619), .B0(new_n19533_), .Y(new_n19534_));
  AND2X1   g17098(.A(new_n19469_), .B(new_n12645_), .Y(new_n19535_));
  AND2X1   g17099(.A(new_n19535_), .B(new_n19534_), .Y(new_n19536_));
  NOR4X1   g17100(.A(new_n19484_), .B(new_n12764_), .C(new_n12762_), .D(pi0619), .Y(new_n19537_));
  NOR2X1   g17101(.A(new_n19537_), .B(new_n12638_), .Y(new_n19538_));
  OAI21X1  g17102(.A0(new_n19531_), .A1(new_n12637_), .B0(new_n19538_), .Y(new_n19539_));
  AND2X1   g17103(.A(new_n19471_), .B(pi0648), .Y(new_n19540_));
  AOI21X1  g17104(.A0(new_n19540_), .A1(new_n19539_), .B0(new_n11886_), .Y(new_n19541_));
  INVX1    g17105(.A(new_n19541_), .Y(new_n19542_));
  AOI21X1  g17106(.A0(new_n19531_), .A1(new_n11886_), .B0(new_n14264_), .Y(new_n19543_));
  OAI21X1  g17107(.A0(new_n19542_), .A1(new_n19536_), .B0(new_n19543_), .Y(new_n19544_));
  AOI21X1  g17108(.A0(new_n19544_), .A1(new_n19501_), .B0(new_n14273_), .Y(new_n19545_));
  INVX1    g17109(.A(new_n19475_), .Y(new_n19546_));
  AND2X1   g17110(.A(new_n19485_), .B(new_n12852_), .Y(new_n19547_));
  AOI22X1  g17111(.A0(new_n19547_), .A1(new_n14564_), .B0(new_n19546_), .B1(new_n12867_), .Y(new_n19548_));
  AOI22X1  g17112(.A0(new_n19547_), .A1(new_n14566_), .B0(new_n19546_), .B1(new_n12865_), .Y(new_n19549_));
  MX2X1    g17113(.A(new_n19549_), .B(new_n19548_), .S0(new_n12689_), .Y(new_n19550_));
  OAI21X1  g17114(.A0(new_n19550_), .A1(new_n11884_), .B0(new_n14562_), .Y(new_n19551_));
  OAI22X1  g17115(.A0(new_n19551_), .A1(new_n19545_), .B0(new_n19493_), .B1(new_n11883_), .Y(new_n19552_));
  INVX1    g17116(.A(new_n19552_), .Y(new_n19553_));
  OAI21X1  g17117(.A0(new_n19491_), .A1(new_n12706_), .B0(new_n19490_), .Y(new_n19554_));
  MX2X1    g17118(.A(new_n19554_), .B(new_n19488_), .S0(new_n11883_), .Y(new_n19555_));
  OAI21X1  g17119(.A0(new_n19555_), .A1(pi0644), .B0(pi0715), .Y(new_n19556_));
  AOI21X1  g17120(.A0(new_n19553_), .A1(pi0644), .B0(new_n19556_), .Y(new_n19557_));
  OR4X1    g17121(.A(new_n12734_), .B(new_n2739_), .C(new_n11883_), .D(pi0186), .Y(new_n19558_));
  OAI21X1  g17122(.A0(new_n19476_), .A1(new_n12735_), .B0(new_n19558_), .Y(new_n19559_));
  OAI21X1  g17123(.A0(new_n19454_), .A1(pi0644), .B0(new_n12739_), .Y(new_n19560_));
  AOI21X1  g17124(.A0(new_n19559_), .A1(pi0644), .B0(new_n19560_), .Y(new_n19561_));
  OR2X1    g17125(.A(new_n19561_), .B(new_n11882_), .Y(new_n19562_));
  OAI21X1  g17126(.A0(new_n19555_), .A1(new_n12743_), .B0(new_n12739_), .Y(new_n19563_));
  AOI21X1  g17127(.A0(new_n19553_), .A1(new_n12743_), .B0(new_n19563_), .Y(new_n19564_));
  OAI21X1  g17128(.A0(new_n19454_), .A1(new_n12743_), .B0(pi0715), .Y(new_n19565_));
  AOI21X1  g17129(.A0(new_n19559_), .A1(new_n12743_), .B0(new_n19565_), .Y(new_n19566_));
  OR2X1    g17130(.A(new_n19566_), .B(pi1160), .Y(new_n19567_));
  OAI22X1  g17131(.A0(new_n19567_), .A1(new_n19564_), .B0(new_n19562_), .B1(new_n19557_), .Y(new_n19568_));
  OAI21X1  g17132(.A0(new_n19552_), .A1(pi0790), .B0(pi0832), .Y(new_n19569_));
  AOI21X1  g17133(.A0(new_n19568_), .A1(pi0790), .B0(new_n19569_), .Y(new_n19570_));
  AOI21X1  g17134(.A0(new_n19452_), .A1(new_n19451_), .B0(new_n19570_), .Y(po0343));
  NOR2X1   g17135(.A(new_n3129_), .B(new_n8729_), .Y(new_n19572_));
  MX2X1    g17136(.A(new_n13704_), .B(new_n13699_), .S0(pi0770), .Y(new_n19573_));
  AOI21X1  g17137(.A0(new_n16745_), .A1(new_n8729_), .B0(pi0770), .Y(new_n19574_));
  NAND2X1  g17138(.A(new_n19574_), .B(new_n16746_), .Y(new_n19575_));
  OAI21X1  g17139(.A0(new_n19573_), .A1(pi0187), .B0(new_n19575_), .Y(new_n19576_));
  NOR2X1   g17140(.A(new_n13676_), .B(new_n14707_), .Y(new_n19577_));
  OAI21X1  g17141(.A0(new_n13674_), .A1(new_n8729_), .B0(new_n19577_), .Y(new_n19578_));
  AOI21X1  g17142(.A0(new_n13672_), .A1(new_n8729_), .B0(new_n19578_), .Y(new_n19579_));
  OAI21X1  g17143(.A0(new_n13694_), .A1(pi0187), .B0(new_n14707_), .Y(new_n19580_));
  AOI21X1  g17144(.A0(new_n13688_), .A1(pi0187), .B0(new_n19580_), .Y(new_n19581_));
  OR2X1    g17145(.A(new_n19581_), .B(new_n14637_), .Y(new_n19582_));
  OAI21X1  g17146(.A0(new_n19582_), .A1(new_n19579_), .B0(new_n3129_), .Y(new_n19583_));
  AOI21X1  g17147(.A0(new_n19576_), .A1(new_n14637_), .B0(new_n19583_), .Y(new_n19584_));
  NOR3X1   g17148(.A(new_n19584_), .B(new_n19572_), .C(pi0625), .Y(new_n19585_));
  INVX1    g17149(.A(new_n19572_), .Y(new_n19586_));
  OAI21X1  g17150(.A0(new_n19576_), .A1(new_n3810_), .B0(new_n19586_), .Y(new_n19587_));
  OAI21X1  g17151(.A0(new_n19587_), .A1(new_n12493_), .B0(new_n12494_), .Y(new_n19588_));
  OAI21X1  g17152(.A0(new_n16436_), .A1(new_n8729_), .B0(new_n2996_), .Y(new_n19589_));
  AOI21X1  g17153(.A0(new_n16435_), .A1(new_n8729_), .B0(new_n19589_), .Y(new_n19590_));
  AOI21X1  g17154(.A0(new_n12901_), .A1(new_n8729_), .B0(new_n12568_), .Y(new_n19591_));
  NOR3X1   g17155(.A(new_n19591_), .B(new_n19590_), .C(new_n14637_), .Y(new_n19592_));
  NOR2X1   g17156(.A(pi0726), .B(pi0187), .Y(new_n19593_));
  INVX1    g17157(.A(new_n19593_), .Y(new_n19594_));
  OAI21X1  g17158(.A0(new_n19594_), .A1(new_n13699_), .B0(new_n3129_), .Y(new_n19595_));
  OAI21X1  g17159(.A0(new_n19595_), .A1(new_n19592_), .B0(new_n19586_), .Y(new_n19596_));
  OR2X1    g17160(.A(new_n19596_), .B(new_n12493_), .Y(new_n19597_));
  AOI21X1  g17161(.A0(new_n13699_), .A1(new_n3129_), .B0(pi0187), .Y(new_n19598_));
  AOI21X1  g17162(.A0(new_n19598_), .A1(new_n12493_), .B0(new_n12494_), .Y(new_n19599_));
  AOI21X1  g17163(.A0(new_n19599_), .A1(new_n19597_), .B0(pi0608), .Y(new_n19600_));
  OAI21X1  g17164(.A0(new_n19588_), .A1(new_n19585_), .B0(new_n19600_), .Y(new_n19601_));
  NOR3X1   g17165(.A(new_n19584_), .B(new_n19572_), .C(new_n12493_), .Y(new_n19602_));
  OAI21X1  g17166(.A0(new_n19587_), .A1(pi0625), .B0(pi1153), .Y(new_n19603_));
  OR2X1    g17167(.A(new_n19596_), .B(pi0625), .Y(new_n19604_));
  AOI21X1  g17168(.A0(new_n19598_), .A1(pi0625), .B0(pi1153), .Y(new_n19605_));
  AOI21X1  g17169(.A0(new_n19605_), .A1(new_n19604_), .B0(new_n12584_), .Y(new_n19606_));
  OAI21X1  g17170(.A0(new_n19603_), .A1(new_n19602_), .B0(new_n19606_), .Y(new_n19607_));
  AOI21X1  g17171(.A0(new_n19607_), .A1(new_n19601_), .B0(new_n11889_), .Y(new_n19608_));
  NOR3X1   g17172(.A(new_n19584_), .B(new_n19572_), .C(pi0778), .Y(new_n19609_));
  NOR2X1   g17173(.A(new_n19609_), .B(new_n19608_), .Y(new_n19610_));
  NAND2X1  g17174(.A(new_n19596_), .B(new_n11889_), .Y(new_n19611_));
  AOI22X1  g17175(.A0(new_n19605_), .A1(new_n19604_), .B0(new_n19599_), .B1(new_n19597_), .Y(new_n19612_));
  OR2X1    g17176(.A(new_n19612_), .B(new_n11889_), .Y(new_n19613_));
  AND2X1   g17177(.A(new_n19613_), .B(new_n19611_), .Y(new_n19614_));
  AOI21X1  g17178(.A0(new_n19614_), .A1(pi0609), .B0(pi1155), .Y(new_n19615_));
  OAI21X1  g17179(.A0(new_n19610_), .A1(pi0609), .B0(new_n19615_), .Y(new_n19616_));
  NAND2X1  g17180(.A(new_n19587_), .B(new_n12623_), .Y(new_n19617_));
  OAI22X1  g17181(.A0(new_n19617_), .A1(new_n12590_), .B0(new_n19598_), .B1(new_n12599_), .Y(new_n19618_));
  AOI21X1  g17182(.A0(new_n19618_), .A1(pi1155), .B0(pi0660), .Y(new_n19619_));
  AOI21X1  g17183(.A0(new_n19614_), .A1(new_n12590_), .B0(new_n12591_), .Y(new_n19620_));
  OAI21X1  g17184(.A0(new_n19610_), .A1(new_n12590_), .B0(new_n19620_), .Y(new_n19621_));
  OAI22X1  g17185(.A0(new_n19617_), .A1(pi0609), .B0(new_n19598_), .B1(new_n12608_), .Y(new_n19622_));
  AOI21X1  g17186(.A0(new_n19622_), .A1(new_n12591_), .B0(new_n12596_), .Y(new_n19623_));
  AOI22X1  g17187(.A0(new_n19623_), .A1(new_n19621_), .B0(new_n19619_), .B1(new_n19616_), .Y(new_n19624_));
  OAI21X1  g17188(.A0(new_n19609_), .A1(new_n19608_), .B0(new_n11888_), .Y(new_n19625_));
  OAI21X1  g17189(.A0(new_n19624_), .A1(new_n11888_), .B0(new_n19625_), .Y(new_n19626_));
  OR2X1    g17190(.A(new_n19598_), .B(new_n13598_), .Y(new_n19627_));
  OAI21X1  g17191(.A0(new_n19614_), .A1(new_n12618_), .B0(new_n19627_), .Y(new_n19628_));
  OAI21X1  g17192(.A0(new_n19628_), .A1(new_n12614_), .B0(new_n12615_), .Y(new_n19629_));
  AOI21X1  g17193(.A0(new_n19626_), .A1(new_n12614_), .B0(new_n19629_), .Y(new_n19630_));
  INVX1    g17194(.A(new_n19598_), .Y(new_n19631_));
  MX2X1    g17195(.A(new_n19631_), .B(new_n19587_), .S0(new_n12623_), .Y(new_n19632_));
  AND2X1   g17196(.A(new_n19632_), .B(new_n11888_), .Y(new_n19633_));
  MX2X1    g17197(.A(new_n19622_), .B(new_n19618_), .S0(pi1155), .Y(new_n19634_));
  AOI21X1  g17198(.A0(new_n19634_), .A1(pi0785), .B0(new_n19633_), .Y(new_n19635_));
  OAI21X1  g17199(.A0(new_n19631_), .A1(pi0618), .B0(pi1154), .Y(new_n19636_));
  AOI21X1  g17200(.A0(new_n19635_), .A1(pi0618), .B0(new_n19636_), .Y(new_n19637_));
  OR2X1    g17201(.A(new_n19637_), .B(pi0627), .Y(new_n19638_));
  OAI21X1  g17202(.A0(new_n19628_), .A1(pi0618), .B0(pi1154), .Y(new_n19639_));
  AOI21X1  g17203(.A0(new_n19626_), .A1(pi0618), .B0(new_n19639_), .Y(new_n19640_));
  OAI21X1  g17204(.A0(new_n19631_), .A1(new_n12614_), .B0(new_n12615_), .Y(new_n19641_));
  AOI21X1  g17205(.A0(new_n19635_), .A1(new_n12614_), .B0(new_n19641_), .Y(new_n19642_));
  OR2X1    g17206(.A(new_n19642_), .B(new_n12622_), .Y(new_n19643_));
  OAI22X1  g17207(.A0(new_n19643_), .A1(new_n19640_), .B0(new_n19638_), .B1(new_n19630_), .Y(new_n19644_));
  MX2X1    g17208(.A(new_n19644_), .B(new_n19626_), .S0(new_n11887_), .Y(new_n19645_));
  MX2X1    g17209(.A(new_n19628_), .B(new_n19631_), .S0(new_n12641_), .Y(new_n19646_));
  OAI21X1  g17210(.A0(new_n19646_), .A1(new_n12637_), .B0(new_n12638_), .Y(new_n19647_));
  AOI21X1  g17211(.A0(new_n19645_), .A1(new_n12637_), .B0(new_n19647_), .Y(new_n19648_));
  OR2X1    g17212(.A(new_n19635_), .B(pi0781), .Y(new_n19649_));
  OAI21X1  g17213(.A0(new_n19642_), .A1(new_n19637_), .B0(pi0781), .Y(new_n19650_));
  NAND2X1  g17214(.A(new_n19650_), .B(new_n19649_), .Y(new_n19651_));
  AOI21X1  g17215(.A0(new_n19598_), .A1(new_n12637_), .B0(new_n12638_), .Y(new_n19652_));
  OAI21X1  g17216(.A0(new_n19651_), .A1(new_n12637_), .B0(new_n19652_), .Y(new_n19653_));
  NAND2X1  g17217(.A(new_n19653_), .B(new_n12645_), .Y(new_n19654_));
  OAI21X1  g17218(.A0(new_n19646_), .A1(pi0619), .B0(pi1159), .Y(new_n19655_));
  AOI21X1  g17219(.A0(new_n19645_), .A1(pi0619), .B0(new_n19655_), .Y(new_n19656_));
  AOI21X1  g17220(.A0(new_n19598_), .A1(pi0619), .B0(pi1159), .Y(new_n19657_));
  OAI21X1  g17221(.A0(new_n19651_), .A1(pi0619), .B0(new_n19657_), .Y(new_n19658_));
  NAND2X1  g17222(.A(new_n19658_), .B(pi0648), .Y(new_n19659_));
  OAI22X1  g17223(.A0(new_n19659_), .A1(new_n19656_), .B0(new_n19654_), .B1(new_n19648_), .Y(new_n19660_));
  MX2X1    g17224(.A(new_n19660_), .B(new_n19645_), .S0(new_n11886_), .Y(new_n19661_));
  MX2X1    g17225(.A(new_n19646_), .B(new_n19631_), .S0(new_n12659_), .Y(new_n19662_));
  AOI21X1  g17226(.A0(new_n19662_), .A1(pi0626), .B0(pi0641), .Y(new_n19663_));
  OAI21X1  g17227(.A0(new_n19661_), .A1(pi0626), .B0(new_n19663_), .Y(new_n19664_));
  NAND2X1  g17228(.A(new_n19658_), .B(new_n19653_), .Y(new_n19665_));
  MX2X1    g17229(.A(new_n19665_), .B(new_n19651_), .S0(new_n11886_), .Y(new_n19666_));
  OAI21X1  g17230(.A0(new_n19598_), .A1(new_n12664_), .B0(pi0641), .Y(new_n19667_));
  AOI21X1  g17231(.A0(new_n19666_), .A1(new_n12664_), .B0(new_n19667_), .Y(new_n19668_));
  NOR2X1   g17232(.A(new_n19668_), .B(pi1158), .Y(new_n19669_));
  AOI21X1  g17233(.A0(new_n19662_), .A1(new_n12664_), .B0(new_n12672_), .Y(new_n19670_));
  OAI21X1  g17234(.A0(new_n19661_), .A1(new_n12664_), .B0(new_n19670_), .Y(new_n19671_));
  OAI21X1  g17235(.A0(new_n19598_), .A1(pi0626), .B0(new_n12672_), .Y(new_n19672_));
  AOI21X1  g17236(.A0(new_n19666_), .A1(pi0626), .B0(new_n19672_), .Y(new_n19673_));
  NOR2X1   g17237(.A(new_n19673_), .B(new_n12676_), .Y(new_n19674_));
  AOI22X1  g17238(.A0(new_n19674_), .A1(new_n19671_), .B0(new_n19669_), .B1(new_n19664_), .Y(new_n19675_));
  MX2X1    g17239(.A(new_n19675_), .B(new_n19661_), .S0(new_n11885_), .Y(new_n19676_));
  MX2X1    g17240(.A(new_n19666_), .B(new_n19631_), .S0(new_n12841_), .Y(new_n19677_));
  OAI21X1  g17241(.A0(new_n19677_), .A1(new_n12683_), .B0(new_n12684_), .Y(new_n19678_));
  AOI21X1  g17242(.A0(new_n19676_), .A1(new_n12683_), .B0(new_n19678_), .Y(new_n19679_));
  MX2X1    g17243(.A(new_n19662_), .B(new_n19631_), .S0(new_n12691_), .Y(new_n19680_));
  AOI21X1  g17244(.A0(new_n19598_), .A1(new_n12683_), .B0(new_n12684_), .Y(new_n19681_));
  OAI21X1  g17245(.A0(new_n19680_), .A1(new_n12683_), .B0(new_n19681_), .Y(new_n19682_));
  NAND2X1  g17246(.A(new_n19682_), .B(new_n12689_), .Y(new_n19683_));
  OAI21X1  g17247(.A0(new_n19677_), .A1(pi0628), .B0(pi1156), .Y(new_n19684_));
  AOI21X1  g17248(.A0(new_n19676_), .A1(pi0628), .B0(new_n19684_), .Y(new_n19685_));
  AOI21X1  g17249(.A0(new_n19598_), .A1(pi0628), .B0(pi1156), .Y(new_n19686_));
  OAI21X1  g17250(.A0(new_n19680_), .A1(pi0628), .B0(new_n19686_), .Y(new_n19687_));
  NAND2X1  g17251(.A(new_n19687_), .B(pi0629), .Y(new_n19688_));
  OAI22X1  g17252(.A0(new_n19688_), .A1(new_n19685_), .B0(new_n19683_), .B1(new_n19679_), .Y(new_n19689_));
  AND2X1   g17253(.A(new_n19676_), .B(new_n11884_), .Y(new_n19690_));
  AOI21X1  g17254(.A0(new_n19689_), .A1(pi0792), .B0(new_n19690_), .Y(new_n19691_));
  MX2X1    g17255(.A(new_n19677_), .B(new_n19631_), .S0(new_n12711_), .Y(new_n19692_));
  INVX1    g17256(.A(new_n19692_), .Y(new_n19693_));
  AOI21X1  g17257(.A0(new_n19693_), .A1(pi0647), .B0(pi1157), .Y(new_n19694_));
  OAI21X1  g17258(.A0(new_n19691_), .A1(pi0647), .B0(new_n19694_), .Y(new_n19695_));
  INVX1    g17259(.A(new_n19680_), .Y(new_n19696_));
  AND2X1   g17260(.A(new_n19687_), .B(new_n19682_), .Y(new_n19697_));
  MX2X1    g17261(.A(new_n19697_), .B(new_n19696_), .S0(new_n11884_), .Y(new_n19698_));
  INVX1    g17262(.A(new_n19698_), .Y(new_n19699_));
  AOI21X1  g17263(.A0(new_n19598_), .A1(new_n12705_), .B0(new_n12706_), .Y(new_n19700_));
  OAI21X1  g17264(.A0(new_n19699_), .A1(new_n12705_), .B0(new_n19700_), .Y(new_n19701_));
  AND2X1   g17265(.A(new_n19701_), .B(new_n12723_), .Y(new_n19702_));
  AOI21X1  g17266(.A0(new_n19693_), .A1(new_n12705_), .B0(new_n12706_), .Y(new_n19703_));
  OAI21X1  g17267(.A0(new_n19691_), .A1(new_n12705_), .B0(new_n19703_), .Y(new_n19704_));
  AOI21X1  g17268(.A0(new_n19598_), .A1(pi0647), .B0(pi1157), .Y(new_n19705_));
  OAI21X1  g17269(.A0(new_n19699_), .A1(pi0647), .B0(new_n19705_), .Y(new_n19706_));
  AND2X1   g17270(.A(new_n19706_), .B(pi0630), .Y(new_n19707_));
  AOI22X1  g17271(.A0(new_n19707_), .A1(new_n19704_), .B0(new_n19702_), .B1(new_n19695_), .Y(new_n19708_));
  MX2X1    g17272(.A(new_n19708_), .B(new_n19691_), .S0(new_n11883_), .Y(new_n19709_));
  AND2X1   g17273(.A(new_n19706_), .B(new_n19701_), .Y(new_n19710_));
  MX2X1    g17274(.A(new_n19710_), .B(new_n19698_), .S0(new_n11883_), .Y(new_n19711_));
  AOI21X1  g17275(.A0(new_n19711_), .A1(new_n12743_), .B0(new_n12739_), .Y(new_n19712_));
  OAI21X1  g17276(.A0(new_n19709_), .A1(new_n12743_), .B0(new_n19712_), .Y(new_n19713_));
  MX2X1    g17277(.A(new_n19693_), .B(new_n19598_), .S0(new_n12735_), .Y(new_n19714_));
  OAI21X1  g17278(.A0(new_n19631_), .A1(pi0644), .B0(new_n12739_), .Y(new_n19715_));
  AOI21X1  g17279(.A0(new_n19714_), .A1(pi0644), .B0(new_n19715_), .Y(new_n19716_));
  NOR2X1   g17280(.A(new_n19716_), .B(new_n11882_), .Y(new_n19717_));
  AND2X1   g17281(.A(new_n19717_), .B(new_n19713_), .Y(new_n19718_));
  OR2X1    g17282(.A(new_n19691_), .B(pi0787), .Y(new_n19719_));
  OAI21X1  g17283(.A0(new_n19708_), .A1(new_n11883_), .B0(new_n19719_), .Y(new_n19720_));
  AND2X1   g17284(.A(new_n19711_), .B(pi0644), .Y(new_n19721_));
  OR2X1    g17285(.A(new_n19721_), .B(pi0715), .Y(new_n19722_));
  AOI21X1  g17286(.A0(new_n19720_), .A1(new_n12743_), .B0(new_n19722_), .Y(new_n19723_));
  OAI21X1  g17287(.A0(new_n19631_), .A1(new_n12743_), .B0(pi0715), .Y(new_n19724_));
  AOI21X1  g17288(.A0(new_n19714_), .A1(new_n12743_), .B0(new_n19724_), .Y(new_n19725_));
  OR2X1    g17289(.A(new_n19725_), .B(pi1160), .Y(new_n19726_));
  OAI21X1  g17290(.A0(new_n19726_), .A1(new_n19723_), .B0(pi0790), .Y(new_n19727_));
  AOI21X1  g17291(.A0(new_n19709_), .A1(new_n12897_), .B0(po1038), .Y(new_n19728_));
  OAI21X1  g17292(.A0(new_n19727_), .A1(new_n19718_), .B0(new_n19728_), .Y(new_n19729_));
  AOI21X1  g17293(.A0(po1038), .A1(new_n8729_), .B0(pi0832), .Y(new_n19730_));
  AOI21X1  g17294(.A0(pi1093), .A1(pi1092), .B0(pi0187), .Y(new_n19731_));
  INVX1    g17295(.A(new_n19731_), .Y(new_n19732_));
  AOI21X1  g17296(.A0(new_n12178_), .A1(new_n14707_), .B0(new_n19731_), .Y(new_n19733_));
  AOI21X1  g17297(.A0(new_n12601_), .A1(new_n2739_), .B0(new_n19733_), .Y(new_n19734_));
  INVX1    g17298(.A(new_n19733_), .Y(new_n19735_));
  AOI21X1  g17299(.A0(new_n19735_), .A1(new_n12776_), .B0(new_n12591_), .Y(new_n19736_));
  AOI21X1  g17300(.A0(new_n19734_), .A1(new_n12779_), .B0(pi1155), .Y(new_n19737_));
  OAI21X1  g17301(.A0(new_n19737_), .A1(new_n19736_), .B0(pi0785), .Y(new_n19738_));
  OAI21X1  g17302(.A0(new_n19734_), .A1(pi0785), .B0(new_n19738_), .Y(new_n19739_));
  INVX1    g17303(.A(new_n19739_), .Y(new_n19740_));
  AOI21X1  g17304(.A0(new_n19740_), .A1(new_n12785_), .B0(new_n12615_), .Y(new_n19741_));
  AOI21X1  g17305(.A0(new_n19740_), .A1(new_n12788_), .B0(pi1154), .Y(new_n19742_));
  OR2X1    g17306(.A(new_n19742_), .B(new_n19741_), .Y(new_n19743_));
  MX2X1    g17307(.A(new_n19743_), .B(new_n19739_), .S0(new_n11887_), .Y(new_n19744_));
  AND2X1   g17308(.A(new_n19744_), .B(new_n11886_), .Y(new_n19745_));
  AOI21X1  g17309(.A0(new_n19731_), .A1(new_n12637_), .B0(new_n12638_), .Y(new_n19746_));
  OAI21X1  g17310(.A0(new_n19744_), .A1(new_n12637_), .B0(new_n19746_), .Y(new_n19747_));
  AOI21X1  g17311(.A0(new_n19731_), .A1(pi0619), .B0(pi1159), .Y(new_n19748_));
  OAI21X1  g17312(.A0(new_n19744_), .A1(pi0619), .B0(new_n19748_), .Y(new_n19749_));
  AOI21X1  g17313(.A0(new_n19749_), .A1(new_n19747_), .B0(new_n11886_), .Y(new_n19750_));
  NOR2X1   g17314(.A(new_n19750_), .B(new_n19745_), .Y(new_n19751_));
  INVX1    g17315(.A(new_n19751_), .Y(new_n19752_));
  MX2X1    g17316(.A(new_n19752_), .B(new_n19732_), .S0(new_n12841_), .Y(new_n19753_));
  MX2X1    g17317(.A(new_n19753_), .B(new_n19732_), .S0(new_n12711_), .Y(new_n19754_));
  AOI21X1  g17318(.A0(new_n12566_), .A1(pi0726), .B0(new_n19731_), .Y(new_n19755_));
  AND2X1   g17319(.A(new_n12566_), .B(pi0726), .Y(new_n19756_));
  AND2X1   g17320(.A(new_n19756_), .B(new_n12493_), .Y(new_n19757_));
  MX2X1    g17321(.A(new_n19731_), .B(pi0625), .S0(new_n19756_), .Y(new_n19758_));
  NOR2X1   g17322(.A(new_n19731_), .B(pi1153), .Y(new_n19759_));
  INVX1    g17323(.A(new_n19759_), .Y(new_n19760_));
  OAI22X1  g17324(.A0(new_n19760_), .A1(new_n19757_), .B0(new_n19758_), .B1(new_n12494_), .Y(new_n19761_));
  MX2X1    g17325(.A(new_n19761_), .B(new_n19755_), .S0(new_n11889_), .Y(new_n19762_));
  NOR4X1   g17326(.A(new_n19762_), .B(new_n12765_), .C(new_n12764_), .D(new_n12762_), .Y(new_n19763_));
  INVX1    g17327(.A(new_n19763_), .Y(new_n19764_));
  NOR3X1   g17328(.A(new_n19764_), .B(new_n12870_), .C(new_n12851_), .Y(new_n19765_));
  INVX1    g17329(.A(new_n19765_), .Y(new_n19766_));
  AOI21X1  g17330(.A0(new_n19731_), .A1(pi0647), .B0(pi1157), .Y(new_n19767_));
  OAI21X1  g17331(.A0(new_n19766_), .A1(pi0647), .B0(new_n19767_), .Y(new_n19768_));
  MX2X1    g17332(.A(new_n19765_), .B(new_n19731_), .S0(new_n12705_), .Y(new_n19769_));
  OAI22X1  g17333(.A0(new_n19769_), .A1(new_n14387_), .B0(new_n19768_), .B1(new_n12723_), .Y(new_n19770_));
  AOI21X1  g17334(.A0(new_n19754_), .A1(new_n14385_), .B0(new_n19770_), .Y(new_n19771_));
  AOI21X1  g17335(.A0(new_n19732_), .A1(pi0626), .B0(new_n16352_), .Y(new_n19772_));
  OAI21X1  g17336(.A0(new_n19751_), .A1(pi0626), .B0(new_n19772_), .Y(new_n19773_));
  AOI21X1  g17337(.A0(new_n19732_), .A1(new_n12664_), .B0(new_n16356_), .Y(new_n19774_));
  OAI21X1  g17338(.A0(new_n19751_), .A1(new_n12664_), .B0(new_n19774_), .Y(new_n19775_));
  NAND2X1  g17339(.A(new_n19763_), .B(new_n12769_), .Y(new_n19776_));
  NAND3X1  g17340(.A(new_n19776_), .B(new_n19775_), .C(new_n19773_), .Y(new_n19777_));
  AND2X1   g17341(.A(new_n19777_), .B(pi0788), .Y(new_n19778_));
  INVX1    g17342(.A(new_n19778_), .Y(new_n19779_));
  NOR2X1   g17343(.A(new_n19755_), .B(new_n12120_), .Y(new_n19780_));
  NOR2X1   g17344(.A(new_n19780_), .B(new_n19735_), .Y(new_n19781_));
  INVX1    g17345(.A(new_n19781_), .Y(new_n19782_));
  MX2X1    g17346(.A(new_n19735_), .B(new_n12493_), .S0(new_n19780_), .Y(new_n19783_));
  NOR2X1   g17347(.A(new_n19783_), .B(new_n19760_), .Y(new_n19784_));
  OAI21X1  g17348(.A0(new_n19758_), .A1(new_n12494_), .B0(new_n12584_), .Y(new_n19785_));
  NOR3X1   g17349(.A(new_n19755_), .B(new_n12120_), .C(new_n12493_), .Y(new_n19786_));
  NOR3X1   g17350(.A(new_n19786_), .B(new_n19735_), .C(new_n12494_), .Y(new_n19787_));
  OAI21X1  g17351(.A0(new_n19760_), .A1(new_n19757_), .B0(pi0608), .Y(new_n19788_));
  OAI22X1  g17352(.A0(new_n19788_), .A1(new_n19787_), .B0(new_n19785_), .B1(new_n19784_), .Y(new_n19789_));
  MX2X1    g17353(.A(new_n19789_), .B(new_n19782_), .S0(new_n11889_), .Y(new_n19790_));
  OAI21X1  g17354(.A0(new_n19762_), .A1(new_n12590_), .B0(new_n12591_), .Y(new_n19791_));
  AOI21X1  g17355(.A0(new_n19790_), .A1(new_n12590_), .B0(new_n19791_), .Y(new_n19792_));
  NOR3X1   g17356(.A(new_n19792_), .B(new_n19736_), .C(pi0660), .Y(new_n19793_));
  OAI21X1  g17357(.A0(new_n19762_), .A1(pi0609), .B0(pi1155), .Y(new_n19794_));
  AOI21X1  g17358(.A0(new_n19790_), .A1(pi0609), .B0(new_n19794_), .Y(new_n19795_));
  NOR3X1   g17359(.A(new_n19795_), .B(new_n19737_), .C(new_n12596_), .Y(new_n19796_));
  OAI21X1  g17360(.A0(new_n19796_), .A1(new_n19793_), .B0(pi0785), .Y(new_n19797_));
  NAND2X1  g17361(.A(new_n19790_), .B(new_n11888_), .Y(new_n19798_));
  AND2X1   g17362(.A(new_n19798_), .B(new_n19797_), .Y(new_n19799_));
  NOR3X1   g17363(.A(new_n19762_), .B(new_n12762_), .C(new_n12614_), .Y(new_n19800_));
  NOR2X1   g17364(.A(new_n19800_), .B(pi1154), .Y(new_n19801_));
  OAI21X1  g17365(.A0(new_n19799_), .A1(pi0618), .B0(new_n19801_), .Y(new_n19802_));
  NOR2X1   g17366(.A(new_n19741_), .B(pi0627), .Y(new_n19803_));
  NOR3X1   g17367(.A(new_n19762_), .B(new_n12762_), .C(pi0618), .Y(new_n19804_));
  NOR2X1   g17368(.A(new_n19804_), .B(new_n12615_), .Y(new_n19805_));
  OAI21X1  g17369(.A0(new_n19799_), .A1(new_n12614_), .B0(new_n19805_), .Y(new_n19806_));
  NOR2X1   g17370(.A(new_n19742_), .B(new_n12622_), .Y(new_n19807_));
  AOI22X1  g17371(.A0(new_n19807_), .A1(new_n19806_), .B0(new_n19803_), .B1(new_n19802_), .Y(new_n19808_));
  MX2X1    g17372(.A(new_n19808_), .B(new_n19799_), .S0(new_n11887_), .Y(new_n19809_));
  OR4X1    g17373(.A(new_n19762_), .B(new_n12764_), .C(new_n12762_), .D(new_n12637_), .Y(new_n19810_));
  AND2X1   g17374(.A(new_n19810_), .B(new_n12638_), .Y(new_n19811_));
  OAI21X1  g17375(.A0(new_n19809_), .A1(pi0619), .B0(new_n19811_), .Y(new_n19812_));
  AND2X1   g17376(.A(new_n19747_), .B(new_n12645_), .Y(new_n19813_));
  AND2X1   g17377(.A(new_n19813_), .B(new_n19812_), .Y(new_n19814_));
  NOR4X1   g17378(.A(new_n19762_), .B(new_n12764_), .C(new_n12762_), .D(pi0619), .Y(new_n19815_));
  NOR2X1   g17379(.A(new_n19815_), .B(new_n12638_), .Y(new_n19816_));
  OAI21X1  g17380(.A0(new_n19809_), .A1(new_n12637_), .B0(new_n19816_), .Y(new_n19817_));
  AND2X1   g17381(.A(new_n19749_), .B(pi0648), .Y(new_n19818_));
  AOI21X1  g17382(.A0(new_n19818_), .A1(new_n19817_), .B0(new_n11886_), .Y(new_n19819_));
  INVX1    g17383(.A(new_n19819_), .Y(new_n19820_));
  AOI21X1  g17384(.A0(new_n19809_), .A1(new_n11886_), .B0(new_n14264_), .Y(new_n19821_));
  OAI21X1  g17385(.A0(new_n19820_), .A1(new_n19814_), .B0(new_n19821_), .Y(new_n19822_));
  AOI21X1  g17386(.A0(new_n19822_), .A1(new_n19779_), .B0(new_n14273_), .Y(new_n19823_));
  INVX1    g17387(.A(new_n19753_), .Y(new_n19824_));
  AND2X1   g17388(.A(new_n19763_), .B(new_n12852_), .Y(new_n19825_));
  AOI22X1  g17389(.A0(new_n19825_), .A1(new_n14564_), .B0(new_n19824_), .B1(new_n12867_), .Y(new_n19826_));
  AOI22X1  g17390(.A0(new_n19825_), .A1(new_n14566_), .B0(new_n19824_), .B1(new_n12865_), .Y(new_n19827_));
  MX2X1    g17391(.A(new_n19827_), .B(new_n19826_), .S0(new_n12689_), .Y(new_n19828_));
  OAI21X1  g17392(.A0(new_n19828_), .A1(new_n11884_), .B0(new_n14562_), .Y(new_n19829_));
  OAI22X1  g17393(.A0(new_n19829_), .A1(new_n19823_), .B0(new_n19771_), .B1(new_n11883_), .Y(new_n19830_));
  INVX1    g17394(.A(new_n19830_), .Y(new_n19831_));
  OAI21X1  g17395(.A0(new_n19769_), .A1(new_n12706_), .B0(new_n19768_), .Y(new_n19832_));
  MX2X1    g17396(.A(new_n19832_), .B(new_n19766_), .S0(new_n11883_), .Y(new_n19833_));
  OAI21X1  g17397(.A0(new_n19833_), .A1(pi0644), .B0(pi0715), .Y(new_n19834_));
  AOI21X1  g17398(.A0(new_n19831_), .A1(pi0644), .B0(new_n19834_), .Y(new_n19835_));
  OR4X1    g17399(.A(new_n12734_), .B(new_n2739_), .C(new_n11883_), .D(pi0187), .Y(new_n19836_));
  OAI21X1  g17400(.A0(new_n19754_), .A1(new_n12735_), .B0(new_n19836_), .Y(new_n19837_));
  OAI21X1  g17401(.A0(new_n19732_), .A1(pi0644), .B0(new_n12739_), .Y(new_n19838_));
  AOI21X1  g17402(.A0(new_n19837_), .A1(pi0644), .B0(new_n19838_), .Y(new_n19839_));
  OR2X1    g17403(.A(new_n19839_), .B(new_n11882_), .Y(new_n19840_));
  OAI21X1  g17404(.A0(new_n19833_), .A1(new_n12743_), .B0(new_n12739_), .Y(new_n19841_));
  AOI21X1  g17405(.A0(new_n19831_), .A1(new_n12743_), .B0(new_n19841_), .Y(new_n19842_));
  OAI21X1  g17406(.A0(new_n19732_), .A1(new_n12743_), .B0(pi0715), .Y(new_n19843_));
  AOI21X1  g17407(.A0(new_n19837_), .A1(new_n12743_), .B0(new_n19843_), .Y(new_n19844_));
  OR2X1    g17408(.A(new_n19844_), .B(pi1160), .Y(new_n19845_));
  OAI22X1  g17409(.A0(new_n19845_), .A1(new_n19842_), .B0(new_n19840_), .B1(new_n19835_), .Y(new_n19846_));
  OAI21X1  g17410(.A0(new_n19830_), .A1(pi0790), .B0(pi0832), .Y(new_n19847_));
  AOI21X1  g17411(.A0(new_n19846_), .A1(pi0790), .B0(new_n19847_), .Y(new_n19848_));
  AOI21X1  g17412(.A0(new_n19730_), .A1(new_n19729_), .B0(new_n19848_), .Y(po0344));
  NOR2X1   g17413(.A(new_n3129_), .B(new_n7389_), .Y(new_n19850_));
  MX2X1    g17414(.A(new_n13704_), .B(new_n13699_), .S0(pi0768), .Y(new_n19851_));
  AOI21X1  g17415(.A0(new_n16745_), .A1(new_n7389_), .B0(pi0768), .Y(new_n19852_));
  NAND2X1  g17416(.A(new_n19852_), .B(new_n16746_), .Y(new_n19853_));
  OAI21X1  g17417(.A0(new_n19851_), .A1(pi0188), .B0(new_n19853_), .Y(new_n19854_));
  NOR2X1   g17418(.A(new_n13676_), .B(new_n15474_), .Y(new_n19855_));
  OAI21X1  g17419(.A0(new_n13674_), .A1(new_n7389_), .B0(new_n19855_), .Y(new_n19856_));
  AOI21X1  g17420(.A0(new_n13672_), .A1(new_n7389_), .B0(new_n19856_), .Y(new_n19857_));
  OAI21X1  g17421(.A0(new_n13694_), .A1(pi0188), .B0(new_n15474_), .Y(new_n19858_));
  AOI21X1  g17422(.A0(new_n13688_), .A1(pi0188), .B0(new_n19858_), .Y(new_n19859_));
  OR2X1    g17423(.A(new_n19859_), .B(new_n15470_), .Y(new_n19860_));
  OAI21X1  g17424(.A0(new_n19860_), .A1(new_n19857_), .B0(new_n3129_), .Y(new_n19861_));
  AOI21X1  g17425(.A0(new_n19854_), .A1(new_n15470_), .B0(new_n19861_), .Y(new_n19862_));
  NOR3X1   g17426(.A(new_n19862_), .B(new_n19850_), .C(pi0625), .Y(new_n19863_));
  INVX1    g17427(.A(new_n19850_), .Y(new_n19864_));
  OAI21X1  g17428(.A0(new_n19854_), .A1(new_n3810_), .B0(new_n19864_), .Y(new_n19865_));
  OAI21X1  g17429(.A0(new_n19865_), .A1(new_n12493_), .B0(new_n12494_), .Y(new_n19866_));
  OAI21X1  g17430(.A0(new_n16436_), .A1(new_n7389_), .B0(new_n2996_), .Y(new_n19867_));
  AOI21X1  g17431(.A0(new_n16435_), .A1(new_n7389_), .B0(new_n19867_), .Y(new_n19868_));
  AOI21X1  g17432(.A0(new_n12901_), .A1(new_n7389_), .B0(new_n12568_), .Y(new_n19869_));
  NOR3X1   g17433(.A(new_n19869_), .B(new_n19868_), .C(new_n15470_), .Y(new_n19870_));
  NOR2X1   g17434(.A(pi0705), .B(pi0188), .Y(new_n19871_));
  INVX1    g17435(.A(new_n19871_), .Y(new_n19872_));
  OAI21X1  g17436(.A0(new_n19872_), .A1(new_n13699_), .B0(new_n3129_), .Y(new_n19873_));
  OAI21X1  g17437(.A0(new_n19873_), .A1(new_n19870_), .B0(new_n19864_), .Y(new_n19874_));
  OR2X1    g17438(.A(new_n19874_), .B(new_n12493_), .Y(new_n19875_));
  AOI21X1  g17439(.A0(new_n13699_), .A1(new_n3129_), .B0(pi0188), .Y(new_n19876_));
  AOI21X1  g17440(.A0(new_n19876_), .A1(new_n12493_), .B0(new_n12494_), .Y(new_n19877_));
  AOI21X1  g17441(.A0(new_n19877_), .A1(new_n19875_), .B0(pi0608), .Y(new_n19878_));
  OAI21X1  g17442(.A0(new_n19866_), .A1(new_n19863_), .B0(new_n19878_), .Y(new_n19879_));
  NOR3X1   g17443(.A(new_n19862_), .B(new_n19850_), .C(new_n12493_), .Y(new_n19880_));
  OAI21X1  g17444(.A0(new_n19865_), .A1(pi0625), .B0(pi1153), .Y(new_n19881_));
  OR2X1    g17445(.A(new_n19874_), .B(pi0625), .Y(new_n19882_));
  AOI21X1  g17446(.A0(new_n19876_), .A1(pi0625), .B0(pi1153), .Y(new_n19883_));
  AOI21X1  g17447(.A0(new_n19883_), .A1(new_n19882_), .B0(new_n12584_), .Y(new_n19884_));
  OAI21X1  g17448(.A0(new_n19881_), .A1(new_n19880_), .B0(new_n19884_), .Y(new_n19885_));
  AOI21X1  g17449(.A0(new_n19885_), .A1(new_n19879_), .B0(new_n11889_), .Y(new_n19886_));
  NOR3X1   g17450(.A(new_n19862_), .B(new_n19850_), .C(pi0778), .Y(new_n19887_));
  NOR2X1   g17451(.A(new_n19887_), .B(new_n19886_), .Y(new_n19888_));
  NAND2X1  g17452(.A(new_n19874_), .B(new_n11889_), .Y(new_n19889_));
  AOI22X1  g17453(.A0(new_n19883_), .A1(new_n19882_), .B0(new_n19877_), .B1(new_n19875_), .Y(new_n19890_));
  OR2X1    g17454(.A(new_n19890_), .B(new_n11889_), .Y(new_n19891_));
  AND2X1   g17455(.A(new_n19891_), .B(new_n19889_), .Y(new_n19892_));
  AOI21X1  g17456(.A0(new_n19892_), .A1(pi0609), .B0(pi1155), .Y(new_n19893_));
  OAI21X1  g17457(.A0(new_n19888_), .A1(pi0609), .B0(new_n19893_), .Y(new_n19894_));
  NAND2X1  g17458(.A(new_n19865_), .B(new_n12623_), .Y(new_n19895_));
  OAI22X1  g17459(.A0(new_n19895_), .A1(new_n12590_), .B0(new_n19876_), .B1(new_n12599_), .Y(new_n19896_));
  AOI21X1  g17460(.A0(new_n19896_), .A1(pi1155), .B0(pi0660), .Y(new_n19897_));
  AOI21X1  g17461(.A0(new_n19892_), .A1(new_n12590_), .B0(new_n12591_), .Y(new_n19898_));
  OAI21X1  g17462(.A0(new_n19888_), .A1(new_n12590_), .B0(new_n19898_), .Y(new_n19899_));
  OAI22X1  g17463(.A0(new_n19895_), .A1(pi0609), .B0(new_n19876_), .B1(new_n12608_), .Y(new_n19900_));
  AOI21X1  g17464(.A0(new_n19900_), .A1(new_n12591_), .B0(new_n12596_), .Y(new_n19901_));
  AOI22X1  g17465(.A0(new_n19901_), .A1(new_n19899_), .B0(new_n19897_), .B1(new_n19894_), .Y(new_n19902_));
  OAI21X1  g17466(.A0(new_n19887_), .A1(new_n19886_), .B0(new_n11888_), .Y(new_n19903_));
  OAI21X1  g17467(.A0(new_n19902_), .A1(new_n11888_), .B0(new_n19903_), .Y(new_n19904_));
  OR2X1    g17468(.A(new_n19876_), .B(new_n13598_), .Y(new_n19905_));
  OAI21X1  g17469(.A0(new_n19892_), .A1(new_n12618_), .B0(new_n19905_), .Y(new_n19906_));
  OAI21X1  g17470(.A0(new_n19906_), .A1(new_n12614_), .B0(new_n12615_), .Y(new_n19907_));
  AOI21X1  g17471(.A0(new_n19904_), .A1(new_n12614_), .B0(new_n19907_), .Y(new_n19908_));
  INVX1    g17472(.A(new_n19876_), .Y(new_n19909_));
  MX2X1    g17473(.A(new_n19909_), .B(new_n19865_), .S0(new_n12623_), .Y(new_n19910_));
  AND2X1   g17474(.A(new_n19910_), .B(new_n11888_), .Y(new_n19911_));
  MX2X1    g17475(.A(new_n19900_), .B(new_n19896_), .S0(pi1155), .Y(new_n19912_));
  AOI21X1  g17476(.A0(new_n19912_), .A1(pi0785), .B0(new_n19911_), .Y(new_n19913_));
  OAI21X1  g17477(.A0(new_n19909_), .A1(pi0618), .B0(pi1154), .Y(new_n19914_));
  AOI21X1  g17478(.A0(new_n19913_), .A1(pi0618), .B0(new_n19914_), .Y(new_n19915_));
  OR2X1    g17479(.A(new_n19915_), .B(pi0627), .Y(new_n19916_));
  OAI21X1  g17480(.A0(new_n19906_), .A1(pi0618), .B0(pi1154), .Y(new_n19917_));
  AOI21X1  g17481(.A0(new_n19904_), .A1(pi0618), .B0(new_n19917_), .Y(new_n19918_));
  OAI21X1  g17482(.A0(new_n19909_), .A1(new_n12614_), .B0(new_n12615_), .Y(new_n19919_));
  AOI21X1  g17483(.A0(new_n19913_), .A1(new_n12614_), .B0(new_n19919_), .Y(new_n19920_));
  OR2X1    g17484(.A(new_n19920_), .B(new_n12622_), .Y(new_n19921_));
  OAI22X1  g17485(.A0(new_n19921_), .A1(new_n19918_), .B0(new_n19916_), .B1(new_n19908_), .Y(new_n19922_));
  MX2X1    g17486(.A(new_n19922_), .B(new_n19904_), .S0(new_n11887_), .Y(new_n19923_));
  MX2X1    g17487(.A(new_n19906_), .B(new_n19909_), .S0(new_n12641_), .Y(new_n19924_));
  OAI21X1  g17488(.A0(new_n19924_), .A1(new_n12637_), .B0(new_n12638_), .Y(new_n19925_));
  AOI21X1  g17489(.A0(new_n19923_), .A1(new_n12637_), .B0(new_n19925_), .Y(new_n19926_));
  OR2X1    g17490(.A(new_n19913_), .B(pi0781), .Y(new_n19927_));
  OAI21X1  g17491(.A0(new_n19920_), .A1(new_n19915_), .B0(pi0781), .Y(new_n19928_));
  NAND2X1  g17492(.A(new_n19928_), .B(new_n19927_), .Y(new_n19929_));
  AOI21X1  g17493(.A0(new_n19876_), .A1(new_n12637_), .B0(new_n12638_), .Y(new_n19930_));
  OAI21X1  g17494(.A0(new_n19929_), .A1(new_n12637_), .B0(new_n19930_), .Y(new_n19931_));
  NAND2X1  g17495(.A(new_n19931_), .B(new_n12645_), .Y(new_n19932_));
  OAI21X1  g17496(.A0(new_n19924_), .A1(pi0619), .B0(pi1159), .Y(new_n19933_));
  AOI21X1  g17497(.A0(new_n19923_), .A1(pi0619), .B0(new_n19933_), .Y(new_n19934_));
  AOI21X1  g17498(.A0(new_n19876_), .A1(pi0619), .B0(pi1159), .Y(new_n19935_));
  OAI21X1  g17499(.A0(new_n19929_), .A1(pi0619), .B0(new_n19935_), .Y(new_n19936_));
  NAND2X1  g17500(.A(new_n19936_), .B(pi0648), .Y(new_n19937_));
  OAI22X1  g17501(.A0(new_n19937_), .A1(new_n19934_), .B0(new_n19932_), .B1(new_n19926_), .Y(new_n19938_));
  MX2X1    g17502(.A(new_n19938_), .B(new_n19923_), .S0(new_n11886_), .Y(new_n19939_));
  MX2X1    g17503(.A(new_n19924_), .B(new_n19909_), .S0(new_n12659_), .Y(new_n19940_));
  AOI21X1  g17504(.A0(new_n19940_), .A1(pi0626), .B0(pi0641), .Y(new_n19941_));
  OAI21X1  g17505(.A0(new_n19939_), .A1(pi0626), .B0(new_n19941_), .Y(new_n19942_));
  NAND2X1  g17506(.A(new_n19936_), .B(new_n19931_), .Y(new_n19943_));
  MX2X1    g17507(.A(new_n19943_), .B(new_n19929_), .S0(new_n11886_), .Y(new_n19944_));
  OAI21X1  g17508(.A0(new_n19876_), .A1(new_n12664_), .B0(pi0641), .Y(new_n19945_));
  AOI21X1  g17509(.A0(new_n19944_), .A1(new_n12664_), .B0(new_n19945_), .Y(new_n19946_));
  NOR2X1   g17510(.A(new_n19946_), .B(pi1158), .Y(new_n19947_));
  AOI21X1  g17511(.A0(new_n19940_), .A1(new_n12664_), .B0(new_n12672_), .Y(new_n19948_));
  OAI21X1  g17512(.A0(new_n19939_), .A1(new_n12664_), .B0(new_n19948_), .Y(new_n19949_));
  OAI21X1  g17513(.A0(new_n19876_), .A1(pi0626), .B0(new_n12672_), .Y(new_n19950_));
  AOI21X1  g17514(.A0(new_n19944_), .A1(pi0626), .B0(new_n19950_), .Y(new_n19951_));
  NOR2X1   g17515(.A(new_n19951_), .B(new_n12676_), .Y(new_n19952_));
  AOI22X1  g17516(.A0(new_n19952_), .A1(new_n19949_), .B0(new_n19947_), .B1(new_n19942_), .Y(new_n19953_));
  MX2X1    g17517(.A(new_n19953_), .B(new_n19939_), .S0(new_n11885_), .Y(new_n19954_));
  MX2X1    g17518(.A(new_n19944_), .B(new_n19909_), .S0(new_n12841_), .Y(new_n19955_));
  OAI21X1  g17519(.A0(new_n19955_), .A1(new_n12683_), .B0(new_n12684_), .Y(new_n19956_));
  AOI21X1  g17520(.A0(new_n19954_), .A1(new_n12683_), .B0(new_n19956_), .Y(new_n19957_));
  MX2X1    g17521(.A(new_n19940_), .B(new_n19909_), .S0(new_n12691_), .Y(new_n19958_));
  AOI21X1  g17522(.A0(new_n19876_), .A1(new_n12683_), .B0(new_n12684_), .Y(new_n19959_));
  OAI21X1  g17523(.A0(new_n19958_), .A1(new_n12683_), .B0(new_n19959_), .Y(new_n19960_));
  NAND2X1  g17524(.A(new_n19960_), .B(new_n12689_), .Y(new_n19961_));
  OAI21X1  g17525(.A0(new_n19955_), .A1(pi0628), .B0(pi1156), .Y(new_n19962_));
  AOI21X1  g17526(.A0(new_n19954_), .A1(pi0628), .B0(new_n19962_), .Y(new_n19963_));
  AOI21X1  g17527(.A0(new_n19876_), .A1(pi0628), .B0(pi1156), .Y(new_n19964_));
  OAI21X1  g17528(.A0(new_n19958_), .A1(pi0628), .B0(new_n19964_), .Y(new_n19965_));
  NAND2X1  g17529(.A(new_n19965_), .B(pi0629), .Y(new_n19966_));
  OAI22X1  g17530(.A0(new_n19966_), .A1(new_n19963_), .B0(new_n19961_), .B1(new_n19957_), .Y(new_n19967_));
  AND2X1   g17531(.A(new_n19954_), .B(new_n11884_), .Y(new_n19968_));
  AOI21X1  g17532(.A0(new_n19967_), .A1(pi0792), .B0(new_n19968_), .Y(new_n19969_));
  MX2X1    g17533(.A(new_n19955_), .B(new_n19909_), .S0(new_n12711_), .Y(new_n19970_));
  INVX1    g17534(.A(new_n19970_), .Y(new_n19971_));
  AOI21X1  g17535(.A0(new_n19971_), .A1(pi0647), .B0(pi1157), .Y(new_n19972_));
  OAI21X1  g17536(.A0(new_n19969_), .A1(pi0647), .B0(new_n19972_), .Y(new_n19973_));
  INVX1    g17537(.A(new_n19958_), .Y(new_n19974_));
  AND2X1   g17538(.A(new_n19965_), .B(new_n19960_), .Y(new_n19975_));
  MX2X1    g17539(.A(new_n19975_), .B(new_n19974_), .S0(new_n11884_), .Y(new_n19976_));
  INVX1    g17540(.A(new_n19976_), .Y(new_n19977_));
  AOI21X1  g17541(.A0(new_n19876_), .A1(new_n12705_), .B0(new_n12706_), .Y(new_n19978_));
  OAI21X1  g17542(.A0(new_n19977_), .A1(new_n12705_), .B0(new_n19978_), .Y(new_n19979_));
  AND2X1   g17543(.A(new_n19979_), .B(new_n12723_), .Y(new_n19980_));
  AOI21X1  g17544(.A0(new_n19971_), .A1(new_n12705_), .B0(new_n12706_), .Y(new_n19981_));
  OAI21X1  g17545(.A0(new_n19969_), .A1(new_n12705_), .B0(new_n19981_), .Y(new_n19982_));
  AOI21X1  g17546(.A0(new_n19876_), .A1(pi0647), .B0(pi1157), .Y(new_n19983_));
  OAI21X1  g17547(.A0(new_n19977_), .A1(pi0647), .B0(new_n19983_), .Y(new_n19984_));
  AND2X1   g17548(.A(new_n19984_), .B(pi0630), .Y(new_n19985_));
  AOI22X1  g17549(.A0(new_n19985_), .A1(new_n19982_), .B0(new_n19980_), .B1(new_n19973_), .Y(new_n19986_));
  MX2X1    g17550(.A(new_n19986_), .B(new_n19969_), .S0(new_n11883_), .Y(new_n19987_));
  AND2X1   g17551(.A(new_n19984_), .B(new_n19979_), .Y(new_n19988_));
  MX2X1    g17552(.A(new_n19988_), .B(new_n19976_), .S0(new_n11883_), .Y(new_n19989_));
  AOI21X1  g17553(.A0(new_n19989_), .A1(new_n12743_), .B0(new_n12739_), .Y(new_n19990_));
  OAI21X1  g17554(.A0(new_n19987_), .A1(new_n12743_), .B0(new_n19990_), .Y(new_n19991_));
  MX2X1    g17555(.A(new_n19971_), .B(new_n19876_), .S0(new_n12735_), .Y(new_n19992_));
  OAI21X1  g17556(.A0(new_n19909_), .A1(pi0644), .B0(new_n12739_), .Y(new_n19993_));
  AOI21X1  g17557(.A0(new_n19992_), .A1(pi0644), .B0(new_n19993_), .Y(new_n19994_));
  NOR2X1   g17558(.A(new_n19994_), .B(new_n11882_), .Y(new_n19995_));
  AND2X1   g17559(.A(new_n19995_), .B(new_n19991_), .Y(new_n19996_));
  OR2X1    g17560(.A(new_n19969_), .B(pi0787), .Y(new_n19997_));
  OAI21X1  g17561(.A0(new_n19986_), .A1(new_n11883_), .B0(new_n19997_), .Y(new_n19998_));
  AND2X1   g17562(.A(new_n19989_), .B(pi0644), .Y(new_n19999_));
  OR2X1    g17563(.A(new_n19999_), .B(pi0715), .Y(new_n20000_));
  AOI21X1  g17564(.A0(new_n19998_), .A1(new_n12743_), .B0(new_n20000_), .Y(new_n20001_));
  OAI21X1  g17565(.A0(new_n19909_), .A1(new_n12743_), .B0(pi0715), .Y(new_n20002_));
  AOI21X1  g17566(.A0(new_n19992_), .A1(new_n12743_), .B0(new_n20002_), .Y(new_n20003_));
  OR2X1    g17567(.A(new_n20003_), .B(pi1160), .Y(new_n20004_));
  OAI21X1  g17568(.A0(new_n20004_), .A1(new_n20001_), .B0(pi0790), .Y(new_n20005_));
  AOI21X1  g17569(.A0(new_n19987_), .A1(new_n12897_), .B0(po1038), .Y(new_n20006_));
  OAI21X1  g17570(.A0(new_n20005_), .A1(new_n19996_), .B0(new_n20006_), .Y(new_n20007_));
  AOI21X1  g17571(.A0(po1038), .A1(new_n7389_), .B0(pi0832), .Y(new_n20008_));
  AOI21X1  g17572(.A0(pi1093), .A1(pi1092), .B0(pi0188), .Y(new_n20009_));
  INVX1    g17573(.A(new_n20009_), .Y(new_n20010_));
  AOI21X1  g17574(.A0(new_n12178_), .A1(new_n15474_), .B0(new_n20009_), .Y(new_n20011_));
  AOI21X1  g17575(.A0(new_n12601_), .A1(new_n2739_), .B0(new_n20011_), .Y(new_n20012_));
  INVX1    g17576(.A(new_n20011_), .Y(new_n20013_));
  AOI21X1  g17577(.A0(new_n20013_), .A1(new_n12776_), .B0(new_n12591_), .Y(new_n20014_));
  AOI21X1  g17578(.A0(new_n20012_), .A1(new_n12779_), .B0(pi1155), .Y(new_n20015_));
  OAI21X1  g17579(.A0(new_n20015_), .A1(new_n20014_), .B0(pi0785), .Y(new_n20016_));
  OAI21X1  g17580(.A0(new_n20012_), .A1(pi0785), .B0(new_n20016_), .Y(new_n20017_));
  INVX1    g17581(.A(new_n20017_), .Y(new_n20018_));
  AOI21X1  g17582(.A0(new_n20018_), .A1(new_n12785_), .B0(new_n12615_), .Y(new_n20019_));
  AOI21X1  g17583(.A0(new_n20018_), .A1(new_n12788_), .B0(pi1154), .Y(new_n20020_));
  OR2X1    g17584(.A(new_n20020_), .B(new_n20019_), .Y(new_n20021_));
  MX2X1    g17585(.A(new_n20021_), .B(new_n20017_), .S0(new_n11887_), .Y(new_n20022_));
  AND2X1   g17586(.A(new_n20022_), .B(new_n11886_), .Y(new_n20023_));
  AOI21X1  g17587(.A0(new_n20009_), .A1(new_n12637_), .B0(new_n12638_), .Y(new_n20024_));
  OAI21X1  g17588(.A0(new_n20022_), .A1(new_n12637_), .B0(new_n20024_), .Y(new_n20025_));
  AOI21X1  g17589(.A0(new_n20009_), .A1(pi0619), .B0(pi1159), .Y(new_n20026_));
  OAI21X1  g17590(.A0(new_n20022_), .A1(pi0619), .B0(new_n20026_), .Y(new_n20027_));
  AOI21X1  g17591(.A0(new_n20027_), .A1(new_n20025_), .B0(new_n11886_), .Y(new_n20028_));
  NOR2X1   g17592(.A(new_n20028_), .B(new_n20023_), .Y(new_n20029_));
  INVX1    g17593(.A(new_n20029_), .Y(new_n20030_));
  MX2X1    g17594(.A(new_n20030_), .B(new_n20010_), .S0(new_n12841_), .Y(new_n20031_));
  MX2X1    g17595(.A(new_n20031_), .B(new_n20010_), .S0(new_n12711_), .Y(new_n20032_));
  AOI21X1  g17596(.A0(new_n12566_), .A1(pi0705), .B0(new_n20009_), .Y(new_n20033_));
  AND2X1   g17597(.A(new_n12566_), .B(pi0705), .Y(new_n20034_));
  AND2X1   g17598(.A(new_n20034_), .B(new_n12493_), .Y(new_n20035_));
  MX2X1    g17599(.A(new_n20009_), .B(pi0625), .S0(new_n20034_), .Y(new_n20036_));
  NOR2X1   g17600(.A(new_n20009_), .B(pi1153), .Y(new_n20037_));
  INVX1    g17601(.A(new_n20037_), .Y(new_n20038_));
  OAI22X1  g17602(.A0(new_n20038_), .A1(new_n20035_), .B0(new_n20036_), .B1(new_n12494_), .Y(new_n20039_));
  MX2X1    g17603(.A(new_n20039_), .B(new_n20033_), .S0(new_n11889_), .Y(new_n20040_));
  NOR4X1   g17604(.A(new_n20040_), .B(new_n12765_), .C(new_n12764_), .D(new_n12762_), .Y(new_n20041_));
  INVX1    g17605(.A(new_n20041_), .Y(new_n20042_));
  NOR3X1   g17606(.A(new_n20042_), .B(new_n12870_), .C(new_n12851_), .Y(new_n20043_));
  INVX1    g17607(.A(new_n20043_), .Y(new_n20044_));
  AOI21X1  g17608(.A0(new_n20009_), .A1(pi0647), .B0(pi1157), .Y(new_n20045_));
  OAI21X1  g17609(.A0(new_n20044_), .A1(pi0647), .B0(new_n20045_), .Y(new_n20046_));
  MX2X1    g17610(.A(new_n20043_), .B(new_n20009_), .S0(new_n12705_), .Y(new_n20047_));
  OAI22X1  g17611(.A0(new_n20047_), .A1(new_n14387_), .B0(new_n20046_), .B1(new_n12723_), .Y(new_n20048_));
  AOI21X1  g17612(.A0(new_n20032_), .A1(new_n14385_), .B0(new_n20048_), .Y(new_n20049_));
  AOI21X1  g17613(.A0(new_n20010_), .A1(pi0626), .B0(new_n16352_), .Y(new_n20050_));
  OAI21X1  g17614(.A0(new_n20029_), .A1(pi0626), .B0(new_n20050_), .Y(new_n20051_));
  AOI21X1  g17615(.A0(new_n20010_), .A1(new_n12664_), .B0(new_n16356_), .Y(new_n20052_));
  OAI21X1  g17616(.A0(new_n20029_), .A1(new_n12664_), .B0(new_n20052_), .Y(new_n20053_));
  NAND2X1  g17617(.A(new_n20041_), .B(new_n12769_), .Y(new_n20054_));
  NAND3X1  g17618(.A(new_n20054_), .B(new_n20053_), .C(new_n20051_), .Y(new_n20055_));
  AND2X1   g17619(.A(new_n20055_), .B(pi0788), .Y(new_n20056_));
  INVX1    g17620(.A(new_n20056_), .Y(new_n20057_));
  NOR2X1   g17621(.A(new_n20033_), .B(new_n12120_), .Y(new_n20058_));
  NOR2X1   g17622(.A(new_n20058_), .B(new_n20013_), .Y(new_n20059_));
  INVX1    g17623(.A(new_n20059_), .Y(new_n20060_));
  MX2X1    g17624(.A(new_n20013_), .B(new_n12493_), .S0(new_n20058_), .Y(new_n20061_));
  NOR2X1   g17625(.A(new_n20061_), .B(new_n20038_), .Y(new_n20062_));
  OAI21X1  g17626(.A0(new_n20036_), .A1(new_n12494_), .B0(new_n12584_), .Y(new_n20063_));
  NOR3X1   g17627(.A(new_n20033_), .B(new_n12120_), .C(new_n12493_), .Y(new_n20064_));
  NOR3X1   g17628(.A(new_n20064_), .B(new_n20013_), .C(new_n12494_), .Y(new_n20065_));
  OAI21X1  g17629(.A0(new_n20038_), .A1(new_n20035_), .B0(pi0608), .Y(new_n20066_));
  OAI22X1  g17630(.A0(new_n20066_), .A1(new_n20065_), .B0(new_n20063_), .B1(new_n20062_), .Y(new_n20067_));
  MX2X1    g17631(.A(new_n20067_), .B(new_n20060_), .S0(new_n11889_), .Y(new_n20068_));
  OAI21X1  g17632(.A0(new_n20040_), .A1(new_n12590_), .B0(new_n12591_), .Y(new_n20069_));
  AOI21X1  g17633(.A0(new_n20068_), .A1(new_n12590_), .B0(new_n20069_), .Y(new_n20070_));
  NOR3X1   g17634(.A(new_n20070_), .B(new_n20014_), .C(pi0660), .Y(new_n20071_));
  OAI21X1  g17635(.A0(new_n20040_), .A1(pi0609), .B0(pi1155), .Y(new_n20072_));
  AOI21X1  g17636(.A0(new_n20068_), .A1(pi0609), .B0(new_n20072_), .Y(new_n20073_));
  NOR3X1   g17637(.A(new_n20073_), .B(new_n20015_), .C(new_n12596_), .Y(new_n20074_));
  OAI21X1  g17638(.A0(new_n20074_), .A1(new_n20071_), .B0(pi0785), .Y(new_n20075_));
  NAND2X1  g17639(.A(new_n20068_), .B(new_n11888_), .Y(new_n20076_));
  AND2X1   g17640(.A(new_n20076_), .B(new_n20075_), .Y(new_n20077_));
  NOR3X1   g17641(.A(new_n20040_), .B(new_n12762_), .C(new_n12614_), .Y(new_n20078_));
  NOR2X1   g17642(.A(new_n20078_), .B(pi1154), .Y(new_n20079_));
  OAI21X1  g17643(.A0(new_n20077_), .A1(pi0618), .B0(new_n20079_), .Y(new_n20080_));
  NOR2X1   g17644(.A(new_n20019_), .B(pi0627), .Y(new_n20081_));
  NOR3X1   g17645(.A(new_n20040_), .B(new_n12762_), .C(pi0618), .Y(new_n20082_));
  NOR2X1   g17646(.A(new_n20082_), .B(new_n12615_), .Y(new_n20083_));
  OAI21X1  g17647(.A0(new_n20077_), .A1(new_n12614_), .B0(new_n20083_), .Y(new_n20084_));
  NOR2X1   g17648(.A(new_n20020_), .B(new_n12622_), .Y(new_n20085_));
  AOI22X1  g17649(.A0(new_n20085_), .A1(new_n20084_), .B0(new_n20081_), .B1(new_n20080_), .Y(new_n20086_));
  MX2X1    g17650(.A(new_n20086_), .B(new_n20077_), .S0(new_n11887_), .Y(new_n20087_));
  OR4X1    g17651(.A(new_n20040_), .B(new_n12764_), .C(new_n12762_), .D(new_n12637_), .Y(new_n20088_));
  AND2X1   g17652(.A(new_n20088_), .B(new_n12638_), .Y(new_n20089_));
  OAI21X1  g17653(.A0(new_n20087_), .A1(pi0619), .B0(new_n20089_), .Y(new_n20090_));
  AND2X1   g17654(.A(new_n20025_), .B(new_n12645_), .Y(new_n20091_));
  AND2X1   g17655(.A(new_n20091_), .B(new_n20090_), .Y(new_n20092_));
  NOR4X1   g17656(.A(new_n20040_), .B(new_n12764_), .C(new_n12762_), .D(pi0619), .Y(new_n20093_));
  NOR2X1   g17657(.A(new_n20093_), .B(new_n12638_), .Y(new_n20094_));
  OAI21X1  g17658(.A0(new_n20087_), .A1(new_n12637_), .B0(new_n20094_), .Y(new_n20095_));
  AND2X1   g17659(.A(new_n20027_), .B(pi0648), .Y(new_n20096_));
  AOI21X1  g17660(.A0(new_n20096_), .A1(new_n20095_), .B0(new_n11886_), .Y(new_n20097_));
  INVX1    g17661(.A(new_n20097_), .Y(new_n20098_));
  AOI21X1  g17662(.A0(new_n20087_), .A1(new_n11886_), .B0(new_n14264_), .Y(new_n20099_));
  OAI21X1  g17663(.A0(new_n20098_), .A1(new_n20092_), .B0(new_n20099_), .Y(new_n20100_));
  AOI21X1  g17664(.A0(new_n20100_), .A1(new_n20057_), .B0(new_n14273_), .Y(new_n20101_));
  INVX1    g17665(.A(new_n20031_), .Y(new_n20102_));
  AND2X1   g17666(.A(new_n20041_), .B(new_n12852_), .Y(new_n20103_));
  AOI22X1  g17667(.A0(new_n20103_), .A1(new_n14564_), .B0(new_n20102_), .B1(new_n12867_), .Y(new_n20104_));
  AOI22X1  g17668(.A0(new_n20103_), .A1(new_n14566_), .B0(new_n20102_), .B1(new_n12865_), .Y(new_n20105_));
  MX2X1    g17669(.A(new_n20105_), .B(new_n20104_), .S0(new_n12689_), .Y(new_n20106_));
  OAI21X1  g17670(.A0(new_n20106_), .A1(new_n11884_), .B0(new_n14562_), .Y(new_n20107_));
  OAI22X1  g17671(.A0(new_n20107_), .A1(new_n20101_), .B0(new_n20049_), .B1(new_n11883_), .Y(new_n20108_));
  INVX1    g17672(.A(new_n20108_), .Y(new_n20109_));
  OAI21X1  g17673(.A0(new_n20047_), .A1(new_n12706_), .B0(new_n20046_), .Y(new_n20110_));
  MX2X1    g17674(.A(new_n20110_), .B(new_n20044_), .S0(new_n11883_), .Y(new_n20111_));
  OAI21X1  g17675(.A0(new_n20111_), .A1(pi0644), .B0(pi0715), .Y(new_n20112_));
  AOI21X1  g17676(.A0(new_n20109_), .A1(pi0644), .B0(new_n20112_), .Y(new_n20113_));
  OR4X1    g17677(.A(new_n12734_), .B(new_n2739_), .C(new_n11883_), .D(pi0188), .Y(new_n20114_));
  OAI21X1  g17678(.A0(new_n20032_), .A1(new_n12735_), .B0(new_n20114_), .Y(new_n20115_));
  OAI21X1  g17679(.A0(new_n20010_), .A1(pi0644), .B0(new_n12739_), .Y(new_n20116_));
  AOI21X1  g17680(.A0(new_n20115_), .A1(pi0644), .B0(new_n20116_), .Y(new_n20117_));
  OR2X1    g17681(.A(new_n20117_), .B(new_n11882_), .Y(new_n20118_));
  OAI21X1  g17682(.A0(new_n20111_), .A1(new_n12743_), .B0(new_n12739_), .Y(new_n20119_));
  AOI21X1  g17683(.A0(new_n20109_), .A1(new_n12743_), .B0(new_n20119_), .Y(new_n20120_));
  OAI21X1  g17684(.A0(new_n20010_), .A1(new_n12743_), .B0(pi0715), .Y(new_n20121_));
  AOI21X1  g17685(.A0(new_n20115_), .A1(new_n12743_), .B0(new_n20121_), .Y(new_n20122_));
  OR2X1    g17686(.A(new_n20122_), .B(pi1160), .Y(new_n20123_));
  OAI22X1  g17687(.A0(new_n20123_), .A1(new_n20120_), .B0(new_n20118_), .B1(new_n20113_), .Y(new_n20124_));
  OAI21X1  g17688(.A0(new_n20108_), .A1(pi0790), .B0(pi0832), .Y(new_n20125_));
  AOI21X1  g17689(.A0(new_n20124_), .A1(pi0790), .B0(new_n20125_), .Y(new_n20126_));
  AOI21X1  g17690(.A0(new_n20008_), .A1(new_n20007_), .B0(new_n20126_), .Y(po0345));
  AND2X1   g17691(.A(new_n12161_), .B(pi0772), .Y(new_n20128_));
  OAI21X1  g17692(.A0(new_n20128_), .A1(new_n15421_), .B0(pi0039), .Y(new_n20129_));
  AOI21X1  g17693(.A0(new_n11947_), .A1(new_n15465_), .B0(pi0039), .Y(new_n20130_));
  OAI21X1  g17694(.A0(new_n12909_), .A1(new_n15465_), .B0(new_n20130_), .Y(new_n20131_));
  AOI21X1  g17695(.A0(new_n20131_), .A1(new_n20129_), .B0(new_n7942_), .Y(new_n20132_));
  NOR3X1   g17696(.A(new_n13977_), .B(new_n15465_), .C(pi0189), .Y(new_n20133_));
  OAI21X1  g17697(.A0(new_n20133_), .A1(new_n20132_), .B0(new_n2996_), .Y(new_n20134_));
  NOR2X1   g17698(.A(new_n12202_), .B(pi0189), .Y(new_n20135_));
  AOI21X1  g17699(.A0(new_n12120_), .A1(pi0772), .B0(new_n12901_), .Y(new_n20136_));
  NOR3X1   g17700(.A(new_n20136_), .B(new_n20135_), .C(new_n2996_), .Y(new_n20137_));
  INVX1    g17701(.A(new_n20137_), .Y(new_n20138_));
  NAND3X1  g17702(.A(new_n20138_), .B(new_n20134_), .C(new_n15428_), .Y(new_n20139_));
  OAI21X1  g17703(.A0(new_n13989_), .A1(pi0189), .B0(new_n15465_), .Y(new_n20140_));
  AOI21X1  g17704(.A0(new_n13986_), .A1(pi0189), .B0(new_n20140_), .Y(new_n20141_));
  AOI21X1  g17705(.A0(new_n12440_), .A1(pi0189), .B0(new_n15465_), .Y(new_n20142_));
  OAI21X1  g17706(.A0(new_n12401_), .A1(pi0189), .B0(new_n20142_), .Y(new_n20143_));
  NAND2X1  g17707(.A(new_n20143_), .B(pi0039), .Y(new_n20144_));
  AOI21X1  g17708(.A0(new_n13996_), .A1(pi0189), .B0(pi0772), .Y(new_n20145_));
  OAI21X1  g17709(.A0(new_n13995_), .A1(pi0189), .B0(new_n20145_), .Y(new_n20146_));
  NAND3X1  g17710(.A(new_n12453_), .B(new_n12104_), .C(pi0189), .Y(new_n20147_));
  AOI21X1  g17711(.A0(new_n12474_), .A1(new_n7942_), .B0(new_n15465_), .Y(new_n20148_));
  AOI21X1  g17712(.A0(new_n20148_), .A1(new_n20147_), .B0(pi0039), .Y(new_n20149_));
  AOI21X1  g17713(.A0(new_n20149_), .A1(new_n20146_), .B0(pi0038), .Y(new_n20150_));
  OAI21X1  g17714(.A0(new_n20144_), .A1(new_n20141_), .B0(new_n20150_), .Y(new_n20151_));
  NOR3X1   g17715(.A(new_n20137_), .B(new_n13676_), .C(new_n15428_), .Y(new_n20152_));
  AOI21X1  g17716(.A0(new_n20152_), .A1(new_n20151_), .B0(new_n3810_), .Y(new_n20153_));
  AOI22X1  g17717(.A0(new_n20153_), .A1(new_n20139_), .B0(new_n3810_), .B1(pi0189), .Y(new_n20154_));
  AND2X1   g17718(.A(new_n20154_), .B(new_n12493_), .Y(new_n20155_));
  NAND2X1  g17719(.A(new_n20138_), .B(new_n20134_), .Y(new_n20156_));
  MX2X1    g17720(.A(new_n20156_), .B(pi0189), .S0(new_n3810_), .Y(new_n20157_));
  OAI21X1  g17721(.A0(new_n20157_), .A1(new_n12493_), .B0(new_n12494_), .Y(new_n20158_));
  OAI21X1  g17722(.A0(new_n12574_), .A1(new_n3810_), .B0(pi0189), .Y(new_n20159_));
  NOR4X1   g17723(.A(new_n3125_), .B(new_n15428_), .C(pi0100), .D(pi0087), .Y(new_n20160_));
  INVX1    g17724(.A(new_n20160_), .Y(new_n20161_));
  OAI21X1  g17725(.A0(new_n12955_), .A1(pi0189), .B0(new_n2996_), .Y(new_n20162_));
  AOI21X1  g17726(.A0(new_n12953_), .A1(pi0189), .B0(new_n20162_), .Y(new_n20163_));
  OAI21X1  g17727(.A0(new_n20135_), .A1(new_n14017_), .B0(new_n20160_), .Y(new_n20164_));
  NOR2X1   g17728(.A(new_n20164_), .B(new_n20163_), .Y(new_n20165_));
  AOI21X1  g17729(.A0(new_n20161_), .A1(new_n20159_), .B0(new_n20165_), .Y(new_n20166_));
  AOI21X1  g17730(.A0(new_n20159_), .A1(new_n12493_), .B0(new_n12494_), .Y(new_n20167_));
  OAI21X1  g17731(.A0(new_n20166_), .A1(new_n12493_), .B0(new_n20167_), .Y(new_n20168_));
  AND2X1   g17732(.A(new_n20168_), .B(new_n12584_), .Y(new_n20169_));
  OAI21X1  g17733(.A0(new_n20158_), .A1(new_n20155_), .B0(new_n20169_), .Y(new_n20170_));
  AND2X1   g17734(.A(new_n20154_), .B(pi0625), .Y(new_n20171_));
  OAI21X1  g17735(.A0(new_n20157_), .A1(pi0625), .B0(pi1153), .Y(new_n20172_));
  AOI21X1  g17736(.A0(new_n20159_), .A1(pi0625), .B0(pi1153), .Y(new_n20173_));
  OAI21X1  g17737(.A0(new_n20166_), .A1(pi0625), .B0(new_n20173_), .Y(new_n20174_));
  AND2X1   g17738(.A(new_n20174_), .B(pi0608), .Y(new_n20175_));
  OAI21X1  g17739(.A0(new_n20172_), .A1(new_n20171_), .B0(new_n20175_), .Y(new_n20176_));
  AOI21X1  g17740(.A0(new_n20176_), .A1(new_n20170_), .B0(new_n11889_), .Y(new_n20177_));
  AND2X1   g17741(.A(new_n20154_), .B(new_n11889_), .Y(new_n20178_));
  OAI21X1  g17742(.A0(new_n20178_), .A1(new_n20177_), .B0(new_n12590_), .Y(new_n20179_));
  AND2X1   g17743(.A(new_n20166_), .B(new_n11889_), .Y(new_n20180_));
  NAND2X1  g17744(.A(new_n20174_), .B(new_n20168_), .Y(new_n20181_));
  AOI21X1  g17745(.A0(new_n20181_), .A1(pi0778), .B0(new_n20180_), .Y(new_n20182_));
  AOI21X1  g17746(.A0(new_n20182_), .A1(pi0609), .B0(pi1155), .Y(new_n20183_));
  NAND2X1  g17747(.A(new_n20159_), .B(new_n12601_), .Y(new_n20184_));
  OAI21X1  g17748(.A0(new_n20157_), .A1(new_n12601_), .B0(new_n20184_), .Y(new_n20185_));
  INVX1    g17749(.A(new_n20159_), .Y(new_n20186_));
  OAI21X1  g17750(.A0(new_n20186_), .A1(pi0609), .B0(pi1155), .Y(new_n20187_));
  AOI21X1  g17751(.A0(new_n20185_), .A1(pi0609), .B0(new_n20187_), .Y(new_n20188_));
  OR2X1    g17752(.A(new_n20188_), .B(pi0660), .Y(new_n20189_));
  AOI21X1  g17753(.A0(new_n20183_), .A1(new_n20179_), .B0(new_n20189_), .Y(new_n20190_));
  OAI21X1  g17754(.A0(new_n20178_), .A1(new_n20177_), .B0(pi0609), .Y(new_n20191_));
  AOI21X1  g17755(.A0(new_n20182_), .A1(new_n12590_), .B0(new_n12591_), .Y(new_n20192_));
  OAI21X1  g17756(.A0(new_n20186_), .A1(new_n12590_), .B0(new_n12591_), .Y(new_n20193_));
  AOI21X1  g17757(.A0(new_n20185_), .A1(new_n12590_), .B0(new_n20193_), .Y(new_n20194_));
  OR2X1    g17758(.A(new_n20194_), .B(new_n12596_), .Y(new_n20195_));
  AOI21X1  g17759(.A0(new_n20192_), .A1(new_n20191_), .B0(new_n20195_), .Y(new_n20196_));
  OAI21X1  g17760(.A0(new_n20196_), .A1(new_n20190_), .B0(pi0785), .Y(new_n20197_));
  OAI21X1  g17761(.A0(new_n20178_), .A1(new_n20177_), .B0(new_n11888_), .Y(new_n20198_));
  AOI21X1  g17762(.A0(new_n20198_), .A1(new_n20197_), .B0(pi0618), .Y(new_n20199_));
  AND2X1   g17763(.A(new_n20159_), .B(new_n12618_), .Y(new_n20200_));
  AOI21X1  g17764(.A0(new_n20182_), .A1(new_n13598_), .B0(new_n20200_), .Y(new_n20201_));
  OAI21X1  g17765(.A0(new_n20201_), .A1(new_n12614_), .B0(new_n12615_), .Y(new_n20202_));
  OAI21X1  g17766(.A0(new_n20194_), .A1(new_n20188_), .B0(pi0785), .Y(new_n20203_));
  OAI21X1  g17767(.A0(new_n20185_), .A1(pi0785), .B0(new_n20203_), .Y(new_n20204_));
  AOI21X1  g17768(.A0(new_n20159_), .A1(new_n12614_), .B0(new_n12615_), .Y(new_n20205_));
  OAI21X1  g17769(.A0(new_n20204_), .A1(new_n12614_), .B0(new_n20205_), .Y(new_n20206_));
  AND2X1   g17770(.A(new_n20206_), .B(new_n12622_), .Y(new_n20207_));
  OAI21X1  g17771(.A0(new_n20202_), .A1(new_n20199_), .B0(new_n20207_), .Y(new_n20208_));
  AOI21X1  g17772(.A0(new_n20198_), .A1(new_n20197_), .B0(new_n12614_), .Y(new_n20209_));
  OAI21X1  g17773(.A0(new_n20201_), .A1(pi0618), .B0(pi1154), .Y(new_n20210_));
  AOI21X1  g17774(.A0(new_n20159_), .A1(pi0618), .B0(pi1154), .Y(new_n20211_));
  OAI21X1  g17775(.A0(new_n20204_), .A1(pi0618), .B0(new_n20211_), .Y(new_n20212_));
  AND2X1   g17776(.A(new_n20212_), .B(pi0627), .Y(new_n20213_));
  OAI21X1  g17777(.A0(new_n20210_), .A1(new_n20209_), .B0(new_n20213_), .Y(new_n20214_));
  AOI21X1  g17778(.A0(new_n20214_), .A1(new_n20208_), .B0(new_n11887_), .Y(new_n20215_));
  AOI21X1  g17779(.A0(new_n20198_), .A1(new_n20197_), .B0(pi0781), .Y(new_n20216_));
  OAI21X1  g17780(.A0(new_n20216_), .A1(new_n20215_), .B0(new_n12637_), .Y(new_n20217_));
  MX2X1    g17781(.A(new_n20201_), .B(new_n20186_), .S0(new_n12641_), .Y(new_n20218_));
  INVX1    g17782(.A(new_n20218_), .Y(new_n20219_));
  AOI21X1  g17783(.A0(new_n20219_), .A1(pi0619), .B0(pi1159), .Y(new_n20220_));
  AOI21X1  g17784(.A0(new_n20212_), .A1(new_n20206_), .B0(new_n11887_), .Y(new_n20221_));
  AOI21X1  g17785(.A0(new_n20204_), .A1(new_n11887_), .B0(new_n20221_), .Y(new_n20222_));
  OAI21X1  g17786(.A0(new_n20186_), .A1(pi0619), .B0(pi1159), .Y(new_n20223_));
  AOI21X1  g17787(.A0(new_n20222_), .A1(pi0619), .B0(new_n20223_), .Y(new_n20224_));
  OR2X1    g17788(.A(new_n20224_), .B(pi0648), .Y(new_n20225_));
  AOI21X1  g17789(.A0(new_n20220_), .A1(new_n20217_), .B0(new_n20225_), .Y(new_n20226_));
  OAI21X1  g17790(.A0(new_n20216_), .A1(new_n20215_), .B0(pi0619), .Y(new_n20227_));
  AOI21X1  g17791(.A0(new_n20219_), .A1(new_n12637_), .B0(new_n12638_), .Y(new_n20228_));
  OAI21X1  g17792(.A0(new_n20186_), .A1(new_n12637_), .B0(new_n12638_), .Y(new_n20229_));
  AOI21X1  g17793(.A0(new_n20222_), .A1(new_n12637_), .B0(new_n20229_), .Y(new_n20230_));
  OR2X1    g17794(.A(new_n20230_), .B(new_n12645_), .Y(new_n20231_));
  AOI21X1  g17795(.A0(new_n20228_), .A1(new_n20227_), .B0(new_n20231_), .Y(new_n20232_));
  OAI21X1  g17796(.A0(new_n20232_), .A1(new_n20226_), .B0(pi0789), .Y(new_n20233_));
  OAI21X1  g17797(.A0(new_n20216_), .A1(new_n20215_), .B0(new_n11886_), .Y(new_n20234_));
  NAND3X1  g17798(.A(new_n20234_), .B(new_n20233_), .C(new_n11885_), .Y(new_n20235_));
  NAND3X1  g17799(.A(new_n20234_), .B(new_n20233_), .C(new_n12664_), .Y(new_n20236_));
  MX2X1    g17800(.A(new_n20218_), .B(new_n20186_), .S0(new_n12659_), .Y(new_n20237_));
  AOI21X1  g17801(.A0(new_n20237_), .A1(pi0626), .B0(pi0641), .Y(new_n20238_));
  NOR2X1   g17802(.A(new_n20230_), .B(new_n20224_), .Y(new_n20239_));
  MX2X1    g17803(.A(new_n20239_), .B(new_n20222_), .S0(new_n11886_), .Y(new_n20240_));
  AOI21X1  g17804(.A0(new_n20186_), .A1(pi0626), .B0(new_n12672_), .Y(new_n20241_));
  OAI21X1  g17805(.A0(new_n20240_), .A1(pi0626), .B0(new_n20241_), .Y(new_n20242_));
  NAND2X1  g17806(.A(new_n20242_), .B(new_n12676_), .Y(new_n20243_));
  AOI21X1  g17807(.A0(new_n20238_), .A1(new_n20236_), .B0(new_n20243_), .Y(new_n20244_));
  NAND3X1  g17808(.A(new_n20234_), .B(new_n20233_), .C(pi0626), .Y(new_n20245_));
  AOI21X1  g17809(.A0(new_n20237_), .A1(new_n12664_), .B0(new_n12672_), .Y(new_n20246_));
  AOI21X1  g17810(.A0(new_n20186_), .A1(new_n12664_), .B0(pi0641), .Y(new_n20247_));
  OAI21X1  g17811(.A0(new_n20240_), .A1(new_n12664_), .B0(new_n20247_), .Y(new_n20248_));
  NAND2X1  g17812(.A(new_n20248_), .B(pi1158), .Y(new_n20249_));
  AOI21X1  g17813(.A0(new_n20246_), .A1(new_n20245_), .B0(new_n20249_), .Y(new_n20250_));
  OAI21X1  g17814(.A0(new_n20250_), .A1(new_n20244_), .B0(pi0788), .Y(new_n20251_));
  NAND3X1  g17815(.A(new_n20251_), .B(new_n20235_), .C(new_n12683_), .Y(new_n20252_));
  MX2X1    g17816(.A(new_n20240_), .B(new_n20159_), .S0(new_n12841_), .Y(new_n20253_));
  AOI21X1  g17817(.A0(new_n20253_), .A1(pi0628), .B0(pi1156), .Y(new_n20254_));
  MX2X1    g17818(.A(new_n20237_), .B(new_n20186_), .S0(new_n12691_), .Y(new_n20255_));
  AOI21X1  g17819(.A0(new_n20159_), .A1(new_n12683_), .B0(new_n12684_), .Y(new_n20256_));
  OAI21X1  g17820(.A0(new_n20255_), .A1(new_n12683_), .B0(new_n20256_), .Y(new_n20257_));
  NAND2X1  g17821(.A(new_n20257_), .B(new_n12689_), .Y(new_n20258_));
  AOI21X1  g17822(.A0(new_n20254_), .A1(new_n20252_), .B0(new_n20258_), .Y(new_n20259_));
  NAND3X1  g17823(.A(new_n20251_), .B(new_n20235_), .C(pi0628), .Y(new_n20260_));
  AOI21X1  g17824(.A0(new_n20253_), .A1(new_n12683_), .B0(new_n12684_), .Y(new_n20261_));
  AOI21X1  g17825(.A0(new_n20159_), .A1(pi0628), .B0(pi1156), .Y(new_n20262_));
  OAI21X1  g17826(.A0(new_n20255_), .A1(pi0628), .B0(new_n20262_), .Y(new_n20263_));
  NAND2X1  g17827(.A(new_n20263_), .B(pi0629), .Y(new_n20264_));
  AOI21X1  g17828(.A0(new_n20261_), .A1(new_n20260_), .B0(new_n20264_), .Y(new_n20265_));
  OAI21X1  g17829(.A0(new_n20265_), .A1(new_n20259_), .B0(pi0792), .Y(new_n20266_));
  NAND3X1  g17830(.A(new_n20251_), .B(new_n20235_), .C(new_n11884_), .Y(new_n20267_));
  AOI21X1  g17831(.A0(new_n20267_), .A1(new_n20266_), .B0(pi0647), .Y(new_n20268_));
  MX2X1    g17832(.A(new_n20253_), .B(new_n20159_), .S0(new_n12711_), .Y(new_n20269_));
  INVX1    g17833(.A(new_n20269_), .Y(new_n20270_));
  OAI21X1  g17834(.A0(new_n20270_), .A1(new_n12705_), .B0(new_n12706_), .Y(new_n20271_));
  AND2X1   g17835(.A(new_n20255_), .B(new_n11884_), .Y(new_n20272_));
  AOI21X1  g17836(.A0(new_n20263_), .A1(new_n20257_), .B0(new_n11884_), .Y(new_n20273_));
  NOR2X1   g17837(.A(new_n20273_), .B(new_n20272_), .Y(new_n20274_));
  INVX1    g17838(.A(new_n20274_), .Y(new_n20275_));
  AOI21X1  g17839(.A0(new_n20159_), .A1(new_n12705_), .B0(new_n12706_), .Y(new_n20276_));
  OAI21X1  g17840(.A0(new_n20275_), .A1(new_n12705_), .B0(new_n20276_), .Y(new_n20277_));
  AND2X1   g17841(.A(new_n20277_), .B(new_n12723_), .Y(new_n20278_));
  OAI21X1  g17842(.A0(new_n20271_), .A1(new_n20268_), .B0(new_n20278_), .Y(new_n20279_));
  AOI21X1  g17843(.A0(new_n20267_), .A1(new_n20266_), .B0(new_n12705_), .Y(new_n20280_));
  OAI21X1  g17844(.A0(new_n20270_), .A1(pi0647), .B0(pi1157), .Y(new_n20281_));
  AOI21X1  g17845(.A0(new_n20159_), .A1(pi0647), .B0(pi1157), .Y(new_n20282_));
  OAI21X1  g17846(.A0(new_n20275_), .A1(pi0647), .B0(new_n20282_), .Y(new_n20283_));
  AND2X1   g17847(.A(new_n20283_), .B(pi0630), .Y(new_n20284_));
  OAI21X1  g17848(.A0(new_n20281_), .A1(new_n20280_), .B0(new_n20284_), .Y(new_n20285_));
  AOI21X1  g17849(.A0(new_n20285_), .A1(new_n20279_), .B0(new_n11883_), .Y(new_n20286_));
  AOI21X1  g17850(.A0(new_n20267_), .A1(new_n20266_), .B0(pi0787), .Y(new_n20287_));
  OAI21X1  g17851(.A0(new_n20287_), .A1(new_n20286_), .B0(pi0644), .Y(new_n20288_));
  AND2X1   g17852(.A(new_n20283_), .B(new_n20277_), .Y(new_n20289_));
  MX2X1    g17853(.A(new_n20289_), .B(new_n20274_), .S0(new_n11883_), .Y(new_n20290_));
  AOI21X1  g17854(.A0(new_n20290_), .A1(new_n12743_), .B0(new_n12739_), .Y(new_n20291_));
  MX2X1    g17855(.A(new_n20269_), .B(new_n20159_), .S0(new_n12735_), .Y(new_n20292_));
  OAI21X1  g17856(.A0(new_n20186_), .A1(pi0644), .B0(new_n12739_), .Y(new_n20293_));
  AOI21X1  g17857(.A0(new_n20292_), .A1(pi0644), .B0(new_n20293_), .Y(new_n20294_));
  OR2X1    g17858(.A(new_n20294_), .B(new_n11882_), .Y(new_n20295_));
  AOI21X1  g17859(.A0(new_n20291_), .A1(new_n20288_), .B0(new_n20295_), .Y(new_n20296_));
  OAI21X1  g17860(.A0(new_n20287_), .A1(new_n20286_), .B0(new_n12743_), .Y(new_n20297_));
  AOI21X1  g17861(.A0(new_n20290_), .A1(pi0644), .B0(pi0715), .Y(new_n20298_));
  OAI21X1  g17862(.A0(new_n20186_), .A1(new_n12743_), .B0(pi0715), .Y(new_n20299_));
  AOI21X1  g17863(.A0(new_n20292_), .A1(new_n12743_), .B0(new_n20299_), .Y(new_n20300_));
  OR2X1    g17864(.A(new_n20300_), .B(pi1160), .Y(new_n20301_));
  AOI21X1  g17865(.A0(new_n20298_), .A1(new_n20297_), .B0(new_n20301_), .Y(new_n20302_));
  NOR3X1   g17866(.A(new_n20302_), .B(new_n20296_), .C(new_n12897_), .Y(new_n20303_));
  NOR3X1   g17867(.A(new_n20287_), .B(new_n20286_), .C(pi0790), .Y(new_n20304_));
  OR2X1    g17868(.A(new_n20304_), .B(new_n5118_), .Y(new_n20305_));
  AOI21X1  g17869(.A0(new_n5118_), .A1(new_n7942_), .B0(pi0057), .Y(new_n20306_));
  OAI21X1  g17870(.A0(new_n20305_), .A1(new_n20303_), .B0(new_n20306_), .Y(new_n20307_));
  AOI21X1  g17871(.A0(pi0189), .A1(pi0057), .B0(pi0832), .Y(new_n20308_));
  NOR2X1   g17872(.A(new_n2739_), .B(new_n7942_), .Y(new_n20309_));
  AOI21X1  g17873(.A0(new_n12178_), .A1(pi0772), .B0(new_n20309_), .Y(new_n20310_));
  OAI21X1  g17874(.A0(new_n14209_), .A1(new_n15428_), .B0(new_n20310_), .Y(new_n20311_));
  NOR4X1   g17875(.A(new_n13585_), .B(new_n12120_), .C(new_n15428_), .D(new_n12493_), .Y(new_n20312_));
  INVX1    g17876(.A(new_n20312_), .Y(new_n20313_));
  AOI21X1  g17877(.A0(new_n20313_), .A1(new_n20311_), .B0(pi1153), .Y(new_n20314_));
  NOR3X1   g17878(.A(new_n13585_), .B(new_n15428_), .C(new_n12493_), .Y(new_n20315_));
  NOR3X1   g17879(.A(new_n20315_), .B(new_n20309_), .C(new_n12494_), .Y(new_n20316_));
  OR2X1    g17880(.A(new_n20316_), .B(pi0608), .Y(new_n20317_));
  AOI21X1  g17881(.A0(new_n12566_), .A1(pi0727), .B0(new_n20309_), .Y(new_n20318_));
  OR2X1    g17882(.A(new_n20318_), .B(new_n20315_), .Y(new_n20319_));
  AND2X1   g17883(.A(new_n20319_), .B(new_n12494_), .Y(new_n20320_));
  NAND2X1  g17884(.A(new_n20310_), .B(pi1153), .Y(new_n20321_));
  OAI21X1  g17885(.A0(new_n20321_), .A1(new_n20312_), .B0(pi0608), .Y(new_n20322_));
  OAI22X1  g17886(.A0(new_n20322_), .A1(new_n20320_), .B0(new_n20317_), .B1(new_n20314_), .Y(new_n20323_));
  MX2X1    g17887(.A(new_n20323_), .B(new_n20311_), .S0(new_n11889_), .Y(new_n20324_));
  INVX1    g17888(.A(new_n20318_), .Y(new_n20325_));
  AOI21X1  g17889(.A0(new_n20319_), .A1(new_n12494_), .B0(new_n20316_), .Y(new_n20326_));
  MX2X1    g17890(.A(new_n20326_), .B(new_n20325_), .S0(new_n11889_), .Y(new_n20327_));
  INVX1    g17891(.A(new_n20327_), .Y(new_n20328_));
  OAI21X1  g17892(.A0(new_n20328_), .A1(new_n12590_), .B0(new_n12591_), .Y(new_n20329_));
  AOI21X1  g17893(.A0(new_n20324_), .A1(new_n12590_), .B0(new_n20329_), .Y(new_n20330_));
  NOR3X1   g17894(.A(new_n13430_), .B(new_n12204_), .C(new_n15465_), .Y(new_n20331_));
  OAI21X1  g17895(.A0(new_n2739_), .A1(new_n7942_), .B0(pi1155), .Y(new_n20332_));
  OAI21X1  g17896(.A0(new_n20332_), .A1(new_n20331_), .B0(new_n12596_), .Y(new_n20333_));
  OAI21X1  g17897(.A0(new_n20328_), .A1(pi0609), .B0(pi1155), .Y(new_n20334_));
  AOI21X1  g17898(.A0(new_n20324_), .A1(pi0609), .B0(new_n20334_), .Y(new_n20335_));
  NOR3X1   g17899(.A(new_n13436_), .B(new_n12204_), .C(new_n15465_), .Y(new_n20336_));
  OAI21X1  g17900(.A0(new_n2739_), .A1(new_n7942_), .B0(new_n12591_), .Y(new_n20337_));
  OAI21X1  g17901(.A0(new_n20337_), .A1(new_n20336_), .B0(pi0660), .Y(new_n20338_));
  OAI22X1  g17902(.A0(new_n20338_), .A1(new_n20335_), .B0(new_n20333_), .B1(new_n20330_), .Y(new_n20339_));
  MX2X1    g17903(.A(new_n20339_), .B(new_n20324_), .S0(new_n11888_), .Y(new_n20340_));
  NAND2X1  g17904(.A(new_n20340_), .B(pi0618), .Y(new_n20341_));
  OAI22X1  g17905(.A0(new_n20328_), .A1(new_n12618_), .B0(new_n2739_), .B1(new_n7942_), .Y(new_n20342_));
  AOI21X1  g17906(.A0(new_n20342_), .A1(new_n12614_), .B0(new_n12615_), .Y(new_n20343_));
  OR4X1    g17907(.A(new_n14178_), .B(new_n12171_), .C(new_n2740_), .D(new_n15465_), .Y(new_n20344_));
  NOR3X1   g17908(.A(new_n20344_), .B(new_n12601_), .C(pi0618), .Y(new_n20345_));
  OAI21X1  g17909(.A0(new_n2739_), .A1(new_n7942_), .B0(new_n12615_), .Y(new_n20346_));
  OAI21X1  g17910(.A0(new_n20346_), .A1(new_n20345_), .B0(pi0627), .Y(new_n20347_));
  AOI21X1  g17911(.A0(new_n20343_), .A1(new_n20341_), .B0(new_n20347_), .Y(new_n20348_));
  NAND2X1  g17912(.A(new_n20340_), .B(new_n12614_), .Y(new_n20349_));
  AOI21X1  g17913(.A0(new_n20342_), .A1(pi0618), .B0(pi1154), .Y(new_n20350_));
  NOR3X1   g17914(.A(new_n20344_), .B(new_n12601_), .C(new_n12614_), .Y(new_n20351_));
  OAI21X1  g17915(.A0(new_n2739_), .A1(new_n7942_), .B0(pi1154), .Y(new_n20352_));
  OAI21X1  g17916(.A0(new_n20352_), .A1(new_n20351_), .B0(new_n12622_), .Y(new_n20353_));
  AOI21X1  g17917(.A0(new_n20350_), .A1(new_n20349_), .B0(new_n20353_), .Y(new_n20354_));
  OAI21X1  g17918(.A0(new_n20354_), .A1(new_n20348_), .B0(pi0781), .Y(new_n20355_));
  AOI21X1  g17919(.A0(new_n20340_), .A1(new_n11887_), .B0(new_n16248_), .Y(new_n20356_));
  NAND3X1  g17920(.A(new_n20327_), .B(new_n14198_), .C(new_n13598_), .Y(new_n20357_));
  NOR4X1   g17921(.A(new_n20344_), .B(new_n14183_), .C(new_n12601_), .D(pi0619), .Y(new_n20358_));
  NOR4X1   g17922(.A(new_n20344_), .B(new_n14183_), .C(new_n12601_), .D(new_n12637_), .Y(new_n20359_));
  OAI22X1  g17923(.A0(new_n20359_), .A1(new_n16251_), .B0(new_n20358_), .B1(new_n16252_), .Y(new_n20360_));
  AOI21X1  g17924(.A0(new_n20357_), .A1(new_n16246_), .B0(new_n20360_), .Y(new_n20361_));
  OAI21X1  g17925(.A0(new_n2739_), .A1(new_n7942_), .B0(pi0789), .Y(new_n20362_));
  OAI21X1  g17926(.A0(new_n20362_), .A1(new_n20361_), .B0(new_n12842_), .Y(new_n20363_));
  AOI21X1  g17927(.A0(new_n20356_), .A1(new_n20355_), .B0(new_n20363_), .Y(new_n20364_));
  OAI22X1  g17928(.A0(new_n20357_), .A1(new_n12659_), .B0(new_n2739_), .B1(new_n7942_), .Y(new_n20365_));
  NOR2X1   g17929(.A(new_n20344_), .B(new_n14185_), .Y(new_n20366_));
  AOI21X1  g17930(.A0(new_n20366_), .A1(new_n12664_), .B0(new_n20309_), .Y(new_n20367_));
  OAI21X1  g17931(.A0(new_n20367_), .A1(pi1158), .B0(pi0641), .Y(new_n20368_));
  AOI21X1  g17932(.A0(new_n20365_), .A1(new_n14196_), .B0(new_n20368_), .Y(new_n20369_));
  AOI21X1  g17933(.A0(new_n20366_), .A1(pi0626), .B0(new_n20309_), .Y(new_n20370_));
  OAI21X1  g17934(.A0(new_n20370_), .A1(new_n12676_), .B0(new_n12672_), .Y(new_n20371_));
  AOI21X1  g17935(.A0(new_n20365_), .A1(new_n14204_), .B0(new_n20371_), .Y(new_n20372_));
  NOR3X1   g17936(.A(new_n20372_), .B(new_n20369_), .C(new_n11885_), .Y(new_n20373_));
  OR2X1    g17937(.A(new_n20373_), .B(new_n14273_), .Y(new_n20374_));
  NOR4X1   g17938(.A(new_n20344_), .B(new_n14185_), .C(new_n12841_), .D(pi0629), .Y(new_n20375_));
  NOR2X1   g17939(.A(new_n20328_), .B(new_n13624_), .Y(new_n20376_));
  OAI22X1  g17940(.A0(new_n20376_), .A1(new_n12689_), .B0(new_n20375_), .B1(new_n12683_), .Y(new_n20377_));
  AOI21X1  g17941(.A0(new_n20366_), .A1(new_n14175_), .B0(pi0628), .Y(new_n20378_));
  OAI21X1  g17942(.A0(new_n20378_), .A1(new_n12689_), .B0(pi1156), .Y(new_n20379_));
  AOI21X1  g17943(.A0(new_n20376_), .A1(pi0628), .B0(new_n20379_), .Y(new_n20380_));
  AOI21X1  g17944(.A0(new_n20377_), .A1(new_n12684_), .B0(new_n20380_), .Y(new_n20381_));
  OAI21X1  g17945(.A0(new_n2739_), .A1(new_n7942_), .B0(pi0792), .Y(new_n20382_));
  OAI22X1  g17946(.A0(new_n20382_), .A1(new_n20381_), .B0(new_n20374_), .B1(new_n20364_), .Y(new_n20383_));
  OR4X1    g17947(.A(new_n20344_), .B(new_n14185_), .C(new_n12841_), .D(new_n12711_), .Y(new_n20384_));
  OR2X1    g17948(.A(new_n20384_), .B(pi0630), .Y(new_n20385_));
  NOR3X1   g17949(.A(new_n20328_), .B(new_n13639_), .C(new_n13624_), .Y(new_n20386_));
  INVX1    g17950(.A(new_n20386_), .Y(new_n20387_));
  AOI22X1  g17951(.A0(new_n20387_), .A1(pi0630), .B0(new_n20385_), .B1(pi0647), .Y(new_n20388_));
  AOI21X1  g17952(.A0(new_n20387_), .A1(new_n12723_), .B0(new_n12705_), .Y(new_n20389_));
  OAI21X1  g17953(.A0(new_n20384_), .A1(new_n12723_), .B0(pi1157), .Y(new_n20390_));
  OAI22X1  g17954(.A0(new_n20390_), .A1(new_n20389_), .B0(new_n20388_), .B1(pi1157), .Y(new_n20391_));
  NOR2X1   g17955(.A(new_n20309_), .B(new_n11883_), .Y(new_n20392_));
  AOI22X1  g17956(.A0(new_n20392_), .A1(new_n20391_), .B0(new_n20383_), .B1(new_n14562_), .Y(new_n20393_));
  AOI21X1  g17957(.A0(new_n20386_), .A1(new_n14286_), .B0(new_n20309_), .Y(new_n20394_));
  OAI21X1  g17958(.A0(new_n20394_), .A1(pi0644), .B0(pi0715), .Y(new_n20395_));
  AOI21X1  g17959(.A0(new_n20393_), .A1(pi0644), .B0(new_n20395_), .Y(new_n20396_));
  NOR4X1   g17960(.A(new_n20344_), .B(new_n16294_), .C(new_n14185_), .D(new_n12841_), .Y(new_n20397_));
  OAI21X1  g17961(.A0(new_n2739_), .A1(new_n7942_), .B0(new_n12739_), .Y(new_n20398_));
  AOI21X1  g17962(.A0(new_n20397_), .A1(pi0644), .B0(new_n20398_), .Y(new_n20399_));
  NOR3X1   g17963(.A(new_n20399_), .B(new_n20396_), .C(new_n11882_), .Y(new_n20400_));
  OAI21X1  g17964(.A0(new_n20394_), .A1(new_n12743_), .B0(new_n12739_), .Y(new_n20401_));
  AOI21X1  g17965(.A0(new_n20393_), .A1(new_n12743_), .B0(new_n20401_), .Y(new_n20402_));
  OAI21X1  g17966(.A0(new_n2739_), .A1(new_n7942_), .B0(pi0715), .Y(new_n20403_));
  AOI21X1  g17967(.A0(new_n20397_), .A1(new_n12743_), .B0(new_n20403_), .Y(new_n20404_));
  NOR3X1   g17968(.A(new_n20404_), .B(new_n20402_), .C(pi1160), .Y(new_n20405_));
  OAI21X1  g17969(.A0(new_n20405_), .A1(new_n20400_), .B0(pi0790), .Y(new_n20406_));
  AOI21X1  g17970(.A0(new_n20393_), .A1(new_n12897_), .B0(new_n12898_), .Y(new_n20407_));
  AOI22X1  g17971(.A0(new_n20407_), .A1(new_n20406_), .B0(new_n20308_), .B1(new_n20307_), .Y(po0346));
  AOI21X1  g17972(.A0(pi1093), .A1(pi1092), .B0(pi0190), .Y(new_n20409_));
  INVX1    g17973(.A(new_n20409_), .Y(new_n20410_));
  AOI21X1  g17974(.A0(new_n12178_), .A1(pi0763), .B0(new_n20409_), .Y(new_n20411_));
  AOI21X1  g17975(.A0(new_n12601_), .A1(new_n2739_), .B0(new_n20411_), .Y(new_n20412_));
  AND2X1   g17976(.A(new_n12178_), .B(pi0763), .Y(new_n20413_));
  AND2X1   g17977(.A(new_n20413_), .B(new_n12608_), .Y(new_n20414_));
  INVX1    g17978(.A(new_n20414_), .Y(new_n20415_));
  AOI21X1  g17979(.A0(new_n20415_), .A1(new_n20412_), .B0(new_n12591_), .Y(new_n20416_));
  NOR3X1   g17980(.A(new_n20414_), .B(new_n20409_), .C(pi1155), .Y(new_n20417_));
  OAI21X1  g17981(.A0(new_n20417_), .A1(new_n20416_), .B0(pi0785), .Y(new_n20418_));
  OAI21X1  g17982(.A0(new_n20412_), .A1(pi0785), .B0(new_n20418_), .Y(new_n20419_));
  INVX1    g17983(.A(new_n20419_), .Y(new_n20420_));
  AOI21X1  g17984(.A0(new_n20420_), .A1(new_n12785_), .B0(new_n12615_), .Y(new_n20421_));
  AOI21X1  g17985(.A0(new_n20420_), .A1(new_n12788_), .B0(pi1154), .Y(new_n20422_));
  NOR2X1   g17986(.A(new_n20422_), .B(new_n20421_), .Y(new_n20423_));
  MX2X1    g17987(.A(new_n20423_), .B(new_n20420_), .S0(new_n11887_), .Y(new_n20424_));
  OR2X1    g17988(.A(new_n20424_), .B(pi0789), .Y(new_n20425_));
  AOI21X1  g17989(.A0(new_n20424_), .A1(new_n15910_), .B0(new_n12638_), .Y(new_n20426_));
  AOI21X1  g17990(.A0(new_n20424_), .A1(new_n15912_), .B0(pi1159), .Y(new_n20427_));
  OAI21X1  g17991(.A0(new_n20427_), .A1(new_n20426_), .B0(pi0789), .Y(new_n20428_));
  AND2X1   g17992(.A(new_n20428_), .B(new_n20425_), .Y(new_n20429_));
  INVX1    g17993(.A(new_n20429_), .Y(new_n20430_));
  MX2X1    g17994(.A(new_n20430_), .B(new_n20410_), .S0(new_n12841_), .Y(new_n20431_));
  MX2X1    g17995(.A(new_n20431_), .B(new_n20410_), .S0(new_n12711_), .Y(new_n20432_));
  AOI21X1  g17996(.A0(new_n12566_), .A1(pi0699), .B0(new_n20409_), .Y(new_n20433_));
  INVX1    g17997(.A(new_n20433_), .Y(new_n20434_));
  NOR3X1   g17998(.A(new_n13585_), .B(new_n15535_), .C(pi0625), .Y(new_n20435_));
  OR2X1    g17999(.A(new_n20435_), .B(new_n20433_), .Y(new_n20436_));
  NOR2X1   g18000(.A(new_n20409_), .B(pi1153), .Y(new_n20437_));
  INVX1    g18001(.A(new_n20437_), .Y(new_n20438_));
  OAI21X1  g18002(.A0(new_n20438_), .A1(new_n20435_), .B0(pi0778), .Y(new_n20439_));
  AOI21X1  g18003(.A0(new_n20436_), .A1(pi1153), .B0(new_n20439_), .Y(new_n20440_));
  AOI21X1  g18004(.A0(new_n20434_), .A1(new_n11889_), .B0(new_n20440_), .Y(new_n20441_));
  NOR4X1   g18005(.A(new_n20441_), .B(new_n12765_), .C(new_n12764_), .D(new_n12762_), .Y(new_n20442_));
  INVX1    g18006(.A(new_n20442_), .Y(new_n20443_));
  NOR3X1   g18007(.A(new_n20443_), .B(new_n12870_), .C(new_n12851_), .Y(new_n20444_));
  INVX1    g18008(.A(new_n20444_), .Y(new_n20445_));
  AOI21X1  g18009(.A0(new_n20409_), .A1(pi0647), .B0(pi1157), .Y(new_n20446_));
  OAI21X1  g18010(.A0(new_n20445_), .A1(pi0647), .B0(new_n20446_), .Y(new_n20447_));
  MX2X1    g18011(.A(new_n20444_), .B(new_n20409_), .S0(new_n12705_), .Y(new_n20448_));
  OAI22X1  g18012(.A0(new_n20448_), .A1(new_n14387_), .B0(new_n20447_), .B1(new_n12723_), .Y(new_n20449_));
  AOI21X1  g18013(.A0(new_n20432_), .A1(new_n14385_), .B0(new_n20449_), .Y(new_n20450_));
  NOR2X1   g18014(.A(new_n20450_), .B(new_n11883_), .Y(new_n20451_));
  AOI21X1  g18015(.A0(new_n20410_), .A1(pi0626), .B0(new_n16352_), .Y(new_n20452_));
  OAI21X1  g18016(.A0(new_n20429_), .A1(pi0626), .B0(new_n20452_), .Y(new_n20453_));
  AOI21X1  g18017(.A0(new_n20428_), .A1(new_n20425_), .B0(new_n12664_), .Y(new_n20454_));
  NOR2X1   g18018(.A(new_n20409_), .B(pi0626), .Y(new_n20455_));
  NOR3X1   g18019(.A(new_n20455_), .B(new_n20454_), .C(new_n16356_), .Y(new_n20456_));
  AOI21X1  g18020(.A0(new_n20442_), .A1(new_n12769_), .B0(new_n20456_), .Y(new_n20457_));
  AOI21X1  g18021(.A0(new_n20457_), .A1(new_n20453_), .B0(new_n11885_), .Y(new_n20458_));
  INVX1    g18022(.A(new_n20411_), .Y(new_n20459_));
  AOI21X1  g18023(.A0(new_n20434_), .A1(new_n12171_), .B0(new_n20459_), .Y(new_n20460_));
  NOR3X1   g18024(.A(new_n20433_), .B(new_n12120_), .C(new_n12493_), .Y(new_n20461_));
  OR2X1    g18025(.A(new_n20460_), .B(new_n20461_), .Y(new_n20462_));
  NOR2X1   g18026(.A(new_n20435_), .B(new_n20433_), .Y(new_n20463_));
  OAI21X1  g18027(.A0(new_n20463_), .A1(new_n12494_), .B0(new_n12584_), .Y(new_n20464_));
  AOI21X1  g18028(.A0(new_n20462_), .A1(new_n20437_), .B0(new_n20464_), .Y(new_n20465_));
  NOR3X1   g18029(.A(new_n20461_), .B(new_n20459_), .C(new_n12494_), .Y(new_n20466_));
  OAI21X1  g18030(.A0(new_n20438_), .A1(new_n20435_), .B0(pi0608), .Y(new_n20467_));
  NOR2X1   g18031(.A(new_n20467_), .B(new_n20466_), .Y(new_n20468_));
  OAI21X1  g18032(.A0(new_n20468_), .A1(new_n20465_), .B0(pi0778), .Y(new_n20469_));
  OAI21X1  g18033(.A0(new_n20460_), .A1(pi0778), .B0(new_n20469_), .Y(new_n20470_));
  OAI21X1  g18034(.A0(new_n20441_), .A1(new_n12590_), .B0(new_n12591_), .Y(new_n20471_));
  AOI21X1  g18035(.A0(new_n20470_), .A1(new_n12590_), .B0(new_n20471_), .Y(new_n20472_));
  NOR3X1   g18036(.A(new_n20472_), .B(new_n20416_), .C(pi0660), .Y(new_n20473_));
  OAI21X1  g18037(.A0(new_n20441_), .A1(pi0609), .B0(pi1155), .Y(new_n20474_));
  AOI21X1  g18038(.A0(new_n20470_), .A1(pi0609), .B0(new_n20474_), .Y(new_n20475_));
  NOR3X1   g18039(.A(new_n20475_), .B(new_n20417_), .C(new_n12596_), .Y(new_n20476_));
  OAI21X1  g18040(.A0(new_n20476_), .A1(new_n20473_), .B0(pi0785), .Y(new_n20477_));
  NAND2X1  g18041(.A(new_n20470_), .B(new_n11888_), .Y(new_n20478_));
  AND2X1   g18042(.A(new_n20478_), .B(new_n20477_), .Y(new_n20479_));
  NOR3X1   g18043(.A(new_n20441_), .B(new_n12762_), .C(new_n12614_), .Y(new_n20480_));
  NOR2X1   g18044(.A(new_n20480_), .B(pi1154), .Y(new_n20481_));
  OAI21X1  g18045(.A0(new_n20479_), .A1(pi0618), .B0(new_n20481_), .Y(new_n20482_));
  NOR2X1   g18046(.A(new_n20421_), .B(pi0627), .Y(new_n20483_));
  NOR3X1   g18047(.A(new_n20441_), .B(new_n12762_), .C(pi0618), .Y(new_n20484_));
  NOR2X1   g18048(.A(new_n20484_), .B(new_n12615_), .Y(new_n20485_));
  OAI21X1  g18049(.A0(new_n20479_), .A1(new_n12614_), .B0(new_n20485_), .Y(new_n20486_));
  NOR2X1   g18050(.A(new_n20422_), .B(new_n12622_), .Y(new_n20487_));
  AOI22X1  g18051(.A0(new_n20487_), .A1(new_n20486_), .B0(new_n20483_), .B1(new_n20482_), .Y(new_n20488_));
  MX2X1    g18052(.A(new_n20488_), .B(new_n20479_), .S0(new_n11887_), .Y(new_n20489_));
  OR4X1    g18053(.A(new_n20441_), .B(new_n12764_), .C(new_n12762_), .D(new_n12637_), .Y(new_n20490_));
  AND2X1   g18054(.A(new_n20490_), .B(new_n12638_), .Y(new_n20491_));
  OAI21X1  g18055(.A0(new_n20489_), .A1(pi0619), .B0(new_n20491_), .Y(new_n20492_));
  NOR2X1   g18056(.A(new_n20426_), .B(pi0648), .Y(new_n20493_));
  AND2X1   g18057(.A(new_n20493_), .B(new_n20492_), .Y(new_n20494_));
  INVX1    g18058(.A(new_n20494_), .Y(new_n20495_));
  NOR4X1   g18059(.A(new_n20441_), .B(new_n12764_), .C(new_n12762_), .D(pi0619), .Y(new_n20496_));
  NOR2X1   g18060(.A(new_n20496_), .B(new_n12638_), .Y(new_n20497_));
  OAI21X1  g18061(.A0(new_n20489_), .A1(new_n12637_), .B0(new_n20497_), .Y(new_n20498_));
  NOR2X1   g18062(.A(new_n20427_), .B(new_n12645_), .Y(new_n20499_));
  AOI21X1  g18063(.A0(new_n20499_), .A1(new_n20498_), .B0(new_n11886_), .Y(new_n20500_));
  AOI21X1  g18064(.A0(new_n20489_), .A1(new_n11886_), .B0(new_n14264_), .Y(new_n20501_));
  INVX1    g18065(.A(new_n20501_), .Y(new_n20502_));
  AOI21X1  g18066(.A0(new_n20500_), .A1(new_n20495_), .B0(new_n20502_), .Y(new_n20503_));
  OAI21X1  g18067(.A0(new_n20503_), .A1(new_n20458_), .B0(new_n16350_), .Y(new_n20504_));
  INVX1    g18068(.A(new_n20431_), .Y(new_n20505_));
  AND2X1   g18069(.A(new_n20442_), .B(new_n12852_), .Y(new_n20506_));
  AOI22X1  g18070(.A0(new_n20506_), .A1(new_n14564_), .B0(new_n20505_), .B1(new_n12867_), .Y(new_n20507_));
  AOI22X1  g18071(.A0(new_n20506_), .A1(new_n14566_), .B0(new_n20505_), .B1(new_n12865_), .Y(new_n20508_));
  MX2X1    g18072(.A(new_n20508_), .B(new_n20507_), .S0(new_n12689_), .Y(new_n20509_));
  OAI21X1  g18073(.A0(new_n20509_), .A1(new_n11884_), .B0(new_n14562_), .Y(new_n20510_));
  INVX1    g18074(.A(new_n20510_), .Y(new_n20511_));
  AOI21X1  g18075(.A0(new_n20511_), .A1(new_n20504_), .B0(new_n20451_), .Y(new_n20512_));
  OAI21X1  g18076(.A0(new_n20448_), .A1(new_n12706_), .B0(new_n20447_), .Y(new_n20513_));
  MX2X1    g18077(.A(new_n20513_), .B(new_n20445_), .S0(new_n11883_), .Y(new_n20514_));
  OAI21X1  g18078(.A0(new_n20514_), .A1(pi0644), .B0(pi0715), .Y(new_n20515_));
  AOI21X1  g18079(.A0(new_n20512_), .A1(pi0644), .B0(new_n20515_), .Y(new_n20516_));
  OR4X1    g18080(.A(new_n12734_), .B(new_n2739_), .C(new_n11883_), .D(pi0190), .Y(new_n20517_));
  OAI21X1  g18081(.A0(new_n20432_), .A1(new_n12735_), .B0(new_n20517_), .Y(new_n20518_));
  OAI21X1  g18082(.A0(new_n20410_), .A1(pi0644), .B0(new_n12739_), .Y(new_n20519_));
  AOI21X1  g18083(.A0(new_n20518_), .A1(pi0644), .B0(new_n20519_), .Y(new_n20520_));
  OR2X1    g18084(.A(new_n20520_), .B(new_n11882_), .Y(new_n20521_));
  OAI21X1  g18085(.A0(new_n20514_), .A1(new_n12743_), .B0(new_n12739_), .Y(new_n20522_));
  AOI21X1  g18086(.A0(new_n20512_), .A1(new_n12743_), .B0(new_n20522_), .Y(new_n20523_));
  OAI21X1  g18087(.A0(new_n20410_), .A1(new_n12743_), .B0(pi0715), .Y(new_n20524_));
  AOI21X1  g18088(.A0(new_n20518_), .A1(new_n12743_), .B0(new_n20524_), .Y(new_n20525_));
  OR2X1    g18089(.A(new_n20525_), .B(pi1160), .Y(new_n20526_));
  OAI22X1  g18090(.A0(new_n20526_), .A1(new_n20523_), .B0(new_n20521_), .B1(new_n20516_), .Y(new_n20527_));
  NAND2X1  g18091(.A(new_n20527_), .B(pi0790), .Y(new_n20528_));
  AOI21X1  g18092(.A0(new_n20512_), .A1(new_n12897_), .B0(new_n12898_), .Y(new_n20529_));
  AOI21X1  g18093(.A0(new_n13699_), .A1(new_n3129_), .B0(pi0190), .Y(new_n20530_));
  INVX1    g18094(.A(new_n20530_), .Y(new_n20531_));
  OAI21X1  g18095(.A0(new_n16436_), .A1(new_n10004_), .B0(new_n2996_), .Y(new_n20532_));
  AOI21X1  g18096(.A0(new_n16435_), .A1(new_n10004_), .B0(new_n20532_), .Y(new_n20533_));
  AOI21X1  g18097(.A0(new_n12901_), .A1(new_n10004_), .B0(new_n12568_), .Y(new_n20534_));
  NOR3X1   g18098(.A(new_n20534_), .B(new_n20533_), .C(new_n15535_), .Y(new_n20535_));
  OR2X1    g18099(.A(pi0699), .B(pi0190), .Y(new_n20536_));
  OAI21X1  g18100(.A0(new_n20536_), .A1(new_n13699_), .B0(new_n3129_), .Y(new_n20537_));
  OAI22X1  g18101(.A0(new_n20537_), .A1(new_n20535_), .B0(new_n3129_), .B1(new_n10004_), .Y(new_n20538_));
  AND2X1   g18102(.A(new_n20538_), .B(new_n11889_), .Y(new_n20539_));
  AOI21X1  g18103(.A0(new_n20530_), .A1(new_n12493_), .B0(new_n12494_), .Y(new_n20540_));
  OAI21X1  g18104(.A0(new_n20538_), .A1(new_n12493_), .B0(new_n20540_), .Y(new_n20541_));
  AOI21X1  g18105(.A0(new_n20530_), .A1(pi0625), .B0(pi1153), .Y(new_n20542_));
  OAI21X1  g18106(.A0(new_n20538_), .A1(pi0625), .B0(new_n20542_), .Y(new_n20543_));
  AOI21X1  g18107(.A0(new_n20543_), .A1(new_n20541_), .B0(new_n11889_), .Y(new_n20544_));
  NOR2X1   g18108(.A(new_n20544_), .B(new_n20539_), .Y(new_n20545_));
  MX2X1    g18109(.A(new_n20545_), .B(new_n20530_), .S0(new_n12618_), .Y(new_n20546_));
  AND2X1   g18110(.A(new_n20530_), .B(new_n12641_), .Y(new_n20547_));
  AOI21X1  g18111(.A0(new_n20546_), .A1(new_n14198_), .B0(new_n20547_), .Y(new_n20548_));
  MX2X1    g18112(.A(new_n20548_), .B(new_n20531_), .S0(new_n12659_), .Y(new_n20549_));
  MX2X1    g18113(.A(new_n20549_), .B(new_n20531_), .S0(new_n12691_), .Y(new_n20550_));
  MX2X1    g18114(.A(new_n20550_), .B(new_n20531_), .S0(pi0628), .Y(new_n20551_));
  MX2X1    g18115(.A(new_n20550_), .B(new_n20531_), .S0(new_n12683_), .Y(new_n20552_));
  MX2X1    g18116(.A(new_n20552_), .B(new_n20551_), .S0(new_n12684_), .Y(new_n20553_));
  MX2X1    g18117(.A(new_n20553_), .B(new_n20550_), .S0(new_n11884_), .Y(new_n20554_));
  MX2X1    g18118(.A(new_n20554_), .B(new_n20531_), .S0(pi0647), .Y(new_n20555_));
  MX2X1    g18119(.A(new_n20554_), .B(new_n20531_), .S0(new_n12705_), .Y(new_n20556_));
  MX2X1    g18120(.A(new_n20556_), .B(new_n20555_), .S0(new_n12706_), .Y(new_n20557_));
  MX2X1    g18121(.A(new_n20557_), .B(new_n20554_), .S0(new_n11883_), .Y(new_n20558_));
  OAI21X1  g18122(.A0(new_n20558_), .A1(pi0644), .B0(pi0715), .Y(new_n20559_));
  OAI22X1  g18123(.A0(new_n12904_), .A1(new_n10004_), .B0(new_n12089_), .B1(pi0763), .Y(new_n20560_));
  NAND2X1  g18124(.A(new_n20560_), .B(pi0039), .Y(new_n20561_));
  AND2X1   g18125(.A(pi0763), .B(new_n10004_), .Y(new_n20562_));
  AOI21X1  g18126(.A0(new_n13683_), .A1(new_n2959_), .B0(new_n15495_), .Y(new_n20563_));
  OAI21X1  g18127(.A0(new_n20563_), .A1(new_n10004_), .B0(new_n15499_), .Y(new_n20564_));
  AOI21X1  g18128(.A0(new_n20562_), .A1(new_n12162_), .B0(new_n20564_), .Y(new_n20565_));
  AOI21X1  g18129(.A0(new_n20565_), .A1(new_n20561_), .B0(pi0038), .Y(new_n20566_));
  OAI21X1  g18130(.A0(new_n12202_), .A1(pi0190), .B0(pi0038), .Y(new_n20567_));
  AOI21X1  g18131(.A0(new_n12205_), .A1(pi0763), .B0(new_n20567_), .Y(new_n20568_));
  NOR2X1   g18132(.A(new_n20568_), .B(new_n20566_), .Y(new_n20569_));
  MX2X1    g18133(.A(new_n20569_), .B(new_n10004_), .S0(new_n3810_), .Y(new_n20570_));
  MX2X1    g18134(.A(new_n20570_), .B(new_n20530_), .S0(new_n12601_), .Y(new_n20571_));
  NOR2X1   g18135(.A(new_n20570_), .B(new_n12601_), .Y(new_n20572_));
  AOI22X1  g18136(.A0(new_n20572_), .A1(pi0609), .B0(new_n20531_), .B1(new_n13430_), .Y(new_n20573_));
  AOI22X1  g18137(.A0(new_n20572_), .A1(new_n12590_), .B0(new_n20531_), .B1(new_n13436_), .Y(new_n20574_));
  MX2X1    g18138(.A(new_n20574_), .B(new_n20573_), .S0(pi1155), .Y(new_n20575_));
  MX2X1    g18139(.A(new_n20575_), .B(new_n20571_), .S0(new_n11888_), .Y(new_n20576_));
  OAI21X1  g18140(.A0(new_n20531_), .A1(pi0618), .B0(pi1154), .Y(new_n20577_));
  AOI21X1  g18141(.A0(new_n20576_), .A1(pi0618), .B0(new_n20577_), .Y(new_n20578_));
  OAI21X1  g18142(.A0(new_n20531_), .A1(new_n12614_), .B0(new_n12615_), .Y(new_n20579_));
  AOI21X1  g18143(.A0(new_n20576_), .A1(new_n12614_), .B0(new_n20579_), .Y(new_n20580_));
  NOR2X1   g18144(.A(new_n20580_), .B(new_n20578_), .Y(new_n20581_));
  MX2X1    g18145(.A(new_n20581_), .B(new_n20576_), .S0(new_n11887_), .Y(new_n20582_));
  OAI21X1  g18146(.A0(new_n20531_), .A1(pi0619), .B0(pi1159), .Y(new_n20583_));
  AOI21X1  g18147(.A0(new_n20582_), .A1(pi0619), .B0(new_n20583_), .Y(new_n20584_));
  OAI21X1  g18148(.A0(new_n20531_), .A1(new_n12637_), .B0(new_n12638_), .Y(new_n20585_));
  AOI21X1  g18149(.A0(new_n20582_), .A1(new_n12637_), .B0(new_n20585_), .Y(new_n20586_));
  NOR2X1   g18150(.A(new_n20586_), .B(new_n20584_), .Y(new_n20587_));
  MX2X1    g18151(.A(new_n20587_), .B(new_n20582_), .S0(new_n11886_), .Y(new_n20588_));
  MX2X1    g18152(.A(new_n20588_), .B(new_n20530_), .S0(new_n12841_), .Y(new_n20589_));
  MX2X1    g18153(.A(new_n20589_), .B(new_n20530_), .S0(new_n12711_), .Y(new_n20590_));
  MX2X1    g18154(.A(new_n20590_), .B(new_n20530_), .S0(new_n12735_), .Y(new_n20591_));
  OAI21X1  g18155(.A0(new_n20531_), .A1(pi0644), .B0(new_n12739_), .Y(new_n20592_));
  AOI21X1  g18156(.A0(new_n20591_), .A1(pi0644), .B0(new_n20592_), .Y(new_n20593_));
  NOR2X1   g18157(.A(new_n20593_), .B(new_n11882_), .Y(new_n20594_));
  OAI21X1  g18158(.A0(new_n20558_), .A1(new_n12743_), .B0(new_n12739_), .Y(new_n20595_));
  OAI21X1  g18159(.A0(new_n20531_), .A1(new_n12743_), .B0(pi0715), .Y(new_n20596_));
  AOI21X1  g18160(.A0(new_n20591_), .A1(new_n12743_), .B0(new_n20596_), .Y(new_n20597_));
  NOR2X1   g18161(.A(new_n20597_), .B(pi1160), .Y(new_n20598_));
  AOI22X1  g18162(.A0(new_n20598_), .A1(new_n20595_), .B0(new_n20594_), .B1(new_n20559_), .Y(new_n20599_));
  NOR3X1   g18163(.A(new_n20597_), .B(pi1160), .C(pi0644), .Y(new_n20600_));
  NOR3X1   g18164(.A(new_n20593_), .B(new_n11882_), .C(new_n12743_), .Y(new_n20601_));
  NOR3X1   g18165(.A(new_n20601_), .B(new_n20600_), .C(new_n12897_), .Y(new_n20602_));
  AOI22X1  g18166(.A0(new_n20552_), .A1(new_n12707_), .B0(new_n20551_), .B1(new_n12709_), .Y(new_n20603_));
  OAI21X1  g18167(.A0(new_n20589_), .A1(new_n14395_), .B0(new_n20603_), .Y(new_n20604_));
  NOR3X1   g18168(.A(new_n20568_), .B(new_n20566_), .C(pi0699), .Y(new_n20605_));
  INVX1    g18169(.A(new_n20605_), .Y(new_n20606_));
  AOI21X1  g18170(.A0(new_n13989_), .A1(pi0190), .B0(pi0763), .Y(new_n20607_));
  OAI21X1  g18171(.A0(new_n13986_), .A1(pi0190), .B0(new_n20607_), .Y(new_n20608_));
  OAI21X1  g18172(.A0(new_n12440_), .A1(pi0190), .B0(pi0763), .Y(new_n20609_));
  AOI21X1  g18173(.A0(new_n12401_), .A1(pi0190), .B0(new_n20609_), .Y(new_n20610_));
  NOR2X1   g18174(.A(new_n20610_), .B(new_n2959_), .Y(new_n20611_));
  AND2X1   g18175(.A(new_n20611_), .B(new_n20608_), .Y(new_n20612_));
  AOI21X1  g18176(.A0(new_n13995_), .A1(pi0190), .B0(pi0763), .Y(new_n20613_));
  OAI21X1  g18177(.A0(new_n13996_), .A1(pi0190), .B0(new_n20613_), .Y(new_n20614_));
  AOI21X1  g18178(.A0(new_n12453_), .A1(new_n12104_), .B0(pi0190), .Y(new_n20615_));
  INVX1    g18179(.A(new_n20615_), .Y(new_n20616_));
  AOI21X1  g18180(.A0(new_n12929_), .A1(pi0190), .B0(new_n15495_), .Y(new_n20617_));
  AOI21X1  g18181(.A0(new_n20617_), .A1(new_n20616_), .B0(pi0039), .Y(new_n20618_));
  AOI21X1  g18182(.A0(new_n20618_), .A1(new_n20614_), .B0(pi0038), .Y(new_n20619_));
  INVX1    g18183(.A(new_n20619_), .Y(new_n20620_));
  AOI21X1  g18184(.A0(new_n16526_), .A1(new_n15495_), .B0(new_n12478_), .Y(new_n20621_));
  OAI21X1  g18185(.A0(new_n20621_), .A1(pi0039), .B0(new_n10004_), .Y(new_n20622_));
  OAI21X1  g18186(.A0(new_n20413_), .A1(new_n13576_), .B0(pi0190), .Y(new_n20623_));
  OAI21X1  g18187(.A0(new_n20623_), .A1(new_n14411_), .B0(pi0038), .Y(new_n20624_));
  INVX1    g18188(.A(new_n20624_), .Y(new_n20625_));
  AOI21X1  g18189(.A0(new_n20625_), .A1(new_n20622_), .B0(new_n15535_), .Y(new_n20626_));
  OAI21X1  g18190(.A0(new_n20620_), .A1(new_n20612_), .B0(new_n20626_), .Y(new_n20627_));
  AND2X1   g18191(.A(new_n20627_), .B(new_n3129_), .Y(new_n20628_));
  AOI22X1  g18192(.A0(new_n20628_), .A1(new_n20606_), .B0(new_n3810_), .B1(pi0190), .Y(new_n20629_));
  INVX1    g18193(.A(new_n20629_), .Y(new_n20630_));
  AOI21X1  g18194(.A0(new_n20570_), .A1(pi0625), .B0(pi1153), .Y(new_n20631_));
  OAI21X1  g18195(.A0(new_n20630_), .A1(pi0625), .B0(new_n20631_), .Y(new_n20632_));
  AND2X1   g18196(.A(new_n20541_), .B(new_n12584_), .Y(new_n20633_));
  AOI21X1  g18197(.A0(new_n20570_), .A1(new_n12493_), .B0(new_n12494_), .Y(new_n20634_));
  OAI21X1  g18198(.A0(new_n20630_), .A1(new_n12493_), .B0(new_n20634_), .Y(new_n20635_));
  AND2X1   g18199(.A(new_n20543_), .B(pi0608), .Y(new_n20636_));
  AOI22X1  g18200(.A0(new_n20636_), .A1(new_n20635_), .B0(new_n20633_), .B1(new_n20632_), .Y(new_n20637_));
  MX2X1    g18201(.A(new_n20637_), .B(new_n20630_), .S0(new_n11889_), .Y(new_n20638_));
  AOI21X1  g18202(.A0(new_n20545_), .A1(pi0609), .B0(pi1155), .Y(new_n20639_));
  OAI21X1  g18203(.A0(new_n20638_), .A1(pi0609), .B0(new_n20639_), .Y(new_n20640_));
  OAI21X1  g18204(.A0(new_n20573_), .A1(new_n12591_), .B0(new_n12596_), .Y(new_n20641_));
  INVX1    g18205(.A(new_n20641_), .Y(new_n20642_));
  AOI21X1  g18206(.A0(new_n20545_), .A1(new_n12590_), .B0(new_n12591_), .Y(new_n20643_));
  OAI21X1  g18207(.A0(new_n20638_), .A1(new_n12590_), .B0(new_n20643_), .Y(new_n20644_));
  OAI21X1  g18208(.A0(new_n20574_), .A1(pi1155), .B0(pi0660), .Y(new_n20645_));
  INVX1    g18209(.A(new_n20645_), .Y(new_n20646_));
  AOI22X1  g18210(.A0(new_n20646_), .A1(new_n20644_), .B0(new_n20642_), .B1(new_n20640_), .Y(new_n20647_));
  MX2X1    g18211(.A(new_n20647_), .B(new_n20638_), .S0(new_n11888_), .Y(new_n20648_));
  AOI21X1  g18212(.A0(new_n20546_), .A1(pi0618), .B0(pi1154), .Y(new_n20649_));
  OAI21X1  g18213(.A0(new_n20648_), .A1(pi0618), .B0(new_n20649_), .Y(new_n20650_));
  NOR2X1   g18214(.A(new_n20578_), .B(pi0627), .Y(new_n20651_));
  AOI21X1  g18215(.A0(new_n20546_), .A1(new_n12614_), .B0(new_n12615_), .Y(new_n20652_));
  OAI21X1  g18216(.A0(new_n20648_), .A1(new_n12614_), .B0(new_n20652_), .Y(new_n20653_));
  NOR2X1   g18217(.A(new_n20580_), .B(new_n12622_), .Y(new_n20654_));
  AOI22X1  g18218(.A0(new_n20654_), .A1(new_n20653_), .B0(new_n20651_), .B1(new_n20650_), .Y(new_n20655_));
  MX2X1    g18219(.A(new_n20655_), .B(new_n20648_), .S0(new_n11887_), .Y(new_n20656_));
  INVX1    g18220(.A(new_n20656_), .Y(new_n20657_));
  OAI21X1  g18221(.A0(new_n20548_), .A1(new_n12637_), .B0(new_n12638_), .Y(new_n20658_));
  AOI21X1  g18222(.A0(new_n20657_), .A1(new_n12637_), .B0(new_n20658_), .Y(new_n20659_));
  NOR3X1   g18223(.A(new_n20659_), .B(new_n20584_), .C(pi0648), .Y(new_n20660_));
  OAI21X1  g18224(.A0(new_n20548_), .A1(pi0619), .B0(pi1159), .Y(new_n20661_));
  AOI21X1  g18225(.A0(new_n20657_), .A1(pi0619), .B0(new_n20661_), .Y(new_n20662_));
  OR2X1    g18226(.A(new_n20586_), .B(new_n12645_), .Y(new_n20663_));
  OAI21X1  g18227(.A0(new_n20663_), .A1(new_n20662_), .B0(pi0789), .Y(new_n20664_));
  AOI21X1  g18228(.A0(new_n20656_), .A1(new_n11886_), .B0(new_n14264_), .Y(new_n20665_));
  OAI21X1  g18229(.A0(new_n20664_), .A1(new_n20660_), .B0(new_n20665_), .Y(new_n20666_));
  AOI21X1  g18230(.A0(new_n20531_), .A1(pi0626), .B0(new_n16352_), .Y(new_n20667_));
  OAI21X1  g18231(.A0(new_n20588_), .A1(pi0626), .B0(new_n20667_), .Y(new_n20668_));
  AOI21X1  g18232(.A0(new_n20531_), .A1(new_n12664_), .B0(new_n16356_), .Y(new_n20669_));
  OAI21X1  g18233(.A0(new_n20588_), .A1(new_n12664_), .B0(new_n20669_), .Y(new_n20670_));
  OR2X1    g18234(.A(new_n20549_), .B(new_n12770_), .Y(new_n20671_));
  NAND3X1  g18235(.A(new_n20671_), .B(new_n20670_), .C(new_n20668_), .Y(new_n20672_));
  AOI21X1  g18236(.A0(new_n20672_), .A1(pi0788), .B0(new_n14273_), .Y(new_n20673_));
  AOI22X1  g18237(.A0(new_n20673_), .A1(new_n20666_), .B0(new_n20604_), .B1(pi0792), .Y(new_n20674_));
  NOR2X1   g18238(.A(new_n20590_), .B(new_n14384_), .Y(new_n20675_));
  AND2X1   g18239(.A(new_n20556_), .B(new_n14386_), .Y(new_n20676_));
  AND2X1   g18240(.A(new_n20555_), .B(new_n14388_), .Y(new_n20677_));
  OR2X1    g18241(.A(new_n20677_), .B(new_n20676_), .Y(new_n20678_));
  OAI21X1  g18242(.A0(new_n20678_), .A1(new_n20675_), .B0(pi0787), .Y(new_n20679_));
  OAI21X1  g18243(.A0(new_n20674_), .A1(new_n14269_), .B0(new_n20679_), .Y(new_n20680_));
  OAI22X1  g18244(.A0(new_n20680_), .A1(new_n20602_), .B0(new_n20599_), .B1(new_n12897_), .Y(new_n20681_));
  OAI21X1  g18245(.A0(new_n6520_), .A1(pi0190), .B0(new_n12898_), .Y(new_n20682_));
  AOI21X1  g18246(.A0(new_n20681_), .A1(new_n6520_), .B0(new_n20682_), .Y(new_n20683_));
  AOI21X1  g18247(.A0(new_n20529_), .A1(new_n20528_), .B0(new_n20683_), .Y(po0347));
  AOI21X1  g18248(.A0(pi1093), .A1(pi1092), .B0(pi0191), .Y(new_n20685_));
  INVX1    g18249(.A(new_n20685_), .Y(new_n20686_));
  AOI21X1  g18250(.A0(new_n12178_), .A1(pi0746), .B0(new_n20685_), .Y(new_n20687_));
  AOI21X1  g18251(.A0(new_n12601_), .A1(new_n2739_), .B0(new_n20687_), .Y(new_n20688_));
  AND2X1   g18252(.A(new_n12178_), .B(pi0746), .Y(new_n20689_));
  AND2X1   g18253(.A(new_n20689_), .B(new_n12608_), .Y(new_n20690_));
  INVX1    g18254(.A(new_n20690_), .Y(new_n20691_));
  AOI21X1  g18255(.A0(new_n20691_), .A1(new_n20688_), .B0(new_n12591_), .Y(new_n20692_));
  NOR3X1   g18256(.A(new_n20690_), .B(new_n20685_), .C(pi1155), .Y(new_n20693_));
  OAI21X1  g18257(.A0(new_n20693_), .A1(new_n20692_), .B0(pi0785), .Y(new_n20694_));
  OAI21X1  g18258(.A0(new_n20688_), .A1(pi0785), .B0(new_n20694_), .Y(new_n20695_));
  INVX1    g18259(.A(new_n20695_), .Y(new_n20696_));
  AOI21X1  g18260(.A0(new_n20696_), .A1(new_n12785_), .B0(new_n12615_), .Y(new_n20697_));
  AOI21X1  g18261(.A0(new_n20696_), .A1(new_n12788_), .B0(pi1154), .Y(new_n20698_));
  NOR2X1   g18262(.A(new_n20698_), .B(new_n20697_), .Y(new_n20699_));
  MX2X1    g18263(.A(new_n20699_), .B(new_n20696_), .S0(new_n11887_), .Y(new_n20700_));
  OR2X1    g18264(.A(new_n20700_), .B(pi0789), .Y(new_n20701_));
  AOI21X1  g18265(.A0(new_n20700_), .A1(new_n15910_), .B0(new_n12638_), .Y(new_n20702_));
  AOI21X1  g18266(.A0(new_n20700_), .A1(new_n15912_), .B0(pi1159), .Y(new_n20703_));
  OAI21X1  g18267(.A0(new_n20703_), .A1(new_n20702_), .B0(pi0789), .Y(new_n20704_));
  AND2X1   g18268(.A(new_n20704_), .B(new_n20701_), .Y(new_n20705_));
  INVX1    g18269(.A(new_n20705_), .Y(new_n20706_));
  MX2X1    g18270(.A(new_n20706_), .B(new_n20686_), .S0(new_n12841_), .Y(new_n20707_));
  MX2X1    g18271(.A(new_n20707_), .B(new_n20686_), .S0(new_n12711_), .Y(new_n20708_));
  AOI21X1  g18272(.A0(new_n12566_), .A1(pi0729), .B0(new_n20685_), .Y(new_n20709_));
  INVX1    g18273(.A(new_n20709_), .Y(new_n20710_));
  NOR3X1   g18274(.A(new_n13585_), .B(new_n15585_), .C(pi0625), .Y(new_n20711_));
  OR2X1    g18275(.A(new_n20711_), .B(new_n20709_), .Y(new_n20712_));
  NOR2X1   g18276(.A(new_n20685_), .B(pi1153), .Y(new_n20713_));
  INVX1    g18277(.A(new_n20713_), .Y(new_n20714_));
  OAI21X1  g18278(.A0(new_n20714_), .A1(new_n20711_), .B0(pi0778), .Y(new_n20715_));
  AOI21X1  g18279(.A0(new_n20712_), .A1(pi1153), .B0(new_n20715_), .Y(new_n20716_));
  AOI21X1  g18280(.A0(new_n20710_), .A1(new_n11889_), .B0(new_n20716_), .Y(new_n20717_));
  NOR4X1   g18281(.A(new_n20717_), .B(new_n12765_), .C(new_n12764_), .D(new_n12762_), .Y(new_n20718_));
  INVX1    g18282(.A(new_n20718_), .Y(new_n20719_));
  NOR3X1   g18283(.A(new_n20719_), .B(new_n12870_), .C(new_n12851_), .Y(new_n20720_));
  INVX1    g18284(.A(new_n20720_), .Y(new_n20721_));
  AOI21X1  g18285(.A0(new_n20685_), .A1(pi0647), .B0(pi1157), .Y(new_n20722_));
  OAI21X1  g18286(.A0(new_n20721_), .A1(pi0647), .B0(new_n20722_), .Y(new_n20723_));
  MX2X1    g18287(.A(new_n20720_), .B(new_n20685_), .S0(new_n12705_), .Y(new_n20724_));
  OAI22X1  g18288(.A0(new_n20724_), .A1(new_n14387_), .B0(new_n20723_), .B1(new_n12723_), .Y(new_n20725_));
  AOI21X1  g18289(.A0(new_n20708_), .A1(new_n14385_), .B0(new_n20725_), .Y(new_n20726_));
  NOR2X1   g18290(.A(new_n20726_), .B(new_n11883_), .Y(new_n20727_));
  AOI21X1  g18291(.A0(new_n20686_), .A1(pi0626), .B0(new_n16352_), .Y(new_n20728_));
  OAI21X1  g18292(.A0(new_n20705_), .A1(pi0626), .B0(new_n20728_), .Y(new_n20729_));
  AOI21X1  g18293(.A0(new_n20704_), .A1(new_n20701_), .B0(new_n12664_), .Y(new_n20730_));
  NOR2X1   g18294(.A(new_n20685_), .B(pi0626), .Y(new_n20731_));
  NOR3X1   g18295(.A(new_n20731_), .B(new_n20730_), .C(new_n16356_), .Y(new_n20732_));
  AOI21X1  g18296(.A0(new_n20718_), .A1(new_n12769_), .B0(new_n20732_), .Y(new_n20733_));
  AOI21X1  g18297(.A0(new_n20733_), .A1(new_n20729_), .B0(new_n11885_), .Y(new_n20734_));
  INVX1    g18298(.A(new_n20687_), .Y(new_n20735_));
  AOI21X1  g18299(.A0(new_n20710_), .A1(new_n12171_), .B0(new_n20735_), .Y(new_n20736_));
  NOR3X1   g18300(.A(new_n20709_), .B(new_n12120_), .C(new_n12493_), .Y(new_n20737_));
  OR2X1    g18301(.A(new_n20736_), .B(new_n20737_), .Y(new_n20738_));
  NOR2X1   g18302(.A(new_n20711_), .B(new_n20709_), .Y(new_n20739_));
  OAI21X1  g18303(.A0(new_n20739_), .A1(new_n12494_), .B0(new_n12584_), .Y(new_n20740_));
  AOI21X1  g18304(.A0(new_n20738_), .A1(new_n20713_), .B0(new_n20740_), .Y(new_n20741_));
  NOR3X1   g18305(.A(new_n20737_), .B(new_n20735_), .C(new_n12494_), .Y(new_n20742_));
  OAI21X1  g18306(.A0(new_n20714_), .A1(new_n20711_), .B0(pi0608), .Y(new_n20743_));
  NOR2X1   g18307(.A(new_n20743_), .B(new_n20742_), .Y(new_n20744_));
  OAI21X1  g18308(.A0(new_n20744_), .A1(new_n20741_), .B0(pi0778), .Y(new_n20745_));
  OAI21X1  g18309(.A0(new_n20736_), .A1(pi0778), .B0(new_n20745_), .Y(new_n20746_));
  OAI21X1  g18310(.A0(new_n20717_), .A1(new_n12590_), .B0(new_n12591_), .Y(new_n20747_));
  AOI21X1  g18311(.A0(new_n20746_), .A1(new_n12590_), .B0(new_n20747_), .Y(new_n20748_));
  NOR3X1   g18312(.A(new_n20748_), .B(new_n20692_), .C(pi0660), .Y(new_n20749_));
  OAI21X1  g18313(.A0(new_n20717_), .A1(pi0609), .B0(pi1155), .Y(new_n20750_));
  AOI21X1  g18314(.A0(new_n20746_), .A1(pi0609), .B0(new_n20750_), .Y(new_n20751_));
  NOR3X1   g18315(.A(new_n20751_), .B(new_n20693_), .C(new_n12596_), .Y(new_n20752_));
  OAI21X1  g18316(.A0(new_n20752_), .A1(new_n20749_), .B0(pi0785), .Y(new_n20753_));
  NAND2X1  g18317(.A(new_n20746_), .B(new_n11888_), .Y(new_n20754_));
  AND2X1   g18318(.A(new_n20754_), .B(new_n20753_), .Y(new_n20755_));
  NOR3X1   g18319(.A(new_n20717_), .B(new_n12762_), .C(new_n12614_), .Y(new_n20756_));
  NOR2X1   g18320(.A(new_n20756_), .B(pi1154), .Y(new_n20757_));
  OAI21X1  g18321(.A0(new_n20755_), .A1(pi0618), .B0(new_n20757_), .Y(new_n20758_));
  NOR2X1   g18322(.A(new_n20697_), .B(pi0627), .Y(new_n20759_));
  NOR3X1   g18323(.A(new_n20717_), .B(new_n12762_), .C(pi0618), .Y(new_n20760_));
  NOR2X1   g18324(.A(new_n20760_), .B(new_n12615_), .Y(new_n20761_));
  OAI21X1  g18325(.A0(new_n20755_), .A1(new_n12614_), .B0(new_n20761_), .Y(new_n20762_));
  NOR2X1   g18326(.A(new_n20698_), .B(new_n12622_), .Y(new_n20763_));
  AOI22X1  g18327(.A0(new_n20763_), .A1(new_n20762_), .B0(new_n20759_), .B1(new_n20758_), .Y(new_n20764_));
  MX2X1    g18328(.A(new_n20764_), .B(new_n20755_), .S0(new_n11887_), .Y(new_n20765_));
  OR4X1    g18329(.A(new_n20717_), .B(new_n12764_), .C(new_n12762_), .D(new_n12637_), .Y(new_n20766_));
  AND2X1   g18330(.A(new_n20766_), .B(new_n12638_), .Y(new_n20767_));
  OAI21X1  g18331(.A0(new_n20765_), .A1(pi0619), .B0(new_n20767_), .Y(new_n20768_));
  NOR2X1   g18332(.A(new_n20702_), .B(pi0648), .Y(new_n20769_));
  AND2X1   g18333(.A(new_n20769_), .B(new_n20768_), .Y(new_n20770_));
  INVX1    g18334(.A(new_n20770_), .Y(new_n20771_));
  NOR4X1   g18335(.A(new_n20717_), .B(new_n12764_), .C(new_n12762_), .D(pi0619), .Y(new_n20772_));
  NOR2X1   g18336(.A(new_n20772_), .B(new_n12638_), .Y(new_n20773_));
  OAI21X1  g18337(.A0(new_n20765_), .A1(new_n12637_), .B0(new_n20773_), .Y(new_n20774_));
  NOR2X1   g18338(.A(new_n20703_), .B(new_n12645_), .Y(new_n20775_));
  AOI21X1  g18339(.A0(new_n20775_), .A1(new_n20774_), .B0(new_n11886_), .Y(new_n20776_));
  AOI21X1  g18340(.A0(new_n20765_), .A1(new_n11886_), .B0(new_n14264_), .Y(new_n20777_));
  INVX1    g18341(.A(new_n20777_), .Y(new_n20778_));
  AOI21X1  g18342(.A0(new_n20776_), .A1(new_n20771_), .B0(new_n20778_), .Y(new_n20779_));
  OAI21X1  g18343(.A0(new_n20779_), .A1(new_n20734_), .B0(new_n16350_), .Y(new_n20780_));
  INVX1    g18344(.A(new_n20707_), .Y(new_n20781_));
  AND2X1   g18345(.A(new_n20718_), .B(new_n12852_), .Y(new_n20782_));
  AOI22X1  g18346(.A0(new_n20782_), .A1(new_n14564_), .B0(new_n20781_), .B1(new_n12867_), .Y(new_n20783_));
  AOI22X1  g18347(.A0(new_n20782_), .A1(new_n14566_), .B0(new_n20781_), .B1(new_n12865_), .Y(new_n20784_));
  MX2X1    g18348(.A(new_n20784_), .B(new_n20783_), .S0(new_n12689_), .Y(new_n20785_));
  OAI21X1  g18349(.A0(new_n20785_), .A1(new_n11884_), .B0(new_n14562_), .Y(new_n20786_));
  INVX1    g18350(.A(new_n20786_), .Y(new_n20787_));
  AOI21X1  g18351(.A0(new_n20787_), .A1(new_n20780_), .B0(new_n20727_), .Y(new_n20788_));
  OAI21X1  g18352(.A0(new_n20724_), .A1(new_n12706_), .B0(new_n20723_), .Y(new_n20789_));
  MX2X1    g18353(.A(new_n20789_), .B(new_n20721_), .S0(new_n11883_), .Y(new_n20790_));
  OAI21X1  g18354(.A0(new_n20790_), .A1(pi0644), .B0(pi0715), .Y(new_n20791_));
  AOI21X1  g18355(.A0(new_n20788_), .A1(pi0644), .B0(new_n20791_), .Y(new_n20792_));
  OR4X1    g18356(.A(new_n12734_), .B(new_n2739_), .C(new_n11883_), .D(pi0191), .Y(new_n20793_));
  OAI21X1  g18357(.A0(new_n20708_), .A1(new_n12735_), .B0(new_n20793_), .Y(new_n20794_));
  OAI21X1  g18358(.A0(new_n20686_), .A1(pi0644), .B0(new_n12739_), .Y(new_n20795_));
  AOI21X1  g18359(.A0(new_n20794_), .A1(pi0644), .B0(new_n20795_), .Y(new_n20796_));
  OR2X1    g18360(.A(new_n20796_), .B(new_n11882_), .Y(new_n20797_));
  OAI21X1  g18361(.A0(new_n20790_), .A1(new_n12743_), .B0(new_n12739_), .Y(new_n20798_));
  AOI21X1  g18362(.A0(new_n20788_), .A1(new_n12743_), .B0(new_n20798_), .Y(new_n20799_));
  OAI21X1  g18363(.A0(new_n20686_), .A1(new_n12743_), .B0(pi0715), .Y(new_n20800_));
  AOI21X1  g18364(.A0(new_n20794_), .A1(new_n12743_), .B0(new_n20800_), .Y(new_n20801_));
  OR2X1    g18365(.A(new_n20801_), .B(pi1160), .Y(new_n20802_));
  OAI22X1  g18366(.A0(new_n20802_), .A1(new_n20799_), .B0(new_n20797_), .B1(new_n20792_), .Y(new_n20803_));
  NAND2X1  g18367(.A(new_n20803_), .B(pi0790), .Y(new_n20804_));
  AOI21X1  g18368(.A0(new_n20788_), .A1(new_n12897_), .B0(new_n12898_), .Y(new_n20805_));
  AOI21X1  g18369(.A0(new_n13699_), .A1(new_n3129_), .B0(pi0191), .Y(new_n20806_));
  INVX1    g18370(.A(new_n20806_), .Y(new_n20807_));
  OAI21X1  g18371(.A0(new_n16436_), .A1(new_n6844_), .B0(new_n2996_), .Y(new_n20808_));
  AOI21X1  g18372(.A0(new_n16435_), .A1(new_n6844_), .B0(new_n20808_), .Y(new_n20809_));
  AOI21X1  g18373(.A0(new_n12901_), .A1(new_n6844_), .B0(new_n12568_), .Y(new_n20810_));
  NOR3X1   g18374(.A(new_n20810_), .B(new_n20809_), .C(new_n15585_), .Y(new_n20811_));
  OR2X1    g18375(.A(pi0729), .B(pi0191), .Y(new_n20812_));
  OAI21X1  g18376(.A0(new_n20812_), .A1(new_n13699_), .B0(new_n3129_), .Y(new_n20813_));
  OAI22X1  g18377(.A0(new_n20813_), .A1(new_n20811_), .B0(new_n3129_), .B1(new_n6844_), .Y(new_n20814_));
  AND2X1   g18378(.A(new_n20814_), .B(new_n11889_), .Y(new_n20815_));
  AOI21X1  g18379(.A0(new_n20806_), .A1(new_n12493_), .B0(new_n12494_), .Y(new_n20816_));
  OAI21X1  g18380(.A0(new_n20814_), .A1(new_n12493_), .B0(new_n20816_), .Y(new_n20817_));
  AOI21X1  g18381(.A0(new_n20806_), .A1(pi0625), .B0(pi1153), .Y(new_n20818_));
  OAI21X1  g18382(.A0(new_n20814_), .A1(pi0625), .B0(new_n20818_), .Y(new_n20819_));
  AOI21X1  g18383(.A0(new_n20819_), .A1(new_n20817_), .B0(new_n11889_), .Y(new_n20820_));
  NOR2X1   g18384(.A(new_n20820_), .B(new_n20815_), .Y(new_n20821_));
  MX2X1    g18385(.A(new_n20821_), .B(new_n20806_), .S0(new_n12618_), .Y(new_n20822_));
  AND2X1   g18386(.A(new_n20806_), .B(new_n12641_), .Y(new_n20823_));
  AOI21X1  g18387(.A0(new_n20822_), .A1(new_n14198_), .B0(new_n20823_), .Y(new_n20824_));
  MX2X1    g18388(.A(new_n20824_), .B(new_n20807_), .S0(new_n12659_), .Y(new_n20825_));
  MX2X1    g18389(.A(new_n20825_), .B(new_n20807_), .S0(new_n12691_), .Y(new_n20826_));
  MX2X1    g18390(.A(new_n20826_), .B(new_n20807_), .S0(pi0628), .Y(new_n20827_));
  MX2X1    g18391(.A(new_n20826_), .B(new_n20807_), .S0(new_n12683_), .Y(new_n20828_));
  MX2X1    g18392(.A(new_n20828_), .B(new_n20827_), .S0(new_n12684_), .Y(new_n20829_));
  MX2X1    g18393(.A(new_n20829_), .B(new_n20826_), .S0(new_n11884_), .Y(new_n20830_));
  MX2X1    g18394(.A(new_n20830_), .B(new_n20807_), .S0(pi0647), .Y(new_n20831_));
  MX2X1    g18395(.A(new_n20830_), .B(new_n20807_), .S0(new_n12705_), .Y(new_n20832_));
  MX2X1    g18396(.A(new_n20832_), .B(new_n20831_), .S0(new_n12706_), .Y(new_n20833_));
  MX2X1    g18397(.A(new_n20833_), .B(new_n20830_), .S0(new_n11883_), .Y(new_n20834_));
  OAI21X1  g18398(.A0(new_n20834_), .A1(pi0644), .B0(pi0715), .Y(new_n20835_));
  OAI22X1  g18399(.A0(new_n12904_), .A1(new_n6844_), .B0(new_n12089_), .B1(pi0746), .Y(new_n20836_));
  NAND2X1  g18400(.A(new_n20836_), .B(pi0039), .Y(new_n20837_));
  AND2X1   g18401(.A(pi0746), .B(new_n6844_), .Y(new_n20838_));
  AOI21X1  g18402(.A0(new_n13683_), .A1(new_n2959_), .B0(new_n15545_), .Y(new_n20839_));
  OAI21X1  g18403(.A0(new_n20839_), .A1(new_n6844_), .B0(new_n15549_), .Y(new_n20840_));
  AOI21X1  g18404(.A0(new_n20838_), .A1(new_n12162_), .B0(new_n20840_), .Y(new_n20841_));
  AOI21X1  g18405(.A0(new_n20841_), .A1(new_n20837_), .B0(pi0038), .Y(new_n20842_));
  OAI21X1  g18406(.A0(new_n12202_), .A1(pi0191), .B0(pi0038), .Y(new_n20843_));
  AOI21X1  g18407(.A0(new_n12205_), .A1(pi0746), .B0(new_n20843_), .Y(new_n20844_));
  NOR2X1   g18408(.A(new_n20844_), .B(new_n20842_), .Y(new_n20845_));
  MX2X1    g18409(.A(new_n20845_), .B(new_n6844_), .S0(new_n3810_), .Y(new_n20846_));
  MX2X1    g18410(.A(new_n20846_), .B(new_n20806_), .S0(new_n12601_), .Y(new_n20847_));
  NOR2X1   g18411(.A(new_n20846_), .B(new_n12601_), .Y(new_n20848_));
  AOI22X1  g18412(.A0(new_n20848_), .A1(pi0609), .B0(new_n20807_), .B1(new_n13430_), .Y(new_n20849_));
  AOI22X1  g18413(.A0(new_n20848_), .A1(new_n12590_), .B0(new_n20807_), .B1(new_n13436_), .Y(new_n20850_));
  MX2X1    g18414(.A(new_n20850_), .B(new_n20849_), .S0(pi1155), .Y(new_n20851_));
  MX2X1    g18415(.A(new_n20851_), .B(new_n20847_), .S0(new_n11888_), .Y(new_n20852_));
  OAI21X1  g18416(.A0(new_n20807_), .A1(pi0618), .B0(pi1154), .Y(new_n20853_));
  AOI21X1  g18417(.A0(new_n20852_), .A1(pi0618), .B0(new_n20853_), .Y(new_n20854_));
  OAI21X1  g18418(.A0(new_n20807_), .A1(new_n12614_), .B0(new_n12615_), .Y(new_n20855_));
  AOI21X1  g18419(.A0(new_n20852_), .A1(new_n12614_), .B0(new_n20855_), .Y(new_n20856_));
  NOR2X1   g18420(.A(new_n20856_), .B(new_n20854_), .Y(new_n20857_));
  MX2X1    g18421(.A(new_n20857_), .B(new_n20852_), .S0(new_n11887_), .Y(new_n20858_));
  OAI21X1  g18422(.A0(new_n20807_), .A1(pi0619), .B0(pi1159), .Y(new_n20859_));
  AOI21X1  g18423(.A0(new_n20858_), .A1(pi0619), .B0(new_n20859_), .Y(new_n20860_));
  OAI21X1  g18424(.A0(new_n20807_), .A1(new_n12637_), .B0(new_n12638_), .Y(new_n20861_));
  AOI21X1  g18425(.A0(new_n20858_), .A1(new_n12637_), .B0(new_n20861_), .Y(new_n20862_));
  NOR2X1   g18426(.A(new_n20862_), .B(new_n20860_), .Y(new_n20863_));
  MX2X1    g18427(.A(new_n20863_), .B(new_n20858_), .S0(new_n11886_), .Y(new_n20864_));
  MX2X1    g18428(.A(new_n20864_), .B(new_n20806_), .S0(new_n12841_), .Y(new_n20865_));
  MX2X1    g18429(.A(new_n20865_), .B(new_n20806_), .S0(new_n12711_), .Y(new_n20866_));
  MX2X1    g18430(.A(new_n20866_), .B(new_n20806_), .S0(new_n12735_), .Y(new_n20867_));
  OAI21X1  g18431(.A0(new_n20807_), .A1(pi0644), .B0(new_n12739_), .Y(new_n20868_));
  AOI21X1  g18432(.A0(new_n20867_), .A1(pi0644), .B0(new_n20868_), .Y(new_n20869_));
  NOR2X1   g18433(.A(new_n20869_), .B(new_n11882_), .Y(new_n20870_));
  OAI21X1  g18434(.A0(new_n20834_), .A1(new_n12743_), .B0(new_n12739_), .Y(new_n20871_));
  OAI21X1  g18435(.A0(new_n20807_), .A1(new_n12743_), .B0(pi0715), .Y(new_n20872_));
  AOI21X1  g18436(.A0(new_n20867_), .A1(new_n12743_), .B0(new_n20872_), .Y(new_n20873_));
  NOR2X1   g18437(.A(new_n20873_), .B(pi1160), .Y(new_n20874_));
  AOI22X1  g18438(.A0(new_n20874_), .A1(new_n20871_), .B0(new_n20870_), .B1(new_n20835_), .Y(new_n20875_));
  NOR3X1   g18439(.A(new_n20873_), .B(pi1160), .C(pi0644), .Y(new_n20876_));
  NOR3X1   g18440(.A(new_n20869_), .B(new_n11882_), .C(new_n12743_), .Y(new_n20877_));
  NOR3X1   g18441(.A(new_n20877_), .B(new_n20876_), .C(new_n12897_), .Y(new_n20878_));
  AOI22X1  g18442(.A0(new_n20828_), .A1(new_n12707_), .B0(new_n20827_), .B1(new_n12709_), .Y(new_n20879_));
  OAI21X1  g18443(.A0(new_n20865_), .A1(new_n14395_), .B0(new_n20879_), .Y(new_n20880_));
  NOR3X1   g18444(.A(new_n20844_), .B(new_n20842_), .C(pi0729), .Y(new_n20881_));
  INVX1    g18445(.A(new_n20881_), .Y(new_n20882_));
  AOI21X1  g18446(.A0(new_n13989_), .A1(pi0191), .B0(pi0746), .Y(new_n20883_));
  OAI21X1  g18447(.A0(new_n13986_), .A1(pi0191), .B0(new_n20883_), .Y(new_n20884_));
  OAI21X1  g18448(.A0(new_n12440_), .A1(pi0191), .B0(pi0746), .Y(new_n20885_));
  AOI21X1  g18449(.A0(new_n12401_), .A1(pi0191), .B0(new_n20885_), .Y(new_n20886_));
  NOR2X1   g18450(.A(new_n20886_), .B(new_n2959_), .Y(new_n20887_));
  AND2X1   g18451(.A(new_n20887_), .B(new_n20884_), .Y(new_n20888_));
  AOI21X1  g18452(.A0(new_n13995_), .A1(pi0191), .B0(pi0746), .Y(new_n20889_));
  OAI21X1  g18453(.A0(new_n13996_), .A1(pi0191), .B0(new_n20889_), .Y(new_n20890_));
  AOI21X1  g18454(.A0(new_n12453_), .A1(new_n12104_), .B0(pi0191), .Y(new_n20891_));
  INVX1    g18455(.A(new_n20891_), .Y(new_n20892_));
  AOI21X1  g18456(.A0(new_n12929_), .A1(pi0191), .B0(new_n15545_), .Y(new_n20893_));
  AOI21X1  g18457(.A0(new_n20893_), .A1(new_n20892_), .B0(pi0039), .Y(new_n20894_));
  AOI21X1  g18458(.A0(new_n20894_), .A1(new_n20890_), .B0(pi0038), .Y(new_n20895_));
  INVX1    g18459(.A(new_n20895_), .Y(new_n20896_));
  AOI21X1  g18460(.A0(new_n16526_), .A1(new_n15545_), .B0(new_n12478_), .Y(new_n20897_));
  OAI21X1  g18461(.A0(new_n20897_), .A1(pi0039), .B0(new_n6844_), .Y(new_n20898_));
  OAI21X1  g18462(.A0(new_n20689_), .A1(new_n13576_), .B0(pi0191), .Y(new_n20899_));
  OAI21X1  g18463(.A0(new_n20899_), .A1(new_n14411_), .B0(pi0038), .Y(new_n20900_));
  INVX1    g18464(.A(new_n20900_), .Y(new_n20901_));
  AOI21X1  g18465(.A0(new_n20901_), .A1(new_n20898_), .B0(new_n15585_), .Y(new_n20902_));
  OAI21X1  g18466(.A0(new_n20896_), .A1(new_n20888_), .B0(new_n20902_), .Y(new_n20903_));
  AND2X1   g18467(.A(new_n20903_), .B(new_n3129_), .Y(new_n20904_));
  AOI22X1  g18468(.A0(new_n20904_), .A1(new_n20882_), .B0(new_n3810_), .B1(pi0191), .Y(new_n20905_));
  INVX1    g18469(.A(new_n20905_), .Y(new_n20906_));
  AOI21X1  g18470(.A0(new_n20846_), .A1(pi0625), .B0(pi1153), .Y(new_n20907_));
  OAI21X1  g18471(.A0(new_n20906_), .A1(pi0625), .B0(new_n20907_), .Y(new_n20908_));
  AND2X1   g18472(.A(new_n20817_), .B(new_n12584_), .Y(new_n20909_));
  AOI21X1  g18473(.A0(new_n20846_), .A1(new_n12493_), .B0(new_n12494_), .Y(new_n20910_));
  OAI21X1  g18474(.A0(new_n20906_), .A1(new_n12493_), .B0(new_n20910_), .Y(new_n20911_));
  AND2X1   g18475(.A(new_n20819_), .B(pi0608), .Y(new_n20912_));
  AOI22X1  g18476(.A0(new_n20912_), .A1(new_n20911_), .B0(new_n20909_), .B1(new_n20908_), .Y(new_n20913_));
  MX2X1    g18477(.A(new_n20913_), .B(new_n20906_), .S0(new_n11889_), .Y(new_n20914_));
  AOI21X1  g18478(.A0(new_n20821_), .A1(pi0609), .B0(pi1155), .Y(new_n20915_));
  OAI21X1  g18479(.A0(new_n20914_), .A1(pi0609), .B0(new_n20915_), .Y(new_n20916_));
  OAI21X1  g18480(.A0(new_n20849_), .A1(new_n12591_), .B0(new_n12596_), .Y(new_n20917_));
  INVX1    g18481(.A(new_n20917_), .Y(new_n20918_));
  AOI21X1  g18482(.A0(new_n20821_), .A1(new_n12590_), .B0(new_n12591_), .Y(new_n20919_));
  OAI21X1  g18483(.A0(new_n20914_), .A1(new_n12590_), .B0(new_n20919_), .Y(new_n20920_));
  OAI21X1  g18484(.A0(new_n20850_), .A1(pi1155), .B0(pi0660), .Y(new_n20921_));
  INVX1    g18485(.A(new_n20921_), .Y(new_n20922_));
  AOI22X1  g18486(.A0(new_n20922_), .A1(new_n20920_), .B0(new_n20918_), .B1(new_n20916_), .Y(new_n20923_));
  MX2X1    g18487(.A(new_n20923_), .B(new_n20914_), .S0(new_n11888_), .Y(new_n20924_));
  AOI21X1  g18488(.A0(new_n20822_), .A1(pi0618), .B0(pi1154), .Y(new_n20925_));
  OAI21X1  g18489(.A0(new_n20924_), .A1(pi0618), .B0(new_n20925_), .Y(new_n20926_));
  NOR2X1   g18490(.A(new_n20854_), .B(pi0627), .Y(new_n20927_));
  AOI21X1  g18491(.A0(new_n20822_), .A1(new_n12614_), .B0(new_n12615_), .Y(new_n20928_));
  OAI21X1  g18492(.A0(new_n20924_), .A1(new_n12614_), .B0(new_n20928_), .Y(new_n20929_));
  NOR2X1   g18493(.A(new_n20856_), .B(new_n12622_), .Y(new_n20930_));
  AOI22X1  g18494(.A0(new_n20930_), .A1(new_n20929_), .B0(new_n20927_), .B1(new_n20926_), .Y(new_n20931_));
  MX2X1    g18495(.A(new_n20931_), .B(new_n20924_), .S0(new_n11887_), .Y(new_n20932_));
  INVX1    g18496(.A(new_n20932_), .Y(new_n20933_));
  OAI21X1  g18497(.A0(new_n20824_), .A1(new_n12637_), .B0(new_n12638_), .Y(new_n20934_));
  AOI21X1  g18498(.A0(new_n20933_), .A1(new_n12637_), .B0(new_n20934_), .Y(new_n20935_));
  NOR3X1   g18499(.A(new_n20935_), .B(new_n20860_), .C(pi0648), .Y(new_n20936_));
  OAI21X1  g18500(.A0(new_n20824_), .A1(pi0619), .B0(pi1159), .Y(new_n20937_));
  AOI21X1  g18501(.A0(new_n20933_), .A1(pi0619), .B0(new_n20937_), .Y(new_n20938_));
  OR2X1    g18502(.A(new_n20862_), .B(new_n12645_), .Y(new_n20939_));
  OAI21X1  g18503(.A0(new_n20939_), .A1(new_n20938_), .B0(pi0789), .Y(new_n20940_));
  AOI21X1  g18504(.A0(new_n20932_), .A1(new_n11886_), .B0(new_n14264_), .Y(new_n20941_));
  OAI21X1  g18505(.A0(new_n20940_), .A1(new_n20936_), .B0(new_n20941_), .Y(new_n20942_));
  AOI21X1  g18506(.A0(new_n20807_), .A1(pi0626), .B0(new_n16352_), .Y(new_n20943_));
  OAI21X1  g18507(.A0(new_n20864_), .A1(pi0626), .B0(new_n20943_), .Y(new_n20944_));
  AOI21X1  g18508(.A0(new_n20807_), .A1(new_n12664_), .B0(new_n16356_), .Y(new_n20945_));
  OAI21X1  g18509(.A0(new_n20864_), .A1(new_n12664_), .B0(new_n20945_), .Y(new_n20946_));
  OR2X1    g18510(.A(new_n20825_), .B(new_n12770_), .Y(new_n20947_));
  NAND3X1  g18511(.A(new_n20947_), .B(new_n20946_), .C(new_n20944_), .Y(new_n20948_));
  AOI21X1  g18512(.A0(new_n20948_), .A1(pi0788), .B0(new_n14273_), .Y(new_n20949_));
  AOI22X1  g18513(.A0(new_n20949_), .A1(new_n20942_), .B0(new_n20880_), .B1(pi0792), .Y(new_n20950_));
  NOR2X1   g18514(.A(new_n20866_), .B(new_n14384_), .Y(new_n20951_));
  AND2X1   g18515(.A(new_n20832_), .B(new_n14386_), .Y(new_n20952_));
  AND2X1   g18516(.A(new_n20831_), .B(new_n14388_), .Y(new_n20953_));
  OR2X1    g18517(.A(new_n20953_), .B(new_n20952_), .Y(new_n20954_));
  OAI21X1  g18518(.A0(new_n20954_), .A1(new_n20951_), .B0(pi0787), .Y(new_n20955_));
  OAI21X1  g18519(.A0(new_n20950_), .A1(new_n14269_), .B0(new_n20955_), .Y(new_n20956_));
  OAI22X1  g18520(.A0(new_n20956_), .A1(new_n20878_), .B0(new_n20875_), .B1(new_n12897_), .Y(new_n20957_));
  OAI21X1  g18521(.A0(new_n6520_), .A1(pi0191), .B0(new_n12898_), .Y(new_n20958_));
  AOI21X1  g18522(.A0(new_n20957_), .A1(new_n6520_), .B0(new_n20958_), .Y(new_n20959_));
  AOI21X1  g18523(.A0(new_n20805_), .A1(new_n20804_), .B0(new_n20959_), .Y(po0348));
  AOI21X1  g18524(.A0(pi1093), .A1(pi1092), .B0(pi0192), .Y(new_n20961_));
  INVX1    g18525(.A(new_n20961_), .Y(new_n20962_));
  AOI21X1  g18526(.A0(new_n12178_), .A1(pi0764), .B0(new_n20961_), .Y(new_n20963_));
  AOI21X1  g18527(.A0(new_n12601_), .A1(new_n2739_), .B0(new_n20963_), .Y(new_n20964_));
  AND2X1   g18528(.A(new_n12178_), .B(pi0764), .Y(new_n20965_));
  AND2X1   g18529(.A(new_n20965_), .B(new_n12608_), .Y(new_n20966_));
  INVX1    g18530(.A(new_n20966_), .Y(new_n20967_));
  AOI21X1  g18531(.A0(new_n20967_), .A1(new_n20964_), .B0(new_n12591_), .Y(new_n20968_));
  NOR3X1   g18532(.A(new_n20966_), .B(new_n20961_), .C(pi1155), .Y(new_n20969_));
  OAI21X1  g18533(.A0(new_n20969_), .A1(new_n20968_), .B0(pi0785), .Y(new_n20970_));
  OAI21X1  g18534(.A0(new_n20964_), .A1(pi0785), .B0(new_n20970_), .Y(new_n20971_));
  INVX1    g18535(.A(new_n20971_), .Y(new_n20972_));
  AOI21X1  g18536(.A0(new_n20972_), .A1(new_n12785_), .B0(new_n12615_), .Y(new_n20973_));
  AOI21X1  g18537(.A0(new_n20972_), .A1(new_n12788_), .B0(pi1154), .Y(new_n20974_));
  NOR2X1   g18538(.A(new_n20974_), .B(new_n20973_), .Y(new_n20975_));
  MX2X1    g18539(.A(new_n20975_), .B(new_n20972_), .S0(new_n11887_), .Y(new_n20976_));
  OR2X1    g18540(.A(new_n20976_), .B(pi0789), .Y(new_n20977_));
  AOI21X1  g18541(.A0(new_n20976_), .A1(new_n15910_), .B0(new_n12638_), .Y(new_n20978_));
  AOI21X1  g18542(.A0(new_n20976_), .A1(new_n15912_), .B0(pi1159), .Y(new_n20979_));
  OAI21X1  g18543(.A0(new_n20979_), .A1(new_n20978_), .B0(pi0789), .Y(new_n20980_));
  AND2X1   g18544(.A(new_n20980_), .B(new_n20977_), .Y(new_n20981_));
  INVX1    g18545(.A(new_n20981_), .Y(new_n20982_));
  MX2X1    g18546(.A(new_n20982_), .B(new_n20962_), .S0(new_n12841_), .Y(new_n20983_));
  MX2X1    g18547(.A(new_n20983_), .B(new_n20962_), .S0(new_n12711_), .Y(new_n20984_));
  AOI21X1  g18548(.A0(new_n12566_), .A1(pi0691), .B0(new_n20961_), .Y(new_n20985_));
  INVX1    g18549(.A(new_n20985_), .Y(new_n20986_));
  NOR3X1   g18550(.A(new_n13585_), .B(new_n15681_), .C(pi0625), .Y(new_n20987_));
  OR2X1    g18551(.A(new_n20987_), .B(new_n20985_), .Y(new_n20988_));
  NOR2X1   g18552(.A(new_n20961_), .B(pi1153), .Y(new_n20989_));
  INVX1    g18553(.A(new_n20989_), .Y(new_n20990_));
  OAI21X1  g18554(.A0(new_n20990_), .A1(new_n20987_), .B0(pi0778), .Y(new_n20991_));
  AOI21X1  g18555(.A0(new_n20988_), .A1(pi1153), .B0(new_n20991_), .Y(new_n20992_));
  AOI21X1  g18556(.A0(new_n20986_), .A1(new_n11889_), .B0(new_n20992_), .Y(new_n20993_));
  NOR4X1   g18557(.A(new_n20993_), .B(new_n12765_), .C(new_n12764_), .D(new_n12762_), .Y(new_n20994_));
  INVX1    g18558(.A(new_n20994_), .Y(new_n20995_));
  NOR3X1   g18559(.A(new_n20995_), .B(new_n12870_), .C(new_n12851_), .Y(new_n20996_));
  INVX1    g18560(.A(new_n20996_), .Y(new_n20997_));
  AOI21X1  g18561(.A0(new_n20961_), .A1(pi0647), .B0(pi1157), .Y(new_n20998_));
  OAI21X1  g18562(.A0(new_n20997_), .A1(pi0647), .B0(new_n20998_), .Y(new_n20999_));
  MX2X1    g18563(.A(new_n20996_), .B(new_n20961_), .S0(new_n12705_), .Y(new_n21000_));
  OAI22X1  g18564(.A0(new_n21000_), .A1(new_n14387_), .B0(new_n20999_), .B1(new_n12723_), .Y(new_n21001_));
  AOI21X1  g18565(.A0(new_n20984_), .A1(new_n14385_), .B0(new_n21001_), .Y(new_n21002_));
  NOR2X1   g18566(.A(new_n21002_), .B(new_n11883_), .Y(new_n21003_));
  AOI21X1  g18567(.A0(new_n20962_), .A1(pi0626), .B0(new_n16352_), .Y(new_n21004_));
  OAI21X1  g18568(.A0(new_n20981_), .A1(pi0626), .B0(new_n21004_), .Y(new_n21005_));
  AOI21X1  g18569(.A0(new_n20980_), .A1(new_n20977_), .B0(new_n12664_), .Y(new_n21006_));
  NOR2X1   g18570(.A(new_n20961_), .B(pi0626), .Y(new_n21007_));
  NOR3X1   g18571(.A(new_n21007_), .B(new_n21006_), .C(new_n16356_), .Y(new_n21008_));
  AOI21X1  g18572(.A0(new_n20994_), .A1(new_n12769_), .B0(new_n21008_), .Y(new_n21009_));
  AOI21X1  g18573(.A0(new_n21009_), .A1(new_n21005_), .B0(new_n11885_), .Y(new_n21010_));
  INVX1    g18574(.A(new_n20963_), .Y(new_n21011_));
  AOI21X1  g18575(.A0(new_n20986_), .A1(new_n12171_), .B0(new_n21011_), .Y(new_n21012_));
  NOR3X1   g18576(.A(new_n20985_), .B(new_n12120_), .C(new_n12493_), .Y(new_n21013_));
  OR2X1    g18577(.A(new_n21012_), .B(new_n21013_), .Y(new_n21014_));
  NOR2X1   g18578(.A(new_n20987_), .B(new_n20985_), .Y(new_n21015_));
  OAI21X1  g18579(.A0(new_n21015_), .A1(new_n12494_), .B0(new_n12584_), .Y(new_n21016_));
  AOI21X1  g18580(.A0(new_n21014_), .A1(new_n20989_), .B0(new_n21016_), .Y(new_n21017_));
  NOR3X1   g18581(.A(new_n21013_), .B(new_n21011_), .C(new_n12494_), .Y(new_n21018_));
  OAI21X1  g18582(.A0(new_n20990_), .A1(new_n20987_), .B0(pi0608), .Y(new_n21019_));
  NOR2X1   g18583(.A(new_n21019_), .B(new_n21018_), .Y(new_n21020_));
  OAI21X1  g18584(.A0(new_n21020_), .A1(new_n21017_), .B0(pi0778), .Y(new_n21021_));
  OAI21X1  g18585(.A0(new_n21012_), .A1(pi0778), .B0(new_n21021_), .Y(new_n21022_));
  OAI21X1  g18586(.A0(new_n20993_), .A1(new_n12590_), .B0(new_n12591_), .Y(new_n21023_));
  AOI21X1  g18587(.A0(new_n21022_), .A1(new_n12590_), .B0(new_n21023_), .Y(new_n21024_));
  NOR3X1   g18588(.A(new_n21024_), .B(new_n20968_), .C(pi0660), .Y(new_n21025_));
  OAI21X1  g18589(.A0(new_n20993_), .A1(pi0609), .B0(pi1155), .Y(new_n21026_));
  AOI21X1  g18590(.A0(new_n21022_), .A1(pi0609), .B0(new_n21026_), .Y(new_n21027_));
  NOR3X1   g18591(.A(new_n21027_), .B(new_n20969_), .C(new_n12596_), .Y(new_n21028_));
  OAI21X1  g18592(.A0(new_n21028_), .A1(new_n21025_), .B0(pi0785), .Y(new_n21029_));
  NAND2X1  g18593(.A(new_n21022_), .B(new_n11888_), .Y(new_n21030_));
  AND2X1   g18594(.A(new_n21030_), .B(new_n21029_), .Y(new_n21031_));
  NOR3X1   g18595(.A(new_n20993_), .B(new_n12762_), .C(new_n12614_), .Y(new_n21032_));
  NOR2X1   g18596(.A(new_n21032_), .B(pi1154), .Y(new_n21033_));
  OAI21X1  g18597(.A0(new_n21031_), .A1(pi0618), .B0(new_n21033_), .Y(new_n21034_));
  NOR2X1   g18598(.A(new_n20973_), .B(pi0627), .Y(new_n21035_));
  NOR3X1   g18599(.A(new_n20993_), .B(new_n12762_), .C(pi0618), .Y(new_n21036_));
  NOR2X1   g18600(.A(new_n21036_), .B(new_n12615_), .Y(new_n21037_));
  OAI21X1  g18601(.A0(new_n21031_), .A1(new_n12614_), .B0(new_n21037_), .Y(new_n21038_));
  NOR2X1   g18602(.A(new_n20974_), .B(new_n12622_), .Y(new_n21039_));
  AOI22X1  g18603(.A0(new_n21039_), .A1(new_n21038_), .B0(new_n21035_), .B1(new_n21034_), .Y(new_n21040_));
  MX2X1    g18604(.A(new_n21040_), .B(new_n21031_), .S0(new_n11887_), .Y(new_n21041_));
  OR4X1    g18605(.A(new_n20993_), .B(new_n12764_), .C(new_n12762_), .D(new_n12637_), .Y(new_n21042_));
  AND2X1   g18606(.A(new_n21042_), .B(new_n12638_), .Y(new_n21043_));
  OAI21X1  g18607(.A0(new_n21041_), .A1(pi0619), .B0(new_n21043_), .Y(new_n21044_));
  NOR2X1   g18608(.A(new_n20978_), .B(pi0648), .Y(new_n21045_));
  AND2X1   g18609(.A(new_n21045_), .B(new_n21044_), .Y(new_n21046_));
  INVX1    g18610(.A(new_n21046_), .Y(new_n21047_));
  NOR4X1   g18611(.A(new_n20993_), .B(new_n12764_), .C(new_n12762_), .D(pi0619), .Y(new_n21048_));
  NOR2X1   g18612(.A(new_n21048_), .B(new_n12638_), .Y(new_n21049_));
  OAI21X1  g18613(.A0(new_n21041_), .A1(new_n12637_), .B0(new_n21049_), .Y(new_n21050_));
  NOR2X1   g18614(.A(new_n20979_), .B(new_n12645_), .Y(new_n21051_));
  AOI21X1  g18615(.A0(new_n21051_), .A1(new_n21050_), .B0(new_n11886_), .Y(new_n21052_));
  AOI21X1  g18616(.A0(new_n21041_), .A1(new_n11886_), .B0(new_n14264_), .Y(new_n21053_));
  INVX1    g18617(.A(new_n21053_), .Y(new_n21054_));
  AOI21X1  g18618(.A0(new_n21052_), .A1(new_n21047_), .B0(new_n21054_), .Y(new_n21055_));
  OAI21X1  g18619(.A0(new_n21055_), .A1(new_n21010_), .B0(new_n16350_), .Y(new_n21056_));
  INVX1    g18620(.A(new_n20983_), .Y(new_n21057_));
  AND2X1   g18621(.A(new_n20994_), .B(new_n12852_), .Y(new_n21058_));
  AOI22X1  g18622(.A0(new_n21058_), .A1(new_n14564_), .B0(new_n21057_), .B1(new_n12867_), .Y(new_n21059_));
  AOI22X1  g18623(.A0(new_n21058_), .A1(new_n14566_), .B0(new_n21057_), .B1(new_n12865_), .Y(new_n21060_));
  MX2X1    g18624(.A(new_n21060_), .B(new_n21059_), .S0(new_n12689_), .Y(new_n21061_));
  OAI21X1  g18625(.A0(new_n21061_), .A1(new_n11884_), .B0(new_n14562_), .Y(new_n21062_));
  INVX1    g18626(.A(new_n21062_), .Y(new_n21063_));
  AOI21X1  g18627(.A0(new_n21063_), .A1(new_n21056_), .B0(new_n21003_), .Y(new_n21064_));
  OAI21X1  g18628(.A0(new_n21000_), .A1(new_n12706_), .B0(new_n20999_), .Y(new_n21065_));
  MX2X1    g18629(.A(new_n21065_), .B(new_n20997_), .S0(new_n11883_), .Y(new_n21066_));
  OAI21X1  g18630(.A0(new_n21066_), .A1(pi0644), .B0(pi0715), .Y(new_n21067_));
  AOI21X1  g18631(.A0(new_n21064_), .A1(pi0644), .B0(new_n21067_), .Y(new_n21068_));
  OR4X1    g18632(.A(new_n12734_), .B(new_n2739_), .C(new_n11883_), .D(pi0192), .Y(new_n21069_));
  OAI21X1  g18633(.A0(new_n20984_), .A1(new_n12735_), .B0(new_n21069_), .Y(new_n21070_));
  OAI21X1  g18634(.A0(new_n20962_), .A1(pi0644), .B0(new_n12739_), .Y(new_n21071_));
  AOI21X1  g18635(.A0(new_n21070_), .A1(pi0644), .B0(new_n21071_), .Y(new_n21072_));
  OR2X1    g18636(.A(new_n21072_), .B(new_n11882_), .Y(new_n21073_));
  OAI21X1  g18637(.A0(new_n21066_), .A1(new_n12743_), .B0(new_n12739_), .Y(new_n21074_));
  AOI21X1  g18638(.A0(new_n21064_), .A1(new_n12743_), .B0(new_n21074_), .Y(new_n21075_));
  OAI21X1  g18639(.A0(new_n20962_), .A1(new_n12743_), .B0(pi0715), .Y(new_n21076_));
  AOI21X1  g18640(.A0(new_n21070_), .A1(new_n12743_), .B0(new_n21076_), .Y(new_n21077_));
  OR2X1    g18641(.A(new_n21077_), .B(pi1160), .Y(new_n21078_));
  OAI22X1  g18642(.A0(new_n21078_), .A1(new_n21075_), .B0(new_n21073_), .B1(new_n21068_), .Y(new_n21079_));
  NAND2X1  g18643(.A(new_n21079_), .B(pi0790), .Y(new_n21080_));
  AOI21X1  g18644(.A0(new_n21064_), .A1(new_n12897_), .B0(new_n12898_), .Y(new_n21081_));
  AOI21X1  g18645(.A0(new_n13699_), .A1(new_n3129_), .B0(pi0192), .Y(new_n21082_));
  INVX1    g18646(.A(new_n21082_), .Y(new_n21083_));
  OAI21X1  g18647(.A0(new_n16436_), .A1(new_n11594_), .B0(new_n2996_), .Y(new_n21084_));
  AOI21X1  g18648(.A0(new_n16435_), .A1(new_n11594_), .B0(new_n21084_), .Y(new_n21085_));
  AOI21X1  g18649(.A0(new_n12901_), .A1(new_n11594_), .B0(new_n12568_), .Y(new_n21086_));
  NOR3X1   g18650(.A(new_n21086_), .B(new_n21085_), .C(new_n15681_), .Y(new_n21087_));
  OR2X1    g18651(.A(pi0691), .B(pi0192), .Y(new_n21088_));
  OAI21X1  g18652(.A0(new_n21088_), .A1(new_n13699_), .B0(new_n3129_), .Y(new_n21089_));
  OAI22X1  g18653(.A0(new_n21089_), .A1(new_n21087_), .B0(new_n3129_), .B1(new_n11594_), .Y(new_n21090_));
  AND2X1   g18654(.A(new_n21090_), .B(new_n11889_), .Y(new_n21091_));
  AOI21X1  g18655(.A0(new_n21082_), .A1(new_n12493_), .B0(new_n12494_), .Y(new_n21092_));
  OAI21X1  g18656(.A0(new_n21090_), .A1(new_n12493_), .B0(new_n21092_), .Y(new_n21093_));
  AOI21X1  g18657(.A0(new_n21082_), .A1(pi0625), .B0(pi1153), .Y(new_n21094_));
  OAI21X1  g18658(.A0(new_n21090_), .A1(pi0625), .B0(new_n21094_), .Y(new_n21095_));
  AOI21X1  g18659(.A0(new_n21095_), .A1(new_n21093_), .B0(new_n11889_), .Y(new_n21096_));
  NOR2X1   g18660(.A(new_n21096_), .B(new_n21091_), .Y(new_n21097_));
  MX2X1    g18661(.A(new_n21097_), .B(new_n21082_), .S0(new_n12618_), .Y(new_n21098_));
  AND2X1   g18662(.A(new_n21082_), .B(new_n12641_), .Y(new_n21099_));
  AOI21X1  g18663(.A0(new_n21098_), .A1(new_n14198_), .B0(new_n21099_), .Y(new_n21100_));
  MX2X1    g18664(.A(new_n21100_), .B(new_n21083_), .S0(new_n12659_), .Y(new_n21101_));
  MX2X1    g18665(.A(new_n21101_), .B(new_n21083_), .S0(new_n12691_), .Y(new_n21102_));
  MX2X1    g18666(.A(new_n21102_), .B(new_n21083_), .S0(pi0628), .Y(new_n21103_));
  MX2X1    g18667(.A(new_n21102_), .B(new_n21083_), .S0(new_n12683_), .Y(new_n21104_));
  MX2X1    g18668(.A(new_n21104_), .B(new_n21103_), .S0(new_n12684_), .Y(new_n21105_));
  MX2X1    g18669(.A(new_n21105_), .B(new_n21102_), .S0(new_n11884_), .Y(new_n21106_));
  MX2X1    g18670(.A(new_n21106_), .B(new_n21083_), .S0(pi0647), .Y(new_n21107_));
  MX2X1    g18671(.A(new_n21106_), .B(new_n21083_), .S0(new_n12705_), .Y(new_n21108_));
  MX2X1    g18672(.A(new_n21108_), .B(new_n21107_), .S0(new_n12706_), .Y(new_n21109_));
  MX2X1    g18673(.A(new_n21109_), .B(new_n21106_), .S0(new_n11883_), .Y(new_n21110_));
  OAI21X1  g18674(.A0(new_n21110_), .A1(pi0644), .B0(pi0715), .Y(new_n21111_));
  OAI22X1  g18675(.A0(new_n12904_), .A1(new_n11594_), .B0(new_n12089_), .B1(pi0764), .Y(new_n21112_));
  NAND2X1  g18676(.A(new_n21112_), .B(pi0039), .Y(new_n21113_));
  AND2X1   g18677(.A(pi0764), .B(new_n11594_), .Y(new_n21114_));
  AOI21X1  g18678(.A0(new_n13683_), .A1(new_n2959_), .B0(new_n15641_), .Y(new_n21115_));
  OAI21X1  g18679(.A0(new_n21115_), .A1(new_n11594_), .B0(new_n15645_), .Y(new_n21116_));
  AOI21X1  g18680(.A0(new_n21114_), .A1(new_n12162_), .B0(new_n21116_), .Y(new_n21117_));
  AOI21X1  g18681(.A0(new_n21117_), .A1(new_n21113_), .B0(pi0038), .Y(new_n21118_));
  OAI21X1  g18682(.A0(new_n12202_), .A1(pi0192), .B0(pi0038), .Y(new_n21119_));
  AOI21X1  g18683(.A0(new_n12205_), .A1(pi0764), .B0(new_n21119_), .Y(new_n21120_));
  NOR2X1   g18684(.A(new_n21120_), .B(new_n21118_), .Y(new_n21121_));
  MX2X1    g18685(.A(new_n21121_), .B(new_n11594_), .S0(new_n3810_), .Y(new_n21122_));
  MX2X1    g18686(.A(new_n21122_), .B(new_n21082_), .S0(new_n12601_), .Y(new_n21123_));
  NOR2X1   g18687(.A(new_n21122_), .B(new_n12601_), .Y(new_n21124_));
  AOI22X1  g18688(.A0(new_n21124_), .A1(pi0609), .B0(new_n21083_), .B1(new_n13430_), .Y(new_n21125_));
  AOI22X1  g18689(.A0(new_n21124_), .A1(new_n12590_), .B0(new_n21083_), .B1(new_n13436_), .Y(new_n21126_));
  MX2X1    g18690(.A(new_n21126_), .B(new_n21125_), .S0(pi1155), .Y(new_n21127_));
  MX2X1    g18691(.A(new_n21127_), .B(new_n21123_), .S0(new_n11888_), .Y(new_n21128_));
  OAI21X1  g18692(.A0(new_n21083_), .A1(pi0618), .B0(pi1154), .Y(new_n21129_));
  AOI21X1  g18693(.A0(new_n21128_), .A1(pi0618), .B0(new_n21129_), .Y(new_n21130_));
  OAI21X1  g18694(.A0(new_n21083_), .A1(new_n12614_), .B0(new_n12615_), .Y(new_n21131_));
  AOI21X1  g18695(.A0(new_n21128_), .A1(new_n12614_), .B0(new_n21131_), .Y(new_n21132_));
  NOR2X1   g18696(.A(new_n21132_), .B(new_n21130_), .Y(new_n21133_));
  MX2X1    g18697(.A(new_n21133_), .B(new_n21128_), .S0(new_n11887_), .Y(new_n21134_));
  OAI21X1  g18698(.A0(new_n21083_), .A1(pi0619), .B0(pi1159), .Y(new_n21135_));
  AOI21X1  g18699(.A0(new_n21134_), .A1(pi0619), .B0(new_n21135_), .Y(new_n21136_));
  OAI21X1  g18700(.A0(new_n21083_), .A1(new_n12637_), .B0(new_n12638_), .Y(new_n21137_));
  AOI21X1  g18701(.A0(new_n21134_), .A1(new_n12637_), .B0(new_n21137_), .Y(new_n21138_));
  NOR2X1   g18702(.A(new_n21138_), .B(new_n21136_), .Y(new_n21139_));
  MX2X1    g18703(.A(new_n21139_), .B(new_n21134_), .S0(new_n11886_), .Y(new_n21140_));
  MX2X1    g18704(.A(new_n21140_), .B(new_n21082_), .S0(new_n12841_), .Y(new_n21141_));
  MX2X1    g18705(.A(new_n21141_), .B(new_n21082_), .S0(new_n12711_), .Y(new_n21142_));
  MX2X1    g18706(.A(new_n21142_), .B(new_n21082_), .S0(new_n12735_), .Y(new_n21143_));
  OAI21X1  g18707(.A0(new_n21083_), .A1(pi0644), .B0(new_n12739_), .Y(new_n21144_));
  AOI21X1  g18708(.A0(new_n21143_), .A1(pi0644), .B0(new_n21144_), .Y(new_n21145_));
  NOR2X1   g18709(.A(new_n21145_), .B(new_n11882_), .Y(new_n21146_));
  OAI21X1  g18710(.A0(new_n21110_), .A1(new_n12743_), .B0(new_n12739_), .Y(new_n21147_));
  OAI21X1  g18711(.A0(new_n21083_), .A1(new_n12743_), .B0(pi0715), .Y(new_n21148_));
  AOI21X1  g18712(.A0(new_n21143_), .A1(new_n12743_), .B0(new_n21148_), .Y(new_n21149_));
  NOR2X1   g18713(.A(new_n21149_), .B(pi1160), .Y(new_n21150_));
  AOI22X1  g18714(.A0(new_n21150_), .A1(new_n21147_), .B0(new_n21146_), .B1(new_n21111_), .Y(new_n21151_));
  NOR3X1   g18715(.A(new_n21149_), .B(pi1160), .C(pi0644), .Y(new_n21152_));
  NOR3X1   g18716(.A(new_n21145_), .B(new_n11882_), .C(new_n12743_), .Y(new_n21153_));
  NOR3X1   g18717(.A(new_n21153_), .B(new_n21152_), .C(new_n12897_), .Y(new_n21154_));
  AOI22X1  g18718(.A0(new_n21104_), .A1(new_n12707_), .B0(new_n21103_), .B1(new_n12709_), .Y(new_n21155_));
  OAI21X1  g18719(.A0(new_n21141_), .A1(new_n14395_), .B0(new_n21155_), .Y(new_n21156_));
  NOR3X1   g18720(.A(new_n21120_), .B(new_n21118_), .C(pi0691), .Y(new_n21157_));
  INVX1    g18721(.A(new_n21157_), .Y(new_n21158_));
  AOI21X1  g18722(.A0(new_n13989_), .A1(pi0192), .B0(pi0764), .Y(new_n21159_));
  OAI21X1  g18723(.A0(new_n13986_), .A1(pi0192), .B0(new_n21159_), .Y(new_n21160_));
  OAI21X1  g18724(.A0(new_n12440_), .A1(pi0192), .B0(pi0764), .Y(new_n21161_));
  AOI21X1  g18725(.A0(new_n12401_), .A1(pi0192), .B0(new_n21161_), .Y(new_n21162_));
  NOR2X1   g18726(.A(new_n21162_), .B(new_n2959_), .Y(new_n21163_));
  AND2X1   g18727(.A(new_n21163_), .B(new_n21160_), .Y(new_n21164_));
  AOI21X1  g18728(.A0(new_n13995_), .A1(pi0192), .B0(pi0764), .Y(new_n21165_));
  OAI21X1  g18729(.A0(new_n13996_), .A1(pi0192), .B0(new_n21165_), .Y(new_n21166_));
  AOI21X1  g18730(.A0(new_n12453_), .A1(new_n12104_), .B0(pi0192), .Y(new_n21167_));
  INVX1    g18731(.A(new_n21167_), .Y(new_n21168_));
  AOI21X1  g18732(.A0(new_n12929_), .A1(pi0192), .B0(new_n15641_), .Y(new_n21169_));
  AOI21X1  g18733(.A0(new_n21169_), .A1(new_n21168_), .B0(pi0039), .Y(new_n21170_));
  AOI21X1  g18734(.A0(new_n21170_), .A1(new_n21166_), .B0(pi0038), .Y(new_n21171_));
  INVX1    g18735(.A(new_n21171_), .Y(new_n21172_));
  AOI21X1  g18736(.A0(new_n16526_), .A1(new_n15641_), .B0(new_n12478_), .Y(new_n21173_));
  OAI21X1  g18737(.A0(new_n21173_), .A1(pi0039), .B0(new_n11594_), .Y(new_n21174_));
  OAI21X1  g18738(.A0(new_n20965_), .A1(new_n13576_), .B0(pi0192), .Y(new_n21175_));
  OAI21X1  g18739(.A0(new_n21175_), .A1(new_n14411_), .B0(pi0038), .Y(new_n21176_));
  INVX1    g18740(.A(new_n21176_), .Y(new_n21177_));
  AOI21X1  g18741(.A0(new_n21177_), .A1(new_n21174_), .B0(new_n15681_), .Y(new_n21178_));
  OAI21X1  g18742(.A0(new_n21172_), .A1(new_n21164_), .B0(new_n21178_), .Y(new_n21179_));
  AND2X1   g18743(.A(new_n21179_), .B(new_n3129_), .Y(new_n21180_));
  AOI22X1  g18744(.A0(new_n21180_), .A1(new_n21158_), .B0(new_n3810_), .B1(pi0192), .Y(new_n21181_));
  INVX1    g18745(.A(new_n21181_), .Y(new_n21182_));
  AOI21X1  g18746(.A0(new_n21122_), .A1(pi0625), .B0(pi1153), .Y(new_n21183_));
  OAI21X1  g18747(.A0(new_n21182_), .A1(pi0625), .B0(new_n21183_), .Y(new_n21184_));
  AND2X1   g18748(.A(new_n21093_), .B(new_n12584_), .Y(new_n21185_));
  AOI21X1  g18749(.A0(new_n21122_), .A1(new_n12493_), .B0(new_n12494_), .Y(new_n21186_));
  OAI21X1  g18750(.A0(new_n21182_), .A1(new_n12493_), .B0(new_n21186_), .Y(new_n21187_));
  AND2X1   g18751(.A(new_n21095_), .B(pi0608), .Y(new_n21188_));
  AOI22X1  g18752(.A0(new_n21188_), .A1(new_n21187_), .B0(new_n21185_), .B1(new_n21184_), .Y(new_n21189_));
  MX2X1    g18753(.A(new_n21189_), .B(new_n21182_), .S0(new_n11889_), .Y(new_n21190_));
  AOI21X1  g18754(.A0(new_n21097_), .A1(pi0609), .B0(pi1155), .Y(new_n21191_));
  OAI21X1  g18755(.A0(new_n21190_), .A1(pi0609), .B0(new_n21191_), .Y(new_n21192_));
  OAI21X1  g18756(.A0(new_n21125_), .A1(new_n12591_), .B0(new_n12596_), .Y(new_n21193_));
  INVX1    g18757(.A(new_n21193_), .Y(new_n21194_));
  AOI21X1  g18758(.A0(new_n21097_), .A1(new_n12590_), .B0(new_n12591_), .Y(new_n21195_));
  OAI21X1  g18759(.A0(new_n21190_), .A1(new_n12590_), .B0(new_n21195_), .Y(new_n21196_));
  OAI21X1  g18760(.A0(new_n21126_), .A1(pi1155), .B0(pi0660), .Y(new_n21197_));
  INVX1    g18761(.A(new_n21197_), .Y(new_n21198_));
  AOI22X1  g18762(.A0(new_n21198_), .A1(new_n21196_), .B0(new_n21194_), .B1(new_n21192_), .Y(new_n21199_));
  MX2X1    g18763(.A(new_n21199_), .B(new_n21190_), .S0(new_n11888_), .Y(new_n21200_));
  AOI21X1  g18764(.A0(new_n21098_), .A1(pi0618), .B0(pi1154), .Y(new_n21201_));
  OAI21X1  g18765(.A0(new_n21200_), .A1(pi0618), .B0(new_n21201_), .Y(new_n21202_));
  NOR2X1   g18766(.A(new_n21130_), .B(pi0627), .Y(new_n21203_));
  AOI21X1  g18767(.A0(new_n21098_), .A1(new_n12614_), .B0(new_n12615_), .Y(new_n21204_));
  OAI21X1  g18768(.A0(new_n21200_), .A1(new_n12614_), .B0(new_n21204_), .Y(new_n21205_));
  NOR2X1   g18769(.A(new_n21132_), .B(new_n12622_), .Y(new_n21206_));
  AOI22X1  g18770(.A0(new_n21206_), .A1(new_n21205_), .B0(new_n21203_), .B1(new_n21202_), .Y(new_n21207_));
  MX2X1    g18771(.A(new_n21207_), .B(new_n21200_), .S0(new_n11887_), .Y(new_n21208_));
  INVX1    g18772(.A(new_n21208_), .Y(new_n21209_));
  OAI21X1  g18773(.A0(new_n21100_), .A1(new_n12637_), .B0(new_n12638_), .Y(new_n21210_));
  AOI21X1  g18774(.A0(new_n21209_), .A1(new_n12637_), .B0(new_n21210_), .Y(new_n21211_));
  NOR3X1   g18775(.A(new_n21211_), .B(new_n21136_), .C(pi0648), .Y(new_n21212_));
  OAI21X1  g18776(.A0(new_n21100_), .A1(pi0619), .B0(pi1159), .Y(new_n21213_));
  AOI21X1  g18777(.A0(new_n21209_), .A1(pi0619), .B0(new_n21213_), .Y(new_n21214_));
  OR2X1    g18778(.A(new_n21138_), .B(new_n12645_), .Y(new_n21215_));
  OAI21X1  g18779(.A0(new_n21215_), .A1(new_n21214_), .B0(pi0789), .Y(new_n21216_));
  AOI21X1  g18780(.A0(new_n21208_), .A1(new_n11886_), .B0(new_n14264_), .Y(new_n21217_));
  OAI21X1  g18781(.A0(new_n21216_), .A1(new_n21212_), .B0(new_n21217_), .Y(new_n21218_));
  AOI21X1  g18782(.A0(new_n21083_), .A1(pi0626), .B0(new_n16352_), .Y(new_n21219_));
  OAI21X1  g18783(.A0(new_n21140_), .A1(pi0626), .B0(new_n21219_), .Y(new_n21220_));
  AOI21X1  g18784(.A0(new_n21083_), .A1(new_n12664_), .B0(new_n16356_), .Y(new_n21221_));
  OAI21X1  g18785(.A0(new_n21140_), .A1(new_n12664_), .B0(new_n21221_), .Y(new_n21222_));
  OR2X1    g18786(.A(new_n21101_), .B(new_n12770_), .Y(new_n21223_));
  NAND3X1  g18787(.A(new_n21223_), .B(new_n21222_), .C(new_n21220_), .Y(new_n21224_));
  AOI21X1  g18788(.A0(new_n21224_), .A1(pi0788), .B0(new_n14273_), .Y(new_n21225_));
  AOI22X1  g18789(.A0(new_n21225_), .A1(new_n21218_), .B0(new_n21156_), .B1(pi0792), .Y(new_n21226_));
  NOR2X1   g18790(.A(new_n21142_), .B(new_n14384_), .Y(new_n21227_));
  AND2X1   g18791(.A(new_n21108_), .B(new_n14386_), .Y(new_n21228_));
  AND2X1   g18792(.A(new_n21107_), .B(new_n14388_), .Y(new_n21229_));
  OR2X1    g18793(.A(new_n21229_), .B(new_n21228_), .Y(new_n21230_));
  OAI21X1  g18794(.A0(new_n21230_), .A1(new_n21227_), .B0(pi0787), .Y(new_n21231_));
  OAI21X1  g18795(.A0(new_n21226_), .A1(new_n14269_), .B0(new_n21231_), .Y(new_n21232_));
  OAI22X1  g18796(.A0(new_n21232_), .A1(new_n21154_), .B0(new_n21151_), .B1(new_n12897_), .Y(new_n21233_));
  OAI21X1  g18797(.A0(new_n6520_), .A1(pi0192), .B0(new_n12898_), .Y(new_n21234_));
  AOI21X1  g18798(.A0(new_n21233_), .A1(new_n6520_), .B0(new_n21234_), .Y(new_n21235_));
  AOI21X1  g18799(.A0(new_n21081_), .A1(new_n21080_), .B0(new_n21235_), .Y(po0349));
  AOI21X1  g18800(.A0(pi1093), .A1(pi1092), .B0(pi0193), .Y(new_n21237_));
  INVX1    g18801(.A(new_n21237_), .Y(new_n21238_));
  AOI21X1  g18802(.A0(new_n12178_), .A1(pi0739), .B0(new_n21237_), .Y(new_n21239_));
  AOI21X1  g18803(.A0(new_n12601_), .A1(new_n2739_), .B0(new_n21239_), .Y(new_n21240_));
  NAND2X1  g18804(.A(new_n12178_), .B(pi0739), .Y(new_n21241_));
  OAI21X1  g18805(.A0(new_n21241_), .A1(new_n13436_), .B0(new_n21240_), .Y(new_n21242_));
  AND2X1   g18806(.A(new_n21242_), .B(pi1155), .Y(new_n21243_));
  NOR2X1   g18807(.A(new_n21241_), .B(new_n13436_), .Y(new_n21244_));
  NOR3X1   g18808(.A(new_n21244_), .B(new_n21237_), .C(pi1155), .Y(new_n21245_));
  OAI21X1  g18809(.A0(new_n21245_), .A1(new_n21243_), .B0(pi0785), .Y(new_n21246_));
  OAI21X1  g18810(.A0(new_n21240_), .A1(pi0785), .B0(new_n21246_), .Y(new_n21247_));
  INVX1    g18811(.A(new_n21247_), .Y(new_n21248_));
  AOI21X1  g18812(.A0(new_n21248_), .A1(new_n12785_), .B0(new_n12615_), .Y(new_n21249_));
  AOI21X1  g18813(.A0(new_n21248_), .A1(new_n12788_), .B0(pi1154), .Y(new_n21250_));
  NOR2X1   g18814(.A(new_n21250_), .B(new_n21249_), .Y(new_n21251_));
  MX2X1    g18815(.A(new_n21251_), .B(new_n21248_), .S0(new_n11887_), .Y(new_n21252_));
  OR2X1    g18816(.A(new_n21252_), .B(pi0789), .Y(new_n21253_));
  AOI21X1  g18817(.A0(new_n21252_), .A1(new_n15910_), .B0(new_n12638_), .Y(new_n21254_));
  AOI21X1  g18818(.A0(new_n21252_), .A1(new_n15912_), .B0(pi1159), .Y(new_n21255_));
  OAI21X1  g18819(.A0(new_n21255_), .A1(new_n21254_), .B0(pi0789), .Y(new_n21256_));
  AND2X1   g18820(.A(new_n21256_), .B(new_n21253_), .Y(new_n21257_));
  INVX1    g18821(.A(new_n21257_), .Y(new_n21258_));
  MX2X1    g18822(.A(new_n21258_), .B(new_n21238_), .S0(new_n12841_), .Y(new_n21259_));
  MX2X1    g18823(.A(new_n21259_), .B(new_n21238_), .S0(new_n12711_), .Y(new_n21260_));
  AOI21X1  g18824(.A0(new_n12566_), .A1(pi0690), .B0(new_n21237_), .Y(new_n21261_));
  INVX1    g18825(.A(new_n21261_), .Y(new_n21262_));
  NOR3X1   g18826(.A(new_n13585_), .B(new_n15732_), .C(pi0625), .Y(new_n21263_));
  OR2X1    g18827(.A(new_n21263_), .B(new_n21261_), .Y(new_n21264_));
  NOR2X1   g18828(.A(new_n21237_), .B(pi1153), .Y(new_n21265_));
  INVX1    g18829(.A(new_n21265_), .Y(new_n21266_));
  OAI21X1  g18830(.A0(new_n21266_), .A1(new_n21263_), .B0(pi0778), .Y(new_n21267_));
  AOI21X1  g18831(.A0(new_n21264_), .A1(pi1153), .B0(new_n21267_), .Y(new_n21268_));
  AOI21X1  g18832(.A0(new_n21262_), .A1(new_n11889_), .B0(new_n21268_), .Y(new_n21269_));
  NOR4X1   g18833(.A(new_n21269_), .B(new_n12765_), .C(new_n12764_), .D(new_n12762_), .Y(new_n21270_));
  INVX1    g18834(.A(new_n21270_), .Y(new_n21271_));
  NOR3X1   g18835(.A(new_n21271_), .B(new_n12870_), .C(new_n12851_), .Y(new_n21272_));
  INVX1    g18836(.A(new_n21272_), .Y(new_n21273_));
  AOI21X1  g18837(.A0(new_n21237_), .A1(pi0647), .B0(pi1157), .Y(new_n21274_));
  OAI21X1  g18838(.A0(new_n21273_), .A1(pi0647), .B0(new_n21274_), .Y(new_n21275_));
  MX2X1    g18839(.A(new_n21272_), .B(new_n21237_), .S0(new_n12705_), .Y(new_n21276_));
  OAI22X1  g18840(.A0(new_n21276_), .A1(new_n14387_), .B0(new_n21275_), .B1(new_n12723_), .Y(new_n21277_));
  AOI21X1  g18841(.A0(new_n21260_), .A1(new_n14385_), .B0(new_n21277_), .Y(new_n21278_));
  NOR2X1   g18842(.A(new_n21278_), .B(new_n11883_), .Y(new_n21279_));
  AOI21X1  g18843(.A0(new_n21238_), .A1(pi0626), .B0(new_n16352_), .Y(new_n21280_));
  OAI21X1  g18844(.A0(new_n21257_), .A1(pi0626), .B0(new_n21280_), .Y(new_n21281_));
  AOI21X1  g18845(.A0(new_n21256_), .A1(new_n21253_), .B0(new_n12664_), .Y(new_n21282_));
  NOR2X1   g18846(.A(new_n21237_), .B(pi0626), .Y(new_n21283_));
  NOR3X1   g18847(.A(new_n21283_), .B(new_n21282_), .C(new_n16356_), .Y(new_n21284_));
  AOI21X1  g18848(.A0(new_n21270_), .A1(new_n12769_), .B0(new_n21284_), .Y(new_n21285_));
  AOI21X1  g18849(.A0(new_n21285_), .A1(new_n21281_), .B0(new_n11885_), .Y(new_n21286_));
  INVX1    g18850(.A(new_n21239_), .Y(new_n21287_));
  AOI21X1  g18851(.A0(new_n21262_), .A1(new_n12171_), .B0(new_n21287_), .Y(new_n21288_));
  NOR3X1   g18852(.A(new_n21261_), .B(new_n12120_), .C(new_n12493_), .Y(new_n21289_));
  OR2X1    g18853(.A(new_n21288_), .B(new_n21289_), .Y(new_n21290_));
  NOR2X1   g18854(.A(new_n21263_), .B(new_n21261_), .Y(new_n21291_));
  OAI21X1  g18855(.A0(new_n21291_), .A1(new_n12494_), .B0(new_n12584_), .Y(new_n21292_));
  AOI21X1  g18856(.A0(new_n21290_), .A1(new_n21265_), .B0(new_n21292_), .Y(new_n21293_));
  NOR3X1   g18857(.A(new_n21289_), .B(new_n21287_), .C(new_n12494_), .Y(new_n21294_));
  OAI21X1  g18858(.A0(new_n21266_), .A1(new_n21263_), .B0(pi0608), .Y(new_n21295_));
  NOR2X1   g18859(.A(new_n21295_), .B(new_n21294_), .Y(new_n21296_));
  OAI21X1  g18860(.A0(new_n21296_), .A1(new_n21293_), .B0(pi0778), .Y(new_n21297_));
  OAI21X1  g18861(.A0(new_n21288_), .A1(pi0778), .B0(new_n21297_), .Y(new_n21298_));
  OAI21X1  g18862(.A0(new_n21269_), .A1(new_n12590_), .B0(new_n12591_), .Y(new_n21299_));
  AOI21X1  g18863(.A0(new_n21298_), .A1(new_n12590_), .B0(new_n21299_), .Y(new_n21300_));
  NOR3X1   g18864(.A(new_n21300_), .B(new_n21243_), .C(pi0660), .Y(new_n21301_));
  OAI21X1  g18865(.A0(new_n21269_), .A1(pi0609), .B0(pi1155), .Y(new_n21302_));
  AOI21X1  g18866(.A0(new_n21298_), .A1(pi0609), .B0(new_n21302_), .Y(new_n21303_));
  NOR3X1   g18867(.A(new_n21303_), .B(new_n21245_), .C(new_n12596_), .Y(new_n21304_));
  OAI21X1  g18868(.A0(new_n21304_), .A1(new_n21301_), .B0(pi0785), .Y(new_n21305_));
  NAND2X1  g18869(.A(new_n21298_), .B(new_n11888_), .Y(new_n21306_));
  AND2X1   g18870(.A(new_n21306_), .B(new_n21305_), .Y(new_n21307_));
  NOR3X1   g18871(.A(new_n21269_), .B(new_n12762_), .C(new_n12614_), .Y(new_n21308_));
  NOR2X1   g18872(.A(new_n21308_), .B(pi1154), .Y(new_n21309_));
  OAI21X1  g18873(.A0(new_n21307_), .A1(pi0618), .B0(new_n21309_), .Y(new_n21310_));
  NOR2X1   g18874(.A(new_n21249_), .B(pi0627), .Y(new_n21311_));
  NOR3X1   g18875(.A(new_n21269_), .B(new_n12762_), .C(pi0618), .Y(new_n21312_));
  NOR2X1   g18876(.A(new_n21312_), .B(new_n12615_), .Y(new_n21313_));
  OAI21X1  g18877(.A0(new_n21307_), .A1(new_n12614_), .B0(new_n21313_), .Y(new_n21314_));
  NOR2X1   g18878(.A(new_n21250_), .B(new_n12622_), .Y(new_n21315_));
  AOI22X1  g18879(.A0(new_n21315_), .A1(new_n21314_), .B0(new_n21311_), .B1(new_n21310_), .Y(new_n21316_));
  MX2X1    g18880(.A(new_n21316_), .B(new_n21307_), .S0(new_n11887_), .Y(new_n21317_));
  OR4X1    g18881(.A(new_n21269_), .B(new_n12764_), .C(new_n12762_), .D(new_n12637_), .Y(new_n21318_));
  AND2X1   g18882(.A(new_n21318_), .B(new_n12638_), .Y(new_n21319_));
  OAI21X1  g18883(.A0(new_n21317_), .A1(pi0619), .B0(new_n21319_), .Y(new_n21320_));
  NOR2X1   g18884(.A(new_n21254_), .B(pi0648), .Y(new_n21321_));
  AND2X1   g18885(.A(new_n21321_), .B(new_n21320_), .Y(new_n21322_));
  INVX1    g18886(.A(new_n21322_), .Y(new_n21323_));
  NOR4X1   g18887(.A(new_n21269_), .B(new_n12764_), .C(new_n12762_), .D(pi0619), .Y(new_n21324_));
  NOR2X1   g18888(.A(new_n21324_), .B(new_n12638_), .Y(new_n21325_));
  OAI21X1  g18889(.A0(new_n21317_), .A1(new_n12637_), .B0(new_n21325_), .Y(new_n21326_));
  NOR2X1   g18890(.A(new_n21255_), .B(new_n12645_), .Y(new_n21327_));
  AOI21X1  g18891(.A0(new_n21327_), .A1(new_n21326_), .B0(new_n11886_), .Y(new_n21328_));
  AOI21X1  g18892(.A0(new_n21317_), .A1(new_n11886_), .B0(new_n14264_), .Y(new_n21329_));
  INVX1    g18893(.A(new_n21329_), .Y(new_n21330_));
  AOI21X1  g18894(.A0(new_n21328_), .A1(new_n21323_), .B0(new_n21330_), .Y(new_n21331_));
  OAI21X1  g18895(.A0(new_n21331_), .A1(new_n21286_), .B0(new_n16350_), .Y(new_n21332_));
  INVX1    g18896(.A(new_n21259_), .Y(new_n21333_));
  AND2X1   g18897(.A(new_n21270_), .B(new_n12852_), .Y(new_n21334_));
  AOI22X1  g18898(.A0(new_n21334_), .A1(new_n14564_), .B0(new_n21333_), .B1(new_n12867_), .Y(new_n21335_));
  AOI22X1  g18899(.A0(new_n21334_), .A1(new_n14566_), .B0(new_n21333_), .B1(new_n12865_), .Y(new_n21336_));
  MX2X1    g18900(.A(new_n21336_), .B(new_n21335_), .S0(new_n12689_), .Y(new_n21337_));
  OAI21X1  g18901(.A0(new_n21337_), .A1(new_n11884_), .B0(new_n14562_), .Y(new_n21338_));
  INVX1    g18902(.A(new_n21338_), .Y(new_n21339_));
  AOI21X1  g18903(.A0(new_n21339_), .A1(new_n21332_), .B0(new_n21279_), .Y(new_n21340_));
  OAI21X1  g18904(.A0(new_n21276_), .A1(new_n12706_), .B0(new_n21275_), .Y(new_n21341_));
  MX2X1    g18905(.A(new_n21341_), .B(new_n21273_), .S0(new_n11883_), .Y(new_n21342_));
  OAI21X1  g18906(.A0(new_n21342_), .A1(pi0644), .B0(pi0715), .Y(new_n21343_));
  AOI21X1  g18907(.A0(new_n21340_), .A1(pi0644), .B0(new_n21343_), .Y(new_n21344_));
  OR4X1    g18908(.A(new_n12734_), .B(new_n2739_), .C(new_n11883_), .D(pi0193), .Y(new_n21345_));
  OAI21X1  g18909(.A0(new_n21260_), .A1(new_n12735_), .B0(new_n21345_), .Y(new_n21346_));
  OAI21X1  g18910(.A0(new_n21238_), .A1(pi0644), .B0(new_n12739_), .Y(new_n21347_));
  AOI21X1  g18911(.A0(new_n21346_), .A1(pi0644), .B0(new_n21347_), .Y(new_n21348_));
  OR2X1    g18912(.A(new_n21348_), .B(new_n11882_), .Y(new_n21349_));
  OAI21X1  g18913(.A0(new_n21342_), .A1(new_n12743_), .B0(new_n12739_), .Y(new_n21350_));
  AOI21X1  g18914(.A0(new_n21340_), .A1(new_n12743_), .B0(new_n21350_), .Y(new_n21351_));
  OAI21X1  g18915(.A0(new_n21238_), .A1(new_n12743_), .B0(pi0715), .Y(new_n21352_));
  AOI21X1  g18916(.A0(new_n21346_), .A1(new_n12743_), .B0(new_n21352_), .Y(new_n21353_));
  OR2X1    g18917(.A(new_n21353_), .B(pi1160), .Y(new_n21354_));
  OAI22X1  g18918(.A0(new_n21354_), .A1(new_n21351_), .B0(new_n21349_), .B1(new_n21344_), .Y(new_n21355_));
  NAND2X1  g18919(.A(new_n21355_), .B(pi0790), .Y(new_n21356_));
  AOI21X1  g18920(.A0(new_n21340_), .A1(new_n12897_), .B0(new_n12898_), .Y(new_n21357_));
  AOI21X1  g18921(.A0(new_n13699_), .A1(new_n3129_), .B0(pi0193), .Y(new_n21358_));
  INVX1    g18922(.A(new_n21358_), .Y(new_n21359_));
  OAI21X1  g18923(.A0(new_n3810_), .A1(new_n15732_), .B0(new_n21358_), .Y(new_n21360_));
  AOI21X1  g18924(.A0(new_n12955_), .A1(pi0193), .B0(pi0038), .Y(new_n21361_));
  OAI22X1  g18925(.A0(new_n21361_), .A1(new_n3810_), .B0(new_n12953_), .B1(pi0193), .Y(new_n21362_));
  OAI21X1  g18926(.A0(new_n12202_), .A1(pi0193), .B0(new_n12567_), .Y(new_n21363_));
  NAND3X1  g18927(.A(new_n21363_), .B(new_n21362_), .C(pi0690), .Y(new_n21364_));
  AND2X1   g18928(.A(new_n21364_), .B(new_n21360_), .Y(new_n21365_));
  INVX1    g18929(.A(new_n21365_), .Y(new_n21366_));
  AOI21X1  g18930(.A0(new_n21358_), .A1(new_n12493_), .B0(new_n12494_), .Y(new_n21367_));
  OAI21X1  g18931(.A0(new_n21365_), .A1(new_n12493_), .B0(new_n21367_), .Y(new_n21368_));
  AOI21X1  g18932(.A0(new_n21358_), .A1(pi0625), .B0(pi1153), .Y(new_n21369_));
  OAI21X1  g18933(.A0(new_n21365_), .A1(pi0625), .B0(new_n21369_), .Y(new_n21370_));
  AND2X1   g18934(.A(new_n21370_), .B(new_n21368_), .Y(new_n21371_));
  MX2X1    g18935(.A(new_n21371_), .B(new_n21366_), .S0(new_n11889_), .Y(new_n21372_));
  MX2X1    g18936(.A(new_n21372_), .B(new_n21358_), .S0(new_n12618_), .Y(new_n21373_));
  INVX1    g18937(.A(new_n21373_), .Y(new_n21374_));
  MX2X1    g18938(.A(new_n21374_), .B(new_n21359_), .S0(new_n12641_), .Y(new_n21375_));
  INVX1    g18939(.A(new_n21375_), .Y(new_n21376_));
  MX2X1    g18940(.A(new_n21376_), .B(new_n21358_), .S0(new_n12659_), .Y(new_n21377_));
  AND2X1   g18941(.A(new_n21358_), .B(new_n12691_), .Y(new_n21378_));
  AOI21X1  g18942(.A0(new_n21377_), .A1(new_n17252_), .B0(new_n21378_), .Y(new_n21379_));
  AOI21X1  g18943(.A0(new_n21358_), .A1(new_n12683_), .B0(new_n12684_), .Y(new_n21380_));
  OAI21X1  g18944(.A0(new_n21379_), .A1(new_n12683_), .B0(new_n21380_), .Y(new_n21381_));
  AOI21X1  g18945(.A0(new_n21358_), .A1(pi0628), .B0(pi1156), .Y(new_n21382_));
  OAI21X1  g18946(.A0(new_n21379_), .A1(pi0628), .B0(new_n21382_), .Y(new_n21383_));
  AOI21X1  g18947(.A0(new_n21383_), .A1(new_n21381_), .B0(new_n11884_), .Y(new_n21384_));
  AOI21X1  g18948(.A0(new_n21379_), .A1(new_n11884_), .B0(new_n21384_), .Y(new_n21385_));
  MX2X1    g18949(.A(new_n21385_), .B(new_n21358_), .S0(pi0647), .Y(new_n21386_));
  MX2X1    g18950(.A(new_n21385_), .B(new_n21358_), .S0(new_n12705_), .Y(new_n21387_));
  MX2X1    g18951(.A(new_n21387_), .B(new_n21386_), .S0(new_n12706_), .Y(new_n21388_));
  MX2X1    g18952(.A(new_n21388_), .B(new_n21385_), .S0(new_n11883_), .Y(new_n21389_));
  AOI21X1  g18953(.A0(new_n21389_), .A1(new_n12743_), .B0(new_n12739_), .Y(new_n21390_));
  OAI22X1  g18954(.A0(new_n14342_), .A1(new_n15697_), .B0(new_n12202_), .B1(pi0193), .Y(new_n21391_));
  AOI21X1  g18955(.A0(new_n13977_), .A1(pi0193), .B0(new_n15697_), .Y(new_n21392_));
  OAI21X1  g18956(.A0(new_n12910_), .A1(pi0193), .B0(new_n21392_), .Y(new_n21393_));
  NAND3X1  g18957(.A(new_n12090_), .B(new_n15697_), .C(new_n7083_), .Y(new_n21394_));
  AOI21X1  g18958(.A0(new_n21394_), .A1(new_n21393_), .B0(pi0038), .Y(new_n21395_));
  AOI21X1  g18959(.A0(new_n21391_), .A1(pi0038), .B0(new_n21395_), .Y(new_n21396_));
  MX2X1    g18960(.A(new_n21396_), .B(pi0193), .S0(new_n3810_), .Y(new_n21397_));
  AND2X1   g18961(.A(new_n21397_), .B(new_n12623_), .Y(new_n21398_));
  AOI21X1  g18962(.A0(new_n21359_), .A1(new_n12601_), .B0(new_n21398_), .Y(new_n21399_));
  AOI22X1  g18963(.A0(new_n21398_), .A1(pi0609), .B0(new_n21359_), .B1(new_n13430_), .Y(new_n21400_));
  AOI22X1  g18964(.A0(new_n21398_), .A1(new_n12590_), .B0(new_n21359_), .B1(new_n13436_), .Y(new_n21401_));
  MX2X1    g18965(.A(new_n21401_), .B(new_n21400_), .S0(pi1155), .Y(new_n21402_));
  MX2X1    g18966(.A(new_n21402_), .B(new_n21399_), .S0(new_n11888_), .Y(new_n21403_));
  OAI21X1  g18967(.A0(new_n21359_), .A1(pi0618), .B0(pi1154), .Y(new_n21404_));
  AOI21X1  g18968(.A0(new_n21403_), .A1(pi0618), .B0(new_n21404_), .Y(new_n21405_));
  OAI21X1  g18969(.A0(new_n21359_), .A1(new_n12614_), .B0(new_n12615_), .Y(new_n21406_));
  AOI21X1  g18970(.A0(new_n21403_), .A1(new_n12614_), .B0(new_n21406_), .Y(new_n21407_));
  NOR2X1   g18971(.A(new_n21407_), .B(new_n21405_), .Y(new_n21408_));
  MX2X1    g18972(.A(new_n21408_), .B(new_n21403_), .S0(new_n11887_), .Y(new_n21409_));
  OAI21X1  g18973(.A0(new_n21359_), .A1(pi0619), .B0(pi1159), .Y(new_n21410_));
  AOI21X1  g18974(.A0(new_n21409_), .A1(pi0619), .B0(new_n21410_), .Y(new_n21411_));
  OAI21X1  g18975(.A0(new_n21359_), .A1(new_n12637_), .B0(new_n12638_), .Y(new_n21412_));
  AOI21X1  g18976(.A0(new_n21409_), .A1(new_n12637_), .B0(new_n21412_), .Y(new_n21413_));
  NOR2X1   g18977(.A(new_n21413_), .B(new_n21411_), .Y(new_n21414_));
  MX2X1    g18978(.A(new_n21414_), .B(new_n21409_), .S0(new_n11886_), .Y(new_n21415_));
  MX2X1    g18979(.A(new_n21415_), .B(new_n21358_), .S0(new_n12841_), .Y(new_n21416_));
  MX2X1    g18980(.A(new_n21416_), .B(new_n21358_), .S0(new_n12711_), .Y(new_n21417_));
  MX2X1    g18981(.A(new_n21417_), .B(new_n21358_), .S0(new_n12735_), .Y(new_n21418_));
  OAI21X1  g18982(.A0(new_n21359_), .A1(pi0644), .B0(new_n12739_), .Y(new_n21419_));
  AOI21X1  g18983(.A0(new_n21418_), .A1(pi0644), .B0(new_n21419_), .Y(new_n21420_));
  OR2X1    g18984(.A(new_n21420_), .B(new_n11882_), .Y(new_n21421_));
  AOI21X1  g18985(.A0(new_n21389_), .A1(pi0644), .B0(pi0715), .Y(new_n21422_));
  OAI21X1  g18986(.A0(new_n21359_), .A1(new_n12743_), .B0(pi0715), .Y(new_n21423_));
  AOI21X1  g18987(.A0(new_n21418_), .A1(new_n12743_), .B0(new_n21423_), .Y(new_n21424_));
  OR2X1    g18988(.A(new_n21424_), .B(pi1160), .Y(new_n21425_));
  OAI22X1  g18989(.A0(new_n21425_), .A1(new_n21422_), .B0(new_n21421_), .B1(new_n21390_), .Y(new_n21426_));
  NOR3X1   g18990(.A(new_n21424_), .B(pi1160), .C(pi0644), .Y(new_n21427_));
  NOR3X1   g18991(.A(new_n21420_), .B(new_n11882_), .C(new_n12743_), .Y(new_n21428_));
  NOR3X1   g18992(.A(new_n21428_), .B(new_n21427_), .C(new_n12897_), .Y(new_n21429_));
  MX2X1    g18993(.A(new_n21383_), .B(new_n21381_), .S0(new_n12689_), .Y(new_n21430_));
  OAI21X1  g18994(.A0(new_n21416_), .A1(new_n14395_), .B0(new_n21430_), .Y(new_n21431_));
  NAND2X1  g18995(.A(new_n21431_), .B(pi0792), .Y(new_n21432_));
  OR2X1    g18996(.A(new_n21396_), .B(pi0690), .Y(new_n21433_));
  OAI21X1  g18997(.A0(new_n12349_), .A1(new_n7083_), .B0(new_n15697_), .Y(new_n21434_));
  AOI21X1  g18998(.A0(new_n12289_), .A1(new_n7083_), .B0(new_n21434_), .Y(new_n21435_));
  OAI21X1  g18999(.A0(new_n12440_), .A1(pi0193), .B0(pi0739), .Y(new_n21436_));
  AOI21X1  g19000(.A0(new_n12401_), .A1(pi0193), .B0(new_n21436_), .Y(new_n21437_));
  OR2X1    g19001(.A(new_n21437_), .B(new_n2959_), .Y(new_n21438_));
  NOR4X1   g19002(.A(new_n13391_), .B(new_n12908_), .C(new_n12907_), .D(pi0193), .Y(new_n21439_));
  OAI21X1  g19003(.A0(new_n12929_), .A1(new_n7083_), .B0(pi0739), .Y(new_n21440_));
  AND2X1   g19004(.A(new_n12467_), .B(pi0193), .Y(new_n21441_));
  OAI21X1  g19005(.A0(new_n12454_), .A1(pi0193), .B0(new_n15697_), .Y(new_n21442_));
  OAI22X1  g19006(.A0(new_n21442_), .A1(new_n21441_), .B0(new_n21440_), .B1(new_n21439_), .Y(new_n21443_));
  AOI21X1  g19007(.A0(new_n21443_), .A1(new_n2959_), .B0(pi0038), .Y(new_n21444_));
  OAI21X1  g19008(.A0(new_n21438_), .A1(new_n21435_), .B0(new_n21444_), .Y(new_n21445_));
  AOI21X1  g19009(.A0(new_n16526_), .A1(new_n15697_), .B0(new_n12478_), .Y(new_n21446_));
  OAI21X1  g19010(.A0(new_n21446_), .A1(pi0039), .B0(new_n7083_), .Y(new_n21447_));
  AOI21X1  g19011(.A0(new_n21241_), .A1(new_n14209_), .B0(new_n7083_), .Y(new_n21448_));
  AOI21X1  g19012(.A0(new_n21448_), .A1(new_n6857_), .B0(new_n2996_), .Y(new_n21449_));
  AOI21X1  g19013(.A0(new_n21449_), .A1(new_n21447_), .B0(new_n15732_), .Y(new_n21450_));
  AOI21X1  g19014(.A0(new_n21450_), .A1(new_n21445_), .B0(new_n3810_), .Y(new_n21451_));
  AOI22X1  g19015(.A0(new_n21451_), .A1(new_n21433_), .B0(new_n3810_), .B1(pi0193), .Y(new_n21452_));
  OAI21X1  g19016(.A0(new_n21397_), .A1(new_n12493_), .B0(new_n12494_), .Y(new_n21453_));
  AOI21X1  g19017(.A0(new_n21452_), .A1(new_n12493_), .B0(new_n21453_), .Y(new_n21454_));
  NAND2X1  g19018(.A(new_n21368_), .B(new_n12584_), .Y(new_n21455_));
  OAI21X1  g19019(.A0(new_n21397_), .A1(pi0625), .B0(pi1153), .Y(new_n21456_));
  AOI21X1  g19020(.A0(new_n21452_), .A1(pi0625), .B0(new_n21456_), .Y(new_n21457_));
  NAND2X1  g19021(.A(new_n21370_), .B(pi0608), .Y(new_n21458_));
  OAI22X1  g19022(.A0(new_n21458_), .A1(new_n21457_), .B0(new_n21455_), .B1(new_n21454_), .Y(new_n21459_));
  MX2X1    g19023(.A(new_n21459_), .B(new_n21452_), .S0(new_n11889_), .Y(new_n21460_));
  INVX1    g19024(.A(new_n21372_), .Y(new_n21461_));
  OAI21X1  g19025(.A0(new_n21461_), .A1(new_n12590_), .B0(new_n12591_), .Y(new_n21462_));
  AOI21X1  g19026(.A0(new_n21460_), .A1(new_n12590_), .B0(new_n21462_), .Y(new_n21463_));
  OAI21X1  g19027(.A0(new_n21400_), .A1(new_n12591_), .B0(new_n12596_), .Y(new_n21464_));
  OAI21X1  g19028(.A0(new_n21461_), .A1(pi0609), .B0(pi1155), .Y(new_n21465_));
  AOI21X1  g19029(.A0(new_n21460_), .A1(pi0609), .B0(new_n21465_), .Y(new_n21466_));
  OAI21X1  g19030(.A0(new_n21401_), .A1(pi1155), .B0(pi0660), .Y(new_n21467_));
  OAI22X1  g19031(.A0(new_n21467_), .A1(new_n21466_), .B0(new_n21464_), .B1(new_n21463_), .Y(new_n21468_));
  MX2X1    g19032(.A(new_n21468_), .B(new_n21460_), .S0(new_n11888_), .Y(new_n21469_));
  OAI21X1  g19033(.A0(new_n21374_), .A1(new_n12614_), .B0(new_n12615_), .Y(new_n21470_));
  AOI21X1  g19034(.A0(new_n21469_), .A1(new_n12614_), .B0(new_n21470_), .Y(new_n21471_));
  OR2X1    g19035(.A(new_n21405_), .B(pi0627), .Y(new_n21472_));
  OAI21X1  g19036(.A0(new_n21374_), .A1(pi0618), .B0(pi1154), .Y(new_n21473_));
  AOI21X1  g19037(.A0(new_n21469_), .A1(pi0618), .B0(new_n21473_), .Y(new_n21474_));
  OR2X1    g19038(.A(new_n21407_), .B(new_n12622_), .Y(new_n21475_));
  OAI22X1  g19039(.A0(new_n21475_), .A1(new_n21474_), .B0(new_n21472_), .B1(new_n21471_), .Y(new_n21476_));
  MX2X1    g19040(.A(new_n21476_), .B(new_n21469_), .S0(new_n11887_), .Y(new_n21477_));
  NAND2X1  g19041(.A(new_n21477_), .B(new_n12637_), .Y(new_n21478_));
  AOI21X1  g19042(.A0(new_n21376_), .A1(pi0619), .B0(pi1159), .Y(new_n21479_));
  OR2X1    g19043(.A(new_n21411_), .B(pi0648), .Y(new_n21480_));
  AOI21X1  g19044(.A0(new_n21479_), .A1(new_n21478_), .B0(new_n21480_), .Y(new_n21481_));
  NAND2X1  g19045(.A(new_n21477_), .B(pi0619), .Y(new_n21482_));
  AOI21X1  g19046(.A0(new_n21376_), .A1(new_n12637_), .B0(new_n12638_), .Y(new_n21483_));
  OR2X1    g19047(.A(new_n21413_), .B(new_n12645_), .Y(new_n21484_));
  AOI21X1  g19048(.A0(new_n21483_), .A1(new_n21482_), .B0(new_n21484_), .Y(new_n21485_));
  NOR3X1   g19049(.A(new_n21485_), .B(new_n21481_), .C(new_n11886_), .Y(new_n21486_));
  OAI21X1  g19050(.A0(new_n21477_), .A1(pi0789), .B0(new_n12842_), .Y(new_n21487_));
  AOI21X1  g19051(.A0(new_n21359_), .A1(pi0626), .B0(new_n16352_), .Y(new_n21488_));
  OAI21X1  g19052(.A0(new_n21415_), .A1(pi0626), .B0(new_n21488_), .Y(new_n21489_));
  AOI21X1  g19053(.A0(new_n21359_), .A1(new_n12664_), .B0(new_n16356_), .Y(new_n21490_));
  OAI21X1  g19054(.A0(new_n21415_), .A1(new_n12664_), .B0(new_n21490_), .Y(new_n21491_));
  NAND2X1  g19055(.A(new_n21377_), .B(new_n12769_), .Y(new_n21492_));
  NAND3X1  g19056(.A(new_n21492_), .B(new_n21491_), .C(new_n21489_), .Y(new_n21493_));
  AOI21X1  g19057(.A0(new_n21493_), .A1(pi0788), .B0(new_n14273_), .Y(new_n21494_));
  OAI21X1  g19058(.A0(new_n21487_), .A1(new_n21486_), .B0(new_n21494_), .Y(new_n21495_));
  AOI21X1  g19059(.A0(new_n21495_), .A1(new_n21432_), .B0(new_n14269_), .Y(new_n21496_));
  OR2X1    g19060(.A(new_n21417_), .B(new_n14384_), .Y(new_n21497_));
  OR2X1    g19061(.A(new_n21386_), .B(new_n14389_), .Y(new_n21498_));
  OR2X1    g19062(.A(new_n21387_), .B(new_n14387_), .Y(new_n21499_));
  NAND3X1  g19063(.A(new_n21499_), .B(new_n21498_), .C(new_n21497_), .Y(new_n21500_));
  AND2X1   g19064(.A(new_n21500_), .B(pi0787), .Y(new_n21501_));
  NOR3X1   g19065(.A(new_n21501_), .B(new_n21496_), .C(new_n21429_), .Y(new_n21502_));
  AOI21X1  g19066(.A0(new_n21426_), .A1(pi0790), .B0(new_n21502_), .Y(new_n21503_));
  OR2X1    g19067(.A(new_n21503_), .B(po1038), .Y(new_n21504_));
  AOI21X1  g19068(.A0(po1038), .A1(new_n7083_), .B0(pi0832), .Y(new_n21505_));
  AOI22X1  g19069(.A0(new_n21505_), .A1(new_n21504_), .B0(new_n21357_), .B1(new_n21356_), .Y(po0350));
  MX2X1    g19070(.A(new_n16746_), .B(new_n16744_), .S0(new_n11641_), .Y(new_n21507_));
  OAI21X1  g19071(.A0(new_n13699_), .A1(pi0194), .B0(new_n15595_), .Y(new_n21508_));
  OAI21X1  g19072(.A0(new_n21507_), .A1(new_n15595_), .B0(new_n21508_), .Y(new_n21509_));
  OR2X1    g19073(.A(new_n21509_), .B(pi0730), .Y(new_n21510_));
  AND2X1   g19074(.A(new_n13672_), .B(new_n11641_), .Y(new_n21511_));
  OAI21X1  g19075(.A0(new_n13676_), .A1(new_n16792_), .B0(pi0194), .Y(new_n21512_));
  NAND2X1  g19076(.A(new_n21512_), .B(new_n15595_), .Y(new_n21513_));
  INVX1    g19077(.A(pi0730), .Y(new_n21514_));
  OAI21X1  g19078(.A0(new_n13694_), .A1(pi0194), .B0(pi0748), .Y(new_n21515_));
  AOI21X1  g19079(.A0(new_n13688_), .A1(pi0194), .B0(new_n21515_), .Y(new_n21516_));
  NOR2X1   g19080(.A(new_n21516_), .B(new_n21514_), .Y(new_n21517_));
  OAI21X1  g19081(.A0(new_n21513_), .A1(new_n21511_), .B0(new_n21517_), .Y(new_n21518_));
  AND2X1   g19082(.A(new_n21518_), .B(new_n3129_), .Y(new_n21519_));
  AOI22X1  g19083(.A0(new_n21519_), .A1(new_n21510_), .B0(new_n3810_), .B1(pi0194), .Y(new_n21520_));
  MX2X1    g19084(.A(new_n21509_), .B(pi0194), .S0(new_n3810_), .Y(new_n21521_));
  OAI21X1  g19085(.A0(new_n21521_), .A1(new_n12493_), .B0(new_n12494_), .Y(new_n21522_));
  AOI21X1  g19086(.A0(new_n21520_), .A1(new_n12493_), .B0(new_n21522_), .Y(new_n21523_));
  OAI21X1  g19087(.A0(new_n16716_), .A1(pi0194), .B0(pi0730), .Y(new_n21524_));
  NAND3X1  g19088(.A(new_n12574_), .B(new_n21514_), .C(new_n11641_), .Y(new_n21525_));
  AND2X1   g19089(.A(new_n21525_), .B(new_n3129_), .Y(new_n21526_));
  AOI22X1  g19090(.A0(new_n21526_), .A1(new_n21524_), .B0(new_n16715_), .B1(pi0194), .Y(new_n21527_));
  OAI21X1  g19091(.A0(new_n12574_), .A1(new_n3810_), .B0(new_n11641_), .Y(new_n21528_));
  OAI21X1  g19092(.A0(new_n21528_), .A1(pi0625), .B0(pi1153), .Y(new_n21529_));
  AOI21X1  g19093(.A0(new_n21527_), .A1(pi0625), .B0(new_n21529_), .Y(new_n21530_));
  OR2X1    g19094(.A(new_n21530_), .B(pi0608), .Y(new_n21531_));
  OAI21X1  g19095(.A0(new_n21521_), .A1(pi0625), .B0(pi1153), .Y(new_n21532_));
  AOI21X1  g19096(.A0(new_n21520_), .A1(pi0625), .B0(new_n21532_), .Y(new_n21533_));
  OAI21X1  g19097(.A0(new_n21528_), .A1(new_n12493_), .B0(new_n12494_), .Y(new_n21534_));
  AOI21X1  g19098(.A0(new_n21527_), .A1(new_n12493_), .B0(new_n21534_), .Y(new_n21535_));
  OR2X1    g19099(.A(new_n21535_), .B(new_n12584_), .Y(new_n21536_));
  OAI22X1  g19100(.A0(new_n21536_), .A1(new_n21533_), .B0(new_n21531_), .B1(new_n21523_), .Y(new_n21537_));
  MX2X1    g19101(.A(new_n21537_), .B(new_n21520_), .S0(new_n11889_), .Y(new_n21538_));
  OAI21X1  g19102(.A0(new_n21535_), .A1(new_n21530_), .B0(pi0778), .Y(new_n21539_));
  OAI21X1  g19103(.A0(new_n21527_), .A1(pi0778), .B0(new_n21539_), .Y(new_n21540_));
  OAI21X1  g19104(.A0(new_n21540_), .A1(new_n12590_), .B0(new_n12591_), .Y(new_n21541_));
  AOI21X1  g19105(.A0(new_n21538_), .A1(new_n12590_), .B0(new_n21541_), .Y(new_n21542_));
  AND2X1   g19106(.A(new_n21521_), .B(new_n12623_), .Y(new_n21543_));
  AOI22X1  g19107(.A0(new_n21543_), .A1(pi0609), .B0(new_n21528_), .B1(new_n13430_), .Y(new_n21544_));
  OAI21X1  g19108(.A0(new_n21544_), .A1(new_n12591_), .B0(new_n12596_), .Y(new_n21545_));
  OAI21X1  g19109(.A0(new_n21540_), .A1(pi0609), .B0(pi1155), .Y(new_n21546_));
  AOI21X1  g19110(.A0(new_n21538_), .A1(pi0609), .B0(new_n21546_), .Y(new_n21547_));
  AOI22X1  g19111(.A0(new_n21543_), .A1(new_n12590_), .B0(new_n21528_), .B1(new_n13436_), .Y(new_n21548_));
  OAI21X1  g19112(.A0(new_n21548_), .A1(pi1155), .B0(pi0660), .Y(new_n21549_));
  OAI22X1  g19113(.A0(new_n21549_), .A1(new_n21547_), .B0(new_n21545_), .B1(new_n21542_), .Y(new_n21550_));
  MX2X1    g19114(.A(new_n21550_), .B(new_n21538_), .S0(new_n11888_), .Y(new_n21551_));
  MX2X1    g19115(.A(new_n21540_), .B(new_n21528_), .S0(new_n12618_), .Y(new_n21552_));
  OAI21X1  g19116(.A0(new_n21552_), .A1(new_n12614_), .B0(new_n12615_), .Y(new_n21553_));
  AOI21X1  g19117(.A0(new_n21551_), .A1(new_n12614_), .B0(new_n21553_), .Y(new_n21554_));
  AOI21X1  g19118(.A0(new_n21528_), .A1(new_n12601_), .B0(new_n21543_), .Y(new_n21555_));
  MX2X1    g19119(.A(new_n21548_), .B(new_n21544_), .S0(pi1155), .Y(new_n21556_));
  MX2X1    g19120(.A(new_n21556_), .B(new_n21555_), .S0(new_n11888_), .Y(new_n21557_));
  OAI21X1  g19121(.A0(new_n21528_), .A1(pi0618), .B0(pi1154), .Y(new_n21558_));
  AOI21X1  g19122(.A0(new_n21557_), .A1(pi0618), .B0(new_n21558_), .Y(new_n21559_));
  OR2X1    g19123(.A(new_n21559_), .B(pi0627), .Y(new_n21560_));
  OAI21X1  g19124(.A0(new_n21552_), .A1(pi0618), .B0(pi1154), .Y(new_n21561_));
  AOI21X1  g19125(.A0(new_n21551_), .A1(pi0618), .B0(new_n21561_), .Y(new_n21562_));
  OAI21X1  g19126(.A0(new_n21528_), .A1(new_n12614_), .B0(new_n12615_), .Y(new_n21563_));
  AOI21X1  g19127(.A0(new_n21557_), .A1(new_n12614_), .B0(new_n21563_), .Y(new_n21564_));
  OR2X1    g19128(.A(new_n21564_), .B(new_n12622_), .Y(new_n21565_));
  OAI22X1  g19129(.A0(new_n21565_), .A1(new_n21562_), .B0(new_n21560_), .B1(new_n21554_), .Y(new_n21566_));
  MX2X1    g19130(.A(new_n21566_), .B(new_n21551_), .S0(new_n11887_), .Y(new_n21567_));
  MX2X1    g19131(.A(new_n21552_), .B(new_n21528_), .S0(new_n12641_), .Y(new_n21568_));
  OAI21X1  g19132(.A0(new_n21568_), .A1(new_n12637_), .B0(new_n12638_), .Y(new_n21569_));
  AOI21X1  g19133(.A0(new_n21567_), .A1(new_n12637_), .B0(new_n21569_), .Y(new_n21570_));
  NOR2X1   g19134(.A(new_n21564_), .B(new_n21559_), .Y(new_n21571_));
  MX2X1    g19135(.A(new_n21571_), .B(new_n21557_), .S0(new_n11887_), .Y(new_n21572_));
  OAI21X1  g19136(.A0(new_n21528_), .A1(pi0619), .B0(pi1159), .Y(new_n21573_));
  AOI21X1  g19137(.A0(new_n21572_), .A1(pi0619), .B0(new_n21573_), .Y(new_n21574_));
  OR2X1    g19138(.A(new_n21574_), .B(pi0648), .Y(new_n21575_));
  OAI21X1  g19139(.A0(new_n21568_), .A1(pi0619), .B0(pi1159), .Y(new_n21576_));
  AOI21X1  g19140(.A0(new_n21567_), .A1(pi0619), .B0(new_n21576_), .Y(new_n21577_));
  OAI21X1  g19141(.A0(new_n21528_), .A1(new_n12637_), .B0(new_n12638_), .Y(new_n21578_));
  AOI21X1  g19142(.A0(new_n21572_), .A1(new_n12637_), .B0(new_n21578_), .Y(new_n21579_));
  OR2X1    g19143(.A(new_n21579_), .B(new_n12645_), .Y(new_n21580_));
  OAI22X1  g19144(.A0(new_n21580_), .A1(new_n21577_), .B0(new_n21575_), .B1(new_n21570_), .Y(new_n21581_));
  MX2X1    g19145(.A(new_n21581_), .B(new_n21567_), .S0(new_n11886_), .Y(new_n21582_));
  MX2X1    g19146(.A(new_n21568_), .B(new_n21528_), .S0(new_n12659_), .Y(new_n21583_));
  AOI21X1  g19147(.A0(new_n21583_), .A1(pi0626), .B0(pi0641), .Y(new_n21584_));
  OAI21X1  g19148(.A0(new_n21582_), .A1(pi0626), .B0(new_n21584_), .Y(new_n21585_));
  OR2X1    g19149(.A(new_n21572_), .B(pi0789), .Y(new_n21586_));
  OAI21X1  g19150(.A0(new_n21579_), .A1(new_n21574_), .B0(pi0789), .Y(new_n21587_));
  NAND2X1  g19151(.A(new_n21587_), .B(new_n21586_), .Y(new_n21588_));
  NAND2X1  g19152(.A(new_n21588_), .B(new_n12664_), .Y(new_n21589_));
  AOI21X1  g19153(.A0(new_n21528_), .A1(pi0626), .B0(new_n12672_), .Y(new_n21590_));
  AOI21X1  g19154(.A0(new_n21590_), .A1(new_n21589_), .B0(pi1158), .Y(new_n21591_));
  AOI21X1  g19155(.A0(new_n21583_), .A1(new_n12664_), .B0(new_n12672_), .Y(new_n21592_));
  OAI21X1  g19156(.A0(new_n21582_), .A1(new_n12664_), .B0(new_n21592_), .Y(new_n21593_));
  NAND2X1  g19157(.A(new_n21588_), .B(pi0626), .Y(new_n21594_));
  AOI21X1  g19158(.A0(new_n21528_), .A1(new_n12664_), .B0(pi0641), .Y(new_n21595_));
  AOI21X1  g19159(.A0(new_n21595_), .A1(new_n21594_), .B0(new_n12676_), .Y(new_n21596_));
  AOI22X1  g19160(.A0(new_n21596_), .A1(new_n21593_), .B0(new_n21591_), .B1(new_n21585_), .Y(new_n21597_));
  MX2X1    g19161(.A(new_n21597_), .B(new_n21582_), .S0(new_n11885_), .Y(new_n21598_));
  MX2X1    g19162(.A(new_n21588_), .B(new_n21528_), .S0(new_n12841_), .Y(new_n21599_));
  OAI21X1  g19163(.A0(new_n21599_), .A1(new_n12683_), .B0(new_n12684_), .Y(new_n21600_));
  AOI21X1  g19164(.A0(new_n21598_), .A1(new_n12683_), .B0(new_n21600_), .Y(new_n21601_));
  MX2X1    g19165(.A(new_n21583_), .B(new_n21528_), .S0(new_n12691_), .Y(new_n21602_));
  INVX1    g19166(.A(new_n21528_), .Y(new_n21603_));
  AOI21X1  g19167(.A0(new_n21603_), .A1(new_n12683_), .B0(new_n12684_), .Y(new_n21604_));
  OAI21X1  g19168(.A0(new_n21602_), .A1(new_n12683_), .B0(new_n21604_), .Y(new_n21605_));
  AND2X1   g19169(.A(new_n21605_), .B(new_n12689_), .Y(new_n21606_));
  INVX1    g19170(.A(new_n21606_), .Y(new_n21607_));
  OAI21X1  g19171(.A0(new_n21599_), .A1(pi0628), .B0(pi1156), .Y(new_n21608_));
  AOI21X1  g19172(.A0(new_n21598_), .A1(pi0628), .B0(new_n21608_), .Y(new_n21609_));
  AOI21X1  g19173(.A0(new_n21603_), .A1(pi0628), .B0(pi1156), .Y(new_n21610_));
  OAI21X1  g19174(.A0(new_n21602_), .A1(pi0628), .B0(new_n21610_), .Y(new_n21611_));
  AND2X1   g19175(.A(new_n21611_), .B(pi0629), .Y(new_n21612_));
  INVX1    g19176(.A(new_n21612_), .Y(new_n21613_));
  OAI22X1  g19177(.A0(new_n21613_), .A1(new_n21609_), .B0(new_n21607_), .B1(new_n21601_), .Y(new_n21614_));
  MX2X1    g19178(.A(new_n21614_), .B(new_n21598_), .S0(new_n11884_), .Y(new_n21615_));
  MX2X1    g19179(.A(new_n21599_), .B(new_n21528_), .S0(new_n12711_), .Y(new_n21616_));
  OAI21X1  g19180(.A0(new_n21616_), .A1(new_n12705_), .B0(new_n12706_), .Y(new_n21617_));
  AOI21X1  g19181(.A0(new_n21615_), .A1(new_n12705_), .B0(new_n21617_), .Y(new_n21618_));
  AOI21X1  g19182(.A0(new_n21611_), .A1(new_n21605_), .B0(new_n11884_), .Y(new_n21619_));
  AOI21X1  g19183(.A0(new_n21602_), .A1(new_n11884_), .B0(new_n21619_), .Y(new_n21620_));
  OAI21X1  g19184(.A0(new_n21528_), .A1(pi0647), .B0(pi1157), .Y(new_n21621_));
  AOI21X1  g19185(.A0(new_n21620_), .A1(pi0647), .B0(new_n21621_), .Y(new_n21622_));
  NOR2X1   g19186(.A(new_n21622_), .B(pi0630), .Y(new_n21623_));
  INVX1    g19187(.A(new_n21623_), .Y(new_n21624_));
  OAI21X1  g19188(.A0(new_n21616_), .A1(pi0647), .B0(pi1157), .Y(new_n21625_));
  AOI21X1  g19189(.A0(new_n21615_), .A1(pi0647), .B0(new_n21625_), .Y(new_n21626_));
  OAI21X1  g19190(.A0(new_n21528_), .A1(new_n12705_), .B0(new_n12706_), .Y(new_n21627_));
  AOI21X1  g19191(.A0(new_n21620_), .A1(new_n12705_), .B0(new_n21627_), .Y(new_n21628_));
  NOR2X1   g19192(.A(new_n21628_), .B(new_n12723_), .Y(new_n21629_));
  INVX1    g19193(.A(new_n21629_), .Y(new_n21630_));
  OAI22X1  g19194(.A0(new_n21630_), .A1(new_n21626_), .B0(new_n21624_), .B1(new_n21618_), .Y(new_n21631_));
  MX2X1    g19195(.A(new_n21631_), .B(new_n21615_), .S0(new_n11883_), .Y(new_n21632_));
  OAI21X1  g19196(.A0(new_n21628_), .A1(new_n21622_), .B0(pi0787), .Y(new_n21633_));
  OAI21X1  g19197(.A0(new_n21620_), .A1(pi0787), .B0(new_n21633_), .Y(new_n21634_));
  OAI21X1  g19198(.A0(new_n21634_), .A1(pi0644), .B0(pi0715), .Y(new_n21635_));
  AOI21X1  g19199(.A0(new_n21632_), .A1(pi0644), .B0(new_n21635_), .Y(new_n21636_));
  AND2X1   g19200(.A(new_n21528_), .B(new_n12735_), .Y(new_n21637_));
  AOI21X1  g19201(.A0(new_n21616_), .A1(new_n12736_), .B0(new_n21637_), .Y(new_n21638_));
  OAI21X1  g19202(.A0(new_n21528_), .A1(pi0644), .B0(new_n12739_), .Y(new_n21639_));
  AOI21X1  g19203(.A0(new_n21638_), .A1(pi0644), .B0(new_n21639_), .Y(new_n21640_));
  NOR3X1   g19204(.A(new_n21640_), .B(new_n21636_), .C(new_n11882_), .Y(new_n21641_));
  OAI21X1  g19205(.A0(new_n21634_), .A1(new_n12743_), .B0(new_n12739_), .Y(new_n21642_));
  AOI21X1  g19206(.A0(new_n21632_), .A1(new_n12743_), .B0(new_n21642_), .Y(new_n21643_));
  OAI21X1  g19207(.A0(new_n21528_), .A1(new_n12743_), .B0(pi0715), .Y(new_n21644_));
  AOI21X1  g19208(.A0(new_n21638_), .A1(new_n12743_), .B0(new_n21644_), .Y(new_n21645_));
  OR2X1    g19209(.A(new_n21645_), .B(pi1160), .Y(new_n21646_));
  OAI21X1  g19210(.A0(new_n21646_), .A1(new_n21643_), .B0(pi0790), .Y(new_n21647_));
  OR2X1    g19211(.A(new_n21632_), .B(pi0790), .Y(new_n21648_));
  AND2X1   g19212(.A(new_n21648_), .B(new_n6520_), .Y(new_n21649_));
  OAI21X1  g19213(.A0(new_n21647_), .A1(new_n21641_), .B0(new_n21649_), .Y(new_n21650_));
  AOI21X1  g19214(.A0(po1038), .A1(new_n11641_), .B0(pi0832), .Y(new_n21651_));
  AOI21X1  g19215(.A0(pi1093), .A1(pi1092), .B0(pi0194), .Y(new_n21652_));
  INVX1    g19216(.A(new_n21652_), .Y(new_n21653_));
  AOI21X1  g19217(.A0(new_n12178_), .A1(pi0748), .B0(new_n21652_), .Y(new_n21654_));
  AOI21X1  g19218(.A0(new_n12601_), .A1(new_n2739_), .B0(new_n21654_), .Y(new_n21655_));
  INVX1    g19219(.A(new_n21654_), .Y(new_n21656_));
  AOI21X1  g19220(.A0(new_n21656_), .A1(new_n12776_), .B0(new_n12591_), .Y(new_n21657_));
  AOI21X1  g19221(.A0(new_n21655_), .A1(new_n12779_), .B0(pi1155), .Y(new_n21658_));
  OAI21X1  g19222(.A0(new_n21658_), .A1(new_n21657_), .B0(pi0785), .Y(new_n21659_));
  OAI21X1  g19223(.A0(new_n21655_), .A1(pi0785), .B0(new_n21659_), .Y(new_n21660_));
  INVX1    g19224(.A(new_n21660_), .Y(new_n21661_));
  AOI21X1  g19225(.A0(new_n21661_), .A1(new_n12785_), .B0(new_n12615_), .Y(new_n21662_));
  AOI21X1  g19226(.A0(new_n21661_), .A1(new_n12788_), .B0(pi1154), .Y(new_n21663_));
  OR2X1    g19227(.A(new_n21663_), .B(new_n21662_), .Y(new_n21664_));
  MX2X1    g19228(.A(new_n21664_), .B(new_n21660_), .S0(new_n11887_), .Y(new_n21665_));
  AND2X1   g19229(.A(new_n21665_), .B(new_n11886_), .Y(new_n21666_));
  AOI21X1  g19230(.A0(new_n21652_), .A1(new_n12637_), .B0(new_n12638_), .Y(new_n21667_));
  OAI21X1  g19231(.A0(new_n21665_), .A1(new_n12637_), .B0(new_n21667_), .Y(new_n21668_));
  AOI21X1  g19232(.A0(new_n21652_), .A1(pi0619), .B0(pi1159), .Y(new_n21669_));
  OAI21X1  g19233(.A0(new_n21665_), .A1(pi0619), .B0(new_n21669_), .Y(new_n21670_));
  AOI21X1  g19234(.A0(new_n21670_), .A1(new_n21668_), .B0(new_n11886_), .Y(new_n21671_));
  NOR2X1   g19235(.A(new_n21671_), .B(new_n21666_), .Y(new_n21672_));
  INVX1    g19236(.A(new_n21672_), .Y(new_n21673_));
  MX2X1    g19237(.A(new_n21673_), .B(new_n21653_), .S0(new_n12841_), .Y(new_n21674_));
  MX2X1    g19238(.A(new_n21674_), .B(new_n21653_), .S0(new_n12711_), .Y(new_n21675_));
  AOI21X1  g19239(.A0(new_n12566_), .A1(pi0730), .B0(new_n21652_), .Y(new_n21676_));
  AND2X1   g19240(.A(new_n12566_), .B(pi0730), .Y(new_n21677_));
  AND2X1   g19241(.A(new_n21677_), .B(new_n12493_), .Y(new_n21678_));
  MX2X1    g19242(.A(new_n21652_), .B(pi0625), .S0(new_n21677_), .Y(new_n21679_));
  NOR2X1   g19243(.A(new_n21652_), .B(pi1153), .Y(new_n21680_));
  INVX1    g19244(.A(new_n21680_), .Y(new_n21681_));
  OAI22X1  g19245(.A0(new_n21681_), .A1(new_n21678_), .B0(new_n21679_), .B1(new_n12494_), .Y(new_n21682_));
  MX2X1    g19246(.A(new_n21682_), .B(new_n21676_), .S0(new_n11889_), .Y(new_n21683_));
  NOR4X1   g19247(.A(new_n21683_), .B(new_n12765_), .C(new_n12764_), .D(new_n12762_), .Y(new_n21684_));
  INVX1    g19248(.A(new_n21684_), .Y(new_n21685_));
  NOR3X1   g19249(.A(new_n21685_), .B(new_n12870_), .C(new_n12851_), .Y(new_n21686_));
  INVX1    g19250(.A(new_n21686_), .Y(new_n21687_));
  AOI21X1  g19251(.A0(new_n21652_), .A1(pi0647), .B0(pi1157), .Y(new_n21688_));
  OAI21X1  g19252(.A0(new_n21687_), .A1(pi0647), .B0(new_n21688_), .Y(new_n21689_));
  MX2X1    g19253(.A(new_n21686_), .B(new_n21652_), .S0(new_n12705_), .Y(new_n21690_));
  OAI22X1  g19254(.A0(new_n21690_), .A1(new_n14387_), .B0(new_n21689_), .B1(new_n12723_), .Y(new_n21691_));
  AOI21X1  g19255(.A0(new_n21675_), .A1(new_n14385_), .B0(new_n21691_), .Y(new_n21692_));
  AOI21X1  g19256(.A0(new_n21653_), .A1(pi0626), .B0(new_n16352_), .Y(new_n21693_));
  OAI21X1  g19257(.A0(new_n21672_), .A1(pi0626), .B0(new_n21693_), .Y(new_n21694_));
  AOI21X1  g19258(.A0(new_n21653_), .A1(new_n12664_), .B0(new_n16356_), .Y(new_n21695_));
  OAI21X1  g19259(.A0(new_n21672_), .A1(new_n12664_), .B0(new_n21695_), .Y(new_n21696_));
  NAND2X1  g19260(.A(new_n21684_), .B(new_n12769_), .Y(new_n21697_));
  NAND3X1  g19261(.A(new_n21697_), .B(new_n21696_), .C(new_n21694_), .Y(new_n21698_));
  AND2X1   g19262(.A(new_n21698_), .B(pi0788), .Y(new_n21699_));
  INVX1    g19263(.A(new_n21699_), .Y(new_n21700_));
  NOR2X1   g19264(.A(new_n21676_), .B(new_n12120_), .Y(new_n21701_));
  NOR2X1   g19265(.A(new_n21701_), .B(new_n21656_), .Y(new_n21702_));
  INVX1    g19266(.A(new_n21702_), .Y(new_n21703_));
  MX2X1    g19267(.A(new_n21656_), .B(new_n12493_), .S0(new_n21701_), .Y(new_n21704_));
  NOR2X1   g19268(.A(new_n21704_), .B(new_n21681_), .Y(new_n21705_));
  OAI21X1  g19269(.A0(new_n21679_), .A1(new_n12494_), .B0(new_n12584_), .Y(new_n21706_));
  NOR3X1   g19270(.A(new_n21676_), .B(new_n12120_), .C(new_n12493_), .Y(new_n21707_));
  NOR3X1   g19271(.A(new_n21707_), .B(new_n21656_), .C(new_n12494_), .Y(new_n21708_));
  OAI21X1  g19272(.A0(new_n21681_), .A1(new_n21678_), .B0(pi0608), .Y(new_n21709_));
  OAI22X1  g19273(.A0(new_n21709_), .A1(new_n21708_), .B0(new_n21706_), .B1(new_n21705_), .Y(new_n21710_));
  MX2X1    g19274(.A(new_n21710_), .B(new_n21703_), .S0(new_n11889_), .Y(new_n21711_));
  OAI21X1  g19275(.A0(new_n21683_), .A1(new_n12590_), .B0(new_n12591_), .Y(new_n21712_));
  AOI21X1  g19276(.A0(new_n21711_), .A1(new_n12590_), .B0(new_n21712_), .Y(new_n21713_));
  NOR3X1   g19277(.A(new_n21713_), .B(new_n21657_), .C(pi0660), .Y(new_n21714_));
  OAI21X1  g19278(.A0(new_n21683_), .A1(pi0609), .B0(pi1155), .Y(new_n21715_));
  AOI21X1  g19279(.A0(new_n21711_), .A1(pi0609), .B0(new_n21715_), .Y(new_n21716_));
  NOR3X1   g19280(.A(new_n21716_), .B(new_n21658_), .C(new_n12596_), .Y(new_n21717_));
  OAI21X1  g19281(.A0(new_n21717_), .A1(new_n21714_), .B0(pi0785), .Y(new_n21718_));
  NAND2X1  g19282(.A(new_n21711_), .B(new_n11888_), .Y(new_n21719_));
  AND2X1   g19283(.A(new_n21719_), .B(new_n21718_), .Y(new_n21720_));
  NOR3X1   g19284(.A(new_n21683_), .B(new_n12762_), .C(new_n12614_), .Y(new_n21721_));
  NOR2X1   g19285(.A(new_n21721_), .B(pi1154), .Y(new_n21722_));
  OAI21X1  g19286(.A0(new_n21720_), .A1(pi0618), .B0(new_n21722_), .Y(new_n21723_));
  NOR2X1   g19287(.A(new_n21662_), .B(pi0627), .Y(new_n21724_));
  NOR3X1   g19288(.A(new_n21683_), .B(new_n12762_), .C(pi0618), .Y(new_n21725_));
  NOR2X1   g19289(.A(new_n21725_), .B(new_n12615_), .Y(new_n21726_));
  OAI21X1  g19290(.A0(new_n21720_), .A1(new_n12614_), .B0(new_n21726_), .Y(new_n21727_));
  NOR2X1   g19291(.A(new_n21663_), .B(new_n12622_), .Y(new_n21728_));
  AOI22X1  g19292(.A0(new_n21728_), .A1(new_n21727_), .B0(new_n21724_), .B1(new_n21723_), .Y(new_n21729_));
  MX2X1    g19293(.A(new_n21729_), .B(new_n21720_), .S0(new_n11887_), .Y(new_n21730_));
  OR4X1    g19294(.A(new_n21683_), .B(new_n12764_), .C(new_n12762_), .D(new_n12637_), .Y(new_n21731_));
  AND2X1   g19295(.A(new_n21731_), .B(new_n12638_), .Y(new_n21732_));
  OAI21X1  g19296(.A0(new_n21730_), .A1(pi0619), .B0(new_n21732_), .Y(new_n21733_));
  AND2X1   g19297(.A(new_n21668_), .B(new_n12645_), .Y(new_n21734_));
  AND2X1   g19298(.A(new_n21734_), .B(new_n21733_), .Y(new_n21735_));
  NOR4X1   g19299(.A(new_n21683_), .B(new_n12764_), .C(new_n12762_), .D(pi0619), .Y(new_n21736_));
  NOR2X1   g19300(.A(new_n21736_), .B(new_n12638_), .Y(new_n21737_));
  OAI21X1  g19301(.A0(new_n21730_), .A1(new_n12637_), .B0(new_n21737_), .Y(new_n21738_));
  AND2X1   g19302(.A(new_n21670_), .B(pi0648), .Y(new_n21739_));
  AOI21X1  g19303(.A0(new_n21739_), .A1(new_n21738_), .B0(new_n11886_), .Y(new_n21740_));
  INVX1    g19304(.A(new_n21740_), .Y(new_n21741_));
  AOI21X1  g19305(.A0(new_n21730_), .A1(new_n11886_), .B0(new_n14264_), .Y(new_n21742_));
  OAI21X1  g19306(.A0(new_n21741_), .A1(new_n21735_), .B0(new_n21742_), .Y(new_n21743_));
  AOI21X1  g19307(.A0(new_n21743_), .A1(new_n21700_), .B0(new_n14273_), .Y(new_n21744_));
  INVX1    g19308(.A(new_n21674_), .Y(new_n21745_));
  AND2X1   g19309(.A(new_n21684_), .B(new_n12852_), .Y(new_n21746_));
  AOI22X1  g19310(.A0(new_n21746_), .A1(new_n14564_), .B0(new_n21745_), .B1(new_n12867_), .Y(new_n21747_));
  AOI22X1  g19311(.A0(new_n21746_), .A1(new_n14566_), .B0(new_n21745_), .B1(new_n12865_), .Y(new_n21748_));
  MX2X1    g19312(.A(new_n21748_), .B(new_n21747_), .S0(new_n12689_), .Y(new_n21749_));
  OAI21X1  g19313(.A0(new_n21749_), .A1(new_n11884_), .B0(new_n14562_), .Y(new_n21750_));
  OAI22X1  g19314(.A0(new_n21750_), .A1(new_n21744_), .B0(new_n21692_), .B1(new_n11883_), .Y(new_n21751_));
  INVX1    g19315(.A(new_n21751_), .Y(new_n21752_));
  OAI21X1  g19316(.A0(new_n21690_), .A1(new_n12706_), .B0(new_n21689_), .Y(new_n21753_));
  MX2X1    g19317(.A(new_n21753_), .B(new_n21687_), .S0(new_n11883_), .Y(new_n21754_));
  OAI21X1  g19318(.A0(new_n21754_), .A1(pi0644), .B0(pi0715), .Y(new_n21755_));
  AOI21X1  g19319(.A0(new_n21752_), .A1(pi0644), .B0(new_n21755_), .Y(new_n21756_));
  OR4X1    g19320(.A(new_n12734_), .B(new_n2739_), .C(new_n11883_), .D(pi0194), .Y(new_n21757_));
  OAI21X1  g19321(.A0(new_n21675_), .A1(new_n12735_), .B0(new_n21757_), .Y(new_n21758_));
  OAI21X1  g19322(.A0(new_n21653_), .A1(pi0644), .B0(new_n12739_), .Y(new_n21759_));
  AOI21X1  g19323(.A0(new_n21758_), .A1(pi0644), .B0(new_n21759_), .Y(new_n21760_));
  OR2X1    g19324(.A(new_n21760_), .B(new_n11882_), .Y(new_n21761_));
  OAI21X1  g19325(.A0(new_n21754_), .A1(new_n12743_), .B0(new_n12739_), .Y(new_n21762_));
  AOI21X1  g19326(.A0(new_n21752_), .A1(new_n12743_), .B0(new_n21762_), .Y(new_n21763_));
  OAI21X1  g19327(.A0(new_n21653_), .A1(new_n12743_), .B0(pi0715), .Y(new_n21764_));
  AOI21X1  g19328(.A0(new_n21758_), .A1(new_n12743_), .B0(new_n21764_), .Y(new_n21765_));
  OR2X1    g19329(.A(new_n21765_), .B(pi1160), .Y(new_n21766_));
  OAI22X1  g19330(.A0(new_n21766_), .A1(new_n21763_), .B0(new_n21761_), .B1(new_n21756_), .Y(new_n21767_));
  OAI21X1  g19331(.A0(new_n21751_), .A1(pi0790), .B0(pi0832), .Y(new_n21768_));
  AOI21X1  g19332(.A0(new_n21767_), .A1(pi0790), .B0(new_n21768_), .Y(new_n21769_));
  AOI21X1  g19333(.A0(new_n21651_), .A1(new_n21650_), .B0(new_n21769_), .Y(po0351));
  NAND2X1  g19334(.A(pi0299), .B(pi0171), .Y(new_n21771_));
  OAI21X1  g19335(.A0(new_n21771_), .A1(new_n6269_), .B0(new_n8574_), .Y(new_n21772_));
  OAI22X1  g19336(.A0(new_n11831_), .A1(new_n11589_), .B0(new_n11576_), .B1(new_n8571_), .Y(new_n21773_));
  OAI21X1  g19337(.A0(new_n21773_), .A1(new_n21772_), .B0(pi0232), .Y(new_n21774_));
  AOI21X1  g19338(.A0(new_n21774_), .A1(new_n11828_), .B0(new_n2959_), .Y(new_n21775_));
  AOI21X1  g19339(.A0(new_n11596_), .A1(new_n5930_), .B0(new_n10092_), .Y(new_n21776_));
  NOR3X1   g19340(.A(new_n11838_), .B(pi0139), .C(pi0138), .Y(new_n21777_));
  AOI21X1  g19341(.A0(new_n21777_), .A1(new_n11843_), .B0(new_n11842_), .Y(new_n21778_));
  NOR3X1   g19342(.A(new_n21778_), .B(new_n9580_), .C(pi0038), .Y(new_n21779_));
  OAI21X1  g19343(.A0(new_n21776_), .A1(pi0039), .B0(new_n21779_), .Y(new_n21780_));
  OR2X1    g19344(.A(new_n11793_), .B(pi0299), .Y(new_n21781_));
  OR2X1    g19345(.A(new_n21781_), .B(new_n11594_), .Y(new_n21782_));
  OR4X1    g19346(.A(new_n7114_), .B(pi0468), .C(pi0332), .D(new_n3774_), .Y(new_n21783_));
  OAI21X1  g19347(.A0(new_n11579_), .A1(new_n11788_), .B0(new_n21783_), .Y(new_n21784_));
  NOR3X1   g19348(.A(new_n7419_), .B(pi0299), .C(pi0192), .Y(new_n21785_));
  OR2X1    g19349(.A(new_n21785_), .B(new_n5237_), .Y(new_n21786_));
  AOI21X1  g19350(.A0(new_n21784_), .A1(pi0299), .B0(new_n21786_), .Y(new_n21787_));
  NAND2X1  g19351(.A(new_n21787_), .B(new_n21782_), .Y(new_n21788_));
  INVX1    g19352(.A(new_n11808_), .Y(new_n21789_));
  AOI21X1  g19353(.A0(new_n6902_), .A1(new_n3774_), .B0(new_n11809_), .Y(new_n21790_));
  OAI21X1  g19354(.A0(new_n21790_), .A1(new_n6905_), .B0(new_n6895_), .Y(new_n21791_));
  OR4X1    g19355(.A(new_n11814_), .B(new_n6887_), .C(pi0299), .D(new_n11594_), .Y(new_n21792_));
  OR4X1    g19356(.A(new_n11803_), .B(new_n6887_), .C(pi0299), .D(pi0192), .Y(new_n21793_));
  NAND3X1  g19357(.A(new_n21793_), .B(new_n21792_), .C(new_n21791_), .Y(new_n21794_));
  AOI21X1  g19358(.A0(new_n21794_), .A1(pi0232), .B0(new_n21789_), .Y(new_n21795_));
  OAI21X1  g19359(.A0(new_n21795_), .A1(new_n2959_), .B0(new_n3277_), .Y(new_n21796_));
  AOI21X1  g19360(.A0(new_n21788_), .A1(new_n11792_), .B0(new_n21796_), .Y(new_n21797_));
  OAI21X1  g19361(.A0(new_n21797_), .A1(pi0087), .B0(new_n11786_), .Y(new_n21798_));
  AOI21X1  g19362(.A0(new_n21798_), .A1(new_n3100_), .B0(new_n11784_), .Y(new_n21799_));
  OAI21X1  g19363(.A0(new_n21799_), .A1(pi0055), .B0(new_n11823_), .Y(new_n21800_));
  AND2X1   g19364(.A(new_n21800_), .B(new_n3148_), .Y(new_n21801_));
  NAND2X1  g19365(.A(new_n21778_), .B(new_n7369_), .Y(new_n21802_));
  OAI22X1  g19366(.A0(new_n21802_), .A1(new_n21801_), .B0(new_n21780_), .B1(new_n21775_), .Y(po0352));
  OAI21X1  g19367(.A0(new_n7474_), .A1(pi0170), .B0(new_n11810_), .Y(new_n21804_));
  AOI21X1  g19368(.A0(new_n21804_), .A1(new_n6893_), .B0(new_n6922_), .Y(new_n21805_));
  OAI21X1  g19369(.A0(new_n21805_), .A1(new_n11804_), .B0(pi0232), .Y(new_n21806_));
  AND2X1   g19370(.A(new_n21806_), .B(new_n11808_), .Y(new_n21807_));
  OR4X1    g19371(.A(new_n11814_), .B(new_n6887_), .C(pi0299), .D(new_n5237_), .Y(new_n21808_));
  AND2X1   g19372(.A(new_n21808_), .B(new_n21807_), .Y(new_n21809_));
  AND2X1   g19373(.A(pi0194), .B(new_n2996_), .Y(new_n21810_));
  OAI21X1  g19374(.A0(new_n21809_), .A1(new_n2959_), .B0(new_n21810_), .Y(new_n21811_));
  NOR2X1   g19375(.A(pi0194), .B(pi0038), .Y(new_n21812_));
  OAI21X1  g19376(.A0(new_n21807_), .A1(new_n2959_), .B0(new_n21812_), .Y(new_n21813_));
  AND2X1   g19377(.A(new_n21813_), .B(new_n21811_), .Y(new_n21814_));
  INVX1    g19378(.A(new_n21811_), .Y(new_n21815_));
  NOR2X1   g19379(.A(new_n21813_), .B(new_n11790_), .Y(new_n21816_));
  AOI21X1  g19380(.A0(new_n21815_), .A1(new_n21781_), .B0(new_n21816_), .Y(new_n21817_));
  AOI22X1  g19381(.A0(new_n11706_), .A1(new_n11850_), .B0(new_n11795_), .B1(pi0170), .Y(new_n21818_));
  OAI21X1  g19382(.A0(new_n21818_), .A1(new_n2953_), .B0(pi0232), .Y(new_n21819_));
  OAI22X1  g19383(.A0(new_n21819_), .A1(new_n21817_), .B0(new_n21814_), .B1(new_n11792_), .Y(new_n21820_));
  AOI21X1  g19384(.A0(new_n21820_), .A1(new_n3026_), .B0(pi0087), .Y(new_n21821_));
  OAI21X1  g19385(.A0(new_n21821_), .A1(new_n11787_), .B0(new_n3100_), .Y(new_n21822_));
  AOI21X1  g19386(.A0(new_n21822_), .A1(new_n11785_), .B0(pi0055), .Y(new_n21823_));
  OAI21X1  g19387(.A0(new_n21823_), .A1(new_n11824_), .B0(new_n3148_), .Y(new_n21824_));
  AOI21X1  g19388(.A0(new_n21824_), .A1(new_n7369_), .B0(new_n11843_), .Y(new_n21825_));
  AOI21X1  g19389(.A0(new_n7237_), .A1(new_n3917_), .B0(new_n11830_), .Y(new_n21826_));
  NOR4X1   g19390(.A(new_n21826_), .B(new_n7713_), .C(new_n2437_), .D(new_n2438_), .Y(new_n21827_));
  AND2X1   g19391(.A(new_n11830_), .B(new_n9592_), .Y(new_n21828_));
  NOR3X1   g19392(.A(new_n21828_), .B(new_n21827_), .C(new_n5237_), .Y(new_n21829_));
  AOI21X1  g19393(.A0(new_n8575_), .A1(new_n5237_), .B0(new_n21829_), .Y(new_n21830_));
  MX2X1    g19394(.A(new_n21830_), .B(new_n8571_), .S0(new_n2953_), .Y(new_n21831_));
  OR4X1    g19395(.A(new_n11644_), .B(new_n7291_), .C(new_n2900_), .D(pi0095), .Y(new_n21832_));
  AOI21X1  g19396(.A0(new_n21832_), .A1(new_n2959_), .B0(pi0038), .Y(new_n21833_));
  OAI21X1  g19397(.A0(new_n21831_), .A1(new_n2959_), .B0(new_n21833_), .Y(new_n21834_));
  NOR2X1   g19398(.A(new_n21830_), .B(new_n2959_), .Y(new_n21835_));
  AOI21X1  g19399(.A0(new_n11679_), .A1(new_n10091_), .B0(pi0039), .Y(new_n21836_));
  NOR3X1   g19400(.A(new_n21836_), .B(new_n21835_), .C(pi0038), .Y(new_n21837_));
  OAI21X1  g19401(.A0(new_n21837_), .A1(new_n11641_), .B0(new_n7686_), .Y(new_n21838_));
  AOI21X1  g19402(.A0(new_n21834_), .A1(new_n11641_), .B0(new_n21838_), .Y(new_n21839_));
  OAI22X1  g19403(.A0(new_n21839_), .A1(pi0196), .B0(new_n11840_), .B1(pi0138), .Y(new_n21840_));
  AND2X1   g19404(.A(new_n11843_), .B(pi0195), .Y(new_n21841_));
  INVX1    g19405(.A(new_n21841_), .Y(new_n21842_));
  AOI21X1  g19406(.A0(new_n21824_), .A1(new_n7369_), .B0(new_n21842_), .Y(new_n21843_));
  OAI21X1  g19407(.A0(new_n21841_), .A1(new_n21839_), .B0(new_n21777_), .Y(new_n21844_));
  OAI22X1  g19408(.A0(new_n21844_), .A1(new_n21843_), .B0(new_n21840_), .B1(new_n21825_), .Y(po0353));
  AND2X1   g19409(.A(pi0947), .B(new_n14336_), .Y(new_n21846_));
  INVX1    g19410(.A(new_n21846_), .Y(new_n21847_));
  OAI21X1  g19411(.A0(new_n14638_), .A1(pi0698), .B0(new_n21847_), .Y(new_n21848_));
  OAI21X1  g19412(.A0(new_n2739_), .A1(pi0197), .B0(pi0832), .Y(new_n21849_));
  AOI21X1  g19413(.A0(new_n21848_), .A1(new_n2739_), .B0(new_n21849_), .Y(new_n21850_));
  AOI21X1  g19414(.A0(new_n21847_), .A1(new_n12202_), .B0(new_n2996_), .Y(new_n21851_));
  OAI21X1  g19415(.A0(new_n12572_), .A1(new_n7347_), .B0(new_n21851_), .Y(new_n21852_));
  OAI21X1  g19416(.A0(new_n14760_), .A1(new_n7347_), .B0(pi0299), .Y(new_n21853_));
  AOI21X1  g19417(.A0(new_n14759_), .A1(new_n7347_), .B0(new_n21853_), .Y(new_n21854_));
  NOR2X1   g19418(.A(new_n14740_), .B(pi0197), .Y(new_n21855_));
  OAI21X1  g19419(.A0(new_n21855_), .A1(new_n14664_), .B0(new_n14336_), .Y(new_n21856_));
  AND2X1   g19420(.A(pi0767), .B(new_n7347_), .Y(new_n21857_));
  AOI21X1  g19421(.A0(new_n21857_), .A1(new_n12089_), .B0(new_n2959_), .Y(new_n21858_));
  OAI21X1  g19422(.A0(new_n21856_), .A1(new_n21854_), .B0(new_n21858_), .Y(new_n21859_));
  AOI21X1  g19423(.A0(new_n21846_), .A1(new_n11947_), .B0(pi0039), .Y(new_n21860_));
  OAI21X1  g19424(.A0(new_n11947_), .A1(pi0197), .B0(new_n21860_), .Y(new_n21861_));
  NAND3X1  g19425(.A(new_n21861_), .B(new_n21859_), .C(new_n2996_), .Y(new_n21862_));
  AOI21X1  g19426(.A0(new_n21862_), .A1(new_n21852_), .B0(new_n14306_), .Y(new_n21863_));
  OAI21X1  g19427(.A0(new_n14703_), .A1(new_n7347_), .B0(new_n14336_), .Y(new_n21864_));
  AOI21X1  g19428(.A0(new_n14693_), .A1(new_n7347_), .B0(new_n21864_), .Y(new_n21865_));
  NAND3X1  g19429(.A(new_n14722_), .B(new_n14718_), .C(pi0197), .Y(new_n21866_));
  NAND2X1  g19430(.A(new_n21866_), .B(pi0299), .Y(new_n21867_));
  AOI21X1  g19431(.A0(new_n14712_), .A1(new_n7347_), .B0(new_n21867_), .Y(new_n21868_));
  NOR3X1   g19432(.A(new_n21855_), .B(new_n14724_), .C(pi0299), .Y(new_n21869_));
  OR2X1    g19433(.A(new_n21869_), .B(new_n14336_), .Y(new_n21870_));
  OAI21X1  g19434(.A0(new_n21870_), .A1(new_n21868_), .B0(pi0039), .Y(new_n21871_));
  OAI22X1  g19435(.A0(new_n21871_), .A1(new_n21865_), .B0(new_n21861_), .B1(new_n14727_), .Y(new_n21872_));
  NOR2X1   g19436(.A(new_n12202_), .B(pi0197), .Y(new_n21873_));
  OAI21X1  g19437(.A0(new_n14590_), .A1(new_n14336_), .B0(new_n2959_), .Y(new_n21874_));
  OAI21X1  g19438(.A0(new_n21874_), .A1(new_n14811_), .B0(pi0038), .Y(new_n21875_));
  OAI21X1  g19439(.A0(new_n21875_), .A1(new_n21873_), .B0(new_n14306_), .Y(new_n21876_));
  AOI21X1  g19440(.A0(new_n21872_), .A1(new_n2996_), .B0(new_n21876_), .Y(new_n21877_));
  OAI21X1  g19441(.A0(new_n21877_), .A1(new_n21863_), .B0(new_n7686_), .Y(new_n21878_));
  AOI21X1  g19442(.A0(new_n9580_), .A1(new_n7347_), .B0(pi0832), .Y(new_n21879_));
  AOI21X1  g19443(.A0(new_n21879_), .A1(new_n21878_), .B0(new_n21850_), .Y(po0354));
  INVX1    g19444(.A(new_n13403_), .Y(new_n21881_));
  AOI21X1  g19445(.A0(new_n11948_), .A1(new_n3065_), .B0(new_n21881_), .Y(new_n21882_));
  INVX1    g19446(.A(new_n12106_), .Y(new_n21883_));
  NAND3X1  g19447(.A(new_n21883_), .B(new_n5071_), .C(pi0198), .Y(new_n21884_));
  AND2X1   g19448(.A(new_n11953_), .B(pi0198), .Y(new_n21885_));
  NOR2X1   g19449(.A(new_n12029_), .B(new_n2973_), .Y(new_n21886_));
  MX2X1    g19450(.A(new_n21886_), .B(new_n21885_), .S0(new_n5031_), .Y(new_n21887_));
  AOI21X1  g19451(.A0(new_n21887_), .A1(new_n5070_), .B0(new_n10136_), .Y(new_n21888_));
  INVX1    g19452(.A(new_n21885_), .Y(new_n21889_));
  AOI21X1  g19453(.A0(new_n21889_), .A1(new_n10136_), .B0(pi0215), .Y(new_n21890_));
  INVX1    g19454(.A(new_n21890_), .Y(new_n21891_));
  AOI21X1  g19455(.A0(new_n21888_), .A1(new_n21884_), .B0(new_n21891_), .Y(new_n21892_));
  AOI21X1  g19456(.A0(new_n11953_), .A1(pi0198), .B0(po1101), .Y(new_n21893_));
  NOR3X1   g19457(.A(new_n21893_), .B(new_n12135_), .C(new_n2973_), .Y(new_n21894_));
  OR2X1    g19458(.A(new_n11966_), .B(new_n5028_), .Y(new_n21895_));
  AOI21X1  g19459(.A0(new_n12144_), .A1(new_n5028_), .B0(new_n2973_), .Y(new_n21896_));
  AND2X1   g19460(.A(new_n21896_), .B(new_n21895_), .Y(new_n21897_));
  AOI21X1  g19461(.A0(new_n21897_), .A1(new_n5071_), .B0(new_n21894_), .Y(new_n21898_));
  OAI21X1  g19462(.A0(new_n21898_), .A1(new_n2954_), .B0(pi0299), .Y(new_n21899_));
  NOR2X1   g19463(.A(new_n21899_), .B(new_n21892_), .Y(new_n21900_));
  NOR3X1   g19464(.A(new_n12106_), .B(new_n5050_), .C(new_n2973_), .Y(new_n21901_));
  INVX1    g19465(.A(new_n21901_), .Y(new_n21902_));
  AOI21X1  g19466(.A0(new_n21887_), .A1(new_n5050_), .B0(new_n2970_), .Y(new_n21903_));
  AOI21X1  g19467(.A0(new_n21889_), .A1(new_n2970_), .B0(pi0223), .Y(new_n21904_));
  INVX1    g19468(.A(new_n21904_), .Y(new_n21905_));
  AOI21X1  g19469(.A0(new_n21903_), .A1(new_n21902_), .B0(new_n21905_), .Y(new_n21906_));
  AOI21X1  g19470(.A0(new_n21897_), .A1(new_n5051_), .B0(new_n21894_), .Y(new_n21907_));
  OAI21X1  g19471(.A0(new_n21907_), .A1(new_n2964_), .B0(new_n2953_), .Y(new_n21908_));
  AND2X1   g19472(.A(new_n8244_), .B(new_n3129_), .Y(new_n21909_));
  OAI21X1  g19473(.A0(new_n21908_), .A1(new_n21906_), .B0(new_n21909_), .Y(new_n21910_));
  OAI22X1  g19474(.A0(new_n21910_), .A1(new_n21900_), .B0(new_n21882_), .B1(new_n2973_), .Y(new_n21911_));
  INVX1    g19475(.A(new_n21911_), .Y(new_n21912_));
  AOI21X1  g19476(.A0(new_n11942_), .A1(new_n11929_), .B0(new_n2973_), .Y(new_n21913_));
  NAND2X1  g19477(.A(pi0633), .B(pi0603), .Y(new_n21914_));
  MX2X1    g19478(.A(new_n12166_), .B(new_n12096_), .S0(pi0198), .Y(new_n21915_));
  MX2X1    g19479(.A(new_n21915_), .B(new_n21913_), .S0(new_n21914_), .Y(new_n21916_));
  INVX1    g19480(.A(pi0633), .Y(new_n21917_));
  AOI21X1  g19481(.A0(new_n12095_), .A1(pi0198), .B0(new_n12100_), .Y(new_n21918_));
  OAI21X1  g19482(.A0(new_n21918_), .A1(new_n21917_), .B0(new_n11945_), .Y(new_n21919_));
  OAI21X1  g19483(.A0(new_n12102_), .A1(pi0603), .B0(new_n21919_), .Y(new_n21920_));
  OAI21X1  g19484(.A0(new_n21920_), .A1(pi0299), .B0(new_n2959_), .Y(new_n21921_));
  AOI21X1  g19485(.A0(new_n21916_), .A1(pi0299), .B0(new_n21921_), .Y(new_n21922_));
  NOR4X1   g19486(.A(new_n12108_), .B(new_n11952_), .C(new_n2740_), .D(new_n21917_), .Y(new_n21923_));
  AOI22X1  g19487(.A0(new_n21923_), .A1(pi0603), .B0(new_n11953_), .B1(pi0198), .Y(new_n21924_));
  AND2X1   g19488(.A(new_n21885_), .B(new_n5027_), .Y(new_n21925_));
  AOI21X1  g19489(.A0(new_n11953_), .A1(pi0198), .B0(new_n21923_), .Y(new_n21926_));
  NOR2X1   g19490(.A(new_n21926_), .B(new_n5057_), .Y(new_n21927_));
  INVX1    g19491(.A(new_n21927_), .Y(new_n21928_));
  NOR2X1   g19492(.A(new_n12135_), .B(new_n2973_), .Y(new_n21929_));
  AOI21X1  g19493(.A0(new_n21923_), .A1(new_n12144_), .B0(new_n21929_), .Y(new_n21930_));
  AOI21X1  g19494(.A0(new_n21930_), .A1(new_n21928_), .B0(new_n5027_), .Y(new_n21931_));
  NOR3X1   g19495(.A(new_n21931_), .B(new_n21925_), .C(new_n12127_), .Y(new_n21932_));
  AOI21X1  g19496(.A0(new_n21924_), .A1(new_n12127_), .B0(new_n21932_), .Y(new_n21933_));
  OR2X1    g19497(.A(new_n21931_), .B(new_n21929_), .Y(new_n21934_));
  MX2X1    g19498(.A(new_n21934_), .B(new_n21933_), .S0(new_n5282_), .Y(new_n21935_));
  AND2X1   g19499(.A(new_n12172_), .B(new_n12145_), .Y(new_n21936_));
  AND2X1   g19500(.A(new_n12184_), .B(new_n21936_), .Y(new_n21937_));
  AOI21X1  g19501(.A0(new_n21937_), .A1(pi0633), .B0(new_n21897_), .Y(new_n21938_));
  NOR2X1   g19502(.A(new_n21938_), .B(new_n5030_), .Y(new_n21939_));
  MX2X1    g19503(.A(new_n21923_), .B(pi0198), .S0(new_n11965_), .Y(new_n21940_));
  AOI21X1  g19504(.A0(new_n21940_), .A1(new_n12150_), .B0(new_n21939_), .Y(new_n21941_));
  AOI21X1  g19505(.A0(new_n21941_), .A1(new_n5051_), .B0(new_n2964_), .Y(new_n21942_));
  OAI21X1  g19506(.A0(new_n21935_), .A1(new_n5051_), .B0(new_n21942_), .Y(new_n21943_));
  INVX1    g19507(.A(new_n12116_), .Y(new_n21944_));
  NOR2X1   g19508(.A(new_n12028_), .B(new_n2973_), .Y(new_n21945_));
  AOI21X1  g19509(.A0(new_n21944_), .A1(pi0633), .B0(new_n21945_), .Y(new_n21946_));
  MX2X1    g19510(.A(new_n21946_), .B(new_n21926_), .S0(new_n5033_), .Y(new_n21947_));
  OR2X1    g19511(.A(new_n21947_), .B(new_n5027_), .Y(new_n21948_));
  NOR2X1   g19512(.A(new_n21926_), .B(new_n5027_), .Y(new_n21949_));
  OAI21X1  g19513(.A0(new_n21949_), .A1(new_n11968_), .B0(new_n12323_), .Y(new_n21950_));
  AOI21X1  g19514(.A0(new_n21948_), .A1(new_n11968_), .B0(new_n21950_), .Y(new_n21951_));
  NOR3X1   g19515(.A(new_n21926_), .B(new_n12323_), .C(new_n5027_), .Y(new_n21952_));
  OR2X1    g19516(.A(new_n21952_), .B(new_n21925_), .Y(new_n21953_));
  NOR2X1   g19517(.A(new_n21953_), .B(new_n21951_), .Y(new_n21954_));
  AOI21X1  g19518(.A0(new_n21886_), .A1(new_n5027_), .B0(new_n5282_), .Y(new_n21955_));
  AOI22X1  g19519(.A0(new_n21955_), .A1(new_n21948_), .B0(new_n21954_), .B1(new_n5282_), .Y(new_n21956_));
  AND2X1   g19520(.A(new_n21956_), .B(new_n5050_), .Y(new_n21957_));
  NOR2X1   g19521(.A(new_n21946_), .B(new_n5027_), .Y(new_n21958_));
  NOR3X1   g19522(.A(new_n21946_), .B(new_n12127_), .C(new_n5027_), .Y(new_n21959_));
  NOR2X1   g19523(.A(new_n12125_), .B(new_n5027_), .Y(new_n21960_));
  INVX1    g19524(.A(new_n21960_), .Y(new_n21961_));
  AOI21X1  g19525(.A0(new_n21926_), .A1(new_n5057_), .B0(new_n21961_), .Y(new_n21962_));
  INVX1    g19526(.A(new_n21962_), .Y(new_n21963_));
  AOI21X1  g19527(.A0(new_n21946_), .A1(new_n5033_), .B0(new_n21963_), .Y(new_n21964_));
  NOR3X1   g19528(.A(new_n12056_), .B(pi0603), .C(new_n2973_), .Y(new_n21965_));
  OR4X1    g19529(.A(new_n21965_), .B(new_n21964_), .C(new_n21959_), .D(new_n5030_), .Y(new_n21966_));
  OAI21X1  g19530(.A0(new_n12028_), .A1(new_n2973_), .B0(new_n5030_), .Y(new_n21967_));
  OAI21X1  g19531(.A0(new_n21967_), .A1(new_n21958_), .B0(new_n21966_), .Y(new_n21968_));
  OAI21X1  g19532(.A0(new_n21968_), .A1(new_n5050_), .B0(new_n2971_), .Y(new_n21969_));
  AOI21X1  g19533(.A0(new_n21924_), .A1(new_n2970_), .B0(pi0223), .Y(new_n21970_));
  OAI21X1  g19534(.A0(new_n21969_), .A1(new_n21957_), .B0(new_n21970_), .Y(new_n21971_));
  AOI21X1  g19535(.A0(new_n21971_), .A1(new_n21943_), .B0(pi0299), .Y(new_n21972_));
  AOI21X1  g19536(.A0(new_n21941_), .A1(new_n5071_), .B0(new_n2954_), .Y(new_n21973_));
  OAI21X1  g19537(.A0(new_n21935_), .A1(new_n5071_), .B0(new_n21973_), .Y(new_n21974_));
  AND2X1   g19538(.A(new_n21956_), .B(new_n5070_), .Y(new_n21975_));
  OAI21X1  g19539(.A0(new_n21968_), .A1(new_n5070_), .B0(new_n10137_), .Y(new_n21976_));
  AOI21X1  g19540(.A0(new_n21924_), .A1(new_n10136_), .B0(pi0215), .Y(new_n21977_));
  OAI21X1  g19541(.A0(new_n21976_), .A1(new_n21975_), .B0(new_n21977_), .Y(new_n21978_));
  AOI21X1  g19542(.A0(new_n21978_), .A1(new_n21974_), .B0(new_n2953_), .Y(new_n21979_));
  NOR3X1   g19543(.A(new_n21979_), .B(new_n21972_), .C(new_n2959_), .Y(new_n21980_));
  OAI21X1  g19544(.A0(new_n21980_), .A1(new_n21922_), .B0(new_n2996_), .Y(new_n21981_));
  AOI21X1  g19545(.A0(pi0198), .A1(pi0039), .B0(new_n2996_), .Y(new_n21982_));
  INVX1    g19546(.A(new_n21982_), .Y(new_n21983_));
  NOR3X1   g19547(.A(new_n12108_), .B(new_n21917_), .C(new_n5027_), .Y(new_n21984_));
  MX2X1    g19548(.A(pi0198), .B(new_n21984_), .S0(new_n11961_), .Y(new_n21985_));
  AOI21X1  g19549(.A0(new_n21985_), .A1(new_n2959_), .B0(new_n21983_), .Y(new_n21986_));
  NOR2X1   g19550(.A(new_n21986_), .B(new_n3810_), .Y(new_n21987_));
  AOI22X1  g19551(.A0(new_n21987_), .A1(new_n21981_), .B0(new_n3810_), .B1(pi0198), .Y(new_n21988_));
  MX2X1    g19552(.A(new_n21988_), .B(new_n21912_), .S0(new_n12601_), .Y(new_n21989_));
  NOR2X1   g19553(.A(new_n21988_), .B(new_n12601_), .Y(new_n21990_));
  AOI22X1  g19554(.A0(new_n21990_), .A1(pi0609), .B0(new_n21911_), .B1(new_n13430_), .Y(new_n21991_));
  AOI22X1  g19555(.A0(new_n21990_), .A1(new_n12590_), .B0(new_n21911_), .B1(new_n13436_), .Y(new_n21992_));
  MX2X1    g19556(.A(new_n21992_), .B(new_n21991_), .S0(pi1155), .Y(new_n21993_));
  MX2X1    g19557(.A(new_n21993_), .B(new_n21989_), .S0(new_n11888_), .Y(new_n21994_));
  OAI21X1  g19558(.A0(new_n21911_), .A1(pi0618), .B0(pi1154), .Y(new_n21995_));
  AOI21X1  g19559(.A0(new_n21994_), .A1(pi0618), .B0(new_n21995_), .Y(new_n21996_));
  OAI21X1  g19560(.A0(new_n21911_), .A1(new_n12614_), .B0(new_n12615_), .Y(new_n21997_));
  AOI21X1  g19561(.A0(new_n21994_), .A1(new_n12614_), .B0(new_n21997_), .Y(new_n21998_));
  OAI21X1  g19562(.A0(new_n21998_), .A1(new_n21996_), .B0(pi0781), .Y(new_n21999_));
  OAI21X1  g19563(.A0(new_n21994_), .A1(pi0781), .B0(new_n21999_), .Y(new_n22000_));
  AOI21X1  g19564(.A0(new_n21912_), .A1(new_n12637_), .B0(new_n12638_), .Y(new_n22001_));
  OAI21X1  g19565(.A0(new_n22000_), .A1(new_n12637_), .B0(new_n22001_), .Y(new_n22002_));
  AOI21X1  g19566(.A0(new_n21912_), .A1(pi0619), .B0(pi1159), .Y(new_n22003_));
  OAI21X1  g19567(.A0(new_n22000_), .A1(pi0619), .B0(new_n22003_), .Y(new_n22004_));
  AOI21X1  g19568(.A0(new_n22004_), .A1(new_n22002_), .B0(new_n11886_), .Y(new_n22005_));
  AOI21X1  g19569(.A0(new_n22000_), .A1(new_n11886_), .B0(new_n22005_), .Y(new_n22006_));
  MX2X1    g19570(.A(new_n22006_), .B(new_n21912_), .S0(new_n12841_), .Y(new_n22007_));
  MX2X1    g19571(.A(new_n22007_), .B(new_n21912_), .S0(new_n12711_), .Y(new_n22008_));
  NOR2X1   g19572(.A(new_n12691_), .B(new_n12659_), .Y(new_n22009_));
  INVX1    g19573(.A(new_n22009_), .Y(new_n22010_));
  INVX1    g19574(.A(new_n12659_), .Y(new_n22011_));
  AOI22X1  g19575(.A0(new_n12292_), .A1(pi0634), .B0(new_n11953_), .B1(pi0198), .Y(new_n22012_));
  AOI21X1  g19576(.A0(new_n22012_), .A1(new_n5367_), .B0(new_n12235_), .Y(new_n22013_));
  INVX1    g19577(.A(new_n22012_), .Y(new_n22014_));
  NAND2X1  g19578(.A(new_n12293_), .B(new_n12028_), .Y(new_n22015_));
  INVX1    g19579(.A(new_n22015_), .Y(new_n22016_));
  AOI21X1  g19580(.A0(new_n22016_), .A1(pi0634), .B0(new_n21945_), .Y(new_n22017_));
  INVX1    g19581(.A(new_n22017_), .Y(new_n22018_));
  MX2X1    g19582(.A(new_n22018_), .B(new_n22014_), .S0(new_n5033_), .Y(new_n22019_));
  OAI21X1  g19583(.A0(new_n22019_), .A1(new_n5367_), .B0(new_n22013_), .Y(new_n22020_));
  OAI21X1  g19584(.A0(new_n12029_), .A1(new_n2973_), .B0(new_n5028_), .Y(new_n22021_));
  AOI21X1  g19585(.A0(new_n21889_), .A1(new_n5367_), .B0(pi0680), .Y(new_n22022_));
  AOI22X1  g19586(.A0(new_n22022_), .A1(new_n22021_), .B0(new_n22019_), .B1(new_n5030_), .Y(new_n22023_));
  AOI21X1  g19587(.A0(new_n22023_), .A1(new_n22020_), .B0(new_n5051_), .Y(new_n22024_));
  MX2X1    g19588(.A(new_n22017_), .B(new_n22012_), .S0(new_n5057_), .Y(new_n22025_));
  OAI21X1  g19589(.A0(new_n22018_), .A1(new_n5367_), .B0(new_n12209_), .Y(new_n22026_));
  AOI21X1  g19590(.A0(new_n22025_), .A1(new_n5367_), .B0(new_n22026_), .Y(new_n22027_));
  NAND3X1  g19591(.A(new_n12260_), .B(new_n5029_), .C(pi0198), .Y(new_n22028_));
  OAI21X1  g19592(.A0(new_n22017_), .A1(new_n5282_), .B0(new_n22028_), .Y(new_n22029_));
  OR2X1    g19593(.A(new_n22029_), .B(new_n22027_), .Y(new_n22030_));
  AND2X1   g19594(.A(new_n22030_), .B(new_n5051_), .Y(new_n22031_));
  NOR3X1   g19595(.A(new_n22031_), .B(new_n22024_), .C(new_n2970_), .Y(new_n22032_));
  OAI21X1  g19596(.A0(new_n21885_), .A1(new_n12292_), .B0(pi0634), .Y(new_n22033_));
  OAI21X1  g19597(.A0(new_n22033_), .A1(new_n5029_), .B0(new_n21889_), .Y(new_n22034_));
  OAI21X1  g19598(.A0(new_n22034_), .A1(new_n2971_), .B0(new_n2964_), .Y(new_n22035_));
  NAND2X1  g19599(.A(new_n11965_), .B(pi0198), .Y(new_n22036_));
  NAND3X1  g19600(.A(new_n12292_), .B(new_n12144_), .C(pi0634), .Y(new_n22037_));
  AND2X1   g19601(.A(new_n22037_), .B(new_n22036_), .Y(new_n22038_));
  INVX1    g19602(.A(new_n22038_), .Y(new_n22039_));
  MX2X1    g19603(.A(new_n22039_), .B(new_n22014_), .S0(new_n5057_), .Y(new_n22040_));
  AOI21X1  g19604(.A0(new_n22038_), .A1(new_n5028_), .B0(new_n12235_), .Y(new_n22041_));
  OAI21X1  g19605(.A0(new_n22040_), .A1(new_n5028_), .B0(new_n22041_), .Y(new_n22042_));
  AOI22X1  g19606(.A0(new_n22039_), .A1(new_n5030_), .B0(new_n21897_), .B1(new_n5029_), .Y(new_n22043_));
  NAND3X1  g19607(.A(new_n22043_), .B(new_n22042_), .C(new_n5051_), .Y(new_n22044_));
  MX2X1    g19608(.A(new_n22038_), .B(new_n22012_), .S0(new_n5033_), .Y(new_n22045_));
  NAND2X1  g19609(.A(new_n22045_), .B(new_n5028_), .Y(new_n22046_));
  NAND4X1  g19610(.A(new_n21896_), .B(new_n21895_), .C(new_n21929_), .D(new_n5029_), .Y(new_n22047_));
  OAI21X1  g19611(.A0(new_n22045_), .A1(new_n5282_), .B0(new_n22047_), .Y(new_n22048_));
  AOI21X1  g19612(.A0(new_n22046_), .A1(new_n22013_), .B0(new_n22048_), .Y(new_n22049_));
  AOI21X1  g19613(.A0(new_n22049_), .A1(new_n5050_), .B0(new_n2964_), .Y(new_n22050_));
  AOI21X1  g19614(.A0(new_n22050_), .A1(new_n22044_), .B0(pi0299), .Y(new_n22051_));
  OAI21X1  g19615(.A0(new_n22035_), .A1(new_n22032_), .B0(new_n22051_), .Y(new_n22052_));
  AND2X1   g19616(.A(new_n22030_), .B(new_n5071_), .Y(new_n22053_));
  AOI21X1  g19617(.A0(new_n22023_), .A1(new_n22020_), .B0(new_n5071_), .Y(new_n22054_));
  NOR3X1   g19618(.A(new_n22054_), .B(new_n22053_), .C(new_n10136_), .Y(new_n22055_));
  OAI21X1  g19619(.A0(new_n22034_), .A1(new_n10137_), .B0(new_n2954_), .Y(new_n22056_));
  NAND3X1  g19620(.A(new_n22043_), .B(new_n22042_), .C(new_n5071_), .Y(new_n22057_));
  AOI21X1  g19621(.A0(new_n22049_), .A1(new_n5070_), .B0(new_n2954_), .Y(new_n22058_));
  AOI21X1  g19622(.A0(new_n22058_), .A1(new_n22057_), .B0(new_n2953_), .Y(new_n22059_));
  OAI21X1  g19623(.A0(new_n22056_), .A1(new_n22055_), .B0(new_n22059_), .Y(new_n22060_));
  AOI21X1  g19624(.A0(new_n22060_), .A1(new_n22052_), .B0(new_n2959_), .Y(new_n22061_));
  NAND2X1  g19625(.A(pi0680), .B(pi0634), .Y(new_n22062_));
  MX2X1    g19626(.A(new_n12463_), .B(new_n12451_), .S0(pi0198), .Y(new_n22063_));
  MX2X1    g19627(.A(new_n22063_), .B(new_n21913_), .S0(new_n22062_), .Y(new_n22064_));
  INVX1    g19628(.A(new_n11945_), .Y(new_n22065_));
  NAND3X1  g19629(.A(new_n12456_), .B(pi0680), .C(pi0634), .Y(new_n22066_));
  AOI21X1  g19630(.A0(new_n13227_), .A1(pi0198), .B0(new_n22066_), .Y(new_n22067_));
  OAI21X1  g19631(.A0(new_n22067_), .A1(new_n22065_), .B0(new_n2953_), .Y(new_n22068_));
  NAND2X1  g19632(.A(new_n22068_), .B(new_n2959_), .Y(new_n22069_));
  AOI21X1  g19633(.A0(new_n22064_), .A1(pi0299), .B0(new_n22069_), .Y(new_n22070_));
  OAI21X1  g19634(.A0(new_n22070_), .A1(new_n22061_), .B0(new_n2996_), .Y(new_n22071_));
  INVX1    g19635(.A(pi0634), .Y(new_n22072_));
  NOR3X1   g19636(.A(new_n12210_), .B(new_n5029_), .C(new_n22072_), .Y(new_n22073_));
  MX2X1    g19637(.A(pi0198), .B(new_n22073_), .S0(new_n11961_), .Y(new_n22074_));
  AOI21X1  g19638(.A0(new_n22074_), .A1(new_n2959_), .B0(new_n21983_), .Y(new_n22075_));
  NOR2X1   g19639(.A(new_n22075_), .B(new_n3810_), .Y(new_n22076_));
  AOI22X1  g19640(.A0(new_n22076_), .A1(new_n22071_), .B0(new_n3810_), .B1(pi0198), .Y(new_n22077_));
  OAI21X1  g19641(.A0(new_n21911_), .A1(pi0625), .B0(pi1153), .Y(new_n22078_));
  AOI21X1  g19642(.A0(new_n22077_), .A1(pi0625), .B0(new_n22078_), .Y(new_n22079_));
  OAI21X1  g19643(.A0(new_n21911_), .A1(new_n12493_), .B0(new_n12494_), .Y(new_n22080_));
  AOI21X1  g19644(.A0(new_n22077_), .A1(new_n12493_), .B0(new_n22080_), .Y(new_n22081_));
  NOR2X1   g19645(.A(new_n22081_), .B(new_n22079_), .Y(new_n22082_));
  MX2X1    g19646(.A(new_n22082_), .B(new_n22077_), .S0(new_n11889_), .Y(new_n22083_));
  INVX1    g19647(.A(new_n22083_), .Y(new_n22084_));
  MX2X1    g19648(.A(new_n22084_), .B(new_n21911_), .S0(new_n12618_), .Y(new_n22085_));
  INVX1    g19649(.A(new_n22085_), .Y(new_n22086_));
  MX2X1    g19650(.A(new_n22086_), .B(new_n21912_), .S0(new_n12641_), .Y(new_n22087_));
  AND2X1   g19651(.A(new_n22087_), .B(new_n22011_), .Y(new_n22088_));
  AOI22X1  g19652(.A0(new_n22088_), .A1(new_n17252_), .B0(new_n21912_), .B1(new_n22010_), .Y(new_n22089_));
  MX2X1    g19653(.A(new_n22089_), .B(new_n21911_), .S0(new_n12683_), .Y(new_n22090_));
  INVX1    g19654(.A(new_n22090_), .Y(new_n22091_));
  AOI21X1  g19655(.A0(new_n21912_), .A1(pi0628), .B0(pi1156), .Y(new_n22092_));
  OAI21X1  g19656(.A0(new_n22089_), .A1(pi0628), .B0(new_n22092_), .Y(new_n22093_));
  OAI21X1  g19657(.A0(new_n22091_), .A1(new_n12684_), .B0(new_n22093_), .Y(new_n22094_));
  MX2X1    g19658(.A(new_n22094_), .B(new_n22089_), .S0(new_n11884_), .Y(new_n22095_));
  AOI21X1  g19659(.A0(new_n21912_), .A1(pi0647), .B0(pi1157), .Y(new_n22096_));
  OAI21X1  g19660(.A0(new_n22095_), .A1(pi0647), .B0(new_n22096_), .Y(new_n22097_));
  INVX1    g19661(.A(new_n22097_), .Y(new_n22098_));
  INVX1    g19662(.A(new_n22095_), .Y(new_n22099_));
  MX2X1    g19663(.A(new_n22099_), .B(new_n21912_), .S0(new_n12705_), .Y(new_n22100_));
  INVX1    g19664(.A(new_n22100_), .Y(new_n22101_));
  AOI22X1  g19665(.A0(new_n22101_), .A1(new_n14386_), .B0(new_n22098_), .B1(pi0630), .Y(new_n22102_));
  OAI21X1  g19666(.A0(new_n22008_), .A1(new_n14384_), .B0(new_n22102_), .Y(new_n22103_));
  NOR2X1   g19667(.A(new_n22007_), .B(new_n14395_), .Y(new_n22104_));
  OAI22X1  g19668(.A0(new_n22093_), .A1(new_n12689_), .B0(new_n22091_), .B1(new_n12708_), .Y(new_n22105_));
  NOR2X1   g19669(.A(new_n22105_), .B(new_n22104_), .Y(new_n22106_));
  AOI21X1  g19670(.A0(new_n21911_), .A1(pi0626), .B0(new_n16352_), .Y(new_n22107_));
  OAI21X1  g19671(.A0(new_n22006_), .A1(pi0626), .B0(new_n22107_), .Y(new_n22108_));
  OR2X1    g19672(.A(new_n22006_), .B(new_n12664_), .Y(new_n22109_));
  AOI21X1  g19673(.A0(new_n21911_), .A1(new_n12664_), .B0(new_n16356_), .Y(new_n22110_));
  MX2X1    g19674(.A(new_n22087_), .B(new_n21912_), .S0(new_n12659_), .Y(new_n22111_));
  AOI22X1  g19675(.A0(new_n22111_), .A1(new_n12769_), .B0(new_n22110_), .B1(new_n22109_), .Y(new_n22112_));
  AOI21X1  g19676(.A0(new_n22112_), .A1(new_n22108_), .B0(new_n11885_), .Y(new_n22113_));
  AND2X1   g19677(.A(new_n12463_), .B(new_n2973_), .Y(new_n22114_));
  OAI21X1  g19678(.A0(pi0665), .A1(new_n2973_), .B0(pi0633), .Y(new_n22115_));
  NOR3X1   g19679(.A(new_n22115_), .B(new_n22114_), .C(new_n21915_), .Y(new_n22116_));
  NOR3X1   g19680(.A(new_n13240_), .B(new_n12166_), .C(new_n2973_), .Y(new_n22117_));
  OR2X1    g19681(.A(pi0665), .B(pi0198), .Y(new_n22118_));
  OAI21X1  g19682(.A0(new_n22118_), .A1(new_n12096_), .B0(new_n21917_), .Y(new_n22119_));
  OAI21X1  g19683(.A0(new_n22119_), .A1(new_n22117_), .B0(pi0603), .Y(new_n22120_));
  NOR2X1   g19684(.A(new_n22120_), .B(new_n22116_), .Y(new_n22121_));
  AOI21X1  g19685(.A0(new_n22063_), .A1(new_n5027_), .B0(new_n22121_), .Y(new_n22122_));
  AOI21X1  g19686(.A0(new_n22062_), .A1(new_n21916_), .B0(new_n2953_), .Y(new_n22123_));
  OAI21X1  g19687(.A0(new_n22122_), .A1(new_n22062_), .B0(new_n22123_), .Y(new_n22124_));
  OR4X1    g19688(.A(new_n13227_), .B(new_n12101_), .C(new_n22072_), .D(new_n2973_), .Y(new_n22125_));
  OAI21X1  g19689(.A0(new_n11945_), .A1(pi0634), .B0(new_n22125_), .Y(new_n22126_));
  OR2X1    g19690(.A(pi0665), .B(new_n22072_), .Y(new_n22127_));
  AOI21X1  g19691(.A0(new_n21917_), .A1(pi0198), .B0(new_n22127_), .Y(new_n22128_));
  OAI21X1  g19692(.A0(new_n12093_), .A1(pi0198), .B0(new_n22128_), .Y(new_n22129_));
  AND2X1   g19693(.A(new_n22129_), .B(pi0603), .Y(new_n22130_));
  OAI21X1  g19694(.A0(new_n21918_), .A1(new_n21917_), .B0(new_n22130_), .Y(new_n22131_));
  AOI21X1  g19695(.A0(new_n22126_), .A1(new_n21917_), .B0(new_n22131_), .Y(new_n22132_));
  NOR3X1   g19696(.A(new_n22067_), .B(new_n22065_), .C(pi0603), .Y(new_n22133_));
  NOR3X1   g19697(.A(new_n22133_), .B(new_n22132_), .C(new_n5029_), .Y(new_n22134_));
  OAI21X1  g19698(.A0(new_n21920_), .A1(pi0680), .B0(new_n2953_), .Y(new_n22135_));
  OR2X1    g19699(.A(new_n22135_), .B(new_n22134_), .Y(new_n22136_));
  AOI21X1  g19700(.A0(new_n22136_), .A1(new_n22124_), .B0(pi0039), .Y(new_n22137_));
  INVX1    g19701(.A(new_n21954_), .Y(new_n22138_));
  OAI21X1  g19702(.A0(new_n22127_), .A1(new_n12122_), .B0(new_n21926_), .Y(new_n22139_));
  AND2X1   g19703(.A(new_n22139_), .B(new_n5033_), .Y(new_n22140_));
  NAND2X1  g19704(.A(new_n12297_), .B(pi0634), .Y(new_n22141_));
  NAND2X1  g19705(.A(new_n22141_), .B(new_n21946_), .Y(new_n22142_));
  AOI21X1  g19706(.A0(new_n22142_), .A1(new_n5057_), .B0(new_n22140_), .Y(new_n22143_));
  NOR2X1   g19707(.A(new_n22143_), .B(new_n5027_), .Y(new_n22144_));
  INVX1    g19708(.A(new_n22144_), .Y(new_n22145_));
  NOR3X1   g19709(.A(new_n22143_), .B(pi0642), .C(new_n5027_), .Y(new_n22146_));
  OR2X1    g19710(.A(new_n22012_), .B(pi0603), .Y(new_n22147_));
  NAND3X1  g19711(.A(new_n22139_), .B(pi0642), .C(pi0603), .Y(new_n22148_));
  NAND2X1  g19712(.A(new_n22148_), .B(new_n22147_), .Y(new_n22149_));
  OAI21X1  g19713(.A0(new_n22149_), .A1(new_n22146_), .B0(new_n12323_), .Y(new_n22150_));
  AND2X1   g19714(.A(new_n22139_), .B(pi0603), .Y(new_n22151_));
  AOI21X1  g19715(.A0(new_n22014_), .A1(new_n5027_), .B0(new_n22151_), .Y(new_n22152_));
  OR2X1    g19716(.A(new_n22152_), .B(new_n12323_), .Y(new_n22153_));
  AND2X1   g19717(.A(new_n22153_), .B(new_n12290_), .Y(new_n22154_));
  AOI21X1  g19718(.A0(new_n22019_), .A1(new_n5027_), .B0(new_n12290_), .Y(new_n22155_));
  AOI22X1  g19719(.A0(new_n22155_), .A1(new_n22145_), .B0(new_n22154_), .B1(new_n22150_), .Y(new_n22156_));
  MX2X1    g19720(.A(new_n22156_), .B(new_n22138_), .S0(new_n5029_), .Y(new_n22157_));
  NOR3X1   g19721(.A(new_n21965_), .B(new_n21964_), .C(new_n21959_), .Y(new_n22158_));
  OR2X1    g19722(.A(new_n22158_), .B(pi0680), .Y(new_n22159_));
  AOI21X1  g19723(.A0(new_n22151_), .A1(new_n12127_), .B0(new_n21962_), .Y(new_n22160_));
  NAND2X1  g19724(.A(new_n22160_), .B(new_n5367_), .Y(new_n22161_));
  NOR2X1   g19725(.A(new_n22160_), .B(new_n5033_), .Y(new_n22162_));
  OAI21X1  g19726(.A0(new_n22162_), .A1(new_n22142_), .B0(new_n22161_), .Y(new_n22163_));
  OAI21X1  g19727(.A0(new_n22025_), .A1(pi0603), .B0(new_n22163_), .Y(new_n22164_));
  OAI22X1  g19728(.A0(new_n22017_), .A1(new_n12120_), .B0(new_n21946_), .B1(new_n5027_), .Y(new_n22165_));
  AOI22X1  g19729(.A0(new_n22165_), .A1(new_n5030_), .B0(new_n22164_), .B1(new_n12209_), .Y(new_n22166_));
  AND2X1   g19730(.A(new_n22166_), .B(new_n22159_), .Y(new_n22167_));
  OAI21X1  g19731(.A0(new_n22167_), .A1(new_n5050_), .B0(new_n2971_), .Y(new_n22168_));
  AOI21X1  g19732(.A0(new_n22157_), .A1(new_n5050_), .B0(new_n22168_), .Y(new_n22169_));
  OAI21X1  g19733(.A0(new_n22033_), .A1(new_n12482_), .B0(new_n21924_), .Y(new_n22170_));
  OAI21X1  g19734(.A0(new_n22170_), .A1(new_n2971_), .B0(new_n2964_), .Y(new_n22171_));
  NOR2X1   g19735(.A(new_n22171_), .B(new_n22169_), .Y(new_n22172_));
  OR2X1    g19736(.A(new_n22118_), .B(new_n12137_), .Y(new_n22173_));
  NAND3X1  g19737(.A(new_n12108_), .B(new_n12255_), .C(pi0198), .Y(new_n22174_));
  NAND3X1  g19738(.A(new_n22174_), .B(new_n22173_), .C(new_n22036_), .Y(new_n22175_));
  OAI21X1  g19739(.A0(new_n11964_), .A1(new_n11958_), .B0(new_n21923_), .Y(new_n22176_));
  OAI21X1  g19740(.A0(new_n22036_), .A1(pi0634), .B0(new_n22176_), .Y(new_n22177_));
  AOI21X1  g19741(.A0(new_n22175_), .A1(pi0634), .B0(new_n22177_), .Y(new_n22178_));
  NOR2X1   g19742(.A(new_n22178_), .B(new_n5033_), .Y(new_n22179_));
  OAI21X1  g19743(.A0(new_n22179_), .A1(new_n22140_), .B0(pi0603), .Y(new_n22180_));
  OAI21X1  g19744(.A0(new_n22045_), .A1(pi0603), .B0(new_n22180_), .Y(new_n22181_));
  NAND2X1  g19745(.A(new_n22181_), .B(new_n5030_), .Y(new_n22182_));
  NAND3X1  g19746(.A(new_n22180_), .B(new_n22147_), .C(new_n12125_), .Y(new_n22183_));
  AOI21X1  g19747(.A0(new_n22152_), .A1(new_n12127_), .B0(new_n12235_), .Y(new_n22184_));
  AOI22X1  g19748(.A0(new_n22184_), .A1(new_n22183_), .B0(new_n21933_), .B1(new_n5029_), .Y(new_n22185_));
  AND2X1   g19749(.A(new_n22185_), .B(new_n22182_), .Y(new_n22186_));
  AOI21X1  g19750(.A0(new_n22040_), .A1(new_n5027_), .B0(new_n22162_), .Y(new_n22187_));
  NOR3X1   g19751(.A(new_n22178_), .B(new_n12127_), .C(new_n5027_), .Y(new_n22188_));
  NOR2X1   g19752(.A(new_n22178_), .B(new_n22160_), .Y(new_n22189_));
  NOR2X1   g19753(.A(new_n22189_), .B(new_n22188_), .Y(new_n22190_));
  AOI21X1  g19754(.A0(new_n22190_), .A1(new_n22187_), .B0(new_n12235_), .Y(new_n22191_));
  MX2X1    g19755(.A(new_n22178_), .B(new_n22038_), .S0(new_n5027_), .Y(new_n22192_));
  OAI22X1  g19756(.A0(new_n22192_), .A1(new_n5282_), .B0(new_n21938_), .B1(pi0680), .Y(new_n22193_));
  NOR3X1   g19757(.A(new_n22193_), .B(new_n22191_), .C(new_n5050_), .Y(new_n22194_));
  OR2X1    g19758(.A(new_n22194_), .B(new_n2964_), .Y(new_n22195_));
  AOI21X1  g19759(.A0(new_n22186_), .A1(new_n5050_), .B0(new_n22195_), .Y(new_n22196_));
  OAI21X1  g19760(.A0(new_n22196_), .A1(new_n22172_), .B0(new_n2953_), .Y(new_n22197_));
  OAI21X1  g19761(.A0(new_n22167_), .A1(new_n5070_), .B0(new_n10137_), .Y(new_n22198_));
  AOI21X1  g19762(.A0(new_n22157_), .A1(new_n5070_), .B0(new_n22198_), .Y(new_n22199_));
  OAI21X1  g19763(.A0(new_n22170_), .A1(new_n10137_), .B0(new_n2954_), .Y(new_n22200_));
  AND2X1   g19764(.A(new_n22186_), .B(new_n5070_), .Y(new_n22201_));
  NOR3X1   g19765(.A(new_n22193_), .B(new_n22191_), .C(new_n5070_), .Y(new_n22202_));
  OR2X1    g19766(.A(new_n22202_), .B(new_n2954_), .Y(new_n22203_));
  OAI22X1  g19767(.A0(new_n22203_), .A1(new_n22201_), .B0(new_n22200_), .B1(new_n22199_), .Y(new_n22204_));
  AOI21X1  g19768(.A0(new_n22204_), .A1(pi0299), .B0(new_n2959_), .Y(new_n22205_));
  AOI21X1  g19769(.A0(new_n22205_), .A1(new_n22197_), .B0(new_n22137_), .Y(new_n22206_));
  AND2X1   g19770(.A(new_n12483_), .B(pi0634), .Y(new_n22207_));
  OAI21X1  g19771(.A0(new_n22207_), .A1(new_n21985_), .B0(new_n2959_), .Y(new_n22208_));
  AOI21X1  g19772(.A0(new_n22208_), .A1(new_n21982_), .B0(new_n3810_), .Y(new_n22209_));
  OAI21X1  g19773(.A0(new_n22206_), .A1(pi0038), .B0(new_n22209_), .Y(new_n22210_));
  OAI21X1  g19774(.A0(new_n3129_), .A1(new_n2973_), .B0(new_n22210_), .Y(new_n22211_));
  AOI21X1  g19775(.A0(new_n21988_), .A1(pi0625), .B0(pi1153), .Y(new_n22212_));
  OAI21X1  g19776(.A0(new_n22211_), .A1(pi0625), .B0(new_n22212_), .Y(new_n22213_));
  NOR2X1   g19777(.A(new_n22079_), .B(pi0608), .Y(new_n22214_));
  AOI21X1  g19778(.A0(new_n21988_), .A1(new_n12493_), .B0(new_n12494_), .Y(new_n22215_));
  OAI21X1  g19779(.A0(new_n22211_), .A1(new_n12493_), .B0(new_n22215_), .Y(new_n22216_));
  NOR2X1   g19780(.A(new_n22081_), .B(new_n12584_), .Y(new_n22217_));
  AOI22X1  g19781(.A0(new_n22217_), .A1(new_n22216_), .B0(new_n22214_), .B1(new_n22213_), .Y(new_n22218_));
  OR2X1    g19782(.A(new_n22211_), .B(pi0778), .Y(new_n22219_));
  OAI21X1  g19783(.A0(new_n22218_), .A1(new_n11889_), .B0(new_n22219_), .Y(new_n22220_));
  OAI21X1  g19784(.A0(new_n22084_), .A1(new_n12590_), .B0(new_n12591_), .Y(new_n22221_));
  AOI21X1  g19785(.A0(new_n22220_), .A1(new_n12590_), .B0(new_n22221_), .Y(new_n22222_));
  OAI21X1  g19786(.A0(new_n21991_), .A1(new_n12591_), .B0(new_n12596_), .Y(new_n22223_));
  OAI21X1  g19787(.A0(new_n22084_), .A1(pi0609), .B0(pi1155), .Y(new_n22224_));
  AOI21X1  g19788(.A0(new_n22220_), .A1(pi0609), .B0(new_n22224_), .Y(new_n22225_));
  OAI21X1  g19789(.A0(new_n21992_), .A1(pi1155), .B0(pi0660), .Y(new_n22226_));
  OAI22X1  g19790(.A0(new_n22226_), .A1(new_n22225_), .B0(new_n22223_), .B1(new_n22222_), .Y(new_n22227_));
  AND2X1   g19791(.A(new_n22220_), .B(new_n11888_), .Y(new_n22228_));
  AOI21X1  g19792(.A0(new_n22227_), .A1(pi0785), .B0(new_n22228_), .Y(new_n22229_));
  AOI21X1  g19793(.A0(new_n22086_), .A1(pi0618), .B0(pi1154), .Y(new_n22230_));
  OAI21X1  g19794(.A0(new_n22229_), .A1(pi0618), .B0(new_n22230_), .Y(new_n22231_));
  NOR2X1   g19795(.A(new_n21996_), .B(pi0627), .Y(new_n22232_));
  AOI21X1  g19796(.A0(new_n22086_), .A1(new_n12614_), .B0(new_n12615_), .Y(new_n22233_));
  OAI21X1  g19797(.A0(new_n22229_), .A1(new_n12614_), .B0(new_n22233_), .Y(new_n22234_));
  NOR2X1   g19798(.A(new_n21998_), .B(new_n12622_), .Y(new_n22235_));
  AOI22X1  g19799(.A0(new_n22235_), .A1(new_n22234_), .B0(new_n22232_), .B1(new_n22231_), .Y(new_n22236_));
  MX2X1    g19800(.A(new_n22236_), .B(new_n22229_), .S0(new_n11887_), .Y(new_n22237_));
  NOR2X1   g19801(.A(new_n22237_), .B(pi0619), .Y(new_n22238_));
  AND2X1   g19802(.A(new_n22087_), .B(pi0619), .Y(new_n22239_));
  OR2X1    g19803(.A(new_n22239_), .B(pi1159), .Y(new_n22240_));
  AND2X1   g19804(.A(new_n22002_), .B(new_n12645_), .Y(new_n22241_));
  OAI21X1  g19805(.A0(new_n22240_), .A1(new_n22238_), .B0(new_n22241_), .Y(new_n22242_));
  AOI21X1  g19806(.A0(new_n22087_), .A1(new_n12637_), .B0(new_n12638_), .Y(new_n22243_));
  OAI21X1  g19807(.A0(new_n22237_), .A1(new_n12637_), .B0(new_n22243_), .Y(new_n22244_));
  NAND3X1  g19808(.A(new_n22244_), .B(new_n22004_), .C(pi0648), .Y(new_n22245_));
  NAND3X1  g19809(.A(new_n22245_), .B(new_n22242_), .C(pi0789), .Y(new_n22246_));
  AOI21X1  g19810(.A0(new_n22237_), .A1(new_n11886_), .B0(new_n14264_), .Y(new_n22247_));
  AND2X1   g19811(.A(new_n22247_), .B(new_n22246_), .Y(new_n22248_));
  OAI22X1  g19812(.A0(new_n22248_), .A1(new_n22113_), .B0(new_n22106_), .B1(new_n11884_), .Y(new_n22249_));
  AOI21X1  g19813(.A0(new_n22106_), .A1(new_n14273_), .B0(new_n14269_), .Y(new_n22250_));
  AOI22X1  g19814(.A0(new_n22250_), .A1(new_n22249_), .B0(new_n22103_), .B1(pi0787), .Y(new_n22251_));
  NAND2X1  g19815(.A(new_n22251_), .B(pi0644), .Y(new_n22252_));
  AOI21X1  g19816(.A0(new_n22101_), .A1(pi1157), .B0(new_n22098_), .Y(new_n22253_));
  MX2X1    g19817(.A(new_n22253_), .B(new_n22099_), .S0(new_n11883_), .Y(new_n22254_));
  AOI21X1  g19818(.A0(new_n22254_), .A1(new_n12743_), .B0(new_n12739_), .Y(new_n22255_));
  MX2X1    g19819(.A(new_n22008_), .B(new_n21912_), .S0(new_n12735_), .Y(new_n22256_));
  OAI21X1  g19820(.A0(new_n21911_), .A1(pi0644), .B0(new_n12739_), .Y(new_n22257_));
  AOI21X1  g19821(.A0(new_n22256_), .A1(pi0644), .B0(new_n22257_), .Y(new_n22258_));
  OR2X1    g19822(.A(new_n22258_), .B(new_n11882_), .Y(new_n22259_));
  AOI21X1  g19823(.A0(new_n22255_), .A1(new_n22252_), .B0(new_n22259_), .Y(new_n22260_));
  NAND2X1  g19824(.A(new_n22251_), .B(new_n12743_), .Y(new_n22261_));
  AOI21X1  g19825(.A0(new_n22254_), .A1(pi0644), .B0(pi0715), .Y(new_n22262_));
  OAI21X1  g19826(.A0(new_n21911_), .A1(new_n12743_), .B0(pi0715), .Y(new_n22263_));
  AOI21X1  g19827(.A0(new_n22256_), .A1(new_n12743_), .B0(new_n22263_), .Y(new_n22264_));
  OR2X1    g19828(.A(new_n22264_), .B(pi1160), .Y(new_n22265_));
  AOI21X1  g19829(.A0(new_n22262_), .A1(new_n22261_), .B0(new_n22265_), .Y(new_n22266_));
  OR2X1    g19830(.A(new_n22266_), .B(new_n12897_), .Y(new_n22267_));
  OAI22X1  g19831(.A0(new_n22267_), .A1(new_n22260_), .B0(new_n22251_), .B1(pi0790), .Y(new_n22268_));
  MX2X1    g19832(.A(new_n22268_), .B(pi0198), .S0(po1038), .Y(po0355));
  INVX1    g19833(.A(pi0637), .Y(new_n22270_));
  INVX1    g19834(.A(pi0617), .Y(new_n22271_));
  OAI21X1  g19835(.A0(new_n12574_), .A1(new_n3810_), .B0(pi0199), .Y(new_n22272_));
  AND2X1   g19836(.A(new_n12178_), .B(new_n4995_), .Y(new_n22273_));
  INVX1    g19837(.A(new_n22273_), .Y(new_n22274_));
  INVX1    g19838(.A(new_n13703_), .Y(new_n22275_));
  AOI21X1  g19839(.A0(new_n22274_), .A1(new_n7941_), .B0(new_n22275_), .Y(new_n22276_));
  OAI21X1  g19840(.A0(new_n12199_), .A1(pi0199), .B0(new_n2996_), .Y(new_n22277_));
  AOI21X1  g19841(.A0(new_n12162_), .A1(pi0199), .B0(new_n22277_), .Y(new_n22278_));
  OAI21X1  g19842(.A0(new_n22278_), .A1(new_n22276_), .B0(new_n3129_), .Y(new_n22279_));
  NOR2X1   g19843(.A(new_n3129_), .B(new_n7941_), .Y(new_n22280_));
  NOR2X1   g19844(.A(new_n22280_), .B(new_n22271_), .Y(new_n22281_));
  AOI22X1  g19845(.A0(new_n22281_), .A1(new_n22279_), .B0(new_n22272_), .B1(new_n22271_), .Y(new_n22282_));
  NOR3X1   g19846(.A(new_n13671_), .B(new_n7941_), .C(pi0038), .Y(new_n22283_));
  AND2X1   g19847(.A(new_n16793_), .B(new_n3129_), .Y(new_n22284_));
  AOI21X1  g19848(.A0(new_n13669_), .A1(pi0038), .B0(pi0617), .Y(new_n22285_));
  OAI21X1  g19849(.A0(new_n22284_), .A1(pi0199), .B0(new_n22285_), .Y(new_n22286_));
  OAI21X1  g19850(.A0(new_n16796_), .A1(new_n3810_), .B0(new_n7941_), .Y(new_n22287_));
  AOI21X1  g19851(.A0(new_n13694_), .A1(pi0199), .B0(new_n22271_), .Y(new_n22288_));
  AOI21X1  g19852(.A0(new_n22288_), .A1(new_n22287_), .B0(new_n22280_), .Y(new_n22289_));
  OAI21X1  g19853(.A0(new_n22286_), .A1(new_n22283_), .B0(new_n22289_), .Y(new_n22290_));
  MX2X1    g19854(.A(new_n22290_), .B(new_n22282_), .S0(new_n22270_), .Y(new_n22291_));
  AOI21X1  g19855(.A0(new_n13699_), .A1(new_n3129_), .B0(new_n7941_), .Y(new_n22292_));
  NAND2X1  g19856(.A(new_n22281_), .B(new_n22279_), .Y(new_n22293_));
  OAI21X1  g19857(.A0(new_n22292_), .A1(pi0617), .B0(new_n22293_), .Y(new_n22294_));
  AOI21X1  g19858(.A0(new_n22294_), .A1(pi0625), .B0(pi1153), .Y(new_n22295_));
  OAI21X1  g19859(.A0(new_n22291_), .A1(pi0625), .B0(new_n22295_), .Y(new_n22296_));
  NOR2X1   g19860(.A(new_n12202_), .B(pi0199), .Y(new_n22297_));
  OAI21X1  g19861(.A0(new_n12522_), .A1(pi0199), .B0(pi0039), .Y(new_n22298_));
  AOI21X1  g19862(.A0(new_n12560_), .A1(pi0199), .B0(new_n22298_), .Y(new_n22299_));
  AND2X1   g19863(.A(new_n13391_), .B(pi0199), .Y(new_n22300_));
  OAI21X1  g19864(.A0(new_n13685_), .A1(pi0199), .B0(new_n2959_), .Y(new_n22301_));
  OAI21X1  g19865(.A0(new_n22301_), .A1(new_n22300_), .B0(new_n2996_), .Y(new_n22302_));
  OAI22X1  g19866(.A0(new_n22302_), .A1(new_n22299_), .B0(new_n22297_), .B1(new_n14017_), .Y(new_n22303_));
  OAI21X1  g19867(.A0(new_n3129_), .A1(new_n7941_), .B0(pi0637), .Y(new_n22304_));
  AOI21X1  g19868(.A0(new_n22303_), .A1(new_n3129_), .B0(new_n22304_), .Y(new_n22305_));
  AOI21X1  g19869(.A0(new_n22272_), .A1(new_n22270_), .B0(new_n22305_), .Y(new_n22306_));
  AOI21X1  g19870(.A0(new_n22272_), .A1(new_n12493_), .B0(new_n12494_), .Y(new_n22307_));
  OAI21X1  g19871(.A0(new_n22306_), .A1(new_n12493_), .B0(new_n22307_), .Y(new_n22308_));
  AND2X1   g19872(.A(new_n22308_), .B(new_n12584_), .Y(new_n22309_));
  AOI21X1  g19873(.A0(new_n22294_), .A1(new_n12493_), .B0(new_n12494_), .Y(new_n22310_));
  OAI21X1  g19874(.A0(new_n22291_), .A1(new_n12493_), .B0(new_n22310_), .Y(new_n22311_));
  AOI21X1  g19875(.A0(new_n22272_), .A1(pi0625), .B0(pi1153), .Y(new_n22312_));
  OAI21X1  g19876(.A0(new_n22306_), .A1(pi0625), .B0(new_n22312_), .Y(new_n22313_));
  AND2X1   g19877(.A(new_n22313_), .B(pi0608), .Y(new_n22314_));
  AOI22X1  g19878(.A0(new_n22314_), .A1(new_n22311_), .B0(new_n22309_), .B1(new_n22296_), .Y(new_n22315_));
  MX2X1    g19879(.A(new_n22315_), .B(new_n22291_), .S0(new_n11889_), .Y(new_n22316_));
  AOI21X1  g19880(.A0(new_n22313_), .A1(new_n22308_), .B0(new_n11889_), .Y(new_n22317_));
  AOI21X1  g19881(.A0(new_n22306_), .A1(new_n11889_), .B0(new_n22317_), .Y(new_n22318_));
  AOI21X1  g19882(.A0(new_n22318_), .A1(pi0609), .B0(pi1155), .Y(new_n22319_));
  OAI21X1  g19883(.A0(new_n22316_), .A1(pi0609), .B0(new_n22319_), .Y(new_n22320_));
  MX2X1    g19884(.A(new_n22282_), .B(new_n22292_), .S0(new_n12601_), .Y(new_n22321_));
  AOI21X1  g19885(.A0(new_n22272_), .A1(new_n12590_), .B0(new_n12591_), .Y(new_n22322_));
  OAI21X1  g19886(.A0(new_n22321_), .A1(new_n12590_), .B0(new_n22322_), .Y(new_n22323_));
  AND2X1   g19887(.A(new_n22323_), .B(new_n12596_), .Y(new_n22324_));
  AOI21X1  g19888(.A0(new_n22318_), .A1(new_n12590_), .B0(new_n12591_), .Y(new_n22325_));
  OAI21X1  g19889(.A0(new_n22316_), .A1(new_n12590_), .B0(new_n22325_), .Y(new_n22326_));
  AOI21X1  g19890(.A0(new_n22272_), .A1(pi0609), .B0(pi1155), .Y(new_n22327_));
  OAI21X1  g19891(.A0(new_n22321_), .A1(pi0609), .B0(new_n22327_), .Y(new_n22328_));
  AND2X1   g19892(.A(new_n22328_), .B(pi0660), .Y(new_n22329_));
  AOI22X1  g19893(.A0(new_n22329_), .A1(new_n22326_), .B0(new_n22324_), .B1(new_n22320_), .Y(new_n22330_));
  MX2X1    g19894(.A(new_n22330_), .B(new_n22316_), .S0(new_n11888_), .Y(new_n22331_));
  MX2X1    g19895(.A(new_n22318_), .B(new_n22272_), .S0(new_n12618_), .Y(new_n22332_));
  AOI21X1  g19896(.A0(new_n22332_), .A1(pi0618), .B0(pi1154), .Y(new_n22333_));
  OAI21X1  g19897(.A0(new_n22331_), .A1(pi0618), .B0(new_n22333_), .Y(new_n22334_));
  AOI21X1  g19898(.A0(new_n22328_), .A1(new_n22323_), .B0(new_n11888_), .Y(new_n22335_));
  AOI21X1  g19899(.A0(new_n22321_), .A1(new_n11888_), .B0(new_n22335_), .Y(new_n22336_));
  OAI21X1  g19900(.A0(new_n22292_), .A1(pi0618), .B0(pi1154), .Y(new_n22337_));
  AOI21X1  g19901(.A0(new_n22336_), .A1(pi0618), .B0(new_n22337_), .Y(new_n22338_));
  NOR2X1   g19902(.A(new_n22338_), .B(pi0627), .Y(new_n22339_));
  AOI21X1  g19903(.A0(new_n22332_), .A1(new_n12614_), .B0(new_n12615_), .Y(new_n22340_));
  OAI21X1  g19904(.A0(new_n22331_), .A1(new_n12614_), .B0(new_n22340_), .Y(new_n22341_));
  OAI21X1  g19905(.A0(new_n22292_), .A1(new_n12614_), .B0(new_n12615_), .Y(new_n22342_));
  AOI21X1  g19906(.A0(new_n22336_), .A1(new_n12614_), .B0(new_n22342_), .Y(new_n22343_));
  NOR2X1   g19907(.A(new_n22343_), .B(new_n12622_), .Y(new_n22344_));
  AOI22X1  g19908(.A0(new_n22344_), .A1(new_n22341_), .B0(new_n22339_), .B1(new_n22334_), .Y(new_n22345_));
  MX2X1    g19909(.A(new_n22345_), .B(new_n22331_), .S0(new_n11887_), .Y(new_n22346_));
  MX2X1    g19910(.A(new_n22332_), .B(new_n22272_), .S0(new_n12641_), .Y(new_n22347_));
  AOI21X1  g19911(.A0(new_n22347_), .A1(pi0619), .B0(pi1159), .Y(new_n22348_));
  OAI21X1  g19912(.A0(new_n22346_), .A1(pi0619), .B0(new_n22348_), .Y(new_n22349_));
  OR2X1    g19913(.A(new_n22336_), .B(pi0781), .Y(new_n22350_));
  OAI21X1  g19914(.A0(new_n22343_), .A1(new_n22338_), .B0(pi0781), .Y(new_n22351_));
  NAND2X1  g19915(.A(new_n22351_), .B(new_n22350_), .Y(new_n22352_));
  AOI21X1  g19916(.A0(new_n22272_), .A1(new_n12637_), .B0(new_n12638_), .Y(new_n22353_));
  OAI21X1  g19917(.A0(new_n22352_), .A1(new_n12637_), .B0(new_n22353_), .Y(new_n22354_));
  AND2X1   g19918(.A(new_n22354_), .B(new_n12645_), .Y(new_n22355_));
  AOI21X1  g19919(.A0(new_n22347_), .A1(new_n12637_), .B0(new_n12638_), .Y(new_n22356_));
  OAI21X1  g19920(.A0(new_n22346_), .A1(new_n12637_), .B0(new_n22356_), .Y(new_n22357_));
  AOI21X1  g19921(.A0(new_n22272_), .A1(pi0619), .B0(pi1159), .Y(new_n22358_));
  OAI21X1  g19922(.A0(new_n22352_), .A1(pi0619), .B0(new_n22358_), .Y(new_n22359_));
  AND2X1   g19923(.A(new_n22359_), .B(pi0648), .Y(new_n22360_));
  AOI22X1  g19924(.A0(new_n22360_), .A1(new_n22357_), .B0(new_n22355_), .B1(new_n22349_), .Y(new_n22361_));
  MX2X1    g19925(.A(new_n22361_), .B(new_n22346_), .S0(new_n11886_), .Y(new_n22362_));
  MX2X1    g19926(.A(new_n22347_), .B(new_n22272_), .S0(new_n12659_), .Y(new_n22363_));
  OAI21X1  g19927(.A0(new_n22363_), .A1(new_n12664_), .B0(new_n12672_), .Y(new_n22364_));
  AOI21X1  g19928(.A0(new_n22362_), .A1(new_n12664_), .B0(new_n22364_), .Y(new_n22365_));
  AOI21X1  g19929(.A0(new_n22359_), .A1(new_n22354_), .B0(new_n11886_), .Y(new_n22366_));
  AOI21X1  g19930(.A0(new_n22352_), .A1(new_n11886_), .B0(new_n22366_), .Y(new_n22367_));
  AOI21X1  g19931(.A0(new_n22292_), .A1(pi0626), .B0(new_n12672_), .Y(new_n22368_));
  OAI21X1  g19932(.A0(new_n22367_), .A1(pi0626), .B0(new_n22368_), .Y(new_n22369_));
  NAND2X1  g19933(.A(new_n22369_), .B(new_n12676_), .Y(new_n22370_));
  OAI21X1  g19934(.A0(new_n22363_), .A1(pi0626), .B0(pi0641), .Y(new_n22371_));
  AOI21X1  g19935(.A0(new_n22362_), .A1(pi0626), .B0(new_n22371_), .Y(new_n22372_));
  AOI21X1  g19936(.A0(new_n22292_), .A1(new_n12664_), .B0(pi0641), .Y(new_n22373_));
  OAI21X1  g19937(.A0(new_n22367_), .A1(new_n12664_), .B0(new_n22373_), .Y(new_n22374_));
  NAND2X1  g19938(.A(new_n22374_), .B(pi1158), .Y(new_n22375_));
  OAI22X1  g19939(.A0(new_n22375_), .A1(new_n22372_), .B0(new_n22370_), .B1(new_n22365_), .Y(new_n22376_));
  MX2X1    g19940(.A(new_n22376_), .B(new_n22362_), .S0(new_n11885_), .Y(new_n22377_));
  MX2X1    g19941(.A(new_n22367_), .B(new_n22272_), .S0(new_n12841_), .Y(new_n22378_));
  AOI21X1  g19942(.A0(new_n22378_), .A1(pi0628), .B0(pi1156), .Y(new_n22379_));
  OAI21X1  g19943(.A0(new_n22377_), .A1(pi0628), .B0(new_n22379_), .Y(new_n22380_));
  MX2X1    g19944(.A(new_n22363_), .B(new_n22272_), .S0(new_n12691_), .Y(new_n22381_));
  INVX1    g19945(.A(new_n22381_), .Y(new_n22382_));
  AOI21X1  g19946(.A0(new_n22272_), .A1(new_n12683_), .B0(new_n12684_), .Y(new_n22383_));
  OAI21X1  g19947(.A0(new_n22382_), .A1(new_n12683_), .B0(new_n22383_), .Y(new_n22384_));
  AND2X1   g19948(.A(new_n22384_), .B(new_n12689_), .Y(new_n22385_));
  AOI21X1  g19949(.A0(new_n22378_), .A1(new_n12683_), .B0(new_n12684_), .Y(new_n22386_));
  OAI21X1  g19950(.A0(new_n22377_), .A1(new_n12683_), .B0(new_n22386_), .Y(new_n22387_));
  AOI21X1  g19951(.A0(new_n22272_), .A1(pi0628), .B0(pi1156), .Y(new_n22388_));
  OAI21X1  g19952(.A0(new_n22382_), .A1(pi0628), .B0(new_n22388_), .Y(new_n22389_));
  AND2X1   g19953(.A(new_n22389_), .B(pi0629), .Y(new_n22390_));
  AOI22X1  g19954(.A0(new_n22390_), .A1(new_n22387_), .B0(new_n22385_), .B1(new_n22380_), .Y(new_n22391_));
  MX2X1    g19955(.A(new_n22391_), .B(new_n22377_), .S0(new_n11884_), .Y(new_n22392_));
  MX2X1    g19956(.A(new_n22378_), .B(new_n22272_), .S0(new_n12711_), .Y(new_n22393_));
  AOI21X1  g19957(.A0(new_n22393_), .A1(pi0647), .B0(pi1157), .Y(new_n22394_));
  OAI21X1  g19958(.A0(new_n22392_), .A1(pi0647), .B0(new_n22394_), .Y(new_n22395_));
  NOR2X1   g19959(.A(new_n22381_), .B(pi0792), .Y(new_n22396_));
  AOI21X1  g19960(.A0(new_n22389_), .A1(new_n22384_), .B0(new_n11884_), .Y(new_n22397_));
  NOR2X1   g19961(.A(new_n22397_), .B(new_n22396_), .Y(new_n22398_));
  INVX1    g19962(.A(new_n22398_), .Y(new_n22399_));
  AOI21X1  g19963(.A0(new_n22272_), .A1(new_n12705_), .B0(new_n12706_), .Y(new_n22400_));
  OAI21X1  g19964(.A0(new_n22399_), .A1(new_n12705_), .B0(new_n22400_), .Y(new_n22401_));
  AND2X1   g19965(.A(new_n22401_), .B(new_n12723_), .Y(new_n22402_));
  AOI21X1  g19966(.A0(new_n22393_), .A1(new_n12705_), .B0(new_n12706_), .Y(new_n22403_));
  OAI21X1  g19967(.A0(new_n22392_), .A1(new_n12705_), .B0(new_n22403_), .Y(new_n22404_));
  AOI21X1  g19968(.A0(new_n22272_), .A1(pi0647), .B0(pi1157), .Y(new_n22405_));
  OAI21X1  g19969(.A0(new_n22399_), .A1(pi0647), .B0(new_n22405_), .Y(new_n22406_));
  AND2X1   g19970(.A(new_n22406_), .B(pi0630), .Y(new_n22407_));
  AOI22X1  g19971(.A0(new_n22407_), .A1(new_n22404_), .B0(new_n22402_), .B1(new_n22395_), .Y(new_n22408_));
  MX2X1    g19972(.A(new_n22408_), .B(new_n22392_), .S0(new_n11883_), .Y(new_n22409_));
  NOR2X1   g19973(.A(new_n22409_), .B(new_n12743_), .Y(new_n22410_));
  AND2X1   g19974(.A(new_n22406_), .B(new_n22401_), .Y(new_n22411_));
  MX2X1    g19975(.A(new_n22411_), .B(new_n22398_), .S0(new_n11883_), .Y(new_n22412_));
  AND2X1   g19976(.A(new_n22412_), .B(new_n12743_), .Y(new_n22413_));
  OR2X1    g19977(.A(new_n22413_), .B(new_n12739_), .Y(new_n22414_));
  AND2X1   g19978(.A(new_n22272_), .B(new_n12735_), .Y(new_n22415_));
  AOI21X1  g19979(.A0(new_n22393_), .A1(new_n12736_), .B0(new_n22415_), .Y(new_n22416_));
  AOI21X1  g19980(.A0(new_n22272_), .A1(new_n12743_), .B0(pi0715), .Y(new_n22417_));
  OAI21X1  g19981(.A0(new_n22416_), .A1(new_n12743_), .B0(new_n22417_), .Y(new_n22418_));
  AND2X1   g19982(.A(new_n22418_), .B(pi1160), .Y(new_n22419_));
  OAI21X1  g19983(.A0(new_n22414_), .A1(new_n22410_), .B0(new_n22419_), .Y(new_n22420_));
  AOI21X1  g19984(.A0(new_n22412_), .A1(pi0644), .B0(pi0715), .Y(new_n22421_));
  OAI21X1  g19985(.A0(new_n22409_), .A1(pi0644), .B0(new_n22421_), .Y(new_n22422_));
  AOI21X1  g19986(.A0(new_n22272_), .A1(pi0644), .B0(new_n12739_), .Y(new_n22423_));
  OAI21X1  g19987(.A0(new_n22416_), .A1(pi0644), .B0(new_n22423_), .Y(new_n22424_));
  AND2X1   g19988(.A(new_n22424_), .B(new_n11882_), .Y(new_n22425_));
  AOI21X1  g19989(.A0(new_n22425_), .A1(new_n22422_), .B0(new_n12897_), .Y(new_n22426_));
  AOI22X1  g19990(.A0(new_n22426_), .A1(new_n22420_), .B0(new_n22409_), .B1(new_n12897_), .Y(new_n22427_));
  OR2X1    g19991(.A(new_n6520_), .B(new_n7941_), .Y(new_n22428_));
  OAI21X1  g19992(.A0(new_n22427_), .A1(po1038), .B0(new_n22428_), .Y(po0356));
  AOI21X1  g19993(.A0(new_n13699_), .A1(new_n3129_), .B0(new_n8009_), .Y(new_n22430_));
  INVX1    g19994(.A(new_n22430_), .Y(new_n22431_));
  INVX1    g19995(.A(pi0606), .Y(new_n22432_));
  AOI21X1  g19996(.A0(new_n22274_), .A1(new_n8009_), .B0(new_n22275_), .Y(new_n22433_));
  INVX1    g19997(.A(new_n22433_), .Y(new_n22434_));
  AOI21X1  g19998(.A0(new_n13977_), .A1(new_n8009_), .B0(pi0038), .Y(new_n22435_));
  OAI21X1  g19999(.A0(new_n12910_), .A1(new_n8009_), .B0(new_n22435_), .Y(new_n22436_));
  AOI21X1  g20000(.A0(new_n22436_), .A1(new_n22434_), .B0(new_n3810_), .Y(new_n22437_));
  NOR2X1   g20001(.A(new_n3129_), .B(new_n8009_), .Y(new_n22438_));
  NOR3X1   g20002(.A(new_n22438_), .B(new_n22437_), .C(new_n22432_), .Y(new_n22439_));
  AOI21X1  g20003(.A0(new_n22431_), .A1(new_n22432_), .B0(new_n22439_), .Y(new_n22440_));
  MX2X1    g20004(.A(new_n22440_), .B(new_n22430_), .S0(new_n12601_), .Y(new_n22441_));
  AOI21X1  g20005(.A0(new_n22431_), .A1(new_n12590_), .B0(new_n12591_), .Y(new_n22442_));
  OAI21X1  g20006(.A0(new_n22441_), .A1(new_n12590_), .B0(new_n22442_), .Y(new_n22443_));
  AOI21X1  g20007(.A0(new_n22431_), .A1(pi0609), .B0(pi1155), .Y(new_n22444_));
  OAI21X1  g20008(.A0(new_n22441_), .A1(pi0609), .B0(new_n22444_), .Y(new_n22445_));
  AOI21X1  g20009(.A0(new_n22445_), .A1(new_n22443_), .B0(new_n11888_), .Y(new_n22446_));
  AOI21X1  g20010(.A0(new_n22441_), .A1(new_n11888_), .B0(new_n22446_), .Y(new_n22447_));
  OAI21X1  g20011(.A0(new_n22430_), .A1(pi0618), .B0(pi1154), .Y(new_n22448_));
  AOI21X1  g20012(.A0(new_n22447_), .A1(pi0618), .B0(new_n22448_), .Y(new_n22449_));
  OAI21X1  g20013(.A0(new_n22430_), .A1(new_n12614_), .B0(new_n12615_), .Y(new_n22450_));
  AOI21X1  g20014(.A0(new_n22447_), .A1(new_n12614_), .B0(new_n22450_), .Y(new_n22451_));
  NOR2X1   g20015(.A(new_n22451_), .B(new_n22449_), .Y(new_n22452_));
  MX2X1    g20016(.A(new_n22452_), .B(new_n22447_), .S0(new_n11887_), .Y(new_n22453_));
  OAI21X1  g20017(.A0(new_n22430_), .A1(pi0619), .B0(pi1159), .Y(new_n22454_));
  AOI21X1  g20018(.A0(new_n22453_), .A1(pi0619), .B0(new_n22454_), .Y(new_n22455_));
  OAI21X1  g20019(.A0(new_n22430_), .A1(new_n12637_), .B0(new_n12638_), .Y(new_n22456_));
  AOI21X1  g20020(.A0(new_n22453_), .A1(new_n12637_), .B0(new_n22456_), .Y(new_n22457_));
  NOR2X1   g20021(.A(new_n22457_), .B(new_n22455_), .Y(new_n22458_));
  MX2X1    g20022(.A(new_n22458_), .B(new_n22453_), .S0(new_n11886_), .Y(new_n22459_));
  MX2X1    g20023(.A(new_n22459_), .B(new_n22431_), .S0(new_n12841_), .Y(new_n22460_));
  INVX1    g20024(.A(pi0643), .Y(new_n22461_));
  AOI21X1  g20025(.A0(new_n12901_), .A1(new_n8009_), .B0(new_n14017_), .Y(new_n22462_));
  AND2X1   g20026(.A(new_n12513_), .B(new_n8009_), .Y(new_n22463_));
  OR2X1    g20027(.A(new_n22463_), .B(pi0299), .Y(new_n22464_));
  AOI21X1  g20028(.A0(new_n12948_), .A1(pi0200), .B0(new_n22464_), .Y(new_n22465_));
  AND2X1   g20029(.A(new_n12521_), .B(new_n8009_), .Y(new_n22466_));
  OR2X1    g20030(.A(new_n22466_), .B(new_n2953_), .Y(new_n22467_));
  AOI21X1  g20031(.A0(new_n12951_), .A1(pi0200), .B0(new_n22467_), .Y(new_n22468_));
  OAI21X1  g20032(.A0(new_n22468_), .A1(new_n22465_), .B0(pi0039), .Y(new_n22469_));
  AOI21X1  g20033(.A0(new_n12453_), .A1(pi0200), .B0(pi0039), .Y(new_n22470_));
  OAI21X1  g20034(.A0(new_n12473_), .A1(pi0200), .B0(new_n22470_), .Y(new_n22471_));
  AOI21X1  g20035(.A0(new_n22471_), .A1(new_n22469_), .B0(pi0038), .Y(new_n22472_));
  OAI21X1  g20036(.A0(new_n22472_), .A1(new_n22462_), .B0(new_n3129_), .Y(new_n22473_));
  NOR2X1   g20037(.A(new_n22438_), .B(new_n22461_), .Y(new_n22474_));
  AOI22X1  g20038(.A0(new_n22474_), .A1(new_n22473_), .B0(new_n22431_), .B1(new_n22461_), .Y(new_n22475_));
  AOI21X1  g20039(.A0(new_n22431_), .A1(new_n12493_), .B0(new_n12494_), .Y(new_n22476_));
  OAI21X1  g20040(.A0(new_n22475_), .A1(new_n12493_), .B0(new_n22476_), .Y(new_n22477_));
  AOI21X1  g20041(.A0(new_n22431_), .A1(pi0625), .B0(pi1153), .Y(new_n22478_));
  OAI21X1  g20042(.A0(new_n22475_), .A1(pi0625), .B0(new_n22478_), .Y(new_n22479_));
  AOI21X1  g20043(.A0(new_n22479_), .A1(new_n22477_), .B0(new_n11889_), .Y(new_n22480_));
  AOI21X1  g20044(.A0(new_n22475_), .A1(new_n11889_), .B0(new_n22480_), .Y(new_n22481_));
  INVX1    g20045(.A(new_n22481_), .Y(new_n22482_));
  MX2X1    g20046(.A(new_n22482_), .B(new_n22430_), .S0(new_n12618_), .Y(new_n22483_));
  INVX1    g20047(.A(new_n22483_), .Y(new_n22484_));
  MX2X1    g20048(.A(new_n22484_), .B(new_n22431_), .S0(new_n12641_), .Y(new_n22485_));
  INVX1    g20049(.A(new_n22485_), .Y(new_n22486_));
  MX2X1    g20050(.A(new_n22486_), .B(new_n22430_), .S0(new_n12659_), .Y(new_n22487_));
  MX2X1    g20051(.A(new_n22487_), .B(new_n22430_), .S0(new_n12691_), .Y(new_n22488_));
  AOI21X1  g20052(.A0(new_n22431_), .A1(new_n12683_), .B0(new_n12684_), .Y(new_n22489_));
  OAI21X1  g20053(.A0(new_n22488_), .A1(new_n12683_), .B0(new_n22489_), .Y(new_n22490_));
  AOI21X1  g20054(.A0(new_n22431_), .A1(pi0628), .B0(pi1156), .Y(new_n22491_));
  OAI21X1  g20055(.A0(new_n22488_), .A1(pi0628), .B0(new_n22491_), .Y(new_n22492_));
  MX2X1    g20056(.A(new_n22492_), .B(new_n22490_), .S0(new_n12689_), .Y(new_n22493_));
  OAI21X1  g20057(.A0(new_n22460_), .A1(new_n14395_), .B0(new_n22493_), .Y(new_n22494_));
  OAI21X1  g20058(.A0(new_n12567_), .A1(new_n12269_), .B0(new_n22462_), .Y(new_n22495_));
  AOI21X1  g20059(.A0(new_n13673_), .A1(new_n8009_), .B0(pi0038), .Y(new_n22496_));
  OAI21X1  g20060(.A0(new_n13671_), .A1(new_n8009_), .B0(new_n22496_), .Y(new_n22497_));
  AND2X1   g20061(.A(new_n22497_), .B(new_n22495_), .Y(new_n22498_));
  OR4X1    g20062(.A(new_n22498_), .B(new_n3125_), .C(new_n3124_), .D(pi0606), .Y(new_n22499_));
  NOR2X1   g20063(.A(new_n12401_), .B(new_n2959_), .Y(new_n22500_));
  OAI21X1  g20064(.A0(new_n22500_), .A1(new_n13682_), .B0(new_n8009_), .Y(new_n22501_));
  OAI21X1  g20065(.A0(new_n13691_), .A1(new_n13690_), .B0(pi0200), .Y(new_n22502_));
  AOI21X1  g20066(.A0(new_n13686_), .A1(new_n8009_), .B0(pi0038), .Y(new_n22503_));
  NOR3X1   g20067(.A(new_n13692_), .B(new_n8009_), .C(new_n2996_), .Y(new_n22504_));
  OR4X1    g20068(.A(new_n22504_), .B(new_n3125_), .C(new_n3124_), .D(new_n22432_), .Y(new_n22505_));
  AOI21X1  g20069(.A0(new_n22503_), .A1(new_n22502_), .B0(new_n22505_), .Y(new_n22506_));
  AOI21X1  g20070(.A0(new_n22506_), .A1(new_n22501_), .B0(new_n22438_), .Y(new_n22507_));
  AOI21X1  g20071(.A0(new_n22507_), .A1(new_n22499_), .B0(new_n22461_), .Y(new_n22508_));
  AOI21X1  g20072(.A0(new_n22440_), .A1(new_n22461_), .B0(new_n22508_), .Y(new_n22509_));
  INVX1    g20073(.A(new_n22509_), .Y(new_n22510_));
  INVX1    g20074(.A(new_n22440_), .Y(new_n22511_));
  AOI21X1  g20075(.A0(new_n22511_), .A1(pi0625), .B0(pi1153), .Y(new_n22512_));
  OAI21X1  g20076(.A0(new_n22510_), .A1(pi0625), .B0(new_n22512_), .Y(new_n22513_));
  AND2X1   g20077(.A(new_n22477_), .B(new_n12584_), .Y(new_n22514_));
  AOI21X1  g20078(.A0(new_n22511_), .A1(new_n12493_), .B0(new_n12494_), .Y(new_n22515_));
  OAI21X1  g20079(.A0(new_n22510_), .A1(new_n12493_), .B0(new_n22515_), .Y(new_n22516_));
  AND2X1   g20080(.A(new_n22479_), .B(pi0608), .Y(new_n22517_));
  AOI22X1  g20081(.A0(new_n22517_), .A1(new_n22516_), .B0(new_n22514_), .B1(new_n22513_), .Y(new_n22518_));
  MX2X1    g20082(.A(new_n22518_), .B(new_n22510_), .S0(new_n11889_), .Y(new_n22519_));
  INVX1    g20083(.A(new_n22519_), .Y(new_n22520_));
  OAI21X1  g20084(.A0(new_n22482_), .A1(new_n12590_), .B0(new_n12591_), .Y(new_n22521_));
  AOI21X1  g20085(.A0(new_n22520_), .A1(new_n12590_), .B0(new_n22521_), .Y(new_n22522_));
  NAND2X1  g20086(.A(new_n22443_), .B(new_n12596_), .Y(new_n22523_));
  OAI21X1  g20087(.A0(new_n22482_), .A1(pi0609), .B0(pi1155), .Y(new_n22524_));
  AOI21X1  g20088(.A0(new_n22520_), .A1(pi0609), .B0(new_n22524_), .Y(new_n22525_));
  NAND2X1  g20089(.A(new_n22445_), .B(pi0660), .Y(new_n22526_));
  OAI22X1  g20090(.A0(new_n22526_), .A1(new_n22525_), .B0(new_n22523_), .B1(new_n22522_), .Y(new_n22527_));
  MX2X1    g20091(.A(new_n22527_), .B(new_n22520_), .S0(new_n11888_), .Y(new_n22528_));
  AOI21X1  g20092(.A0(new_n22484_), .A1(pi0618), .B0(pi1154), .Y(new_n22529_));
  INVX1    g20093(.A(new_n22529_), .Y(new_n22530_));
  AOI21X1  g20094(.A0(new_n22528_), .A1(new_n12614_), .B0(new_n22530_), .Y(new_n22531_));
  NOR2X1   g20095(.A(new_n22449_), .B(pi0627), .Y(new_n22532_));
  INVX1    g20096(.A(new_n22532_), .Y(new_n22533_));
  AOI21X1  g20097(.A0(new_n22484_), .A1(new_n12614_), .B0(new_n12615_), .Y(new_n22534_));
  INVX1    g20098(.A(new_n22534_), .Y(new_n22535_));
  AOI21X1  g20099(.A0(new_n22528_), .A1(pi0618), .B0(new_n22535_), .Y(new_n22536_));
  NOR2X1   g20100(.A(new_n22451_), .B(new_n12622_), .Y(new_n22537_));
  INVX1    g20101(.A(new_n22537_), .Y(new_n22538_));
  OAI22X1  g20102(.A0(new_n22538_), .A1(new_n22536_), .B0(new_n22533_), .B1(new_n22531_), .Y(new_n22539_));
  MX2X1    g20103(.A(new_n22539_), .B(new_n22528_), .S0(new_n11887_), .Y(new_n22540_));
  OAI21X1  g20104(.A0(new_n22486_), .A1(new_n12637_), .B0(new_n12638_), .Y(new_n22541_));
  AOI21X1  g20105(.A0(new_n22540_), .A1(new_n12637_), .B0(new_n22541_), .Y(new_n22542_));
  NOR3X1   g20106(.A(new_n22542_), .B(new_n22455_), .C(pi0648), .Y(new_n22543_));
  OAI21X1  g20107(.A0(new_n22486_), .A1(pi0619), .B0(pi1159), .Y(new_n22544_));
  AOI21X1  g20108(.A0(new_n22540_), .A1(pi0619), .B0(new_n22544_), .Y(new_n22545_));
  OR2X1    g20109(.A(new_n22457_), .B(new_n12645_), .Y(new_n22546_));
  OAI21X1  g20110(.A0(new_n22546_), .A1(new_n22545_), .B0(pi0789), .Y(new_n22547_));
  OR2X1    g20111(.A(new_n22540_), .B(pi0789), .Y(new_n22548_));
  AND2X1   g20112(.A(new_n22548_), .B(new_n12842_), .Y(new_n22549_));
  OAI21X1  g20113(.A0(new_n22547_), .A1(new_n22543_), .B0(new_n22549_), .Y(new_n22550_));
  AOI21X1  g20114(.A0(new_n22430_), .A1(pi0626), .B0(new_n16352_), .Y(new_n22551_));
  OAI21X1  g20115(.A0(new_n22459_), .A1(pi0626), .B0(new_n22551_), .Y(new_n22552_));
  AOI21X1  g20116(.A0(new_n22430_), .A1(new_n12664_), .B0(new_n16356_), .Y(new_n22553_));
  OAI21X1  g20117(.A0(new_n22459_), .A1(new_n12664_), .B0(new_n22553_), .Y(new_n22554_));
  OR2X1    g20118(.A(new_n22487_), .B(new_n12770_), .Y(new_n22555_));
  NAND3X1  g20119(.A(new_n22555_), .B(new_n22554_), .C(new_n22552_), .Y(new_n22556_));
  AOI21X1  g20120(.A0(new_n22556_), .A1(pi0788), .B0(new_n14273_), .Y(new_n22557_));
  AOI22X1  g20121(.A0(new_n22557_), .A1(new_n22550_), .B0(new_n22494_), .B1(pi0792), .Y(new_n22558_));
  NAND2X1  g20122(.A(new_n22430_), .B(new_n12711_), .Y(new_n22559_));
  OAI21X1  g20123(.A0(new_n22460_), .A1(new_n12711_), .B0(new_n22559_), .Y(new_n22560_));
  NAND2X1  g20124(.A(new_n22560_), .B(new_n14385_), .Y(new_n22561_));
  AOI21X1  g20125(.A0(new_n22492_), .A1(new_n22490_), .B0(new_n11884_), .Y(new_n22562_));
  AOI21X1  g20126(.A0(new_n22488_), .A1(new_n11884_), .B0(new_n22562_), .Y(new_n22563_));
  MX2X1    g20127(.A(new_n22563_), .B(new_n22431_), .S0(new_n12705_), .Y(new_n22564_));
  INVX1    g20128(.A(new_n22564_), .Y(new_n22565_));
  AOI21X1  g20129(.A0(new_n22431_), .A1(pi0647), .B0(pi1157), .Y(new_n22566_));
  INVX1    g20130(.A(new_n22566_), .Y(new_n22567_));
  AOI21X1  g20131(.A0(new_n22563_), .A1(new_n12705_), .B0(new_n22567_), .Y(new_n22568_));
  AOI22X1  g20132(.A0(new_n22568_), .A1(pi0630), .B0(new_n22565_), .B1(new_n14386_), .Y(new_n22569_));
  AND2X1   g20133(.A(new_n22569_), .B(new_n22561_), .Y(new_n22570_));
  OAI22X1  g20134(.A0(new_n22570_), .A1(new_n11883_), .B0(new_n22558_), .B1(new_n14269_), .Y(new_n22571_));
  AOI21X1  g20135(.A0(new_n22565_), .A1(pi1157), .B0(new_n22568_), .Y(new_n22572_));
  MX2X1    g20136(.A(new_n22572_), .B(new_n22563_), .S0(new_n11883_), .Y(new_n22573_));
  AOI21X1  g20137(.A0(new_n22573_), .A1(pi0644), .B0(pi0715), .Y(new_n22574_));
  OAI21X1  g20138(.A0(new_n22571_), .A1(pi0644), .B0(new_n22574_), .Y(new_n22575_));
  MX2X1    g20139(.A(new_n22560_), .B(new_n22430_), .S0(new_n12735_), .Y(new_n22576_));
  AOI21X1  g20140(.A0(new_n22431_), .A1(pi0644), .B0(new_n12739_), .Y(new_n22577_));
  OAI21X1  g20141(.A0(new_n22576_), .A1(pi0644), .B0(new_n22577_), .Y(new_n22578_));
  AND2X1   g20142(.A(new_n22578_), .B(new_n11882_), .Y(new_n22579_));
  AOI21X1  g20143(.A0(new_n22573_), .A1(new_n12743_), .B0(new_n12739_), .Y(new_n22580_));
  OAI21X1  g20144(.A0(new_n22571_), .A1(new_n12743_), .B0(new_n22580_), .Y(new_n22581_));
  AOI21X1  g20145(.A0(new_n22431_), .A1(new_n12743_), .B0(pi0715), .Y(new_n22582_));
  OAI21X1  g20146(.A0(new_n22576_), .A1(new_n12743_), .B0(new_n22582_), .Y(new_n22583_));
  AND2X1   g20147(.A(new_n22583_), .B(pi1160), .Y(new_n22584_));
  AOI22X1  g20148(.A0(new_n22584_), .A1(new_n22581_), .B0(new_n22579_), .B1(new_n22575_), .Y(new_n22585_));
  MX2X1    g20149(.A(new_n22585_), .B(new_n22571_), .S0(new_n12897_), .Y(new_n22586_));
  MX2X1    g20150(.A(new_n22586_), .B(pi0200), .S0(po1038), .Y(po0357));
  INVX1    g20151(.A(pi0201), .Y(new_n22588_));
  AND2X1   g20152(.A(pi0237), .B(pi0233), .Y(new_n22589_));
  INVX1    g20153(.A(new_n22589_), .Y(new_n22590_));
  AOI21X1  g20154(.A0(new_n5324_), .A1(pi0332), .B0(pi0059), .Y(new_n22591_));
  AOI21X1  g20155(.A0(pi0332), .A1(pi0074), .B0(pi0055), .Y(new_n22592_));
  MX2X1    g20156(.A(pi0587), .B(pi0947), .S0(pi0299), .Y(new_n22593_));
  MX2X1    g20157(.A(new_n22593_), .B(new_n5028_), .S0(pi0468), .Y(new_n22594_));
  NAND3X1  g20158(.A(new_n22594_), .B(new_n8313_), .C(new_n2507_), .Y(new_n22595_));
  AOI21X1  g20159(.A0(new_n22595_), .A1(new_n2445_), .B0(new_n5850_), .Y(new_n22596_));
  AOI21X1  g20160(.A0(new_n5359_), .A1(new_n3630_), .B0(pi0332), .Y(new_n22597_));
  OAI22X1  g20161(.A0(new_n22597_), .A1(new_n11269_), .B0(new_n3106_), .B1(new_n2445_), .Y(new_n22598_));
  OAI21X1  g20162(.A0(new_n22598_), .A1(new_n22596_), .B0(new_n4991_), .Y(new_n22599_));
  AND2X1   g20163(.A(new_n22599_), .B(new_n22592_), .Y(new_n22600_));
  NAND2X1  g20164(.A(new_n5331_), .B(new_n3130_), .Y(new_n22601_));
  OAI21X1  g20165(.A0(new_n22601_), .A1(new_n3074_), .B0(new_n2445_), .Y(new_n22602_));
  OAI21X1  g20166(.A0(new_n22602_), .A1(new_n3128_), .B0(new_n3148_), .Y(new_n22603_));
  OAI21X1  g20167(.A0(new_n22603_), .A1(new_n22600_), .B0(new_n22591_), .Y(new_n22604_));
  NAND2X1  g20168(.A(new_n22602_), .B(new_n5327_), .Y(new_n22605_));
  INVX1    g20169(.A(new_n5327_), .Y(new_n22606_));
  AOI21X1  g20170(.A0(new_n22606_), .A1(pi0332), .B0(new_n3153_), .Y(new_n22607_));
  AOI21X1  g20171(.A0(new_n22607_), .A1(new_n22605_), .B0(pi0057), .Y(new_n22608_));
  AOI22X1  g20172(.A0(new_n22608_), .A1(new_n22604_), .B0(pi0332), .B1(pi0057), .Y(new_n22609_));
  NOR2X1   g20173(.A(new_n5028_), .B(pi0332), .Y(new_n22610_));
  NOR2X1   g20174(.A(new_n22610_), .B(pi0947), .Y(new_n22611_));
  INVX1    g20175(.A(new_n22611_), .Y(new_n22612_));
  NOR3X1   g20176(.A(new_n2445_), .B(new_n2766_), .C(new_n2526_), .Y(new_n22613_));
  NOR2X1   g20177(.A(pi0841), .B(pi0070), .Y(new_n22614_));
  MX2X1    g20178(.A(new_n22614_), .B(pi0070), .S0(new_n2456_), .Y(new_n22615_));
  NOR2X1   g20179(.A(pi0096), .B(pi0032), .Y(new_n22616_));
  AOI21X1  g20180(.A0(new_n22616_), .A1(pi0070), .B0(pi0332), .Y(new_n22617_));
  INVX1    g20181(.A(new_n22617_), .Y(new_n22618_));
  AOI21X1  g20182(.A0(new_n22615_), .A1(new_n2766_), .B0(new_n22618_), .Y(new_n22619_));
  NOR2X1   g20183(.A(new_n22619_), .B(new_n22613_), .Y(new_n22620_));
  AOI21X1  g20184(.A0(new_n22620_), .A1(new_n5057_), .B0(new_n5367_), .Y(new_n22621_));
  NOR2X1   g20185(.A(new_n22621_), .B(new_n22612_), .Y(new_n22622_));
  MX2X1    g20186(.A(new_n22619_), .B(new_n2445_), .S0(pi0468), .Y(new_n22623_));
  AND2X1   g20187(.A(new_n22623_), .B(new_n5367_), .Y(new_n22624_));
  INVX1    g20188(.A(new_n22624_), .Y(new_n22625_));
  INVX1    g20189(.A(new_n22620_), .Y(new_n22626_));
  AOI21X1  g20190(.A0(new_n22626_), .A1(new_n5028_), .B0(new_n14590_), .Y(new_n22627_));
  AOI21X1  g20191(.A0(new_n22627_), .A1(new_n22625_), .B0(new_n22622_), .Y(new_n22628_));
  INVX1    g20192(.A(new_n22616_), .Y(new_n22629_));
  OR4X1    g20193(.A(new_n2710_), .B(new_n2709_), .C(pi0095), .D(pi0040), .Y(new_n22630_));
  AOI21X1  g20194(.A0(new_n22630_), .A1(new_n5134_), .B0(new_n22629_), .Y(new_n22631_));
  NOR2X1   g20195(.A(new_n22614_), .B(new_n2456_), .Y(new_n22632_));
  NOR3X1   g20196(.A(new_n22632_), .B(new_n2768_), .C(pi0095), .Y(new_n22633_));
  NAND3X1  g20197(.A(new_n22633_), .B(new_n2516_), .C(new_n2518_), .Y(new_n22634_));
  NOR4X1   g20198(.A(new_n22634_), .B(new_n2513_), .C(new_n2520_), .D(pi0093), .Y(new_n22635_));
  NOR2X1   g20199(.A(new_n22635_), .B(new_n22615_), .Y(new_n22636_));
  OAI21X1  g20200(.A0(new_n22636_), .A1(pi0210), .B0(new_n2445_), .Y(new_n22637_));
  AOI21X1  g20201(.A0(new_n22631_), .A1(pi0210), .B0(new_n22637_), .Y(new_n22638_));
  NOR2X1   g20202(.A(new_n22638_), .B(new_n22613_), .Y(new_n22639_));
  AOI21X1  g20203(.A0(new_n22639_), .A1(new_n5057_), .B0(new_n5367_), .Y(new_n22640_));
  NOR2X1   g20204(.A(new_n22640_), .B(new_n22612_), .Y(new_n22641_));
  MX2X1    g20205(.A(new_n22638_), .B(new_n2445_), .S0(pi0468), .Y(new_n22642_));
  AND2X1   g20206(.A(new_n22642_), .B(new_n5367_), .Y(new_n22643_));
  INVX1    g20207(.A(new_n22643_), .Y(new_n22644_));
  INVX1    g20208(.A(new_n22639_), .Y(new_n22645_));
  AOI21X1  g20209(.A0(new_n22645_), .A1(new_n5028_), .B0(new_n14590_), .Y(new_n22646_));
  AOI21X1  g20210(.A0(new_n22646_), .A1(new_n22644_), .B0(new_n22641_), .Y(new_n22647_));
  MX2X1    g20211(.A(new_n22647_), .B(new_n22628_), .S0(new_n3131_), .Y(new_n22648_));
  NAND2X1  g20212(.A(new_n22648_), .B(new_n5327_), .Y(new_n22649_));
  AOI21X1  g20213(.A0(new_n22628_), .A1(new_n22606_), .B0(new_n3153_), .Y(new_n22650_));
  AND2X1   g20214(.A(new_n2532_), .B(new_n2507_), .Y(new_n22651_));
  NOR3X1   g20215(.A(pi0095), .B(pi0072), .C(pi0040), .Y(new_n22652_));
  AOI21X1  g20216(.A0(new_n22652_), .A1(new_n22651_), .B0(pi0070), .Y(new_n22653_));
  OR2X1    g20217(.A(new_n22653_), .B(new_n22629_), .Y(new_n22654_));
  AOI21X1  g20218(.A0(new_n22651_), .A1(new_n22633_), .B0(new_n22615_), .Y(new_n22655_));
  INVX1    g20219(.A(new_n22655_), .Y(new_n22656_));
  AOI21X1  g20220(.A0(new_n22656_), .A1(new_n2766_), .B0(pi0332), .Y(new_n22657_));
  OAI21X1  g20221(.A0(new_n22654_), .A1(new_n2766_), .B0(new_n22657_), .Y(new_n22658_));
  INVX1    g20222(.A(new_n22658_), .Y(new_n22659_));
  NOR2X1   g20223(.A(new_n22659_), .B(new_n22613_), .Y(new_n22660_));
  NAND2X1  g20224(.A(new_n22660_), .B(new_n5057_), .Y(new_n22661_));
  AOI21X1  g20225(.A0(new_n22661_), .A1(new_n5028_), .B0(new_n22612_), .Y(new_n22662_));
  MX2X1    g20226(.A(new_n22659_), .B(new_n2445_), .S0(pi0468), .Y(new_n22663_));
  OAI21X1  g20227(.A0(new_n22660_), .A1(new_n5367_), .B0(pi0947), .Y(new_n22664_));
  AOI21X1  g20228(.A0(new_n22663_), .A1(new_n5367_), .B0(new_n22664_), .Y(new_n22665_));
  NOR3X1   g20229(.A(new_n22665_), .B(new_n22662_), .C(new_n2953_), .Y(new_n22666_));
  INVX1    g20230(.A(pi0587), .Y(new_n22667_));
  OAI21X1  g20231(.A0(new_n5028_), .A1(pi0332), .B0(new_n22667_), .Y(new_n22668_));
  AOI21X1  g20232(.A0(new_n22656_), .A1(new_n2973_), .B0(pi0332), .Y(new_n22669_));
  OAI21X1  g20233(.A0(new_n22654_), .A1(new_n2973_), .B0(new_n22669_), .Y(new_n22670_));
  AND2X1   g20234(.A(pi0198), .B(pi0096), .Y(new_n22671_));
  AND2X1   g20235(.A(new_n22671_), .B(pi0332), .Y(new_n22672_));
  INVX1    g20236(.A(new_n22672_), .Y(new_n22673_));
  NAND3X1  g20237(.A(new_n22673_), .B(new_n22670_), .C(new_n5057_), .Y(new_n22674_));
  AOI21X1  g20238(.A0(new_n22674_), .A1(new_n5028_), .B0(new_n22668_), .Y(new_n22675_));
  AOI21X1  g20239(.A0(new_n22673_), .A1(new_n22670_), .B0(new_n5367_), .Y(new_n22676_));
  AOI21X1  g20240(.A0(pi0468), .A1(pi0332), .B0(new_n5028_), .Y(new_n22677_));
  INVX1    g20241(.A(new_n22677_), .Y(new_n22678_));
  AOI21X1  g20242(.A0(new_n22670_), .A1(new_n5860_), .B0(new_n22678_), .Y(new_n22679_));
  NOR3X1   g20243(.A(new_n22679_), .B(new_n22676_), .C(new_n22667_), .Y(new_n22680_));
  NOR3X1   g20244(.A(new_n22680_), .B(new_n22675_), .C(pi0299), .Y(new_n22681_));
  OAI21X1  g20245(.A0(new_n22681_), .A1(new_n22666_), .B0(new_n5849_), .Y(new_n22682_));
  NOR2X1   g20246(.A(new_n22610_), .B(pi0587), .Y(new_n22683_));
  OAI21X1  g20247(.A0(new_n22636_), .A1(pi0198), .B0(new_n2445_), .Y(new_n22684_));
  AOI21X1  g20248(.A0(new_n22631_), .A1(pi0198), .B0(new_n22684_), .Y(new_n22685_));
  NOR3X1   g20249(.A(new_n22685_), .B(new_n22672_), .C(new_n5033_), .Y(new_n22686_));
  OAI21X1  g20250(.A0(new_n22686_), .A1(new_n5367_), .B0(new_n22683_), .Y(new_n22687_));
  OAI21X1  g20251(.A0(new_n22685_), .A1(new_n22672_), .B0(new_n5028_), .Y(new_n22688_));
  OAI21X1  g20252(.A0(new_n22685_), .A1(pi0468), .B0(new_n22677_), .Y(new_n22689_));
  NAND3X1  g20253(.A(new_n22689_), .B(new_n22688_), .C(pi0587), .Y(new_n22690_));
  AOI21X1  g20254(.A0(new_n22690_), .A1(new_n22687_), .B0(pi0299), .Y(new_n22691_));
  NOR2X1   g20255(.A(new_n22691_), .B(new_n11269_), .Y(new_n22692_));
  OAI21X1  g20256(.A0(new_n22647_), .A1(new_n2953_), .B0(new_n22692_), .Y(new_n22693_));
  AOI21X1  g20257(.A0(new_n22693_), .A1(new_n22682_), .B0(pi0074), .Y(new_n22694_));
  NOR2X1   g20258(.A(new_n22628_), .B(new_n2953_), .Y(new_n22695_));
  NAND2X1  g20259(.A(new_n22615_), .B(new_n2973_), .Y(new_n22696_));
  AOI21X1  g20260(.A0(new_n22696_), .A1(new_n22617_), .B0(new_n22672_), .Y(new_n22697_));
  AND2X1   g20261(.A(new_n22615_), .B(new_n2973_), .Y(new_n22698_));
  OAI21X1  g20262(.A0(new_n22698_), .A1(new_n22618_), .B0(new_n5340_), .Y(new_n22699_));
  OR2X1    g20263(.A(new_n5365_), .B(pi0299), .Y(new_n22700_));
  AOI21X1  g20264(.A0(new_n22699_), .A1(new_n22610_), .B0(new_n22700_), .Y(new_n22701_));
  OAI21X1  g20265(.A0(new_n22697_), .A1(new_n5367_), .B0(new_n22701_), .Y(new_n22702_));
  OAI21X1  g20266(.A0(new_n3107_), .A1(pi0074), .B0(new_n22702_), .Y(new_n22703_));
  OAI21X1  g20267(.A0(new_n22703_), .A1(new_n22695_), .B0(new_n3128_), .Y(new_n22704_));
  OR2X1    g20268(.A(new_n22648_), .B(new_n3128_), .Y(new_n22705_));
  AND2X1   g20269(.A(new_n22705_), .B(new_n3148_), .Y(new_n22706_));
  OAI21X1  g20270(.A0(new_n22704_), .A1(new_n22694_), .B0(new_n22706_), .Y(new_n22707_));
  AOI21X1  g20271(.A0(new_n22628_), .A1(new_n5324_), .B0(pi0059), .Y(new_n22708_));
  AOI22X1  g20272(.A0(new_n22708_), .A1(new_n22707_), .B0(new_n22650_), .B1(new_n22649_), .Y(new_n22709_));
  MX2X1    g20273(.A(new_n22709_), .B(new_n22628_), .S0(pi0057), .Y(new_n22710_));
  MX2X1    g20274(.A(new_n22710_), .B(new_n22609_), .S0(new_n22590_), .Y(new_n22711_));
  AOI21X1  g20275(.A0(new_n22671_), .A1(new_n5340_), .B0(new_n11777_), .Y(new_n22712_));
  AOI22X1  g20276(.A0(new_n6520_), .A1(new_n2953_), .B0(pi0210), .B1(pi0096), .Y(new_n22713_));
  NOR2X1   g20277(.A(new_n11776_), .B(new_n5331_), .Y(new_n22714_));
  NOR4X1   g20278(.A(new_n22714_), .B(new_n22713_), .C(new_n22712_), .D(new_n22590_), .Y(new_n22715_));
  MX2X1    g20279(.A(new_n22715_), .B(new_n22711_), .S0(new_n22588_), .Y(po0358));
  INVX1    g20280(.A(pi0202), .Y(new_n22717_));
  INVX1    g20281(.A(pi0233), .Y(new_n22718_));
  AND2X1   g20282(.A(pi0237), .B(new_n22718_), .Y(new_n22719_));
  INVX1    g20283(.A(new_n22719_), .Y(new_n22720_));
  MX2X1    g20284(.A(new_n22710_), .B(new_n22609_), .S0(new_n22720_), .Y(new_n22721_));
  NOR4X1   g20285(.A(new_n22720_), .B(new_n22714_), .C(new_n22713_), .D(new_n22712_), .Y(new_n22722_));
  MX2X1    g20286(.A(new_n22722_), .B(new_n22721_), .S0(new_n22717_), .Y(po0359));
  INVX1    g20287(.A(pi0203), .Y(new_n22724_));
  NOR2X1   g20288(.A(pi0237), .B(pi0233), .Y(new_n22725_));
  INVX1    g20289(.A(new_n22725_), .Y(new_n22726_));
  MX2X1    g20290(.A(new_n22710_), .B(new_n22609_), .S0(new_n22726_), .Y(new_n22727_));
  NOR4X1   g20291(.A(new_n22726_), .B(new_n22714_), .C(new_n22713_), .D(new_n22712_), .Y(new_n22728_));
  MX2X1    g20292(.A(new_n22728_), .B(new_n22727_), .S0(new_n22724_), .Y(po0360));
  MX2X1    g20293(.A(new_n5030_), .B(pi0602), .S0(new_n5860_), .Y(new_n22730_));
  MX2X1    g20294(.A(new_n22730_), .B(new_n5120_), .S0(pi0299), .Y(new_n22731_));
  AOI21X1  g20295(.A0(new_n22731_), .A1(new_n3630_), .B0(pi0332), .Y(new_n22732_));
  NOR2X1   g20296(.A(pi0602), .B(pi0299), .Y(new_n22733_));
  OAI21X1  g20297(.A0(pi0907), .A1(new_n2953_), .B0(new_n5860_), .Y(new_n22734_));
  OAI22X1  g20298(.A0(new_n22734_), .A1(new_n22733_), .B0(new_n5282_), .B1(new_n5860_), .Y(new_n22735_));
  NAND3X1  g20299(.A(new_n22735_), .B(new_n8313_), .C(new_n2507_), .Y(new_n22736_));
  AND2X1   g20300(.A(new_n22736_), .B(new_n2445_), .Y(new_n22737_));
  OAI22X1  g20301(.A0(new_n22737_), .A1(new_n5850_), .B0(new_n22732_), .B1(new_n11269_), .Y(new_n22738_));
  OAI21X1  g20302(.A0(new_n3106_), .A1(new_n2445_), .B0(new_n22592_), .Y(new_n22739_));
  AOI21X1  g20303(.A0(new_n22738_), .A1(new_n4991_), .B0(new_n22739_), .Y(new_n22740_));
  NAND2X1  g20304(.A(new_n5120_), .B(new_n3130_), .Y(new_n22741_));
  OAI21X1  g20305(.A0(new_n22741_), .A1(new_n3074_), .B0(new_n2445_), .Y(new_n22742_));
  OAI21X1  g20306(.A0(new_n22742_), .A1(new_n3128_), .B0(new_n3148_), .Y(new_n22743_));
  OAI21X1  g20307(.A0(new_n22743_), .A1(new_n22740_), .B0(new_n22591_), .Y(new_n22744_));
  NAND2X1  g20308(.A(new_n22742_), .B(new_n5327_), .Y(new_n22745_));
  AOI21X1  g20309(.A0(new_n22745_), .A1(new_n22607_), .B0(pi0057), .Y(new_n22746_));
  AOI22X1  g20310(.A0(new_n22746_), .A1(new_n22744_), .B0(pi0332), .B1(pi0057), .Y(new_n22747_));
  AOI21X1  g20311(.A0(new_n5282_), .A1(new_n2445_), .B0(pi0907), .Y(new_n22748_));
  INVX1    g20312(.A(new_n22748_), .Y(new_n22749_));
  AOI21X1  g20313(.A0(new_n22620_), .A1(new_n5057_), .B0(new_n5282_), .Y(new_n22750_));
  NOR2X1   g20314(.A(new_n22750_), .B(new_n22749_), .Y(new_n22751_));
  AND2X1   g20315(.A(new_n22623_), .B(new_n5282_), .Y(new_n22752_));
  INVX1    g20316(.A(new_n22752_), .Y(new_n22753_));
  AOI21X1  g20317(.A0(new_n22626_), .A1(new_n5030_), .B0(new_n5297_), .Y(new_n22754_));
  AOI21X1  g20318(.A0(new_n22754_), .A1(new_n22753_), .B0(new_n22751_), .Y(new_n22755_));
  AND2X1   g20319(.A(new_n22642_), .B(new_n5282_), .Y(new_n22756_));
  INVX1    g20320(.A(new_n22756_), .Y(new_n22757_));
  AOI21X1  g20321(.A0(new_n22645_), .A1(new_n5030_), .B0(new_n5297_), .Y(new_n22758_));
  AOI21X1  g20322(.A0(new_n12290_), .A1(pi0332), .B0(new_n5029_), .Y(new_n22759_));
  OAI21X1  g20323(.A0(new_n22645_), .A1(new_n5033_), .B0(new_n22759_), .Y(new_n22760_));
  AOI22X1  g20324(.A0(new_n22760_), .A1(new_n22748_), .B0(new_n22758_), .B1(new_n22757_), .Y(new_n22761_));
  MX2X1    g20325(.A(new_n22761_), .B(new_n22755_), .S0(new_n3131_), .Y(new_n22762_));
  NAND2X1  g20326(.A(new_n22762_), .B(new_n5327_), .Y(new_n22763_));
  AOI21X1  g20327(.A0(new_n22755_), .A1(new_n22606_), .B0(new_n3153_), .Y(new_n22764_));
  AOI21X1  g20328(.A0(new_n22671_), .A1(new_n5030_), .B0(new_n2445_), .Y(new_n22765_));
  NOR2X1   g20329(.A(new_n22765_), .B(pi0299), .Y(new_n22766_));
  OR2X1    g20330(.A(new_n22685_), .B(new_n22672_), .Y(new_n22767_));
  OR2X1    g20331(.A(new_n22767_), .B(new_n5275_), .Y(new_n22768_));
  AOI22X1  g20332(.A0(new_n22768_), .A1(new_n22766_), .B0(new_n22761_), .B1(pi0299), .Y(new_n22769_));
  OR2X1    g20333(.A(new_n22769_), .B(new_n11269_), .Y(new_n22770_));
  NAND3X1  g20334(.A(new_n22673_), .B(new_n22670_), .C(new_n5219_), .Y(new_n22771_));
  AND2X1   g20335(.A(new_n22771_), .B(new_n22766_), .Y(new_n22772_));
  AOI21X1  g20336(.A0(new_n22661_), .A1(new_n5030_), .B0(new_n22749_), .Y(new_n22773_));
  OAI21X1  g20337(.A0(new_n22660_), .A1(new_n5282_), .B0(pi0907), .Y(new_n22774_));
  AOI21X1  g20338(.A0(new_n22663_), .A1(new_n5282_), .B0(new_n22774_), .Y(new_n22775_));
  NOR3X1   g20339(.A(new_n22775_), .B(new_n22773_), .C(new_n2953_), .Y(new_n22776_));
  OAI21X1  g20340(.A0(new_n22776_), .A1(new_n22772_), .B0(new_n5849_), .Y(new_n22777_));
  AOI21X1  g20341(.A0(new_n22777_), .A1(new_n22770_), .B0(pi0074), .Y(new_n22778_));
  NOR2X1   g20342(.A(new_n22755_), .B(new_n2953_), .Y(new_n22779_));
  AOI21X1  g20343(.A0(new_n22730_), .A1(new_n22697_), .B0(new_n22765_), .Y(new_n22780_));
  OAI22X1  g20344(.A0(new_n22780_), .A1(pi0299), .B0(new_n3107_), .B1(pi0074), .Y(new_n22781_));
  OAI21X1  g20345(.A0(new_n22781_), .A1(new_n22779_), .B0(new_n3128_), .Y(new_n22782_));
  OR2X1    g20346(.A(new_n22762_), .B(new_n3128_), .Y(new_n22783_));
  AND2X1   g20347(.A(new_n22783_), .B(new_n3148_), .Y(new_n22784_));
  OAI21X1  g20348(.A0(new_n22782_), .A1(new_n22778_), .B0(new_n22784_), .Y(new_n22785_));
  AOI21X1  g20349(.A0(new_n22755_), .A1(new_n5324_), .B0(pi0059), .Y(new_n22786_));
  AOI22X1  g20350(.A0(new_n22786_), .A1(new_n22785_), .B0(new_n22764_), .B1(new_n22763_), .Y(new_n22787_));
  MX2X1    g20351(.A(new_n22787_), .B(new_n22755_), .S0(pi0057), .Y(new_n22788_));
  MX2X1    g20352(.A(new_n22788_), .B(new_n22747_), .S0(new_n22590_), .Y(new_n22789_));
  AOI21X1  g20353(.A0(new_n22671_), .A1(new_n5219_), .B0(new_n11777_), .Y(new_n22790_));
  NOR2X1   g20354(.A(new_n11776_), .B(new_n5120_), .Y(new_n22791_));
  NOR4X1   g20355(.A(new_n22791_), .B(new_n22790_), .C(new_n22713_), .D(new_n22590_), .Y(new_n22792_));
  MX2X1    g20356(.A(new_n22789_), .B(new_n22792_), .S0(pi0204), .Y(po0361));
  MX2X1    g20357(.A(new_n22788_), .B(new_n22747_), .S0(new_n22720_), .Y(new_n22794_));
  NOR4X1   g20358(.A(new_n22791_), .B(new_n22790_), .C(new_n22720_), .D(new_n22713_), .Y(new_n22795_));
  MX2X1    g20359(.A(new_n22794_), .B(new_n22795_), .S0(pi0205), .Y(po0362));
  INVX1    g20360(.A(pi0237), .Y(new_n22797_));
  AND2X1   g20361(.A(new_n22797_), .B(pi0233), .Y(new_n22798_));
  INVX1    g20362(.A(new_n22798_), .Y(new_n22799_));
  MX2X1    g20363(.A(new_n22788_), .B(new_n22747_), .S0(new_n22799_), .Y(new_n22800_));
  NOR4X1   g20364(.A(new_n22799_), .B(new_n22791_), .C(new_n22790_), .D(new_n22713_), .Y(new_n22801_));
  MX2X1    g20365(.A(new_n22800_), .B(new_n22801_), .S0(pi0206), .Y(po0363));
  INVX1    g20366(.A(pi0207), .Y(new_n22803_));
  OR2X1    g20367(.A(new_n12574_), .B(new_n3810_), .Y(new_n22804_));
  AOI21X1  g20368(.A0(new_n13704_), .A1(new_n3129_), .B0(new_n12601_), .Y(new_n22805_));
  AOI21X1  g20369(.A0(new_n12601_), .A1(new_n22804_), .B0(new_n22805_), .Y(new_n22806_));
  AOI22X1  g20370(.A0(new_n22805_), .A1(new_n12590_), .B0(new_n13436_), .B1(new_n22804_), .Y(new_n22807_));
  AOI22X1  g20371(.A0(new_n22805_), .A1(pi0609), .B0(new_n13430_), .B1(new_n22804_), .Y(new_n22808_));
  MX2X1    g20372(.A(new_n22808_), .B(new_n22807_), .S0(new_n12591_), .Y(new_n22809_));
  MX2X1    g20373(.A(new_n22809_), .B(new_n22806_), .S0(new_n11888_), .Y(new_n22810_));
  OR2X1    g20374(.A(new_n22810_), .B(pi0781), .Y(new_n22811_));
  OAI21X1  g20375(.A0(new_n22804_), .A1(new_n12614_), .B0(new_n12615_), .Y(new_n22812_));
  AOI21X1  g20376(.A0(new_n22810_), .A1(new_n12614_), .B0(new_n22812_), .Y(new_n22813_));
  OAI21X1  g20377(.A0(new_n22804_), .A1(pi0618), .B0(pi1154), .Y(new_n22814_));
  AOI21X1  g20378(.A0(new_n22810_), .A1(pi0618), .B0(new_n22814_), .Y(new_n22815_));
  OAI21X1  g20379(.A0(new_n22815_), .A1(new_n22813_), .B0(pi0781), .Y(new_n22816_));
  AND2X1   g20380(.A(new_n22816_), .B(new_n22811_), .Y(new_n22817_));
  INVX1    g20381(.A(new_n22817_), .Y(new_n22818_));
  INVX1    g20382(.A(new_n22804_), .Y(new_n22819_));
  AOI21X1  g20383(.A0(new_n22819_), .A1(pi0619), .B0(pi1159), .Y(new_n22820_));
  OAI21X1  g20384(.A0(new_n22818_), .A1(pi0619), .B0(new_n22820_), .Y(new_n22821_));
  AOI21X1  g20385(.A0(new_n22819_), .A1(new_n12637_), .B0(new_n12638_), .Y(new_n22822_));
  OAI21X1  g20386(.A0(new_n22818_), .A1(new_n12637_), .B0(new_n22822_), .Y(new_n22823_));
  AND2X1   g20387(.A(new_n22823_), .B(new_n22821_), .Y(new_n22824_));
  MX2X1    g20388(.A(new_n22824_), .B(new_n22817_), .S0(new_n11886_), .Y(new_n22825_));
  NOR3X1   g20389(.A(new_n14175_), .B(new_n12574_), .C(new_n3810_), .Y(new_n22826_));
  AOI21X1  g20390(.A0(new_n22825_), .A1(new_n14175_), .B0(new_n22826_), .Y(new_n22827_));
  MX2X1    g20391(.A(new_n22827_), .B(new_n22804_), .S0(new_n12711_), .Y(new_n22828_));
  NOR2X1   g20392(.A(new_n22828_), .B(pi0207), .Y(new_n22829_));
  INVX1    g20393(.A(new_n16746_), .Y(new_n22830_));
  NOR4X1   g20394(.A(new_n22830_), .B(new_n14178_), .C(new_n12601_), .D(new_n3810_), .Y(new_n22831_));
  INVX1    g20395(.A(new_n22831_), .Y(new_n22832_));
  NOR4X1   g20396(.A(new_n22832_), .B(new_n14183_), .C(new_n14180_), .D(new_n12841_), .Y(new_n22833_));
  AND2X1   g20397(.A(new_n22833_), .B(new_n14123_), .Y(new_n22834_));
  OAI21X1  g20398(.A0(new_n22834_), .A1(new_n22803_), .B0(pi0623), .Y(new_n22835_));
  AOI21X1  g20399(.A0(new_n13699_), .A1(new_n3129_), .B0(pi0207), .Y(new_n22836_));
  INVX1    g20400(.A(new_n22836_), .Y(new_n22837_));
  OAI22X1  g20401(.A0(new_n22837_), .A1(pi0623), .B0(new_n22835_), .B1(new_n22829_), .Y(new_n22838_));
  OR2X1    g20402(.A(new_n22838_), .B(new_n14384_), .Y(new_n22839_));
  INVX1    g20403(.A(pi0710), .Y(new_n22840_));
  NOR4X1   g20404(.A(new_n16715_), .B(new_n13639_), .C(new_n13624_), .D(new_n13569_), .Y(new_n22841_));
  INVX1    g20405(.A(new_n12869_), .Y(new_n22842_));
  OAI21X1  g20406(.A0(new_n16716_), .A1(new_n3810_), .B0(new_n11889_), .Y(new_n22843_));
  OAI21X1  g20407(.A0(new_n12574_), .A1(new_n3810_), .B0(new_n12493_), .Y(new_n22844_));
  OAI21X1  g20408(.A0(new_n16716_), .A1(new_n3810_), .B0(pi0625), .Y(new_n22845_));
  AOI21X1  g20409(.A0(new_n22845_), .A1(new_n22844_), .B0(new_n12494_), .Y(new_n22846_));
  OAI21X1  g20410(.A0(new_n12574_), .A1(new_n3810_), .B0(pi0625), .Y(new_n22847_));
  OAI21X1  g20411(.A0(new_n16716_), .A1(new_n3810_), .B0(new_n12493_), .Y(new_n22848_));
  AOI21X1  g20412(.A0(new_n22848_), .A1(new_n22847_), .B0(pi1153), .Y(new_n22849_));
  OAI21X1  g20413(.A0(new_n22849_), .A1(new_n22846_), .B0(pi0778), .Y(new_n22850_));
  NAND2X1  g20414(.A(new_n22850_), .B(new_n22843_), .Y(new_n22851_));
  MX2X1    g20415(.A(new_n22851_), .B(new_n22804_), .S0(new_n12618_), .Y(new_n22852_));
  MX2X1    g20416(.A(new_n22852_), .B(new_n22804_), .S0(new_n12641_), .Y(new_n22853_));
  INVX1    g20417(.A(new_n22853_), .Y(new_n22854_));
  MX2X1    g20418(.A(new_n22854_), .B(new_n22819_), .S0(new_n12659_), .Y(new_n22855_));
  NOR3X1   g20419(.A(new_n17252_), .B(new_n12574_), .C(new_n3810_), .Y(new_n22856_));
  AOI21X1  g20420(.A0(new_n22855_), .A1(new_n17252_), .B0(new_n22856_), .Y(new_n22857_));
  OAI22X1  g20421(.A0(new_n22857_), .A1(new_n13639_), .B0(new_n22842_), .B1(new_n22804_), .Y(new_n22858_));
  INVX1    g20422(.A(new_n22858_), .Y(new_n22859_));
  MX2X1    g20423(.A(new_n22859_), .B(new_n22841_), .S0(pi0207), .Y(new_n22860_));
  MX2X1    g20424(.A(new_n22860_), .B(new_n22836_), .S0(new_n22840_), .Y(new_n22861_));
  INVX1    g20425(.A(new_n22861_), .Y(new_n22862_));
  AOI21X1  g20426(.A0(new_n22836_), .A1(pi0647), .B0(pi1157), .Y(new_n22863_));
  OAI21X1  g20427(.A0(new_n22862_), .A1(pi0647), .B0(new_n22863_), .Y(new_n22864_));
  AOI21X1  g20428(.A0(new_n22836_), .A1(new_n12705_), .B0(new_n12706_), .Y(new_n22865_));
  OAI21X1  g20429(.A0(new_n22862_), .A1(new_n12705_), .B0(new_n22865_), .Y(new_n22866_));
  MX2X1    g20430(.A(new_n22866_), .B(new_n22864_), .S0(pi0630), .Y(new_n22867_));
  AOI21X1  g20431(.A0(new_n22867_), .A1(new_n22839_), .B0(new_n11883_), .Y(new_n22868_));
  AOI21X1  g20432(.A0(new_n13699_), .A1(new_n3129_), .B0(pi0628), .Y(new_n22869_));
  AND2X1   g20433(.A(new_n22857_), .B(pi0628), .Y(new_n22870_));
  AOI21X1  g20434(.A0(new_n22870_), .A1(new_n12689_), .B0(new_n22869_), .Y(new_n22871_));
  NOR2X1   g20435(.A(new_n22871_), .B(new_n12684_), .Y(new_n22872_));
  OAI21X1  g20436(.A0(new_n12574_), .A1(new_n3810_), .B0(pi0628), .Y(new_n22873_));
  MX2X1    g20437(.A(new_n22857_), .B(new_n22804_), .S0(pi0628), .Y(new_n22874_));
  INVX1    g20438(.A(new_n22874_), .Y(new_n22875_));
  OAI22X1  g20439(.A0(new_n22875_), .A1(new_n12710_), .B0(new_n22873_), .B1(pi1156), .Y(new_n22876_));
  OAI21X1  g20440(.A0(new_n22876_), .A1(new_n22872_), .B0(pi0792), .Y(new_n22877_));
  OAI21X1  g20441(.A0(new_n13672_), .A1(new_n3810_), .B0(new_n11889_), .Y(new_n22878_));
  OAI21X1  g20442(.A0(new_n13672_), .A1(new_n3810_), .B0(new_n12493_), .Y(new_n22879_));
  AOI21X1  g20443(.A0(new_n22879_), .A1(new_n22847_), .B0(pi1153), .Y(new_n22880_));
  NOR3X1   g20444(.A(new_n22880_), .B(new_n22846_), .C(pi0608), .Y(new_n22881_));
  OAI21X1  g20445(.A0(new_n13672_), .A1(new_n3810_), .B0(pi0625), .Y(new_n22882_));
  AOI21X1  g20446(.A0(new_n22882_), .A1(new_n22844_), .B0(new_n12494_), .Y(new_n22883_));
  NOR3X1   g20447(.A(new_n22883_), .B(new_n22849_), .C(new_n12584_), .Y(new_n22884_));
  OR2X1    g20448(.A(new_n22884_), .B(new_n11889_), .Y(new_n22885_));
  OAI21X1  g20449(.A0(new_n22885_), .A1(new_n22881_), .B0(new_n22878_), .Y(new_n22886_));
  MX2X1    g20450(.A(new_n22886_), .B(new_n22851_), .S0(pi0609), .Y(new_n22887_));
  AOI21X1  g20451(.A0(new_n22804_), .A1(pi1155), .B0(pi0660), .Y(new_n22888_));
  INVX1    g20452(.A(new_n22888_), .Y(new_n22889_));
  AOI21X1  g20453(.A0(new_n22887_), .A1(new_n12591_), .B0(new_n22889_), .Y(new_n22890_));
  MX2X1    g20454(.A(new_n22886_), .B(new_n22851_), .S0(new_n12590_), .Y(new_n22891_));
  AOI21X1  g20455(.A0(new_n22804_), .A1(new_n12591_), .B0(new_n12596_), .Y(new_n22892_));
  INVX1    g20456(.A(new_n22892_), .Y(new_n22893_));
  AOI21X1  g20457(.A0(new_n22891_), .A1(pi1155), .B0(new_n22893_), .Y(new_n22894_));
  OAI21X1  g20458(.A0(new_n22894_), .A1(new_n22890_), .B0(pi0785), .Y(new_n22895_));
  OAI21X1  g20459(.A0(new_n22886_), .A1(pi0785), .B0(new_n22895_), .Y(new_n22896_));
  INVX1    g20460(.A(new_n22852_), .Y(new_n22897_));
  MX2X1    g20461(.A(new_n22896_), .B(new_n22897_), .S0(pi0618), .Y(new_n22898_));
  AOI21X1  g20462(.A0(new_n22804_), .A1(pi1154), .B0(pi0627), .Y(new_n22899_));
  OAI21X1  g20463(.A0(new_n22898_), .A1(pi1154), .B0(new_n22899_), .Y(new_n22900_));
  MX2X1    g20464(.A(new_n22896_), .B(new_n22897_), .S0(new_n12614_), .Y(new_n22901_));
  AOI21X1  g20465(.A0(new_n22804_), .A1(new_n12615_), .B0(new_n12622_), .Y(new_n22902_));
  OAI21X1  g20466(.A0(new_n22901_), .A1(new_n12615_), .B0(new_n22902_), .Y(new_n22903_));
  NAND2X1  g20467(.A(new_n22903_), .B(new_n22900_), .Y(new_n22904_));
  MX2X1    g20468(.A(new_n22904_), .B(new_n22896_), .S0(new_n11887_), .Y(new_n22905_));
  MX2X1    g20469(.A(new_n22905_), .B(new_n22854_), .S0(pi0619), .Y(new_n22906_));
  AOI21X1  g20470(.A0(new_n22804_), .A1(pi1159), .B0(pi0648), .Y(new_n22907_));
  OAI21X1  g20471(.A0(new_n22906_), .A1(pi1159), .B0(new_n22907_), .Y(new_n22908_));
  MX2X1    g20472(.A(new_n22905_), .B(new_n22854_), .S0(new_n12637_), .Y(new_n22909_));
  AOI21X1  g20473(.A0(new_n22804_), .A1(new_n12638_), .B0(new_n12645_), .Y(new_n22910_));
  OAI21X1  g20474(.A0(new_n22909_), .A1(new_n12638_), .B0(new_n22910_), .Y(new_n22911_));
  AOI21X1  g20475(.A0(new_n22911_), .A1(new_n22908_), .B0(new_n11886_), .Y(new_n22912_));
  AOI21X1  g20476(.A0(new_n22905_), .A1(new_n11886_), .B0(new_n22912_), .Y(new_n22913_));
  AOI21X1  g20477(.A0(new_n22855_), .A1(pi0626), .B0(pi0641), .Y(new_n22914_));
  OAI21X1  g20478(.A0(new_n22913_), .A1(pi0626), .B0(new_n22914_), .Y(new_n22915_));
  AOI21X1  g20479(.A0(new_n22804_), .A1(pi0641), .B0(pi1158), .Y(new_n22916_));
  AOI21X1  g20480(.A0(new_n22855_), .A1(new_n12664_), .B0(new_n12672_), .Y(new_n22917_));
  OAI21X1  g20481(.A0(new_n22913_), .A1(new_n12664_), .B0(new_n22917_), .Y(new_n22918_));
  AOI21X1  g20482(.A0(new_n22804_), .A1(new_n12672_), .B0(new_n12676_), .Y(new_n22919_));
  AOI22X1  g20483(.A0(new_n22919_), .A1(new_n22918_), .B0(new_n22916_), .B1(new_n22915_), .Y(new_n22920_));
  OR2X1    g20484(.A(new_n22913_), .B(pi0788), .Y(new_n22921_));
  AND2X1   g20485(.A(new_n22921_), .B(new_n16350_), .Y(new_n22922_));
  OAI21X1  g20486(.A0(new_n22920_), .A1(new_n11885_), .B0(new_n22922_), .Y(new_n22923_));
  AOI21X1  g20487(.A0(new_n22923_), .A1(new_n22877_), .B0(pi0207), .Y(new_n22924_));
  INVX1    g20488(.A(pi0623), .Y(new_n22925_));
  NOR3X1   g20489(.A(new_n16715_), .B(new_n13624_), .C(new_n13569_), .Y(new_n22926_));
  NAND3X1  g20490(.A(new_n16793_), .B(new_n3129_), .C(new_n12493_), .Y(new_n22927_));
  NOR4X1   g20491(.A(new_n16714_), .B(new_n12567_), .C(new_n3810_), .D(new_n12493_), .Y(new_n22928_));
  OAI21X1  g20492(.A0(new_n22928_), .A1(new_n12494_), .B0(new_n12584_), .Y(new_n22929_));
  AOI21X1  g20493(.A0(new_n22927_), .A1(new_n12494_), .B0(new_n22929_), .Y(new_n22930_));
  AOI21X1  g20494(.A0(new_n22284_), .A1(pi0625), .B0(new_n12494_), .Y(new_n22931_));
  NOR4X1   g20495(.A(new_n16714_), .B(new_n12567_), .C(new_n3810_), .D(pi0625), .Y(new_n22932_));
  OAI21X1  g20496(.A0(new_n22932_), .A1(pi1153), .B0(pi0608), .Y(new_n22933_));
  OAI21X1  g20497(.A0(new_n22933_), .A1(new_n22931_), .B0(pi0778), .Y(new_n22934_));
  OAI22X1  g20498(.A0(new_n22934_), .A1(new_n22930_), .B0(new_n22284_), .B1(pi0778), .Y(new_n22935_));
  NOR4X1   g20499(.A(new_n16714_), .B(new_n13569_), .C(new_n12567_), .D(new_n3810_), .Y(new_n22936_));
  OAI21X1  g20500(.A0(new_n22936_), .A1(new_n12590_), .B0(new_n12617_), .Y(new_n22937_));
  AOI21X1  g20501(.A0(new_n22935_), .A1(new_n12590_), .B0(new_n22937_), .Y(new_n22938_));
  OAI21X1  g20502(.A0(new_n22936_), .A1(pi0609), .B0(new_n12616_), .Y(new_n22939_));
  AOI21X1  g20503(.A0(new_n22935_), .A1(pi0609), .B0(new_n22939_), .Y(new_n22940_));
  OR2X1    g20504(.A(new_n22940_), .B(new_n22938_), .Y(new_n22941_));
  NOR2X1   g20505(.A(new_n22935_), .B(pi0785), .Y(new_n22942_));
  AOI21X1  g20506(.A0(new_n22941_), .A1(pi0785), .B0(new_n22942_), .Y(new_n22943_));
  AND2X1   g20507(.A(new_n22943_), .B(new_n12614_), .Y(new_n22944_));
  AOI21X1  g20508(.A0(new_n22936_), .A1(new_n13598_), .B0(new_n12614_), .Y(new_n22945_));
  OR4X1    g20509(.A(new_n22945_), .B(new_n22944_), .C(pi1154), .D(pi0627), .Y(new_n22946_));
  AND2X1   g20510(.A(new_n22936_), .B(new_n13598_), .Y(new_n22947_));
  OAI21X1  g20511(.A0(new_n22947_), .A1(pi0618), .B0(new_n12639_), .Y(new_n22948_));
  AOI21X1  g20512(.A0(new_n22943_), .A1(pi0618), .B0(new_n22948_), .Y(new_n22949_));
  NOR2X1   g20513(.A(new_n22949_), .B(new_n11887_), .Y(new_n22950_));
  AOI21X1  g20514(.A0(new_n22943_), .A1(new_n11887_), .B0(new_n16248_), .Y(new_n22951_));
  INVX1    g20515(.A(new_n22951_), .Y(new_n22952_));
  AOI21X1  g20516(.A0(new_n22950_), .A1(new_n22946_), .B0(new_n22952_), .Y(new_n22953_));
  NOR4X1   g20517(.A(new_n16715_), .B(new_n13569_), .C(new_n12641_), .D(new_n12618_), .Y(new_n22954_));
  AND2X1   g20518(.A(new_n14180_), .B(new_n12658_), .Y(new_n22955_));
  AOI21X1  g20519(.A0(new_n22955_), .A1(new_n22954_), .B0(new_n22953_), .Y(new_n22956_));
  INVX1    g20520(.A(new_n22956_), .Y(new_n22957_));
  NAND4X1  g20521(.A(new_n22936_), .B(new_n22011_), .C(new_n14198_), .D(new_n13598_), .Y(new_n22958_));
  AOI21X1  g20522(.A0(new_n22958_), .A1(pi0626), .B0(pi0641), .Y(new_n22959_));
  AND2X1   g20523(.A(new_n22959_), .B(new_n12676_), .Y(new_n22960_));
  OAI21X1  g20524(.A0(new_n22957_), .A1(pi0626), .B0(new_n22960_), .Y(new_n22961_));
  AOI21X1  g20525(.A0(new_n22958_), .A1(new_n12664_), .B0(new_n12672_), .Y(new_n22962_));
  AND2X1   g20526(.A(new_n22962_), .B(pi1158), .Y(new_n22963_));
  OAI21X1  g20527(.A0(new_n22957_), .A1(new_n12664_), .B0(new_n22963_), .Y(new_n22964_));
  NAND3X1  g20528(.A(new_n22964_), .B(new_n22961_), .C(pi0788), .Y(new_n22965_));
  AOI21X1  g20529(.A0(new_n22956_), .A1(new_n11885_), .B0(new_n14273_), .Y(new_n22966_));
  NOR3X1   g20530(.A(new_n12867_), .B(new_n12865_), .C(new_n14123_), .Y(new_n22967_));
  AOI22X1  g20531(.A0(new_n22967_), .A1(new_n22926_), .B0(new_n22966_), .B1(new_n22965_), .Y(new_n22968_));
  OAI21X1  g20532(.A0(new_n22968_), .A1(new_n22803_), .B0(new_n22925_), .Y(new_n22969_));
  OR4X1    g20533(.A(new_n13693_), .B(new_n13690_), .C(new_n3125_), .D(new_n3124_), .Y(new_n22970_));
  AND2X1   g20534(.A(new_n13704_), .B(new_n3129_), .Y(new_n22971_));
  OAI21X1  g20535(.A0(new_n22970_), .A1(new_n12493_), .B0(pi1153), .Y(new_n22972_));
  AOI21X1  g20536(.A0(new_n22971_), .A1(new_n12493_), .B0(new_n22972_), .Y(new_n22973_));
  NOR3X1   g20537(.A(new_n22973_), .B(new_n22849_), .C(new_n12584_), .Y(new_n22974_));
  OAI21X1  g20538(.A0(new_n22970_), .A1(pi0625), .B0(new_n12494_), .Y(new_n22975_));
  AOI21X1  g20539(.A0(new_n22971_), .A1(pi0625), .B0(new_n22975_), .Y(new_n22976_));
  NOR3X1   g20540(.A(new_n22976_), .B(new_n22846_), .C(pi0608), .Y(new_n22977_));
  NOR3X1   g20541(.A(new_n22977_), .B(new_n22974_), .C(new_n11889_), .Y(new_n22978_));
  AOI21X1  g20542(.A0(new_n22970_), .A1(new_n11889_), .B0(new_n22978_), .Y(new_n22979_));
  NAND2X1  g20543(.A(new_n22851_), .B(pi0609), .Y(new_n22980_));
  OAI21X1  g20544(.A0(new_n22979_), .A1(pi0609), .B0(new_n22980_), .Y(new_n22981_));
  OAI21X1  g20545(.A0(new_n22808_), .A1(new_n12591_), .B0(new_n12596_), .Y(new_n22982_));
  AOI21X1  g20546(.A0(new_n22981_), .A1(new_n12591_), .B0(new_n22982_), .Y(new_n22983_));
  NAND2X1  g20547(.A(new_n22851_), .B(new_n12590_), .Y(new_n22984_));
  OAI21X1  g20548(.A0(new_n22979_), .A1(new_n12590_), .B0(new_n22984_), .Y(new_n22985_));
  OAI21X1  g20549(.A0(new_n22807_), .A1(pi1155), .B0(pi0660), .Y(new_n22986_));
  AOI21X1  g20550(.A0(new_n22985_), .A1(pi1155), .B0(new_n22986_), .Y(new_n22987_));
  OR2X1    g20551(.A(new_n22987_), .B(new_n22983_), .Y(new_n22988_));
  MX2X1    g20552(.A(new_n22988_), .B(new_n22979_), .S0(new_n11888_), .Y(new_n22989_));
  MX2X1    g20553(.A(new_n22989_), .B(new_n22897_), .S0(pi0618), .Y(new_n22990_));
  NOR2X1   g20554(.A(new_n22815_), .B(pi0627), .Y(new_n22991_));
  OAI21X1  g20555(.A0(new_n22990_), .A1(pi1154), .B0(new_n22991_), .Y(new_n22992_));
  MX2X1    g20556(.A(new_n22989_), .B(new_n22897_), .S0(new_n12614_), .Y(new_n22993_));
  NOR2X1   g20557(.A(new_n22813_), .B(new_n12622_), .Y(new_n22994_));
  OAI21X1  g20558(.A0(new_n22993_), .A1(new_n12615_), .B0(new_n22994_), .Y(new_n22995_));
  AOI21X1  g20559(.A0(new_n22995_), .A1(new_n22992_), .B0(new_n11887_), .Y(new_n22996_));
  AND2X1   g20560(.A(new_n22989_), .B(new_n11887_), .Y(new_n22997_));
  NOR2X1   g20561(.A(new_n22997_), .B(new_n22996_), .Y(new_n22998_));
  MX2X1    g20562(.A(new_n22998_), .B(new_n22853_), .S0(pi0619), .Y(new_n22999_));
  AND2X1   g20563(.A(new_n22999_), .B(new_n12638_), .Y(new_n23000_));
  AND2X1   g20564(.A(new_n22823_), .B(new_n12645_), .Y(new_n23001_));
  INVX1    g20565(.A(new_n23001_), .Y(new_n23002_));
  AND2X1   g20566(.A(new_n22853_), .B(new_n12637_), .Y(new_n23003_));
  NOR3X1   g20567(.A(new_n22997_), .B(new_n22996_), .C(new_n12637_), .Y(new_n23004_));
  OAI21X1  g20568(.A0(new_n23004_), .A1(new_n23003_), .B0(pi1159), .Y(new_n23005_));
  AND2X1   g20569(.A(new_n22821_), .B(pi0648), .Y(new_n23006_));
  AOI21X1  g20570(.A0(new_n23006_), .A1(new_n23005_), .B0(new_n11886_), .Y(new_n23007_));
  OAI21X1  g20571(.A0(new_n23002_), .A1(new_n23000_), .B0(new_n23007_), .Y(new_n23008_));
  AOI21X1  g20572(.A0(new_n22998_), .A1(new_n11886_), .B0(new_n14264_), .Y(new_n23009_));
  NOR2X1   g20573(.A(new_n12767_), .B(new_n12690_), .Y(new_n23010_));
  INVX1    g20574(.A(new_n14196_), .Y(new_n23011_));
  AOI21X1  g20575(.A0(new_n22804_), .A1(new_n12672_), .B0(new_n23011_), .Y(new_n23012_));
  OAI21X1  g20576(.A0(new_n22855_), .A1(new_n12672_), .B0(new_n23012_), .Y(new_n23013_));
  INVX1    g20577(.A(new_n14204_), .Y(new_n23014_));
  AOI21X1  g20578(.A0(new_n22804_), .A1(pi0641), .B0(new_n23014_), .Y(new_n23015_));
  OAI21X1  g20579(.A0(new_n22855_), .A1(pi0641), .B0(new_n23015_), .Y(new_n23016_));
  AND2X1   g20580(.A(new_n23016_), .B(new_n23013_), .Y(new_n23017_));
  INVX1    g20581(.A(new_n23017_), .Y(new_n23018_));
  AOI21X1  g20582(.A0(new_n23010_), .A1(new_n22825_), .B0(new_n23018_), .Y(new_n23019_));
  OAI21X1  g20583(.A0(new_n23019_), .A1(new_n11885_), .B0(new_n16350_), .Y(new_n23020_));
  AOI21X1  g20584(.A0(new_n23009_), .A1(new_n23008_), .B0(new_n23020_), .Y(new_n23021_));
  OAI21X1  g20585(.A0(new_n22870_), .A1(new_n22869_), .B0(new_n12689_), .Y(new_n23022_));
  OAI22X1  g20586(.A0(new_n22875_), .A1(new_n12710_), .B0(new_n23022_), .B1(new_n12684_), .Y(new_n23023_));
  AOI21X1  g20587(.A0(new_n22827_), .A1(new_n14394_), .B0(new_n23023_), .Y(new_n23024_));
  NOR2X1   g20588(.A(new_n23024_), .B(new_n11884_), .Y(new_n23025_));
  OAI21X1  g20589(.A0(new_n23025_), .A1(new_n23021_), .B0(new_n22803_), .Y(new_n23026_));
  INVX1    g20590(.A(new_n22833_), .Y(new_n23027_));
  OAI21X1  g20591(.A0(new_n22926_), .A1(pi1156), .B0(new_n14392_), .Y(new_n23028_));
  AOI21X1  g20592(.A0(new_n23027_), .A1(pi1156), .B0(new_n23028_), .Y(new_n23029_));
  OAI21X1  g20593(.A0(new_n22926_), .A1(new_n12684_), .B0(new_n14393_), .Y(new_n23030_));
  AOI21X1  g20594(.A0(new_n23027_), .A1(new_n12684_), .B0(new_n23030_), .Y(new_n23031_));
  OAI21X1  g20595(.A0(new_n23031_), .A1(new_n23029_), .B0(pi0792), .Y(new_n23032_));
  OR2X1    g20596(.A(new_n22832_), .B(new_n14183_), .Y(new_n23033_));
  AND2X1   g20597(.A(pi0648), .B(new_n12637_), .Y(new_n23034_));
  OAI21X1  g20598(.A0(new_n22954_), .A1(new_n12638_), .B0(new_n23034_), .Y(new_n23035_));
  AOI21X1  g20599(.A0(new_n23033_), .A1(new_n12638_), .B0(new_n23035_), .Y(new_n23036_));
  AND2X1   g20600(.A(new_n12645_), .B(pi0619), .Y(new_n23037_));
  OAI21X1  g20601(.A0(new_n22954_), .A1(pi1159), .B0(new_n23037_), .Y(new_n23038_));
  AOI21X1  g20602(.A0(new_n23033_), .A1(pi1159), .B0(new_n23038_), .Y(new_n23039_));
  OAI21X1  g20603(.A0(new_n23039_), .A1(new_n23036_), .B0(pi0789), .Y(new_n23040_));
  AOI21X1  g20604(.A0(new_n22831_), .A1(new_n14182_), .B0(pi0627), .Y(new_n23041_));
  OAI21X1  g20605(.A0(new_n22945_), .A1(pi1154), .B0(new_n23041_), .Y(new_n23042_));
  OAI21X1  g20606(.A0(new_n16796_), .A1(new_n3810_), .B0(new_n11889_), .Y(new_n23043_));
  NOR3X1   g20607(.A(new_n16796_), .B(new_n3810_), .C(pi0625), .Y(new_n23044_));
  INVX1    g20608(.A(new_n23044_), .Y(new_n23045_));
  AND2X1   g20609(.A(new_n16746_), .B(new_n3129_), .Y(new_n23046_));
  AOI21X1  g20610(.A0(new_n23046_), .A1(pi0625), .B0(pi1153), .Y(new_n23047_));
  AOI21X1  g20611(.A0(new_n23047_), .A1(new_n23045_), .B0(new_n22929_), .Y(new_n23048_));
  NOR3X1   g20612(.A(new_n16796_), .B(new_n3810_), .C(new_n12493_), .Y(new_n23049_));
  AND2X1   g20613(.A(new_n23046_), .B(new_n12493_), .Y(new_n23050_));
  NOR3X1   g20614(.A(new_n23050_), .B(new_n23049_), .C(new_n12494_), .Y(new_n23051_));
  OAI21X1  g20615(.A0(new_n23051_), .A1(new_n22933_), .B0(pi0778), .Y(new_n23052_));
  OAI21X1  g20616(.A0(new_n23052_), .A1(new_n23048_), .B0(new_n23043_), .Y(new_n23053_));
  INVX1    g20617(.A(new_n23053_), .Y(new_n23054_));
  INVX1    g20618(.A(new_n22936_), .Y(new_n23055_));
  AOI21X1  g20619(.A0(new_n23055_), .A1(pi0609), .B0(pi1155), .Y(new_n23056_));
  OAI21X1  g20620(.A0(new_n23054_), .A1(pi0609), .B0(new_n23056_), .Y(new_n23057_));
  NAND4X1  g20621(.A(new_n16746_), .B(new_n14177_), .C(new_n12623_), .D(new_n3129_), .Y(new_n23058_));
  AND2X1   g20622(.A(new_n23058_), .B(new_n12596_), .Y(new_n23059_));
  AOI21X1  g20623(.A0(new_n23055_), .A1(new_n12590_), .B0(new_n12591_), .Y(new_n23060_));
  OAI21X1  g20624(.A0(new_n23054_), .A1(new_n12590_), .B0(new_n23060_), .Y(new_n23061_));
  NAND4X1  g20625(.A(new_n16746_), .B(new_n14176_), .C(new_n12623_), .D(new_n3129_), .Y(new_n23062_));
  AND2X1   g20626(.A(new_n23062_), .B(pi0660), .Y(new_n23063_));
  AOI22X1  g20627(.A0(new_n23063_), .A1(new_n23061_), .B0(new_n23059_), .B1(new_n23057_), .Y(new_n23064_));
  MX2X1    g20628(.A(new_n23064_), .B(new_n23054_), .S0(new_n11888_), .Y(new_n23065_));
  NOR2X1   g20629(.A(new_n23065_), .B(new_n12614_), .Y(new_n23066_));
  OAI21X1  g20630(.A0(new_n22947_), .A1(pi0618), .B0(pi1154), .Y(new_n23067_));
  AOI21X1  g20631(.A0(new_n22831_), .A1(new_n14181_), .B0(new_n12622_), .Y(new_n23068_));
  OAI21X1  g20632(.A0(new_n23067_), .A1(new_n23066_), .B0(new_n23068_), .Y(new_n23069_));
  AOI21X1  g20633(.A0(new_n23069_), .A1(new_n23042_), .B0(new_n11887_), .Y(new_n23070_));
  AOI21X1  g20634(.A0(new_n12622_), .A1(new_n12614_), .B0(new_n11887_), .Y(new_n23071_));
  OR4X1    g20635(.A(new_n23039_), .B(new_n23036_), .C(new_n16247_), .D(new_n11886_), .Y(new_n23072_));
  OAI21X1  g20636(.A0(new_n23071_), .A1(new_n23065_), .B0(new_n23072_), .Y(new_n23073_));
  OAI21X1  g20637(.A0(new_n23073_), .A1(new_n23070_), .B0(new_n23040_), .Y(new_n23074_));
  OAI21X1  g20638(.A0(new_n23074_), .A1(pi0626), .B0(new_n22959_), .Y(new_n23075_));
  AND2X1   g20639(.A(pi0641), .B(new_n12664_), .Y(new_n23076_));
  NOR3X1   g20640(.A(new_n22832_), .B(new_n14183_), .C(new_n14180_), .Y(new_n23077_));
  AOI21X1  g20641(.A0(new_n23077_), .A1(new_n23076_), .B0(pi1158), .Y(new_n23078_));
  OAI21X1  g20642(.A0(new_n23074_), .A1(new_n12664_), .B0(new_n22962_), .Y(new_n23079_));
  AND2X1   g20643(.A(new_n12672_), .B(pi0626), .Y(new_n23080_));
  AOI21X1  g20644(.A0(new_n23077_), .A1(new_n23080_), .B0(new_n12676_), .Y(new_n23081_));
  AOI22X1  g20645(.A0(new_n23081_), .A1(new_n23079_), .B0(new_n23078_), .B1(new_n23075_), .Y(new_n23082_));
  OR2X1    g20646(.A(new_n23074_), .B(pi0788), .Y(new_n23083_));
  AND2X1   g20647(.A(new_n23083_), .B(new_n16350_), .Y(new_n23084_));
  OAI21X1  g20648(.A0(new_n23082_), .A1(new_n11885_), .B0(new_n23084_), .Y(new_n23085_));
  AND2X1   g20649(.A(new_n23085_), .B(new_n23032_), .Y(new_n23086_));
  INVX1    g20650(.A(new_n23086_), .Y(new_n23087_));
  AOI21X1  g20651(.A0(new_n23087_), .A1(pi0207), .B0(new_n22925_), .Y(new_n23088_));
  AOI21X1  g20652(.A0(new_n23088_), .A1(new_n23026_), .B0(new_n22840_), .Y(new_n23089_));
  OAI21X1  g20653(.A0(new_n22969_), .A1(new_n22924_), .B0(new_n23089_), .Y(new_n23090_));
  AOI21X1  g20654(.A0(new_n22838_), .A1(new_n22840_), .B0(new_n14269_), .Y(new_n23091_));
  AOI21X1  g20655(.A0(new_n23091_), .A1(new_n23090_), .B0(new_n22868_), .Y(new_n23092_));
  NAND2X1  g20656(.A(new_n22866_), .B(new_n22864_), .Y(new_n23093_));
  MX2X1    g20657(.A(new_n23093_), .B(new_n22862_), .S0(new_n11883_), .Y(new_n23094_));
  OAI21X1  g20658(.A0(new_n23094_), .A1(pi0644), .B0(pi0715), .Y(new_n23095_));
  AOI21X1  g20659(.A0(new_n23092_), .A1(pi0644), .B0(new_n23095_), .Y(new_n23096_));
  MX2X1    g20660(.A(new_n22838_), .B(new_n22836_), .S0(new_n12735_), .Y(new_n23097_));
  OAI21X1  g20661(.A0(new_n22837_), .A1(pi0644), .B0(new_n12739_), .Y(new_n23098_));
  AOI21X1  g20662(.A0(new_n23097_), .A1(pi0644), .B0(new_n23098_), .Y(new_n23099_));
  OR2X1    g20663(.A(new_n23099_), .B(new_n11882_), .Y(new_n23100_));
  OAI21X1  g20664(.A0(new_n23094_), .A1(new_n12743_), .B0(new_n12739_), .Y(new_n23101_));
  AOI21X1  g20665(.A0(new_n23092_), .A1(new_n12743_), .B0(new_n23101_), .Y(new_n23102_));
  OAI21X1  g20666(.A0(new_n22837_), .A1(new_n12743_), .B0(pi0715), .Y(new_n23103_));
  AOI21X1  g20667(.A0(new_n23097_), .A1(new_n12743_), .B0(new_n23103_), .Y(new_n23104_));
  OR2X1    g20668(.A(new_n23104_), .B(pi1160), .Y(new_n23105_));
  OAI22X1  g20669(.A0(new_n23105_), .A1(new_n23102_), .B0(new_n23100_), .B1(new_n23096_), .Y(new_n23106_));
  MX2X1    g20670(.A(new_n23106_), .B(new_n23092_), .S0(new_n12897_), .Y(new_n23107_));
  MX2X1    g20671(.A(new_n23107_), .B(new_n22803_), .S0(po1038), .Y(po0364));
  INVX1    g20672(.A(pi0208), .Y(new_n23109_));
  NOR2X1   g20673(.A(new_n22828_), .B(pi0208), .Y(new_n23110_));
  OAI21X1  g20674(.A0(new_n22834_), .A1(new_n23109_), .B0(pi0607), .Y(new_n23111_));
  AOI21X1  g20675(.A0(new_n13699_), .A1(new_n3129_), .B0(pi0208), .Y(new_n23112_));
  INVX1    g20676(.A(new_n23112_), .Y(new_n23113_));
  OAI22X1  g20677(.A0(new_n23113_), .A1(pi0607), .B0(new_n23111_), .B1(new_n23110_), .Y(new_n23114_));
  OR2X1    g20678(.A(new_n23114_), .B(new_n14384_), .Y(new_n23115_));
  INVX1    g20679(.A(pi0638), .Y(new_n23116_));
  MX2X1    g20680(.A(new_n22859_), .B(new_n22841_), .S0(pi0208), .Y(new_n23117_));
  MX2X1    g20681(.A(new_n23117_), .B(new_n23112_), .S0(new_n23116_), .Y(new_n23118_));
  INVX1    g20682(.A(new_n23118_), .Y(new_n23119_));
  AOI21X1  g20683(.A0(new_n23112_), .A1(pi0647), .B0(pi1157), .Y(new_n23120_));
  OAI21X1  g20684(.A0(new_n23119_), .A1(pi0647), .B0(new_n23120_), .Y(new_n23121_));
  AOI21X1  g20685(.A0(new_n23112_), .A1(new_n12705_), .B0(new_n12706_), .Y(new_n23122_));
  OAI21X1  g20686(.A0(new_n23119_), .A1(new_n12705_), .B0(new_n23122_), .Y(new_n23123_));
  MX2X1    g20687(.A(new_n23123_), .B(new_n23121_), .S0(pi0630), .Y(new_n23124_));
  AOI21X1  g20688(.A0(new_n23124_), .A1(new_n23115_), .B0(new_n11883_), .Y(new_n23125_));
  AOI21X1  g20689(.A0(new_n22923_), .A1(new_n22877_), .B0(pi0208), .Y(new_n23126_));
  INVX1    g20690(.A(pi0607), .Y(new_n23127_));
  OAI21X1  g20691(.A0(new_n22968_), .A1(new_n23109_), .B0(new_n23127_), .Y(new_n23128_));
  OAI21X1  g20692(.A0(new_n23025_), .A1(new_n23021_), .B0(new_n23109_), .Y(new_n23129_));
  AOI21X1  g20693(.A0(new_n23087_), .A1(pi0208), .B0(new_n23127_), .Y(new_n23130_));
  AOI21X1  g20694(.A0(new_n23130_), .A1(new_n23129_), .B0(new_n23116_), .Y(new_n23131_));
  OAI21X1  g20695(.A0(new_n23128_), .A1(new_n23126_), .B0(new_n23131_), .Y(new_n23132_));
  AOI21X1  g20696(.A0(new_n23114_), .A1(new_n23116_), .B0(new_n14269_), .Y(new_n23133_));
  AOI21X1  g20697(.A0(new_n23133_), .A1(new_n23132_), .B0(new_n23125_), .Y(new_n23134_));
  NAND2X1  g20698(.A(new_n23123_), .B(new_n23121_), .Y(new_n23135_));
  MX2X1    g20699(.A(new_n23135_), .B(new_n23119_), .S0(new_n11883_), .Y(new_n23136_));
  OAI21X1  g20700(.A0(new_n23136_), .A1(pi0644), .B0(pi0715), .Y(new_n23137_));
  AOI21X1  g20701(.A0(new_n23134_), .A1(pi0644), .B0(new_n23137_), .Y(new_n23138_));
  MX2X1    g20702(.A(new_n23114_), .B(new_n23112_), .S0(new_n12735_), .Y(new_n23139_));
  OAI21X1  g20703(.A0(new_n23113_), .A1(pi0644), .B0(new_n12739_), .Y(new_n23140_));
  AOI21X1  g20704(.A0(new_n23139_), .A1(pi0644), .B0(new_n23140_), .Y(new_n23141_));
  OR2X1    g20705(.A(new_n23141_), .B(new_n11882_), .Y(new_n23142_));
  OAI21X1  g20706(.A0(new_n23136_), .A1(new_n12743_), .B0(new_n12739_), .Y(new_n23143_));
  AOI21X1  g20707(.A0(new_n23134_), .A1(new_n12743_), .B0(new_n23143_), .Y(new_n23144_));
  OAI21X1  g20708(.A0(new_n23113_), .A1(new_n12743_), .B0(pi0715), .Y(new_n23145_));
  AOI21X1  g20709(.A0(new_n23139_), .A1(new_n12743_), .B0(new_n23145_), .Y(new_n23146_));
  OR2X1    g20710(.A(new_n23146_), .B(pi1160), .Y(new_n23147_));
  OAI22X1  g20711(.A0(new_n23147_), .A1(new_n23144_), .B0(new_n23142_), .B1(new_n23138_), .Y(new_n23148_));
  MX2X1    g20712(.A(new_n23148_), .B(new_n23134_), .S0(new_n12897_), .Y(new_n23149_));
  MX2X1    g20713(.A(new_n23149_), .B(new_n23109_), .S0(po1038), .Y(po0365));
  INVX1    g20714(.A(pi0639), .Y(new_n23151_));
  AOI21X1  g20715(.A0(new_n22923_), .A1(new_n22877_), .B0(new_n14269_), .Y(new_n23152_));
  MX2X1    g20716(.A(new_n22858_), .B(new_n22819_), .S0(new_n12705_), .Y(new_n23153_));
  OAI22X1  g20717(.A0(new_n23153_), .A1(pi0630), .B0(new_n22819_), .B1(pi0647), .Y(new_n23154_));
  NAND2X1  g20718(.A(new_n23154_), .B(pi1157), .Y(new_n23155_));
  AOI21X1  g20719(.A0(new_n13699_), .A1(new_n3129_), .B0(new_n12705_), .Y(new_n23156_));
  MX2X1    g20720(.A(new_n22858_), .B(new_n22819_), .S0(pi0647), .Y(new_n23157_));
  INVX1    g20721(.A(new_n23157_), .Y(new_n23158_));
  AOI22X1  g20722(.A0(new_n23158_), .A1(new_n14388_), .B0(new_n23156_), .B1(new_n12706_), .Y(new_n23159_));
  AOI21X1  g20723(.A0(new_n23159_), .A1(new_n23155_), .B0(new_n11883_), .Y(new_n23160_));
  OAI21X1  g20724(.A0(new_n23160_), .A1(new_n23152_), .B0(new_n12743_), .Y(new_n23161_));
  MX2X1    g20725(.A(new_n22858_), .B(new_n22819_), .S0(new_n13651_), .Y(new_n23162_));
  INVX1    g20726(.A(new_n23162_), .Y(new_n23163_));
  AOI21X1  g20727(.A0(new_n23163_), .A1(pi0644), .B0(pi0715), .Y(new_n23164_));
  NAND2X1  g20728(.A(new_n23164_), .B(new_n23161_), .Y(new_n23165_));
  AOI21X1  g20729(.A0(new_n22819_), .A1(pi0715), .B0(pi1160), .Y(new_n23166_));
  OAI21X1  g20730(.A0(new_n23160_), .A1(new_n23152_), .B0(pi0644), .Y(new_n23167_));
  AOI21X1  g20731(.A0(new_n23163_), .A1(new_n12743_), .B0(new_n12739_), .Y(new_n23168_));
  NAND2X1  g20732(.A(new_n23168_), .B(new_n23167_), .Y(new_n23169_));
  AOI21X1  g20733(.A0(new_n22819_), .A1(new_n12739_), .B0(new_n11882_), .Y(new_n23170_));
  AOI22X1  g20734(.A0(new_n23170_), .A1(new_n23169_), .B0(new_n23166_), .B1(new_n23165_), .Y(new_n23171_));
  OAI21X1  g20735(.A0(new_n23160_), .A1(new_n23152_), .B0(new_n12897_), .Y(new_n23172_));
  AND2X1   g20736(.A(new_n23172_), .B(new_n6520_), .Y(new_n23173_));
  OAI21X1  g20737(.A0(new_n23171_), .A1(new_n12897_), .B0(new_n23173_), .Y(new_n23174_));
  OR2X1    g20738(.A(new_n23174_), .B(new_n23151_), .Y(new_n23175_));
  AND2X1   g20739(.A(new_n13699_), .B(new_n7686_), .Y(new_n23176_));
  AOI21X1  g20740(.A0(new_n23176_), .A1(new_n23151_), .B0(pi0622), .Y(new_n23177_));
  OR2X1    g20741(.A(new_n23025_), .B(new_n23021_), .Y(new_n23178_));
  INVX1    g20742(.A(new_n22828_), .Y(new_n23179_));
  NOR3X1   g20743(.A(new_n23153_), .B(new_n12706_), .C(pi0630), .Y(new_n23180_));
  AOI21X1  g20744(.A0(new_n23158_), .A1(new_n14388_), .B0(new_n23180_), .Y(new_n23181_));
  OAI21X1  g20745(.A0(new_n23179_), .A1(new_n14384_), .B0(new_n23181_), .Y(new_n23182_));
  AOI22X1  g20746(.A0(new_n23182_), .A1(pi0787), .B0(new_n23178_), .B1(new_n14562_), .Y(new_n23183_));
  OAI21X1  g20747(.A0(new_n23183_), .A1(pi0644), .B0(new_n23164_), .Y(new_n23184_));
  MX2X1    g20748(.A(new_n23179_), .B(new_n22819_), .S0(new_n12735_), .Y(new_n23185_));
  MX2X1    g20749(.A(new_n23185_), .B(new_n22819_), .S0(pi0644), .Y(new_n23186_));
  AOI21X1  g20750(.A0(new_n23186_), .A1(pi0715), .B0(pi1160), .Y(new_n23187_));
  OAI21X1  g20751(.A0(new_n23183_), .A1(new_n12743_), .B0(new_n23168_), .Y(new_n23188_));
  MX2X1    g20752(.A(new_n23185_), .B(new_n22819_), .S0(new_n12743_), .Y(new_n23189_));
  AOI21X1  g20753(.A0(new_n23189_), .A1(new_n12739_), .B0(new_n11882_), .Y(new_n23190_));
  AOI22X1  g20754(.A0(new_n23190_), .A1(new_n23188_), .B0(new_n23187_), .B1(new_n23184_), .Y(new_n23191_));
  OR2X1    g20755(.A(new_n23191_), .B(new_n12897_), .Y(new_n23192_));
  OAI21X1  g20756(.A0(new_n23183_), .A1(pi0790), .B0(new_n6520_), .Y(new_n23193_));
  INVX1    g20757(.A(new_n23193_), .Y(new_n23194_));
  NAND3X1  g20758(.A(new_n23194_), .B(new_n23192_), .C(pi0639), .Y(new_n23195_));
  INVX1    g20759(.A(pi0622), .Y(new_n23196_));
  AND2X1   g20760(.A(new_n23189_), .B(pi1160), .Y(new_n23197_));
  INVX1    g20761(.A(new_n23197_), .Y(new_n23198_));
  AOI21X1  g20762(.A0(new_n23186_), .A1(new_n11882_), .B0(new_n12897_), .Y(new_n23199_));
  OAI21X1  g20763(.A0(new_n23185_), .A1(pi0790), .B0(new_n6520_), .Y(new_n23200_));
  AOI21X1  g20764(.A0(new_n23199_), .A1(new_n23198_), .B0(new_n23200_), .Y(new_n23201_));
  AOI21X1  g20765(.A0(new_n23201_), .A1(new_n23151_), .B0(new_n23196_), .Y(new_n23202_));
  AOI22X1  g20766(.A0(new_n23202_), .A1(new_n23195_), .B0(new_n23177_), .B1(new_n23175_), .Y(new_n23203_));
  AND2X1   g20767(.A(new_n22841_), .B(new_n14286_), .Y(new_n23204_));
  INVX1    g20768(.A(new_n23204_), .Y(new_n23205_));
  AOI21X1  g20769(.A0(new_n23205_), .A1(pi0644), .B0(pi0715), .Y(new_n23206_));
  INVX1    g20770(.A(new_n23206_), .Y(new_n23207_));
  AOI21X1  g20771(.A0(new_n22834_), .A1(pi0647), .B0(pi1157), .Y(new_n23208_));
  OAI21X1  g20772(.A0(new_n23086_), .A1(pi0647), .B0(new_n23208_), .Y(new_n23209_));
  AOI21X1  g20773(.A0(new_n22841_), .A1(pi0647), .B0(new_n12706_), .Y(new_n23210_));
  OR2X1    g20774(.A(new_n23210_), .B(pi0630), .Y(new_n23211_));
  INVX1    g20775(.A(new_n23211_), .Y(new_n23212_));
  AOI21X1  g20776(.A0(new_n22834_), .A1(new_n12705_), .B0(new_n12706_), .Y(new_n23213_));
  OAI21X1  g20777(.A0(new_n23086_), .A1(new_n12705_), .B0(new_n23213_), .Y(new_n23214_));
  AOI21X1  g20778(.A0(new_n22841_), .A1(new_n12705_), .B0(pi1157), .Y(new_n23215_));
  OR2X1    g20779(.A(new_n23215_), .B(new_n12723_), .Y(new_n23216_));
  INVX1    g20780(.A(new_n23216_), .Y(new_n23217_));
  AOI22X1  g20781(.A0(new_n23217_), .A1(new_n23214_), .B0(new_n23212_), .B1(new_n23209_), .Y(new_n23218_));
  MX2X1    g20782(.A(new_n23218_), .B(new_n23086_), .S0(new_n11883_), .Y(new_n23219_));
  AND2X1   g20783(.A(new_n23219_), .B(new_n12743_), .Y(new_n23220_));
  OR4X1    g20784(.A(new_n23027_), .B(new_n16294_), .C(new_n12739_), .D(pi0644), .Y(new_n23221_));
  AND2X1   g20785(.A(new_n23221_), .B(new_n11882_), .Y(new_n23222_));
  OAI21X1  g20786(.A0(new_n23220_), .A1(new_n23207_), .B0(new_n23222_), .Y(new_n23223_));
  AOI21X1  g20787(.A0(new_n23205_), .A1(new_n12743_), .B0(new_n12739_), .Y(new_n23224_));
  INVX1    g20788(.A(new_n23224_), .Y(new_n23225_));
  AND2X1   g20789(.A(new_n23219_), .B(pi0644), .Y(new_n23226_));
  OR4X1    g20790(.A(new_n23027_), .B(new_n16294_), .C(pi0715), .D(new_n12743_), .Y(new_n23227_));
  AND2X1   g20791(.A(new_n23227_), .B(pi1160), .Y(new_n23228_));
  OAI21X1  g20792(.A0(new_n23226_), .A1(new_n23225_), .B0(new_n23228_), .Y(new_n23229_));
  AND2X1   g20793(.A(new_n23229_), .B(new_n23223_), .Y(new_n23230_));
  AOI21X1  g20794(.A0(new_n23219_), .A1(new_n12897_), .B0(po1038), .Y(new_n23231_));
  OAI21X1  g20795(.A0(new_n23230_), .A1(new_n12897_), .B0(new_n23231_), .Y(new_n23232_));
  NAND3X1  g20796(.A(new_n23232_), .B(pi0639), .C(pi0622), .Y(new_n23233_));
  NOR2X1   g20797(.A(new_n22968_), .B(new_n14269_), .Y(new_n23234_));
  AND2X1   g20798(.A(new_n13650_), .B(new_n12735_), .Y(new_n23235_));
  AOI21X1  g20799(.A0(new_n23235_), .A1(new_n22841_), .B0(new_n23234_), .Y(new_n23236_));
  NAND2X1  g20800(.A(new_n23224_), .B(pi1160), .Y(new_n23237_));
  AOI21X1  g20801(.A0(new_n23236_), .A1(pi0644), .B0(new_n23237_), .Y(new_n23238_));
  NAND2X1  g20802(.A(new_n23206_), .B(new_n11882_), .Y(new_n23239_));
  AOI21X1  g20803(.A0(new_n23236_), .A1(new_n12743_), .B0(new_n23239_), .Y(new_n23240_));
  OR2X1    g20804(.A(new_n23240_), .B(new_n12897_), .Y(new_n23241_));
  AOI21X1  g20805(.A0(new_n23236_), .A1(new_n12897_), .B0(po1038), .Y(new_n23242_));
  OAI21X1  g20806(.A0(new_n23241_), .A1(new_n23238_), .B0(new_n23242_), .Y(new_n23243_));
  INVX1    g20807(.A(pi0209), .Y(new_n23244_));
  XOR2X1   g20808(.A(pi1160), .B(pi0644), .Y(new_n23245_));
  AND2X1   g20809(.A(new_n23245_), .B(pi0790), .Y(new_n23246_));
  NOR4X1   g20810(.A(new_n23246_), .B(new_n23027_), .C(new_n16294_), .D(po1038), .Y(new_n23247_));
  AOI21X1  g20811(.A0(new_n23247_), .A1(pi0622), .B0(pi0639), .Y(new_n23248_));
  OR2X1    g20812(.A(new_n23248_), .B(new_n23244_), .Y(new_n23249_));
  AOI21X1  g20813(.A0(new_n23243_), .A1(new_n23196_), .B0(new_n23249_), .Y(new_n23250_));
  NAND2X1  g20814(.A(new_n23250_), .B(new_n23233_), .Y(new_n23251_));
  OAI21X1  g20815(.A0(new_n23203_), .A1(pi0209), .B0(new_n23251_), .Y(po0366));
  AOI22X1  g20816(.A0(new_n14591_), .A1(pi0634), .B0(pi0947), .B1(pi0633), .Y(new_n23253_));
  OAI21X1  g20817(.A0(new_n23253_), .A1(new_n12901_), .B0(pi0038), .Y(new_n23254_));
  AOI21X1  g20818(.A0(new_n12901_), .A1(pi0210), .B0(new_n23254_), .Y(new_n23255_));
  OAI21X1  g20819(.A0(new_n11952_), .A1(new_n2740_), .B0(pi0210), .Y(new_n23256_));
  OAI21X1  g20820(.A0(new_n5030_), .A1(new_n5028_), .B0(pi0210), .Y(new_n23257_));
  OAI22X1  g20821(.A0(new_n23257_), .A1(new_n12029_), .B0(new_n23256_), .B1(po1101), .Y(new_n23258_));
  MX2X1    g20822(.A(new_n22072_), .B(new_n2766_), .S0(new_n11953_), .Y(new_n23259_));
  OR2X1    g20823(.A(new_n23259_), .B(new_n6269_), .Y(new_n23260_));
  AND2X1   g20824(.A(new_n23260_), .B(pi0907), .Y(new_n23261_));
  MX2X1    g20825(.A(new_n2766_), .B(new_n22072_), .S0(new_n12028_), .Y(new_n23262_));
  OAI21X1  g20826(.A0(new_n23262_), .A1(new_n6270_), .B0(new_n23261_), .Y(new_n23263_));
  AND2X1   g20827(.A(new_n23263_), .B(new_n14590_), .Y(new_n23264_));
  OAI21X1  g20828(.A0(new_n23258_), .A1(pi0907), .B0(new_n23264_), .Y(new_n23265_));
  MX2X1    g20829(.A(new_n21917_), .B(new_n2766_), .S0(new_n11953_), .Y(new_n23266_));
  AOI21X1  g20830(.A0(new_n23266_), .A1(new_n5031_), .B0(new_n14590_), .Y(new_n23267_));
  AND2X1   g20831(.A(new_n23266_), .B(po1101), .Y(new_n23268_));
  OR2X1    g20832(.A(new_n23268_), .B(new_n6269_), .Y(new_n23269_));
  MX2X1    g20833(.A(new_n2766_), .B(new_n21917_), .S0(new_n12028_), .Y(new_n23270_));
  OAI21X1  g20834(.A0(new_n23270_), .A1(new_n5033_), .B0(new_n23269_), .Y(new_n23271_));
  AOI21X1  g20835(.A0(new_n23271_), .A1(new_n23267_), .B0(new_n5051_), .Y(new_n23272_));
  AOI21X1  g20836(.A0(new_n23259_), .A1(new_n5052_), .B0(new_n5297_), .Y(new_n23273_));
  INVX1    g20837(.A(new_n23273_), .Y(new_n23274_));
  AOI21X1  g20838(.A0(new_n23262_), .A1(new_n5053_), .B0(new_n23274_), .Y(new_n23275_));
  NOR3X1   g20839(.A(new_n12106_), .B(pi0907), .C(new_n2766_), .Y(new_n23276_));
  OAI21X1  g20840(.A0(new_n23276_), .A1(new_n23275_), .B0(new_n14590_), .Y(new_n23277_));
  AOI21X1  g20841(.A0(new_n23266_), .A1(new_n5052_), .B0(new_n14590_), .Y(new_n23278_));
  INVX1    g20842(.A(new_n23278_), .Y(new_n23279_));
  AOI21X1  g20843(.A0(new_n23270_), .A1(new_n5053_), .B0(new_n23279_), .Y(new_n23280_));
  NOR2X1   g20844(.A(new_n23280_), .B(new_n5050_), .Y(new_n23281_));
  AOI22X1  g20845(.A0(new_n23281_), .A1(new_n23277_), .B0(new_n23272_), .B1(new_n23265_), .Y(new_n23282_));
  MX2X1    g20846(.A(new_n23253_), .B(new_n2766_), .S0(new_n11953_), .Y(new_n23283_));
  AOI21X1  g20847(.A0(new_n23283_), .A1(new_n2970_), .B0(pi0223), .Y(new_n23284_));
  OAI21X1  g20848(.A0(new_n23282_), .A1(new_n2970_), .B0(new_n23284_), .Y(new_n23285_));
  MX2X1    g20849(.A(new_n22072_), .B(new_n2766_), .S0(new_n11965_), .Y(new_n23286_));
  AND2X1   g20850(.A(new_n23286_), .B(new_n5053_), .Y(new_n23287_));
  NOR3X1   g20851(.A(new_n11952_), .B(new_n5053_), .C(new_n2740_), .Y(new_n23288_));
  OR4X1    g20852(.A(new_n23288_), .B(new_n11964_), .C(new_n11958_), .D(new_n2766_), .Y(new_n23289_));
  OAI21X1  g20853(.A0(new_n23287_), .A1(new_n23274_), .B0(new_n23289_), .Y(new_n23290_));
  AND2X1   g20854(.A(new_n23290_), .B(new_n14590_), .Y(new_n23291_));
  MX2X1    g20855(.A(new_n21917_), .B(new_n2766_), .S0(new_n11965_), .Y(new_n23292_));
  AND2X1   g20856(.A(new_n23292_), .B(new_n5053_), .Y(new_n23293_));
  OAI21X1  g20857(.A0(new_n23293_), .A1(new_n23279_), .B0(new_n5051_), .Y(new_n23294_));
  OAI22X1  g20858(.A0(new_n23257_), .A1(new_n12135_), .B0(new_n23256_), .B1(po1101), .Y(new_n23295_));
  OR2X1    g20859(.A(new_n23295_), .B(pi0907), .Y(new_n23296_));
  OAI21X1  g20860(.A0(new_n23286_), .A1(new_n6270_), .B0(new_n23261_), .Y(new_n23297_));
  NAND3X1  g20861(.A(new_n23297_), .B(new_n23296_), .C(new_n14590_), .Y(new_n23298_));
  OAI22X1  g20862(.A0(new_n23292_), .A1(new_n5033_), .B0(new_n23268_), .B1(new_n6269_), .Y(new_n23299_));
  AOI21X1  g20863(.A0(new_n23299_), .A1(new_n23267_), .B0(new_n5051_), .Y(new_n23300_));
  AOI21X1  g20864(.A0(new_n23300_), .A1(new_n23298_), .B0(new_n2964_), .Y(new_n23301_));
  OAI21X1  g20865(.A0(new_n23294_), .A1(new_n23291_), .B0(new_n23301_), .Y(new_n23302_));
  NAND3X1  g20866(.A(new_n23302_), .B(new_n23285_), .C(new_n2953_), .Y(new_n23303_));
  INVX1    g20867(.A(new_n23275_), .Y(new_n23304_));
  AOI21X1  g20868(.A0(new_n21883_), .A1(pi0210), .B0(new_n12069_), .Y(new_n23305_));
  OAI21X1  g20869(.A0(new_n23258_), .A1(new_n5069_), .B0(new_n5297_), .Y(new_n23306_));
  OAI21X1  g20870(.A0(new_n23306_), .A1(new_n23305_), .B0(new_n23304_), .Y(new_n23307_));
  OR2X1    g20871(.A(new_n23280_), .B(new_n10136_), .Y(new_n23308_));
  AOI21X1  g20872(.A0(new_n23307_), .A1(new_n14590_), .B0(new_n23308_), .Y(new_n23309_));
  AND2X1   g20873(.A(new_n23283_), .B(new_n10136_), .Y(new_n23310_));
  OR2X1    g20874(.A(new_n23310_), .B(pi0215), .Y(new_n23311_));
  NOR2X1   g20875(.A(new_n23287_), .B(new_n23274_), .Y(new_n23312_));
  OR2X1    g20876(.A(new_n23295_), .B(new_n5069_), .Y(new_n23313_));
  AOI21X1  g20877(.A0(new_n23289_), .A1(new_n5069_), .B0(pi0907), .Y(new_n23314_));
  AOI21X1  g20878(.A0(new_n23314_), .A1(new_n23313_), .B0(new_n23312_), .Y(new_n23315_));
  OAI22X1  g20879(.A0(new_n23315_), .A1(pi0947), .B0(new_n23293_), .B1(new_n23279_), .Y(new_n23316_));
  AOI21X1  g20880(.A0(new_n23316_), .A1(pi0215), .B0(new_n2953_), .Y(new_n23317_));
  OAI21X1  g20881(.A0(new_n23311_), .A1(new_n23309_), .B0(new_n23317_), .Y(new_n23318_));
  NAND3X1  g20882(.A(new_n23318_), .B(new_n23303_), .C(pi0039), .Y(new_n23319_));
  INVX1    g20883(.A(new_n23253_), .Y(new_n23320_));
  AOI21X1  g20884(.A0(new_n23320_), .A1(new_n11946_), .B0(pi0299), .Y(new_n23321_));
  OAI21X1  g20885(.A0(new_n11946_), .A1(new_n2766_), .B0(new_n23321_), .Y(new_n23322_));
  AOI21X1  g20886(.A0(new_n23320_), .A1(new_n11929_), .B0(new_n2953_), .Y(new_n23323_));
  AOI21X1  g20887(.A0(new_n23323_), .A1(new_n11942_), .B0(pi0039), .Y(new_n23324_));
  AOI21X1  g20888(.A0(new_n23324_), .A1(new_n23322_), .B0(pi0038), .Y(new_n23325_));
  AOI21X1  g20889(.A0(new_n23325_), .A1(new_n23319_), .B0(new_n23255_), .Y(new_n23326_));
  MX2X1    g20890(.A(new_n23326_), .B(pi0210), .S0(new_n9580_), .Y(po0367));
  NOR2X1   g20891(.A(new_n15077_), .B(new_n3810_), .Y(new_n23328_));
  NAND2X1  g20892(.A(new_n15075_), .B(new_n3129_), .Y(new_n23329_));
  OAI21X1  g20893(.A0(new_n23329_), .A1(new_n22432_), .B0(pi0643), .Y(new_n23330_));
  AOI21X1  g20894(.A0(new_n23328_), .A1(new_n22432_), .B0(new_n23330_), .Y(new_n23331_));
  NOR2X1   g20895(.A(new_n14658_), .B(new_n3810_), .Y(new_n23332_));
  OAI21X1  g20896(.A0(new_n22804_), .A1(pi0606), .B0(new_n22461_), .Y(new_n23333_));
  AOI21X1  g20897(.A0(new_n23332_), .A1(pi0606), .B0(new_n23333_), .Y(new_n23334_));
  NOR3X1   g20898(.A(new_n23334_), .B(new_n23331_), .C(po1038), .Y(new_n23335_));
  NAND2X1  g20899(.A(new_n15069_), .B(new_n3129_), .Y(new_n23336_));
  AND2X1   g20900(.A(new_n15067_), .B(new_n3129_), .Y(new_n23337_));
  OAI21X1  g20901(.A0(new_n23337_), .A1(new_n22432_), .B0(pi0643), .Y(new_n23338_));
  AOI21X1  g20902(.A0(new_n23336_), .A1(new_n22432_), .B0(new_n23338_), .Y(new_n23339_));
  NOR4X1   g20903(.A(new_n14675_), .B(new_n3810_), .C(pi0643), .D(new_n22432_), .Y(new_n23340_));
  AND2X1   g20904(.A(new_n6520_), .B(new_n8548_), .Y(new_n23341_));
  OAI21X1  g20905(.A0(new_n23340_), .A1(new_n23339_), .B0(new_n23341_), .Y(new_n23342_));
  OAI21X1  g20906(.A0(new_n23335_), .A1(new_n8548_), .B0(new_n23342_), .Y(po0368));
  OAI21X1  g20907(.A0(new_n23329_), .A1(new_n23127_), .B0(pi0638), .Y(new_n23344_));
  AOI21X1  g20908(.A0(new_n23328_), .A1(new_n23127_), .B0(new_n23344_), .Y(new_n23345_));
  OAI21X1  g20909(.A0(new_n22804_), .A1(pi0607), .B0(new_n23116_), .Y(new_n23346_));
  AOI21X1  g20910(.A0(new_n23332_), .A1(pi0607), .B0(new_n23346_), .Y(new_n23347_));
  NOR3X1   g20911(.A(new_n23347_), .B(new_n23345_), .C(po1038), .Y(new_n23348_));
  OR2X1    g20912(.A(new_n23337_), .B(new_n23127_), .Y(new_n23349_));
  AOI21X1  g20913(.A0(new_n23336_), .A1(new_n23127_), .B0(new_n23116_), .Y(new_n23350_));
  NOR4X1   g20914(.A(new_n14675_), .B(new_n3810_), .C(pi0638), .D(new_n23127_), .Y(new_n23351_));
  AOI21X1  g20915(.A0(new_n23350_), .A1(new_n23349_), .B0(new_n23351_), .Y(new_n23352_));
  NAND3X1  g20916(.A(new_n5117_), .B(pi0212), .C(new_n2436_), .Y(new_n23353_));
  OAI22X1  g20917(.A0(new_n23353_), .A1(new_n23352_), .B0(new_n23348_), .B1(pi0212), .Y(po0369));
  AND2X1   g20918(.A(new_n6520_), .B(pi0213), .Y(new_n23355_));
  INVX1    g20919(.A(new_n23355_), .Y(new_n23356_));
  OR2X1    g20920(.A(new_n23337_), .B(new_n23196_), .Y(new_n23357_));
  AOI21X1  g20921(.A0(new_n23336_), .A1(new_n23196_), .B0(new_n23151_), .Y(new_n23358_));
  NOR4X1   g20922(.A(new_n14675_), .B(new_n3810_), .C(pi0639), .D(new_n23196_), .Y(new_n23359_));
  AOI21X1  g20923(.A0(new_n23358_), .A1(new_n23357_), .B0(new_n23359_), .Y(new_n23360_));
  OAI21X1  g20924(.A0(new_n23329_), .A1(new_n23151_), .B0(pi0622), .Y(new_n23361_));
  AOI21X1  g20925(.A0(new_n23332_), .A1(new_n23151_), .B0(new_n23361_), .Y(new_n23362_));
  OAI21X1  g20926(.A0(new_n22804_), .A1(pi0639), .B0(new_n23196_), .Y(new_n23363_));
  AOI21X1  g20927(.A0(new_n23328_), .A1(pi0639), .B0(new_n23363_), .Y(new_n23364_));
  NOR3X1   g20928(.A(new_n23364_), .B(new_n23362_), .C(po1038), .Y(new_n23365_));
  OAI22X1  g20929(.A0(new_n23365_), .A1(pi0213), .B0(new_n23360_), .B1(new_n23356_), .Y(po0370));
  OAI21X1  g20930(.A0(new_n23329_), .A1(new_n22925_), .B0(pi0710), .Y(new_n23367_));
  AOI21X1  g20931(.A0(new_n23328_), .A1(new_n22925_), .B0(new_n23367_), .Y(new_n23368_));
  OAI21X1  g20932(.A0(new_n22804_), .A1(pi0623), .B0(new_n22840_), .Y(new_n23369_));
  AOI21X1  g20933(.A0(new_n23332_), .A1(pi0623), .B0(new_n23369_), .Y(new_n23370_));
  NOR3X1   g20934(.A(new_n23370_), .B(new_n23368_), .C(po1038), .Y(new_n23371_));
  OR2X1    g20935(.A(new_n23337_), .B(new_n22925_), .Y(new_n23372_));
  AOI21X1  g20936(.A0(new_n23336_), .A1(new_n22925_), .B0(new_n22840_), .Y(new_n23373_));
  NOR4X1   g20937(.A(new_n14675_), .B(new_n3810_), .C(pi0710), .D(new_n22925_), .Y(new_n23374_));
  AOI21X1  g20938(.A0(new_n23373_), .A1(new_n23372_), .B0(new_n23374_), .Y(new_n23375_));
  NAND3X1  g20939(.A(new_n5117_), .B(pi0214), .C(new_n2436_), .Y(new_n23376_));
  OAI22X1  g20940(.A0(new_n23376_), .A1(new_n23375_), .B0(new_n23371_), .B1(pi0214), .Y(po0371));
  AND2X1   g20941(.A(new_n14862_), .B(new_n14590_), .Y(new_n23378_));
  INVX1    g20942(.A(new_n23378_), .Y(new_n23379_));
  AND2X1   g20943(.A(pi0907), .B(pi0681), .Y(new_n23380_));
  AND2X1   g20944(.A(new_n23380_), .B(new_n14590_), .Y(new_n23381_));
  NOR2X1   g20945(.A(pi0681), .B(pi0661), .Y(new_n23382_));
  AOI21X1  g20946(.A0(new_n23382_), .A1(new_n11984_), .B0(pi0642), .Y(new_n23383_));
  OAI21X1  g20947(.A0(new_n11974_), .A1(new_n5030_), .B0(new_n23383_), .Y(new_n23384_));
  AOI21X1  g20948(.A0(new_n23384_), .A1(pi0947), .B0(new_n23381_), .Y(new_n23385_));
  AOI21X1  g20949(.A0(new_n23385_), .A1(new_n23379_), .B0(new_n2953_), .Y(new_n23386_));
  NOR3X1   g20950(.A(new_n23380_), .B(new_n14929_), .C(pi0947), .Y(new_n23387_));
  AOI21X1  g20951(.A0(new_n12106_), .A1(new_n11968_), .B0(new_n5050_), .Y(new_n23388_));
  OAI21X1  g20952(.A0(new_n12047_), .A1(pi0642), .B0(new_n5030_), .Y(new_n23389_));
  NOR3X1   g20953(.A(new_n11952_), .B(new_n12323_), .C(new_n2740_), .Y(new_n23390_));
  AOI21X1  g20954(.A0(new_n23390_), .A1(new_n11968_), .B0(new_n5030_), .Y(new_n23391_));
  OAI21X1  g20955(.A0(new_n12127_), .A1(new_n12246_), .B0(new_n23391_), .Y(new_n23392_));
  AOI21X1  g20956(.A0(new_n23392_), .A1(new_n23389_), .B0(new_n5051_), .Y(new_n23393_));
  NOR3X1   g20957(.A(new_n23393_), .B(new_n23388_), .C(new_n14590_), .Y(new_n23394_));
  OR2X1    g20958(.A(new_n23394_), .B(new_n2970_), .Y(new_n23395_));
  AND2X1   g20959(.A(new_n11953_), .B(new_n2970_), .Y(new_n23396_));
  INVX1    g20960(.A(new_n23380_), .Y(new_n23397_));
  MX2X1    g20961(.A(new_n23397_), .B(new_n11968_), .S0(pi0947), .Y(new_n23398_));
  NOR2X1   g20962(.A(new_n23398_), .B(new_n2971_), .Y(new_n23399_));
  NOR3X1   g20963(.A(new_n23399_), .B(new_n23396_), .C(pi0223), .Y(new_n23400_));
  OAI21X1  g20964(.A0(new_n23395_), .A1(new_n23387_), .B0(new_n23400_), .Y(new_n23401_));
  OAI21X1  g20965(.A0(new_n12135_), .A1(new_n5282_), .B0(new_n11968_), .Y(new_n23402_));
  AOI21X1  g20966(.A0(new_n12230_), .A1(new_n5282_), .B0(new_n23402_), .Y(new_n23403_));
  AOI21X1  g20967(.A0(new_n23384_), .A1(new_n5051_), .B0(new_n14590_), .Y(new_n23404_));
  OAI21X1  g20968(.A0(new_n23403_), .A1(new_n5051_), .B0(new_n23404_), .Y(new_n23405_));
  OAI21X1  g20969(.A0(new_n12010_), .A1(pi0947), .B0(new_n23405_), .Y(new_n23406_));
  AOI21X1  g20970(.A0(new_n23380_), .A1(new_n14590_), .B0(new_n2964_), .Y(new_n23407_));
  AOI21X1  g20971(.A0(new_n23407_), .A1(new_n23406_), .B0(pi0299), .Y(new_n23408_));
  AOI21X1  g20972(.A0(new_n23408_), .A1(new_n23401_), .B0(new_n23386_), .Y(new_n23409_));
  INVX1    g20973(.A(new_n23381_), .Y(new_n23410_));
  NOR2X1   g20974(.A(new_n12029_), .B(new_n5029_), .Y(new_n23411_));
  NOR2X1   g20975(.A(new_n11993_), .B(new_n11968_), .Y(new_n23412_));
  INVX1    g20976(.A(new_n23412_), .Y(new_n23413_));
  NAND3X1  g20977(.A(new_n12004_), .B(new_n11993_), .C(pi0642), .Y(new_n23414_));
  OAI22X1  g20978(.A0(new_n23414_), .A1(new_n23411_), .B0(new_n23413_), .B1(new_n11953_), .Y(new_n23415_));
  AOI21X1  g20979(.A0(new_n23415_), .A1(pi0947), .B0(new_n5051_), .Y(new_n23416_));
  OAI21X1  g20980(.A0(new_n23410_), .A1(new_n12033_), .B0(new_n23416_), .Y(new_n23417_));
  OAI21X1  g20981(.A0(new_n23397_), .A1(new_n12260_), .B0(new_n14590_), .Y(new_n23418_));
  AND2X1   g20982(.A(new_n11993_), .B(pi0642), .Y(new_n23419_));
  MX2X1    g20983(.A(new_n12056_), .B(new_n12028_), .S0(new_n5030_), .Y(new_n23420_));
  AND2X1   g20984(.A(new_n23420_), .B(new_n23419_), .Y(new_n23421_));
  OAI21X1  g20985(.A0(new_n23413_), .A1(new_n12107_), .B0(pi0947), .Y(new_n23422_));
  OAI21X1  g20986(.A0(new_n23422_), .A1(new_n23421_), .B0(new_n23418_), .Y(new_n23423_));
  AOI21X1  g20987(.A0(new_n23423_), .A1(new_n5051_), .B0(new_n2970_), .Y(new_n23424_));
  INVX1    g20988(.A(new_n23399_), .Y(new_n23425_));
  OAI21X1  g20989(.A0(new_n23425_), .A1(new_n11953_), .B0(new_n2964_), .Y(new_n23426_));
  AOI21X1  g20990(.A0(new_n23424_), .A1(new_n23417_), .B0(new_n23426_), .Y(new_n23427_));
  AOI21X1  g20991(.A0(new_n11981_), .A1(new_n11979_), .B0(new_n5051_), .Y(new_n23428_));
  OAI21X1  g20992(.A0(new_n23428_), .A1(new_n23397_), .B0(new_n14590_), .Y(new_n23429_));
  AOI21X1  g20993(.A0(new_n12145_), .A1(pi0947), .B0(new_n11974_), .Y(new_n23430_));
  NAND3X1  g20994(.A(new_n23419_), .B(new_n12004_), .C(new_n11999_), .Y(new_n23431_));
  AOI21X1  g20995(.A0(new_n23412_), .A1(new_n12012_), .B0(new_n14590_), .Y(new_n23432_));
  AOI22X1  g20996(.A0(new_n23432_), .A1(new_n23431_), .B0(new_n23430_), .B1(new_n5051_), .Y(new_n23433_));
  AOI21X1  g20997(.A0(new_n23433_), .A1(new_n23429_), .B0(new_n2964_), .Y(new_n23434_));
  OAI21X1  g20998(.A0(new_n23434_), .A1(new_n23427_), .B0(new_n2953_), .Y(new_n23435_));
  INVX1    g20999(.A(new_n23398_), .Y(new_n23436_));
  AOI21X1  g21000(.A0(new_n23436_), .A1(new_n12077_), .B0(new_n2953_), .Y(new_n23437_));
  OAI21X1  g21001(.A0(new_n23423_), .A1(new_n10136_), .B0(new_n23437_), .Y(new_n23438_));
  NAND3X1  g21002(.A(new_n23438_), .B(new_n23435_), .C(new_n2954_), .Y(new_n23439_));
  OAI21X1  g21003(.A0(new_n23409_), .A1(new_n2954_), .B0(new_n23439_), .Y(new_n23440_));
  OAI21X1  g21004(.A0(new_n23398_), .A1(new_n12091_), .B0(pi0299), .Y(new_n23441_));
  AOI21X1  g21005(.A0(new_n12091_), .A1(pi0215), .B0(new_n23441_), .Y(new_n23442_));
  NOR2X1   g21006(.A(new_n23398_), .B(new_n12445_), .Y(new_n23443_));
  OAI21X1  g21007(.A0(new_n11946_), .A1(new_n2954_), .B0(new_n2953_), .Y(new_n23444_));
  OAI21X1  g21008(.A0(new_n23444_), .A1(new_n23443_), .B0(new_n2959_), .Y(new_n23445_));
  OAI21X1  g21009(.A0(new_n23445_), .A1(new_n23442_), .B0(new_n2996_), .Y(new_n23446_));
  AOI21X1  g21010(.A0(new_n23440_), .A1(pi0039), .B0(new_n23446_), .Y(new_n23447_));
  AND2X1   g21011(.A(new_n23436_), .B(new_n12202_), .Y(new_n23448_));
  OAI21X1  g21012(.A0(new_n12202_), .A1(new_n2954_), .B0(pi0038), .Y(new_n23449_));
  OAI21X1  g21013(.A0(new_n23449_), .A1(new_n23448_), .B0(new_n7686_), .Y(new_n23450_));
  OAI22X1  g21014(.A0(new_n23450_), .A1(new_n23447_), .B0(new_n7686_), .B1(new_n2954_), .Y(po0372));
  NAND2X1  g21015(.A(pi0907), .B(pi0662), .Y(new_n23452_));
  MX2X1    g21016(.A(new_n23452_), .B(new_n12051_), .S0(pi0947), .Y(new_n23453_));
  AOI21X1  g21017(.A0(new_n12901_), .A1(pi0216), .B0(new_n2996_), .Y(new_n23454_));
  OAI21X1  g21018(.A0(new_n23453_), .A1(new_n12901_), .B0(new_n23454_), .Y(new_n23455_));
  NOR2X1   g21019(.A(new_n23452_), .B(pi0947), .Y(new_n23456_));
  AOI21X1  g21020(.A0(new_n12106_), .A1(new_n12051_), .B0(new_n14590_), .Y(new_n23457_));
  OR2X1    g21021(.A(new_n23457_), .B(new_n23456_), .Y(new_n23458_));
  AOI21X1  g21022(.A0(new_n14646_), .A1(new_n14590_), .B0(new_n23458_), .Y(new_n23459_));
  INVX1    g21023(.A(new_n23453_), .Y(new_n23460_));
  AND2X1   g21024(.A(pi0947), .B(pi0614), .Y(new_n23461_));
  AOI22X1  g21025(.A0(new_n23461_), .A1(new_n23420_), .B0(new_n23456_), .B1(new_n12057_), .Y(new_n23462_));
  NOR3X1   g21026(.A(new_n23462_), .B(new_n2437_), .C(pi0216), .Y(new_n23463_));
  AOI21X1  g21027(.A0(new_n23460_), .A1(new_n12077_), .B0(new_n23463_), .Y(new_n23464_));
  OAI21X1  g21028(.A0(new_n23459_), .A1(new_n2438_), .B0(new_n23464_), .Y(new_n23465_));
  AND2X1   g21029(.A(new_n23465_), .B(new_n2954_), .Y(new_n23466_));
  AOI22X1  g21030(.A0(new_n12144_), .A1(new_n5028_), .B0(new_n11950_), .B1(pi0614), .Y(new_n23467_));
  OAI21X1  g21031(.A0(new_n11966_), .A1(new_n5028_), .B0(new_n23467_), .Y(new_n23468_));
  NOR2X1   g21032(.A(new_n11965_), .B(pi0614), .Y(new_n23469_));
  AOI22X1  g21033(.A0(new_n23469_), .A1(new_n5030_), .B0(new_n23468_), .B1(new_n12034_), .Y(new_n23470_));
  OAI21X1  g21034(.A0(new_n23452_), .A1(pi0947), .B0(pi0216), .Y(new_n23471_));
  AOI21X1  g21035(.A0(new_n23470_), .A1(pi0947), .B0(new_n23471_), .Y(new_n23472_));
  NAND3X1  g21036(.A(new_n11974_), .B(pi0907), .C(pi0662), .Y(new_n23473_));
  NOR2X1   g21037(.A(new_n12052_), .B(new_n14590_), .Y(new_n23474_));
  OAI21X1  g21038(.A0(new_n12049_), .A1(new_n12003_), .B0(new_n23474_), .Y(new_n23475_));
  OAI21X1  g21039(.A0(new_n12145_), .A1(new_n14590_), .B0(new_n23475_), .Y(new_n23476_));
  AOI21X1  g21040(.A0(new_n23473_), .A1(new_n14590_), .B0(new_n23476_), .Y(new_n23477_));
  OAI21X1  g21041(.A0(new_n23477_), .A1(pi0216), .B0(pi0215), .Y(new_n23478_));
  AOI21X1  g21042(.A0(new_n23472_), .A1(new_n23379_), .B0(new_n23478_), .Y(new_n23479_));
  NOR3X1   g21043(.A(new_n23479_), .B(new_n23466_), .C(new_n2953_), .Y(new_n23480_));
  OR2X1    g21044(.A(new_n12048_), .B(new_n12036_), .Y(new_n23481_));
  AND2X1   g21045(.A(new_n12055_), .B(new_n14590_), .Y(new_n23482_));
  AOI22X1  g21046(.A0(new_n23482_), .A1(new_n23452_), .B0(new_n23481_), .B1(pi0947), .Y(new_n23483_));
  OAI21X1  g21047(.A0(new_n12062_), .A1(new_n12058_), .B0(new_n14590_), .Y(new_n23484_));
  NOR3X1   g21048(.A(new_n23457_), .B(new_n23456_), .C(new_n5050_), .Y(new_n23485_));
  AOI21X1  g21049(.A0(new_n23485_), .A1(new_n23484_), .B0(new_n2970_), .Y(new_n23486_));
  OAI21X1  g21050(.A0(new_n23483_), .A1(new_n5051_), .B0(new_n23486_), .Y(new_n23487_));
  NOR2X1   g21051(.A(new_n23453_), .B(new_n2971_), .Y(new_n23488_));
  NOR3X1   g21052(.A(new_n23488_), .B(new_n23396_), .C(pi0223), .Y(new_n23489_));
  NAND3X1  g21053(.A(new_n11972_), .B(new_n11967_), .C(new_n11950_), .Y(new_n23490_));
  AND2X1   g21054(.A(new_n12006_), .B(new_n5282_), .Y(new_n23491_));
  OAI21X1  g21055(.A0(new_n12135_), .A1(new_n5282_), .B0(new_n12051_), .Y(new_n23492_));
  AOI21X1  g21056(.A0(new_n23491_), .A1(new_n23490_), .B0(new_n23492_), .Y(new_n23493_));
  OR2X1    g21057(.A(new_n23493_), .B(new_n5051_), .Y(new_n23494_));
  AOI21X1  g21058(.A0(new_n23470_), .A1(new_n5051_), .B0(new_n14590_), .Y(new_n23495_));
  AOI22X1  g21059(.A0(new_n23495_), .A1(new_n23494_), .B0(new_n14686_), .B1(new_n14590_), .Y(new_n23496_));
  OAI21X1  g21060(.A0(new_n23452_), .A1(pi0947), .B0(pi0223), .Y(new_n23497_));
  OAI21X1  g21061(.A0(new_n23497_), .A1(new_n23496_), .B0(pi0216), .Y(new_n23498_));
  AOI21X1  g21062(.A0(new_n23489_), .A1(new_n23487_), .B0(new_n23498_), .Y(new_n23499_));
  INVX1    g21063(.A(new_n23456_), .Y(new_n23500_));
  AOI21X1  g21064(.A0(new_n12053_), .A1(pi0947), .B0(new_n5051_), .Y(new_n23501_));
  OAI21X1  g21065(.A0(new_n23500_), .A1(new_n12033_), .B0(new_n23501_), .Y(new_n23502_));
  AOI21X1  g21066(.A0(new_n23462_), .A1(new_n5051_), .B0(new_n2970_), .Y(new_n23503_));
  INVX1    g21067(.A(new_n23488_), .Y(new_n23504_));
  OAI21X1  g21068(.A0(new_n23504_), .A1(new_n11953_), .B0(new_n2964_), .Y(new_n23505_));
  AOI21X1  g21069(.A0(new_n23503_), .A1(new_n23502_), .B0(new_n23505_), .Y(new_n23506_));
  OR2X1    g21070(.A(new_n23452_), .B(new_n23428_), .Y(new_n23507_));
  INVX1    g21071(.A(new_n23430_), .Y(new_n23508_));
  OAI21X1  g21072(.A0(new_n23508_), .A1(new_n5050_), .B0(new_n23475_), .Y(new_n23509_));
  AOI21X1  g21073(.A0(new_n23507_), .A1(new_n14590_), .B0(new_n23509_), .Y(new_n23510_));
  OAI21X1  g21074(.A0(new_n23510_), .A1(new_n2964_), .B0(new_n2438_), .Y(new_n23511_));
  OAI21X1  g21075(.A0(new_n23511_), .A1(new_n23506_), .B0(new_n2953_), .Y(new_n23512_));
  OAI21X1  g21076(.A0(new_n23512_), .A1(new_n23499_), .B0(pi0039), .Y(new_n23513_));
  AOI21X1  g21077(.A0(new_n23460_), .A1(new_n11943_), .B0(new_n2953_), .Y(new_n23514_));
  OAI21X1  g21078(.A0(new_n11943_), .A1(new_n2438_), .B0(new_n23514_), .Y(new_n23515_));
  NAND3X1  g21079(.A(new_n23460_), .B(new_n11945_), .C(new_n11944_), .Y(new_n23516_));
  AOI21X1  g21080(.A0(new_n12445_), .A1(pi0216), .B0(pi0299), .Y(new_n23517_));
  AOI21X1  g21081(.A0(new_n23517_), .A1(new_n23516_), .B0(pi0039), .Y(new_n23518_));
  AOI21X1  g21082(.A0(new_n23518_), .A1(new_n23515_), .B0(pi0038), .Y(new_n23519_));
  OAI21X1  g21083(.A0(new_n23513_), .A1(new_n23480_), .B0(new_n23519_), .Y(new_n23520_));
  AND2X1   g21084(.A(new_n23520_), .B(new_n23455_), .Y(new_n23521_));
  MX2X1    g21085(.A(new_n23521_), .B(pi0216), .S0(new_n9580_), .Y(po0373));
  INVX1    g21086(.A(pi0695), .Y(new_n23523_));
  OAI21X1  g21087(.A0(new_n23176_), .A1(new_n23523_), .B0(new_n6637_), .Y(new_n23524_));
  AOI21X1  g21088(.A0(new_n23174_), .A1(new_n23523_), .B0(new_n23524_), .Y(new_n23525_));
  INVX1    g21089(.A(pi0612), .Y(new_n23526_));
  OAI21X1  g21090(.A0(new_n23243_), .A1(pi0695), .B0(pi0217), .Y(new_n23527_));
  NAND2X1  g21091(.A(new_n23527_), .B(new_n23526_), .Y(new_n23528_));
  AOI21X1  g21092(.A0(new_n23194_), .A1(new_n23192_), .B0(pi0695), .Y(new_n23529_));
  OAI21X1  g21093(.A0(new_n23201_), .A1(new_n23523_), .B0(new_n6637_), .Y(new_n23530_));
  OR2X1    g21094(.A(new_n23530_), .B(new_n23529_), .Y(new_n23531_));
  AOI21X1  g21095(.A0(new_n23247_), .A1(pi0695), .B0(new_n6637_), .Y(new_n23532_));
  OAI21X1  g21096(.A0(new_n23232_), .A1(pi0695), .B0(new_n23532_), .Y(new_n23533_));
  NAND3X1  g21097(.A(new_n23533_), .B(new_n23531_), .C(pi0612), .Y(new_n23534_));
  OAI21X1  g21098(.A0(new_n23528_), .A1(new_n23525_), .B0(new_n23534_), .Y(po0374));
  MX2X1    g21099(.A(new_n22788_), .B(new_n22747_), .S0(new_n22726_), .Y(new_n23536_));
  NOR4X1   g21100(.A(new_n22791_), .B(new_n22790_), .C(new_n22726_), .D(new_n22713_), .Y(new_n23537_));
  MX2X1    g21101(.A(new_n23536_), .B(new_n23537_), .S0(pi0218), .Y(po0375));
  INVX1    g21102(.A(pi0219), .Y(new_n23539_));
  NAND3X1  g21103(.A(new_n5117_), .B(new_n23539_), .C(new_n2436_), .Y(new_n23540_));
  OR2X1    g21104(.A(new_n23337_), .B(new_n22271_), .Y(new_n23541_));
  AOI21X1  g21105(.A0(new_n23336_), .A1(new_n22271_), .B0(new_n22270_), .Y(new_n23542_));
  NOR4X1   g21106(.A(new_n14675_), .B(new_n3810_), .C(pi0637), .D(new_n22271_), .Y(new_n23543_));
  AOI21X1  g21107(.A0(new_n23542_), .A1(new_n23541_), .B0(new_n23543_), .Y(new_n23544_));
  OAI21X1  g21108(.A0(new_n23329_), .A1(new_n22271_), .B0(pi0637), .Y(new_n23545_));
  AOI21X1  g21109(.A0(new_n23328_), .A1(new_n22271_), .B0(new_n23545_), .Y(new_n23546_));
  OAI21X1  g21110(.A0(new_n22804_), .A1(pi0617), .B0(new_n22270_), .Y(new_n23547_));
  AOI21X1  g21111(.A0(new_n23332_), .A1(pi0617), .B0(new_n23547_), .Y(new_n23548_));
  NOR3X1   g21112(.A(new_n23548_), .B(new_n23546_), .C(po1038), .Y(new_n23549_));
  OAI22X1  g21113(.A0(new_n23549_), .A1(new_n23539_), .B0(new_n23544_), .B1(new_n23540_), .Y(po0376));
  INVX1    g21114(.A(pi0220), .Y(new_n23551_));
  MX2X1    g21115(.A(new_n22710_), .B(new_n22609_), .S0(new_n22799_), .Y(new_n23552_));
  NOR4X1   g21116(.A(new_n22799_), .B(new_n22714_), .C(new_n22713_), .D(new_n22712_), .Y(new_n23553_));
  MX2X1    g21117(.A(new_n23553_), .B(new_n23552_), .S0(new_n23551_), .Y(po0377));
  AND2X1   g21118(.A(pi0907), .B(pi0661), .Y(new_n23555_));
  AND2X1   g21119(.A(pi0947), .B(pi0616), .Y(new_n23556_));
  AOI21X1  g21120(.A0(new_n23555_), .A1(new_n14590_), .B0(new_n23556_), .Y(new_n23557_));
  AOI21X1  g21121(.A0(new_n12901_), .A1(pi0221), .B0(new_n2996_), .Y(new_n23558_));
  OAI21X1  g21122(.A0(new_n23557_), .A1(new_n12901_), .B0(new_n23558_), .Y(new_n23559_));
  AND2X1   g21123(.A(new_n23555_), .B(new_n14590_), .Y(new_n23560_));
  OR2X1    g21124(.A(new_n12032_), .B(new_n11995_), .Y(new_n23561_));
  OAI21X1  g21125(.A0(new_n12050_), .A1(new_n23481_), .B0(new_n12000_), .Y(new_n23562_));
  AOI21X1  g21126(.A0(new_n23562_), .A1(new_n23561_), .B0(new_n14590_), .Y(new_n23563_));
  NOR3X1   g21127(.A(new_n23563_), .B(new_n23482_), .C(new_n5051_), .Y(new_n23564_));
  MX2X1    g21128(.A(new_n12032_), .B(new_n12046_), .S0(new_n5033_), .Y(new_n23565_));
  AND2X1   g21129(.A(new_n12106_), .B(new_n11968_), .Y(new_n23566_));
  OAI21X1  g21130(.A0(new_n23421_), .A1(new_n23566_), .B0(new_n12000_), .Y(new_n23567_));
  AND2X1   g21131(.A(new_n23567_), .B(pi0947), .Y(new_n23568_));
  OAI21X1  g21132(.A0(new_n23565_), .A1(new_n11995_), .B0(new_n23568_), .Y(new_n23569_));
  AOI21X1  g21133(.A0(new_n23569_), .A1(new_n23484_), .B0(new_n5050_), .Y(new_n23570_));
  NOR3X1   g21134(.A(new_n23570_), .B(new_n23564_), .C(new_n23560_), .Y(new_n23571_));
  NOR3X1   g21135(.A(new_n23557_), .B(new_n11952_), .C(new_n2740_), .Y(new_n23572_));
  AOI21X1  g21136(.A0(new_n23572_), .A1(new_n2970_), .B0(pi0223), .Y(new_n23573_));
  INVX1    g21137(.A(new_n23573_), .Y(new_n23574_));
  NOR2X1   g21138(.A(new_n23574_), .B(new_n23396_), .Y(new_n23575_));
  OAI21X1  g21139(.A0(new_n23571_), .A1(new_n2970_), .B0(new_n23575_), .Y(new_n23576_));
  OAI21X1  g21140(.A0(new_n11973_), .A1(new_n11966_), .B0(new_n5282_), .Y(new_n23577_));
  AOI21X1  g21141(.A0(new_n23382_), .A1(new_n11984_), .B0(pi0616), .Y(new_n23578_));
  AOI21X1  g21142(.A0(new_n23578_), .A1(new_n23577_), .B0(new_n14590_), .Y(new_n23579_));
  AOI21X1  g21143(.A0(new_n11991_), .A1(new_n14590_), .B0(new_n23579_), .Y(new_n23580_));
  OR2X1    g21144(.A(new_n23580_), .B(new_n5050_), .Y(new_n23581_));
  OAI21X1  g21145(.A0(new_n12002_), .A1(new_n11996_), .B0(pi0947), .Y(new_n23582_));
  NAND2X1  g21146(.A(new_n23582_), .B(new_n5050_), .Y(new_n23583_));
  AOI21X1  g21147(.A0(new_n12084_), .A1(new_n14590_), .B0(new_n23583_), .Y(new_n23584_));
  NOR3X1   g21148(.A(new_n23584_), .B(new_n23560_), .C(new_n2964_), .Y(new_n23585_));
  AOI21X1  g21149(.A0(new_n23585_), .A1(new_n23581_), .B0(new_n2437_), .Y(new_n23586_));
  INVX1    g21150(.A(new_n23560_), .Y(new_n23587_));
  OAI22X1  g21151(.A0(new_n23411_), .A1(new_n12005_), .B0(new_n12006_), .B1(new_n11993_), .Y(new_n23588_));
  AOI21X1  g21152(.A0(new_n23588_), .A1(pi0947), .B0(new_n5051_), .Y(new_n23589_));
  OAI21X1  g21153(.A0(new_n23587_), .A1(new_n12033_), .B0(new_n23589_), .Y(new_n23590_));
  AOI22X1  g21154(.A0(new_n23556_), .A1(new_n23420_), .B0(new_n23560_), .B1(new_n12057_), .Y(new_n23591_));
  AOI21X1  g21155(.A0(new_n23591_), .A1(new_n5051_), .B0(new_n2970_), .Y(new_n23592_));
  AOI21X1  g21156(.A0(new_n23592_), .A1(new_n23590_), .B0(new_n23574_), .Y(new_n23593_));
  NAND2X1  g21157(.A(new_n12007_), .B(pi0947), .Y(new_n23594_));
  NAND2X1  g21158(.A(new_n23594_), .B(new_n23428_), .Y(new_n23595_));
  AOI22X1  g21159(.A0(new_n23594_), .A1(new_n23587_), .B0(new_n23430_), .B1(new_n5051_), .Y(new_n23596_));
  AOI21X1  g21160(.A0(new_n23596_), .A1(new_n23595_), .B0(new_n2964_), .Y(new_n23597_));
  OR2X1    g21161(.A(new_n23597_), .B(pi0221), .Y(new_n23598_));
  OAI21X1  g21162(.A0(new_n23598_), .A1(new_n23593_), .B0(new_n2953_), .Y(new_n23599_));
  AOI21X1  g21163(.A0(new_n23586_), .A1(new_n23576_), .B0(new_n23599_), .Y(new_n23600_));
  OAI21X1  g21164(.A0(new_n23555_), .A1(new_n14646_), .B0(new_n14590_), .Y(new_n23601_));
  AND2X1   g21165(.A(new_n23569_), .B(pi0221), .Y(new_n23602_));
  AOI21X1  g21166(.A0(new_n23572_), .A1(new_n2438_), .B0(pi0221), .Y(new_n23603_));
  OAI21X1  g21167(.A0(new_n23591_), .A1(new_n2438_), .B0(new_n23603_), .Y(new_n23604_));
  NAND2X1  g21168(.A(new_n23604_), .B(new_n2954_), .Y(new_n23605_));
  AOI21X1  g21169(.A0(new_n23602_), .A1(new_n23601_), .B0(new_n23605_), .Y(new_n23606_));
  NOR4X1   g21170(.A(new_n23579_), .B(new_n23560_), .C(new_n23378_), .D(new_n2437_), .Y(new_n23607_));
  AOI21X1  g21171(.A0(new_n23594_), .A1(new_n23587_), .B0(new_n23430_), .Y(new_n23608_));
  OAI21X1  g21172(.A0(new_n23608_), .A1(pi0221), .B0(pi0215), .Y(new_n23609_));
  OAI21X1  g21173(.A0(new_n23609_), .A1(new_n23607_), .B0(pi0299), .Y(new_n23610_));
  OAI21X1  g21174(.A0(new_n23610_), .A1(new_n23606_), .B0(pi0039), .Y(new_n23611_));
  AOI21X1  g21175(.A0(new_n11942_), .A1(new_n11929_), .B0(new_n2437_), .Y(new_n23612_));
  OAI21X1  g21176(.A0(new_n23557_), .A1(new_n12091_), .B0(pi0299), .Y(new_n23613_));
  OR2X1    g21177(.A(new_n23613_), .B(new_n23612_), .Y(new_n23614_));
  OR2X1    g21178(.A(new_n23557_), .B(new_n12445_), .Y(new_n23615_));
  AOI21X1  g21179(.A0(new_n12445_), .A1(pi0221), .B0(pi0299), .Y(new_n23616_));
  AOI21X1  g21180(.A0(new_n23616_), .A1(new_n23615_), .B0(pi0039), .Y(new_n23617_));
  AOI21X1  g21181(.A0(new_n23617_), .A1(new_n23614_), .B0(pi0038), .Y(new_n23618_));
  OAI21X1  g21182(.A0(new_n23611_), .A1(new_n23600_), .B0(new_n23618_), .Y(new_n23619_));
  AND2X1   g21183(.A(new_n23619_), .B(new_n23559_), .Y(new_n23620_));
  MX2X1    g21184(.A(new_n23620_), .B(pi0221), .S0(new_n9580_), .Y(po0378));
  MX2X1    g21185(.A(new_n14929_), .B(new_n12010_), .S0(pi0223), .Y(new_n23622_));
  AOI21X1  g21186(.A0(new_n23622_), .A1(new_n2953_), .B0(new_n2959_), .Y(new_n23623_));
  NAND2X1  g21187(.A(new_n12914_), .B(new_n2996_), .Y(new_n23624_));
  AOI21X1  g21188(.A0(new_n23623_), .A1(new_n12088_), .B0(new_n23624_), .Y(new_n23625_));
  NOR2X1   g21189(.A(new_n23625_), .B(new_n21881_), .Y(new_n23626_));
  NOR2X1   g21190(.A(new_n23626_), .B(new_n2960_), .Y(new_n23627_));
  INVX1    g21191(.A(new_n23382_), .Y(new_n23628_));
  MX2X1    g21192(.A(new_n23565_), .B(new_n12291_), .S0(pi0616), .Y(new_n23629_));
  NOR3X1   g21193(.A(new_n12108_), .B(new_n11950_), .C(new_n5027_), .Y(new_n23630_));
  OAI21X1  g21194(.A0(new_n23630_), .A1(new_n12116_), .B0(new_n12115_), .Y(new_n23631_));
  AOI21X1  g21195(.A0(new_n23631_), .A1(new_n11978_), .B0(new_n23628_), .Y(new_n23632_));
  OAI21X1  g21196(.A0(new_n23629_), .A1(new_n11978_), .B0(new_n23632_), .Y(new_n23633_));
  INVX1    g21197(.A(new_n23633_), .Y(new_n23634_));
  AOI21X1  g21198(.A0(new_n23629_), .A1(new_n23628_), .B0(new_n23634_), .Y(new_n23635_));
  INVX1    g21199(.A(new_n23635_), .Y(new_n23636_));
  INVX1    g21200(.A(new_n12121_), .Y(new_n23637_));
  MX2X1    g21201(.A(new_n23637_), .B(new_n12070_), .S0(new_n11950_), .Y(new_n23638_));
  INVX1    g21202(.A(new_n23638_), .Y(new_n23639_));
  NOR3X1   g21203(.A(new_n23630_), .B(new_n5029_), .C(pi0662), .Y(new_n23640_));
  AOI21X1  g21204(.A0(new_n23640_), .A1(new_n12029_), .B0(new_n23628_), .Y(new_n23641_));
  OAI21X1  g21205(.A0(new_n23639_), .A1(new_n11978_), .B0(new_n23641_), .Y(new_n23642_));
  OAI21X1  g21206(.A0(new_n23638_), .A1(new_n23382_), .B0(new_n23642_), .Y(new_n23643_));
  OR2X1    g21207(.A(new_n23643_), .B(new_n5071_), .Y(new_n23644_));
  AND2X1   g21208(.A(new_n23644_), .B(pi0222), .Y(new_n23645_));
  OAI21X1  g21209(.A0(new_n23636_), .A1(new_n5070_), .B0(new_n23645_), .Y(new_n23646_));
  MX2X1    g21210(.A(new_n12181_), .B(new_n12364_), .S0(new_n5030_), .Y(new_n23647_));
  NOR2X1   g21211(.A(new_n23647_), .B(new_n11950_), .Y(new_n23648_));
  NOR2X1   g21212(.A(new_n23648_), .B(new_n5071_), .Y(new_n23649_));
  INVX1    g21213(.A(new_n23649_), .Y(new_n23650_));
  AND2X1   g21214(.A(new_n23630_), .B(new_n12056_), .Y(new_n23651_));
  INVX1    g21215(.A(new_n23651_), .Y(new_n23652_));
  NAND3X1  g21216(.A(new_n23630_), .B(new_n12056_), .C(new_n11983_), .Y(new_n23653_));
  OR4X1    g21217(.A(new_n12116_), .B(new_n11983_), .C(new_n11950_), .D(new_n5027_), .Y(new_n23654_));
  NAND3X1  g21218(.A(new_n23654_), .B(new_n23653_), .C(new_n23382_), .Y(new_n23655_));
  INVX1    g21219(.A(new_n23655_), .Y(new_n23656_));
  AOI21X1  g21220(.A0(new_n23652_), .A1(new_n23628_), .B0(new_n23656_), .Y(new_n23657_));
  OR2X1    g21221(.A(new_n23657_), .B(new_n5070_), .Y(new_n23658_));
  AND2X1   g21222(.A(new_n23658_), .B(new_n2960_), .Y(new_n23659_));
  AOI21X1  g21223(.A0(new_n23659_), .A1(new_n23650_), .B0(new_n10136_), .Y(new_n23660_));
  NOR4X1   g21224(.A(new_n12171_), .B(new_n11952_), .C(new_n2740_), .D(new_n11950_), .Y(new_n23661_));
  INVX1    g21225(.A(new_n23661_), .Y(new_n23662_));
  AOI21X1  g21226(.A0(new_n11953_), .A1(pi0222), .B0(new_n10137_), .Y(new_n23663_));
  AOI21X1  g21227(.A0(new_n23663_), .A1(new_n23662_), .B0(pi0215), .Y(new_n23664_));
  INVX1    g21228(.A(new_n23664_), .Y(new_n23665_));
  AOI21X1  g21229(.A0(new_n23660_), .A1(new_n23646_), .B0(new_n23665_), .Y(new_n23666_));
  NOR4X1   g21230(.A(new_n12171_), .B(new_n11952_), .C(new_n5030_), .D(new_n2740_), .Y(new_n23667_));
  OAI21X1  g21231(.A0(new_n23667_), .A1(new_n12182_), .B0(pi0616), .Y(new_n23668_));
  NOR3X1   g21232(.A(new_n23668_), .B(new_n12186_), .C(pi0222), .Y(new_n23669_));
  INVX1    g21233(.A(new_n12146_), .Y(new_n23670_));
  AOI21X1  g21234(.A0(new_n23670_), .A1(pi0616), .B0(new_n11988_), .Y(new_n23671_));
  INVX1    g21235(.A(new_n23671_), .Y(new_n23672_));
  AOI21X1  g21236(.A0(new_n23670_), .A1(pi0616), .B0(new_n11984_), .Y(new_n23673_));
  OAI21X1  g21237(.A0(new_n11974_), .A1(new_n11978_), .B0(new_n23673_), .Y(new_n23674_));
  AND2X1   g21238(.A(new_n23674_), .B(new_n23382_), .Y(new_n23675_));
  AOI21X1  g21239(.A0(new_n23672_), .A1(new_n23628_), .B0(new_n23675_), .Y(new_n23676_));
  AND2X1   g21240(.A(new_n23676_), .B(new_n5071_), .Y(new_n23677_));
  INVX1    g21241(.A(new_n23677_), .Y(new_n23678_));
  AOI21X1  g21242(.A0(new_n12121_), .A1(pi0616), .B0(new_n11998_), .Y(new_n23679_));
  INVX1    g21243(.A(new_n23679_), .Y(new_n23680_));
  AOI21X1  g21244(.A0(new_n23640_), .A1(new_n12135_), .B0(new_n23628_), .Y(new_n23681_));
  OAI21X1  g21245(.A0(new_n23680_), .A1(new_n11978_), .B0(new_n23681_), .Y(new_n23682_));
  INVX1    g21246(.A(new_n23682_), .Y(new_n23683_));
  AOI21X1  g21247(.A0(new_n23680_), .A1(new_n23628_), .B0(new_n23683_), .Y(new_n23684_));
  AOI21X1  g21248(.A0(new_n23684_), .A1(new_n5070_), .B0(new_n2960_), .Y(new_n23685_));
  AOI21X1  g21249(.A0(new_n23685_), .A1(new_n23678_), .B0(new_n23669_), .Y(new_n23686_));
  OAI21X1  g21250(.A0(new_n23686_), .A1(new_n2954_), .B0(pi0299), .Y(new_n23687_));
  OR2X1    g21251(.A(new_n23687_), .B(new_n23666_), .Y(new_n23688_));
  OAI21X1  g21252(.A0(new_n23643_), .A1(new_n5051_), .B0(pi0222), .Y(new_n23689_));
  AOI21X1  g21253(.A0(new_n23635_), .A1(new_n5051_), .B0(new_n23689_), .Y(new_n23690_));
  NAND2X1  g21254(.A(new_n23648_), .B(new_n5050_), .Y(new_n23691_));
  AOI21X1  g21255(.A0(new_n23657_), .A1(new_n5051_), .B0(new_n2961_), .Y(new_n23692_));
  AOI21X1  g21256(.A0(new_n23662_), .A1(new_n2961_), .B0(pi0222), .Y(new_n23693_));
  INVX1    g21257(.A(new_n23693_), .Y(new_n23694_));
  AOI21X1  g21258(.A0(new_n23692_), .A1(new_n23691_), .B0(new_n23694_), .Y(new_n23695_));
  NOR2X1   g21259(.A(new_n23695_), .B(pi0223), .Y(new_n23696_));
  INVX1    g21260(.A(new_n23696_), .Y(new_n23697_));
  NAND2X1  g21261(.A(new_n23676_), .B(new_n5051_), .Y(new_n23698_));
  AOI21X1  g21262(.A0(new_n23684_), .A1(new_n5050_), .B0(new_n2960_), .Y(new_n23699_));
  AND2X1   g21263(.A(new_n23699_), .B(new_n23698_), .Y(new_n23700_));
  NOR3X1   g21264(.A(new_n23668_), .B(new_n12194_), .C(pi0222), .Y(new_n23701_));
  NOR2X1   g21265(.A(new_n23701_), .B(new_n2964_), .Y(new_n23702_));
  INVX1    g21266(.A(new_n23702_), .Y(new_n23703_));
  OAI22X1  g21267(.A0(new_n23703_), .A1(new_n23700_), .B0(new_n23697_), .B1(new_n23690_), .Y(new_n23704_));
  AOI21X1  g21268(.A0(new_n23704_), .A1(new_n2953_), .B0(new_n2959_), .Y(new_n23705_));
  AND2X1   g21269(.A(new_n12104_), .B(pi0222), .Y(new_n23706_));
  AOI21X1  g21270(.A0(new_n13683_), .A1(new_n2960_), .B0(pi0039), .Y(new_n23707_));
  OAI21X1  g21271(.A0(new_n13683_), .A1(pi0616), .B0(new_n23707_), .Y(new_n23708_));
  OAI21X1  g21272(.A0(new_n23708_), .A1(new_n23706_), .B0(new_n2996_), .Y(new_n23709_));
  AOI21X1  g21273(.A0(new_n23705_), .A1(new_n23688_), .B0(new_n23709_), .Y(new_n23710_));
  AOI21X1  g21274(.A0(new_n12901_), .A1(pi0222), .B0(new_n2996_), .Y(new_n23711_));
  INVX1    g21275(.A(new_n23711_), .Y(new_n23712_));
  AND2X1   g21276(.A(new_n12205_), .B(pi0616), .Y(new_n23713_));
  OAI21X1  g21277(.A0(new_n23713_), .A1(new_n23712_), .B0(new_n3129_), .Y(new_n23714_));
  OAI22X1  g21278(.A0(new_n23714_), .A1(new_n23710_), .B0(new_n3129_), .B1(new_n2960_), .Y(new_n23715_));
  MX2X1    g21279(.A(new_n23715_), .B(new_n23627_), .S0(new_n12601_), .Y(new_n23716_));
  INVX1    g21280(.A(new_n23627_), .Y(new_n23717_));
  AOI21X1  g21281(.A0(new_n23717_), .A1(new_n12590_), .B0(new_n12591_), .Y(new_n23718_));
  OAI21X1  g21282(.A0(new_n23716_), .A1(new_n12590_), .B0(new_n23718_), .Y(new_n23719_));
  AOI21X1  g21283(.A0(new_n23717_), .A1(pi0609), .B0(pi1155), .Y(new_n23720_));
  OAI21X1  g21284(.A0(new_n23716_), .A1(pi0609), .B0(new_n23720_), .Y(new_n23721_));
  NAND2X1  g21285(.A(new_n23721_), .B(new_n23719_), .Y(new_n23722_));
  MX2X1    g21286(.A(new_n23722_), .B(new_n23716_), .S0(new_n11888_), .Y(new_n23723_));
  AOI21X1  g21287(.A0(new_n23717_), .A1(new_n12614_), .B0(new_n12615_), .Y(new_n23724_));
  OAI21X1  g21288(.A0(new_n23723_), .A1(new_n12614_), .B0(new_n23724_), .Y(new_n23725_));
  AOI21X1  g21289(.A0(new_n23717_), .A1(pi0618), .B0(pi1154), .Y(new_n23726_));
  OAI21X1  g21290(.A0(new_n23723_), .A1(pi0618), .B0(new_n23726_), .Y(new_n23727_));
  AOI21X1  g21291(.A0(new_n23727_), .A1(new_n23725_), .B0(new_n11887_), .Y(new_n23728_));
  AOI21X1  g21292(.A0(new_n23723_), .A1(new_n11887_), .B0(new_n23728_), .Y(new_n23729_));
  OAI21X1  g21293(.A0(new_n23627_), .A1(pi0619), .B0(pi1159), .Y(new_n23730_));
  AOI21X1  g21294(.A0(new_n23729_), .A1(pi0619), .B0(new_n23730_), .Y(new_n23731_));
  OAI21X1  g21295(.A0(new_n23627_), .A1(new_n12637_), .B0(new_n12638_), .Y(new_n23732_));
  AOI21X1  g21296(.A0(new_n23729_), .A1(new_n12637_), .B0(new_n23732_), .Y(new_n23733_));
  NOR2X1   g21297(.A(new_n23733_), .B(new_n23731_), .Y(new_n23734_));
  MX2X1    g21298(.A(new_n23734_), .B(new_n23729_), .S0(new_n11886_), .Y(new_n23735_));
  INVX1    g21299(.A(new_n23735_), .Y(new_n23736_));
  MX2X1    g21300(.A(new_n23736_), .B(new_n23627_), .S0(new_n12841_), .Y(new_n23737_));
  NAND2X1  g21301(.A(new_n23737_), .B(new_n14394_), .Y(new_n23738_));
  AND2X1   g21302(.A(pi0680), .B(pi0661), .Y(new_n23739_));
  OR2X1    g21303(.A(new_n23739_), .B(new_n12458_), .Y(new_n23740_));
  NAND2X1  g21304(.A(new_n12458_), .B(new_n2960_), .Y(new_n23741_));
  AOI21X1  g21305(.A0(new_n13228_), .A1(pi0222), .B0(pi0299), .Y(new_n23742_));
  NAND3X1  g21306(.A(new_n23742_), .B(new_n23741_), .C(new_n23740_), .Y(new_n23743_));
  INVX1    g21307(.A(new_n23739_), .Y(new_n23744_));
  NAND2X1  g21308(.A(new_n23744_), .B(new_n12463_), .Y(new_n23745_));
  OR2X1    g21309(.A(new_n12463_), .B(pi0222), .Y(new_n23746_));
  AOI21X1  g21310(.A0(new_n13240_), .A1(pi0222), .B0(new_n2953_), .Y(new_n23747_));
  NAND3X1  g21311(.A(new_n23747_), .B(new_n23746_), .C(new_n23745_), .Y(new_n23748_));
  NAND3X1  g21312(.A(new_n23748_), .B(new_n23743_), .C(new_n2959_), .Y(new_n23749_));
  NAND3X1  g21313(.A(new_n12047_), .B(pi0680), .C(new_n11977_), .Y(new_n23750_));
  OAI21X1  g21314(.A0(new_n12071_), .A1(new_n11978_), .B0(new_n23750_), .Y(new_n23751_));
  AND2X1   g21315(.A(new_n12033_), .B(pi0681), .Y(new_n23752_));
  MX2X1    g21316(.A(new_n12943_), .B(new_n23752_), .S0(new_n11976_), .Y(new_n23753_));
  AOI21X1  g21317(.A0(new_n23751_), .A1(new_n23382_), .B0(new_n23753_), .Y(new_n23754_));
  AND2X1   g21318(.A(new_n23754_), .B(new_n5050_), .Y(new_n23755_));
  MX2X1    g21319(.A(new_n12404_), .B(new_n12057_), .S0(new_n5029_), .Y(new_n23756_));
  OR2X1    g21320(.A(new_n23756_), .B(new_n11976_), .Y(new_n23757_));
  OAI21X1  g21321(.A0(new_n12063_), .A1(pi0661), .B0(new_n23757_), .Y(new_n23758_));
  OAI21X1  g21322(.A0(new_n23758_), .A1(new_n5050_), .B0(pi0222), .Y(new_n23759_));
  OR4X1    g21323(.A(new_n12502_), .B(new_n5051_), .C(new_n5029_), .D(new_n11976_), .Y(new_n23760_));
  OR4X1    g21324(.A(new_n12499_), .B(new_n12260_), .C(new_n5050_), .D(new_n11976_), .Y(new_n23761_));
  NAND3X1  g21325(.A(new_n23761_), .B(new_n23760_), .C(pi0224), .Y(new_n23762_));
  OR4X1    g21326(.A(new_n12499_), .B(new_n11952_), .C(new_n2740_), .D(new_n11976_), .Y(new_n23763_));
  AOI21X1  g21327(.A0(new_n23763_), .A1(new_n2961_), .B0(pi0222), .Y(new_n23764_));
  AOI21X1  g21328(.A0(new_n23764_), .A1(new_n23762_), .B0(pi0223), .Y(new_n23765_));
  OAI21X1  g21329(.A0(new_n23759_), .A1(new_n23755_), .B0(new_n23765_), .Y(new_n23766_));
  OAI22X1  g21330(.A0(new_n12526_), .A1(new_n12224_), .B0(new_n12229_), .B1(pi0680), .Y(new_n23767_));
  INVX1    g21331(.A(new_n23767_), .Y(new_n23768_));
  MX2X1    g21332(.A(new_n23768_), .B(new_n12084_), .S0(new_n11976_), .Y(new_n23769_));
  AND2X1   g21333(.A(new_n23769_), .B(new_n5050_), .Y(new_n23770_));
  NOR2X1   g21334(.A(new_n23628_), .B(new_n11986_), .Y(new_n23771_));
  MX2X1    g21335(.A(new_n12545_), .B(new_n11975_), .S0(new_n11976_), .Y(new_n23772_));
  NOR3X1   g21336(.A(new_n23772_), .B(new_n23771_), .C(new_n5050_), .Y(new_n23773_));
  OR2X1    g21337(.A(new_n23773_), .B(new_n2960_), .Y(new_n23774_));
  AND2X1   g21338(.A(pi0661), .B(new_n2960_), .Y(new_n23775_));
  AOI21X1  g21339(.A0(new_n23775_), .A1(new_n12510_), .B0(new_n2964_), .Y(new_n23776_));
  OAI21X1  g21340(.A0(new_n23774_), .A1(new_n23770_), .B0(new_n23776_), .Y(new_n23777_));
  AOI21X1  g21341(.A0(new_n23777_), .A1(new_n23766_), .B0(pi0299), .Y(new_n23778_));
  OAI21X1  g21342(.A0(new_n23758_), .A1(new_n5070_), .B0(pi0222), .Y(new_n23779_));
  AOI21X1  g21343(.A0(new_n23754_), .A1(new_n5070_), .B0(new_n23779_), .Y(new_n23780_));
  OAI21X1  g21344(.A0(new_n12506_), .A1(new_n11976_), .B0(new_n5071_), .Y(new_n23781_));
  OAI21X1  g21345(.A0(new_n23744_), .A1(new_n12502_), .B0(new_n5070_), .Y(new_n23782_));
  NAND3X1  g21346(.A(new_n23782_), .B(new_n23781_), .C(new_n2960_), .Y(new_n23783_));
  NAND2X1  g21347(.A(new_n23783_), .B(new_n10137_), .Y(new_n23784_));
  OR2X1    g21348(.A(new_n23784_), .B(new_n23780_), .Y(new_n23785_));
  AOI21X1  g21349(.A0(new_n23763_), .A1(new_n23663_), .B0(pi0215), .Y(new_n23786_));
  NAND2X1  g21350(.A(new_n23769_), .B(new_n5070_), .Y(new_n23787_));
  NOR3X1   g21351(.A(new_n23772_), .B(new_n23771_), .C(new_n5070_), .Y(new_n23788_));
  NOR2X1   g21352(.A(new_n23788_), .B(new_n2960_), .Y(new_n23789_));
  AOI22X1  g21353(.A0(new_n23789_), .A1(new_n23787_), .B0(new_n23775_), .B1(new_n12518_), .Y(new_n23790_));
  OAI21X1  g21354(.A0(new_n23790_), .A1(new_n2954_), .B0(pi0299), .Y(new_n23791_));
  AOI21X1  g21355(.A0(new_n23786_), .A1(new_n23785_), .B0(new_n23791_), .Y(new_n23792_));
  OAI21X1  g21356(.A0(new_n23792_), .A1(new_n23778_), .B0(pi0039), .Y(new_n23793_));
  AOI21X1  g21357(.A0(new_n23793_), .A1(new_n23749_), .B0(pi0038), .Y(new_n23794_));
  NOR4X1   g21358(.A(new_n13585_), .B(new_n3074_), .C(new_n11976_), .D(pi0039), .Y(new_n23795_));
  OAI21X1  g21359(.A0(new_n23795_), .A1(new_n23712_), .B0(new_n3129_), .Y(new_n23796_));
  OAI22X1  g21360(.A0(new_n23796_), .A1(new_n23794_), .B0(new_n3129_), .B1(new_n2960_), .Y(new_n23797_));
  AND2X1   g21361(.A(new_n23797_), .B(new_n11889_), .Y(new_n23798_));
  AOI21X1  g21362(.A0(new_n23717_), .A1(new_n12493_), .B0(new_n12494_), .Y(new_n23799_));
  OAI21X1  g21363(.A0(new_n23797_), .A1(new_n12493_), .B0(new_n23799_), .Y(new_n23800_));
  AOI21X1  g21364(.A0(new_n23717_), .A1(pi0625), .B0(pi1153), .Y(new_n23801_));
  OAI21X1  g21365(.A0(new_n23797_), .A1(pi0625), .B0(new_n23801_), .Y(new_n23802_));
  AOI21X1  g21366(.A0(new_n23802_), .A1(new_n23800_), .B0(new_n11889_), .Y(new_n23803_));
  NOR2X1   g21367(.A(new_n23803_), .B(new_n23798_), .Y(new_n23804_));
  MX2X1    g21368(.A(new_n23804_), .B(new_n23717_), .S0(new_n12618_), .Y(new_n23805_));
  OR4X1    g21369(.A(new_n23626_), .B(new_n12640_), .C(new_n12639_), .D(new_n2960_), .Y(new_n23806_));
  OAI21X1  g21370(.A0(new_n23805_), .A1(new_n12641_), .B0(new_n23806_), .Y(new_n23807_));
  NOR2X1   g21371(.A(new_n23807_), .B(new_n12659_), .Y(new_n23808_));
  AOI22X1  g21372(.A0(new_n23808_), .A1(new_n17252_), .B0(new_n23717_), .B1(new_n22010_), .Y(new_n23809_));
  AOI21X1  g21373(.A0(new_n23717_), .A1(pi0628), .B0(new_n12710_), .Y(new_n23810_));
  OAI21X1  g21374(.A0(new_n23809_), .A1(pi0628), .B0(new_n23810_), .Y(new_n23811_));
  AOI21X1  g21375(.A0(new_n23717_), .A1(new_n12683_), .B0(new_n12708_), .Y(new_n23812_));
  OAI21X1  g21376(.A0(new_n23809_), .A1(new_n12683_), .B0(new_n23812_), .Y(new_n23813_));
  NAND3X1  g21377(.A(new_n23813_), .B(new_n23811_), .C(new_n23738_), .Y(new_n23814_));
  INVX1    g21378(.A(new_n23629_), .Y(new_n23815_));
  AOI21X1  g21379(.A0(new_n12252_), .A1(new_n5033_), .B0(new_n12220_), .Y(new_n23816_));
  INVX1    g21380(.A(new_n12256_), .Y(new_n23817_));
  OAI22X1  g21381(.A0(new_n23817_), .A1(new_n12109_), .B0(new_n12028_), .B1(new_n5027_), .Y(new_n23818_));
  AOI21X1  g21382(.A0(new_n23816_), .A1(new_n5027_), .B0(new_n23818_), .Y(new_n23819_));
  OAI21X1  g21383(.A0(new_n12171_), .A1(new_n12107_), .B0(new_n23816_), .Y(new_n23820_));
  INVX1    g21384(.A(new_n23820_), .Y(new_n23821_));
  OAI21X1  g21385(.A0(new_n23821_), .A1(new_n11968_), .B0(new_n12323_), .Y(new_n23822_));
  AOI21X1  g21386(.A0(new_n23819_), .A1(new_n11968_), .B0(new_n23822_), .Y(new_n23823_));
  NOR2X1   g21387(.A(new_n23820_), .B(new_n12326_), .Y(new_n23824_));
  INVX1    g21388(.A(new_n12360_), .Y(new_n23825_));
  NOR2X1   g21389(.A(new_n23816_), .B(new_n23825_), .Y(new_n23826_));
  OAI21X1  g21390(.A0(new_n23826_), .A1(new_n11950_), .B0(pi0680), .Y(new_n23827_));
  OR2X1    g21391(.A(new_n23827_), .B(new_n23824_), .Y(new_n23828_));
  OAI21X1  g21392(.A0(new_n23828_), .A1(new_n23823_), .B0(pi0661), .Y(new_n23829_));
  AOI21X1  g21393(.A0(new_n23815_), .A1(new_n5029_), .B0(new_n23829_), .Y(new_n23830_));
  AND2X1   g21394(.A(pi0681), .B(new_n11976_), .Y(new_n23831_));
  INVX1    g21395(.A(new_n23831_), .Y(new_n23832_));
  OAI21X1  g21396(.A0(new_n23832_), .A1(new_n23815_), .B0(new_n23633_), .Y(new_n23833_));
  NOR2X1   g21397(.A(new_n23833_), .B(new_n23830_), .Y(new_n23834_));
  NOR2X1   g21398(.A(new_n23834_), .B(new_n5070_), .Y(new_n23835_));
  OAI21X1  g21399(.A0(new_n12408_), .A1(new_n11950_), .B0(pi0680), .Y(new_n23836_));
  OAI21X1  g21400(.A0(new_n23836_), .A1(new_n12279_), .B0(pi0661), .Y(new_n23837_));
  AOI21X1  g21401(.A0(new_n23638_), .A1(new_n5029_), .B0(new_n23837_), .Y(new_n23838_));
  OAI21X1  g21402(.A0(new_n23832_), .A1(new_n23638_), .B0(new_n23642_), .Y(new_n23839_));
  OAI21X1  g21403(.A0(new_n23839_), .A1(new_n23838_), .B0(new_n5070_), .Y(new_n23840_));
  NAND2X1  g21404(.A(new_n23840_), .B(pi0222), .Y(new_n23841_));
  NOR2X1   g21405(.A(new_n12304_), .B(new_n12301_), .Y(new_n23842_));
  OAI21X1  g21406(.A0(new_n12354_), .A1(new_n11950_), .B0(pi0680), .Y(new_n23843_));
  AOI21X1  g21407(.A0(new_n23651_), .A1(new_n5029_), .B0(new_n11976_), .Y(new_n23844_));
  OAI21X1  g21408(.A0(new_n23843_), .A1(new_n23842_), .B0(new_n23844_), .Y(new_n23845_));
  AOI21X1  g21409(.A0(new_n23831_), .A1(new_n23652_), .B0(new_n23656_), .Y(new_n23846_));
  NAND3X1  g21410(.A(new_n23846_), .B(new_n23845_), .C(new_n5071_), .Y(new_n23847_));
  NOR2X1   g21411(.A(new_n12361_), .B(new_n11950_), .Y(new_n23848_));
  AND2X1   g21412(.A(new_n12316_), .B(pi0680), .Y(new_n23849_));
  INVX1    g21413(.A(new_n23849_), .Y(new_n23850_));
  AOI21X1  g21414(.A0(new_n23661_), .A1(new_n5029_), .B0(new_n11976_), .Y(new_n23851_));
  OAI21X1  g21415(.A0(new_n23850_), .A1(new_n23848_), .B0(new_n23851_), .Y(new_n23852_));
  NOR4X1   g21416(.A(new_n12171_), .B(new_n12047_), .C(new_n11983_), .D(new_n11950_), .Y(new_n23853_));
  AND2X1   g21417(.A(new_n23661_), .B(new_n11983_), .Y(new_n23854_));
  NOR3X1   g21418(.A(new_n23854_), .B(new_n23853_), .C(new_n23628_), .Y(new_n23855_));
  AOI21X1  g21419(.A0(new_n23831_), .A1(new_n23662_), .B0(new_n23855_), .Y(new_n23856_));
  NAND3X1  g21420(.A(new_n23856_), .B(new_n23852_), .C(new_n5070_), .Y(new_n23857_));
  NAND3X1  g21421(.A(new_n23857_), .B(new_n23847_), .C(new_n2960_), .Y(new_n23858_));
  OAI21X1  g21422(.A0(new_n23841_), .A1(new_n23835_), .B0(new_n23858_), .Y(new_n23859_));
  NOR2X1   g21423(.A(new_n23739_), .B(new_n23630_), .Y(new_n23860_));
  MX2X1    g21424(.A(new_n12361_), .B(new_n12308_), .S0(new_n11950_), .Y(new_n23861_));
  INVX1    g21425(.A(new_n23861_), .Y(new_n23862_));
  OAI21X1  g21426(.A0(new_n23862_), .A1(new_n23860_), .B0(new_n23663_), .Y(new_n23863_));
  AND2X1   g21427(.A(new_n23863_), .B(new_n2954_), .Y(new_n23864_));
  INVX1    g21428(.A(new_n23864_), .Y(new_n23865_));
  AOI21X1  g21429(.A0(new_n23859_), .A1(new_n10137_), .B0(new_n23865_), .Y(new_n23866_));
  AOI21X1  g21430(.A0(new_n23679_), .A1(new_n5029_), .B0(new_n11976_), .Y(new_n23867_));
  OAI21X1  g21431(.A0(new_n23836_), .A1(new_n12227_), .B0(new_n23867_), .Y(new_n23868_));
  AOI21X1  g21432(.A0(new_n23831_), .A1(new_n23680_), .B0(new_n23683_), .Y(new_n23869_));
  AND2X1   g21433(.A(new_n23869_), .B(new_n23868_), .Y(new_n23870_));
  NOR2X1   g21434(.A(new_n23825_), .B(new_n12237_), .Y(new_n23871_));
  OAI21X1  g21435(.A0(new_n23871_), .A1(new_n11950_), .B0(pi0680), .Y(new_n23872_));
  INVX1    g21436(.A(new_n23872_), .Y(new_n23873_));
  AOI21X1  g21437(.A0(new_n23873_), .A1(new_n12239_), .B0(new_n11976_), .Y(new_n23874_));
  OAI21X1  g21438(.A0(new_n23672_), .A1(pi0680), .B0(new_n23874_), .Y(new_n23875_));
  AOI21X1  g21439(.A0(new_n23831_), .A1(new_n23672_), .B0(new_n23675_), .Y(new_n23876_));
  AND2X1   g21440(.A(new_n23876_), .B(new_n23875_), .Y(new_n23877_));
  INVX1    g21441(.A(new_n23877_), .Y(new_n23878_));
  AOI21X1  g21442(.A0(new_n23878_), .A1(new_n5071_), .B0(new_n2960_), .Y(new_n23879_));
  OAI21X1  g21443(.A0(new_n23870_), .A1(new_n5071_), .B0(new_n23879_), .Y(new_n23880_));
  AOI21X1  g21444(.A0(new_n12376_), .A1(new_n12181_), .B0(new_n11966_), .Y(new_n23881_));
  OAI21X1  g21445(.A0(new_n23881_), .A1(new_n11950_), .B0(pi0680), .Y(new_n23882_));
  OR2X1    g21446(.A(new_n23882_), .B(new_n12329_), .Y(new_n23883_));
  NOR3X1   g21447(.A(new_n12181_), .B(new_n11966_), .C(new_n11950_), .Y(new_n23884_));
  AOI21X1  g21448(.A0(new_n23884_), .A1(new_n5029_), .B0(new_n11976_), .Y(new_n23885_));
  OAI21X1  g21449(.A0(new_n23662_), .A1(new_n11965_), .B0(new_n5030_), .Y(new_n23886_));
  OAI21X1  g21450(.A0(new_n23884_), .A1(pi0661), .B0(new_n23886_), .Y(new_n23887_));
  AOI21X1  g21451(.A0(new_n23885_), .A1(new_n23883_), .B0(new_n23887_), .Y(new_n23888_));
  OR4X1    g21452(.A(new_n12210_), .B(new_n12141_), .C(new_n5029_), .D(new_n11976_), .Y(new_n23889_));
  AND2X1   g21453(.A(new_n23889_), .B(new_n23668_), .Y(new_n23890_));
  OAI21X1  g21454(.A0(new_n23890_), .A1(new_n5071_), .B0(new_n2960_), .Y(new_n23891_));
  AOI21X1  g21455(.A0(new_n23888_), .A1(new_n5071_), .B0(new_n23891_), .Y(new_n23892_));
  NOR2X1   g21456(.A(new_n23892_), .B(new_n2954_), .Y(new_n23893_));
  AOI21X1  g21457(.A0(new_n23893_), .A1(new_n23880_), .B0(new_n2953_), .Y(new_n23894_));
  INVX1    g21458(.A(new_n23894_), .Y(new_n23895_));
  INVX1    g21459(.A(new_n3163_), .Y(new_n23896_));
  AOI21X1  g21460(.A0(new_n23744_), .A1(new_n23662_), .B0(pi0222), .Y(new_n23897_));
  OAI21X1  g21461(.A0(new_n23861_), .A1(new_n23744_), .B0(new_n23897_), .Y(new_n23898_));
  NAND3X1  g21462(.A(new_n23846_), .B(new_n23845_), .C(new_n5051_), .Y(new_n23899_));
  NAND3X1  g21463(.A(new_n23856_), .B(new_n23852_), .C(new_n5050_), .Y(new_n23900_));
  AND2X1   g21464(.A(new_n23900_), .B(pi0224), .Y(new_n23901_));
  AOI22X1  g21465(.A0(new_n23901_), .A1(new_n23899_), .B0(new_n23898_), .B1(new_n23896_), .Y(new_n23902_));
  NOR3X1   g21466(.A(new_n23833_), .B(new_n23830_), .C(new_n5050_), .Y(new_n23903_));
  NOR3X1   g21467(.A(new_n23839_), .B(new_n23838_), .C(new_n5051_), .Y(new_n23904_));
  NOR3X1   g21468(.A(new_n23904_), .B(new_n23903_), .C(new_n2960_), .Y(new_n23905_));
  OAI21X1  g21469(.A0(new_n23905_), .A1(new_n23902_), .B0(new_n2964_), .Y(new_n23906_));
  AOI21X1  g21470(.A0(new_n23878_), .A1(new_n5051_), .B0(new_n2960_), .Y(new_n23907_));
  OAI21X1  g21471(.A0(new_n23870_), .A1(new_n5051_), .B0(new_n23907_), .Y(new_n23908_));
  OAI21X1  g21472(.A0(new_n23890_), .A1(new_n5051_), .B0(new_n2960_), .Y(new_n23909_));
  AOI21X1  g21473(.A0(new_n23888_), .A1(new_n5051_), .B0(new_n23909_), .Y(new_n23910_));
  NOR2X1   g21474(.A(new_n23910_), .B(new_n2964_), .Y(new_n23911_));
  AOI21X1  g21475(.A0(new_n23911_), .A1(new_n23908_), .B0(pi0299), .Y(new_n23912_));
  AOI21X1  g21476(.A0(new_n23912_), .A1(new_n23906_), .B0(new_n2959_), .Y(new_n23913_));
  OAI21X1  g21477(.A0(new_n23895_), .A1(new_n23866_), .B0(new_n23913_), .Y(new_n23914_));
  NAND4X1  g21478(.A(new_n12461_), .B(new_n12459_), .C(pi0680), .D(pi0661), .Y(new_n23915_));
  AOI21X1  g21479(.A0(new_n12165_), .A1(pi0616), .B0(pi0222), .Y(new_n23916_));
  AND2X1   g21480(.A(new_n12461_), .B(new_n12459_), .Y(new_n23917_));
  INVX1    g21481(.A(new_n23917_), .Y(new_n23918_));
  AND2X1   g21482(.A(new_n12449_), .B(new_n5027_), .Y(new_n23919_));
  NAND2X1  g21483(.A(new_n12098_), .B(pi0603), .Y(new_n23920_));
  NAND2X1  g21484(.A(new_n23920_), .B(new_n23817_), .Y(new_n23921_));
  NOR2X1   g21485(.A(new_n23921_), .B(new_n23919_), .Y(new_n23922_));
  AOI21X1  g21486(.A0(new_n12165_), .A1(new_n11950_), .B0(new_n23922_), .Y(new_n23923_));
  OAI21X1  g21487(.A0(new_n23739_), .A1(new_n23918_), .B0(new_n23923_), .Y(new_n23924_));
  AOI22X1  g21488(.A0(new_n23924_), .A1(pi0222), .B0(new_n23916_), .B1(new_n23915_), .Y(new_n23925_));
  NOR2X1   g21489(.A(new_n23925_), .B(pi0299), .Y(new_n23926_));
  AND2X1   g21490(.A(new_n12465_), .B(new_n12464_), .Y(new_n23927_));
  INVX1    g21491(.A(new_n23927_), .Y(new_n23928_));
  AND2X1   g21492(.A(new_n12451_), .B(new_n5027_), .Y(new_n23929_));
  INVX1    g21493(.A(new_n12096_), .Y(new_n23930_));
  OAI21X1  g21494(.A0(new_n23930_), .A1(new_n5027_), .B0(new_n23817_), .Y(new_n23931_));
  NOR2X1   g21495(.A(new_n23931_), .B(new_n23929_), .Y(new_n23932_));
  AOI21X1  g21496(.A0(new_n12167_), .A1(new_n11950_), .B0(new_n23932_), .Y(new_n23933_));
  OAI21X1  g21497(.A0(new_n23739_), .A1(new_n23928_), .B0(new_n23933_), .Y(new_n23934_));
  NAND4X1  g21498(.A(new_n12465_), .B(new_n12464_), .C(pi0680), .D(pi0661), .Y(new_n23935_));
  AOI21X1  g21499(.A0(new_n12167_), .A1(pi0616), .B0(pi0222), .Y(new_n23936_));
  AOI22X1  g21500(.A0(new_n23936_), .A1(new_n23935_), .B0(new_n23934_), .B1(pi0222), .Y(new_n23937_));
  OAI21X1  g21501(.A0(new_n23937_), .A1(new_n2953_), .B0(new_n2959_), .Y(new_n23938_));
  OAI21X1  g21502(.A0(new_n23938_), .A1(new_n23926_), .B0(new_n2996_), .Y(new_n23939_));
  INVX1    g21503(.A(new_n23939_), .Y(new_n23940_));
  NOR4X1   g21504(.A(new_n23825_), .B(new_n3003_), .C(new_n2740_), .D(new_n2555_), .Y(new_n23941_));
  INVX1    g21505(.A(new_n23941_), .Y(new_n23942_));
  NOR4X1   g21506(.A(new_n5029_), .B(new_n11976_), .C(new_n11950_), .D(pi0039), .Y(new_n23943_));
  AOI21X1  g21507(.A0(new_n11950_), .A1(new_n2960_), .B0(new_n23943_), .Y(new_n23944_));
  AOI21X1  g21508(.A0(new_n12482_), .A1(new_n11950_), .B0(new_n23860_), .Y(new_n23945_));
  MX2X1    g21509(.A(pi0222), .B(new_n23945_), .S0(new_n12202_), .Y(new_n23946_));
  OAI21X1  g21510(.A0(new_n23944_), .A1(new_n23942_), .B0(new_n23946_), .Y(new_n23947_));
  AOI21X1  g21511(.A0(new_n23947_), .A1(pi0038), .B0(new_n3810_), .Y(new_n23948_));
  INVX1    g21512(.A(new_n23948_), .Y(new_n23949_));
  AOI21X1  g21513(.A0(new_n23940_), .A1(new_n23914_), .B0(new_n23949_), .Y(new_n23950_));
  AOI21X1  g21514(.A0(new_n3810_), .A1(pi0222), .B0(new_n23950_), .Y(new_n23951_));
  INVX1    g21515(.A(new_n23951_), .Y(new_n23952_));
  INVX1    g21516(.A(new_n23715_), .Y(new_n23953_));
  AOI21X1  g21517(.A0(new_n23953_), .A1(pi0625), .B0(pi1153), .Y(new_n23954_));
  OAI21X1  g21518(.A0(new_n23952_), .A1(pi0625), .B0(new_n23954_), .Y(new_n23955_));
  AND2X1   g21519(.A(new_n23800_), .B(new_n12584_), .Y(new_n23956_));
  AOI21X1  g21520(.A0(new_n23953_), .A1(new_n12493_), .B0(new_n12494_), .Y(new_n23957_));
  OAI21X1  g21521(.A0(new_n23952_), .A1(new_n12493_), .B0(new_n23957_), .Y(new_n23958_));
  AND2X1   g21522(.A(new_n23802_), .B(pi0608), .Y(new_n23959_));
  AOI22X1  g21523(.A0(new_n23959_), .A1(new_n23958_), .B0(new_n23956_), .B1(new_n23955_), .Y(new_n23960_));
  MX2X1    g21524(.A(new_n23960_), .B(new_n23952_), .S0(new_n11889_), .Y(new_n23961_));
  AOI21X1  g21525(.A0(new_n23804_), .A1(pi0609), .B0(pi1155), .Y(new_n23962_));
  OAI21X1  g21526(.A0(new_n23961_), .A1(pi0609), .B0(new_n23962_), .Y(new_n23963_));
  AND2X1   g21527(.A(new_n23719_), .B(new_n12596_), .Y(new_n23964_));
  AOI21X1  g21528(.A0(new_n23804_), .A1(new_n12590_), .B0(new_n12591_), .Y(new_n23965_));
  OAI21X1  g21529(.A0(new_n23961_), .A1(new_n12590_), .B0(new_n23965_), .Y(new_n23966_));
  AND2X1   g21530(.A(new_n23721_), .B(pi0660), .Y(new_n23967_));
  AOI22X1  g21531(.A0(new_n23967_), .A1(new_n23966_), .B0(new_n23964_), .B1(new_n23963_), .Y(new_n23968_));
  MX2X1    g21532(.A(new_n23968_), .B(new_n23961_), .S0(new_n11888_), .Y(new_n23969_));
  AOI21X1  g21533(.A0(new_n23805_), .A1(pi0618), .B0(pi1154), .Y(new_n23970_));
  OAI21X1  g21534(.A0(new_n23969_), .A1(pi0618), .B0(new_n23970_), .Y(new_n23971_));
  AND2X1   g21535(.A(new_n23725_), .B(new_n12622_), .Y(new_n23972_));
  AOI21X1  g21536(.A0(new_n23805_), .A1(new_n12614_), .B0(new_n12615_), .Y(new_n23973_));
  OAI21X1  g21537(.A0(new_n23969_), .A1(new_n12614_), .B0(new_n23973_), .Y(new_n23974_));
  AND2X1   g21538(.A(new_n23727_), .B(pi0627), .Y(new_n23975_));
  AOI22X1  g21539(.A0(new_n23975_), .A1(new_n23974_), .B0(new_n23972_), .B1(new_n23971_), .Y(new_n23976_));
  MX2X1    g21540(.A(new_n23976_), .B(new_n23969_), .S0(new_n11887_), .Y(new_n23977_));
  INVX1    g21541(.A(new_n23977_), .Y(new_n23978_));
  OAI21X1  g21542(.A0(new_n23807_), .A1(new_n12637_), .B0(new_n12638_), .Y(new_n23979_));
  AOI21X1  g21543(.A0(new_n23978_), .A1(new_n12637_), .B0(new_n23979_), .Y(new_n23980_));
  NOR3X1   g21544(.A(new_n23980_), .B(new_n23731_), .C(pi0648), .Y(new_n23981_));
  OAI21X1  g21545(.A0(new_n23807_), .A1(pi0619), .B0(pi1159), .Y(new_n23982_));
  AOI21X1  g21546(.A0(new_n23978_), .A1(pi0619), .B0(new_n23982_), .Y(new_n23983_));
  OR2X1    g21547(.A(new_n23733_), .B(new_n12645_), .Y(new_n23984_));
  OAI21X1  g21548(.A0(new_n23984_), .A1(new_n23983_), .B0(pi0789), .Y(new_n23985_));
  AOI21X1  g21549(.A0(new_n23717_), .A1(pi0626), .B0(new_n16352_), .Y(new_n23986_));
  OAI21X1  g21550(.A0(new_n23736_), .A1(pi0626), .B0(new_n23986_), .Y(new_n23987_));
  AOI21X1  g21551(.A0(new_n23717_), .A1(new_n12664_), .B0(new_n16356_), .Y(new_n23988_));
  OAI21X1  g21552(.A0(new_n23736_), .A1(new_n12664_), .B0(new_n23988_), .Y(new_n23989_));
  OAI21X1  g21553(.A0(new_n23627_), .A1(new_n22011_), .B0(new_n12769_), .Y(new_n23990_));
  NOR2X1   g21554(.A(new_n23990_), .B(new_n23808_), .Y(new_n23991_));
  INVX1    g21555(.A(new_n23991_), .Y(new_n23992_));
  NAND3X1  g21556(.A(new_n23992_), .B(new_n23989_), .C(new_n23987_), .Y(new_n23993_));
  AOI22X1  g21557(.A0(new_n23993_), .A1(pi0788), .B0(new_n23977_), .B1(new_n11886_), .Y(new_n23994_));
  OAI21X1  g21558(.A0(new_n23985_), .A1(new_n23981_), .B0(new_n23994_), .Y(new_n23995_));
  NAND4X1  g21559(.A(new_n23992_), .B(new_n23989_), .C(new_n23987_), .D(new_n14264_), .Y(new_n23996_));
  AND2X1   g21560(.A(new_n23996_), .B(new_n16350_), .Y(new_n23997_));
  AOI22X1  g21561(.A0(new_n23997_), .A1(new_n23995_), .B0(new_n23814_), .B1(pi0792), .Y(new_n23998_));
  MX2X1    g21562(.A(new_n23737_), .B(new_n23627_), .S0(new_n12711_), .Y(new_n23999_));
  OAI22X1  g21563(.A0(new_n23809_), .A1(new_n13639_), .B0(new_n23627_), .B1(new_n22842_), .Y(new_n24000_));
  OAI21X1  g21564(.A0(new_n23627_), .A1(pi0647), .B0(pi1157), .Y(new_n24001_));
  AOI21X1  g21565(.A0(new_n24000_), .A1(pi0647), .B0(new_n24001_), .Y(new_n24002_));
  OAI21X1  g21566(.A0(new_n23627_), .A1(new_n12705_), .B0(new_n12706_), .Y(new_n24003_));
  AOI21X1  g21567(.A0(new_n24000_), .A1(new_n12705_), .B0(new_n24003_), .Y(new_n24004_));
  MX2X1    g21568(.A(new_n24004_), .B(new_n24002_), .S0(new_n12723_), .Y(new_n24005_));
  AOI21X1  g21569(.A0(new_n23999_), .A1(new_n14385_), .B0(new_n24005_), .Y(new_n24006_));
  OAI22X1  g21570(.A0(new_n24006_), .A1(new_n11883_), .B0(new_n23998_), .B1(new_n14269_), .Y(new_n24007_));
  NOR2X1   g21571(.A(new_n24004_), .B(new_n24002_), .Y(new_n24008_));
  MX2X1    g21572(.A(new_n24008_), .B(new_n24000_), .S0(new_n11883_), .Y(new_n24009_));
  AOI21X1  g21573(.A0(new_n24009_), .A1(new_n12743_), .B0(new_n12739_), .Y(new_n24010_));
  OAI21X1  g21574(.A0(new_n24007_), .A1(new_n12743_), .B0(new_n24010_), .Y(new_n24011_));
  MX2X1    g21575(.A(new_n23999_), .B(new_n23627_), .S0(new_n12735_), .Y(new_n24012_));
  AOI21X1  g21576(.A0(new_n23717_), .A1(new_n12743_), .B0(pi0715), .Y(new_n24013_));
  OAI21X1  g21577(.A0(new_n24012_), .A1(new_n12743_), .B0(new_n24013_), .Y(new_n24014_));
  AND2X1   g21578(.A(new_n24014_), .B(pi1160), .Y(new_n24015_));
  AOI21X1  g21579(.A0(new_n24009_), .A1(pi0644), .B0(pi0715), .Y(new_n24016_));
  OAI21X1  g21580(.A0(new_n24007_), .A1(pi0644), .B0(new_n24016_), .Y(new_n24017_));
  AOI21X1  g21581(.A0(new_n23717_), .A1(pi0644), .B0(new_n12739_), .Y(new_n24018_));
  OAI21X1  g21582(.A0(new_n24012_), .A1(pi0644), .B0(new_n24018_), .Y(new_n24019_));
  AND2X1   g21583(.A(new_n24019_), .B(new_n11882_), .Y(new_n24020_));
  AOI22X1  g21584(.A0(new_n24020_), .A1(new_n24017_), .B0(new_n24015_), .B1(new_n24011_), .Y(new_n24021_));
  MX2X1    g21585(.A(new_n24021_), .B(new_n24007_), .S0(new_n12897_), .Y(new_n24022_));
  MX2X1    g21586(.A(new_n24022_), .B(pi0222), .S0(po1038), .Y(po0379));
  AOI21X1  g21587(.A0(new_n12010_), .A1(new_n2953_), .B0(new_n2959_), .Y(new_n24024_));
  AOI21X1  g21588(.A0(new_n11947_), .A1(new_n2959_), .B0(new_n10761_), .Y(new_n24025_));
  INVX1    g21589(.A(new_n24025_), .Y(new_n24026_));
  AOI21X1  g21590(.A0(new_n24024_), .A1(new_n12088_), .B0(new_n24026_), .Y(new_n24027_));
  OAI21X1  g21591(.A0(new_n24027_), .A1(new_n21881_), .B0(pi0223), .Y(new_n24028_));
  INVX1    g21592(.A(new_n24028_), .Y(new_n24029_));
  NOR3X1   g21593(.A(new_n12108_), .B(new_n11968_), .C(new_n5027_), .Y(new_n24030_));
  OR4X1    g21594(.A(new_n24030_), .B(new_n11952_), .C(new_n12323_), .D(new_n2740_), .Y(new_n24031_));
  AOI21X1  g21595(.A0(new_n12121_), .A1(pi0642), .B0(new_n12324_), .Y(new_n24032_));
  OAI21X1  g21596(.A0(new_n12030_), .A1(pi0642), .B0(new_n24032_), .Y(new_n24033_));
  AND2X1   g21597(.A(new_n24033_), .B(new_n24031_), .Y(new_n24034_));
  AND2X1   g21598(.A(new_n24034_), .B(pi0681), .Y(new_n24035_));
  AOI21X1  g21599(.A0(new_n24033_), .A1(new_n24031_), .B0(new_n12059_), .Y(new_n24036_));
  AOI21X1  g21600(.A0(new_n12029_), .A1(new_n11968_), .B0(new_n12124_), .Y(new_n24037_));
  OAI21X1  g21601(.A0(new_n24037_), .A1(new_n12060_), .B0(new_n11949_), .Y(new_n24038_));
  OAI21X1  g21602(.A0(new_n24038_), .A1(new_n24036_), .B0(new_n5070_), .Y(new_n24039_));
  OR2X1    g21603(.A(new_n24039_), .B(new_n24035_), .Y(new_n24040_));
  MX2X1    g21604(.A(new_n12291_), .B(new_n12260_), .S0(new_n11968_), .Y(new_n24041_));
  AND2X1   g21605(.A(new_n24041_), .B(pi0681), .Y(new_n24042_));
  INVX1    g21606(.A(new_n24042_), .Y(new_n24043_));
  NOR3X1   g21607(.A(new_n24030_), .B(new_n12046_), .C(new_n12060_), .Y(new_n24044_));
  NOR2X1   g21608(.A(new_n24044_), .B(pi0681), .Y(new_n24045_));
  OAI21X1  g21609(.A0(new_n24041_), .A1(new_n12059_), .B0(new_n24045_), .Y(new_n24046_));
  AND2X1   g21610(.A(new_n24046_), .B(new_n5071_), .Y(new_n24047_));
  AOI21X1  g21611(.A0(new_n24047_), .A1(new_n24043_), .B0(new_n2964_), .Y(new_n24048_));
  NOR4X1   g21612(.A(new_n12171_), .B(new_n11952_), .C(new_n2740_), .D(new_n11968_), .Y(new_n24049_));
  INVX1    g21613(.A(new_n24049_), .Y(new_n24050_));
  AOI21X1  g21614(.A0(new_n24049_), .A1(new_n12060_), .B0(pi0681), .Y(new_n24051_));
  INVX1    g21615(.A(new_n24051_), .Y(new_n24052_));
  NOR4X1   g21616(.A(new_n5029_), .B(pi0662), .C(pi0661), .D(new_n11968_), .Y(new_n24053_));
  AOI21X1  g21617(.A0(new_n24053_), .A1(new_n12170_), .B0(new_n24052_), .Y(new_n24054_));
  AOI21X1  g21618(.A0(new_n24050_), .A1(pi0681), .B0(new_n24054_), .Y(new_n24055_));
  AND2X1   g21619(.A(new_n24030_), .B(new_n12056_), .Y(new_n24056_));
  INVX1    g21620(.A(new_n24056_), .Y(new_n24057_));
  AOI21X1  g21621(.A0(new_n24053_), .A1(new_n12352_), .B0(pi0681), .Y(new_n24058_));
  OAI21X1  g21622(.A0(new_n24057_), .A1(new_n12059_), .B0(new_n24058_), .Y(new_n24059_));
  OAI21X1  g21623(.A0(new_n24056_), .A1(new_n11949_), .B0(new_n24059_), .Y(new_n24060_));
  OAI21X1  g21624(.A0(new_n24060_), .A1(new_n14594_), .B0(new_n14590_), .Y(new_n24061_));
  AOI21X1  g21625(.A0(new_n24055_), .A1(new_n14594_), .B0(new_n24061_), .Y(new_n24062_));
  AND2X1   g21626(.A(new_n24060_), .B(pi0947), .Y(new_n24063_));
  OR2X1    g21627(.A(new_n24063_), .B(pi0223), .Y(new_n24064_));
  OAI21X1  g21628(.A0(new_n24064_), .A1(new_n24062_), .B0(new_n10137_), .Y(new_n24065_));
  AOI21X1  g21629(.A0(new_n24048_), .A1(new_n24040_), .B0(new_n24065_), .Y(new_n24066_));
  AOI21X1  g21630(.A0(new_n11953_), .A1(pi0223), .B0(new_n10137_), .Y(new_n24067_));
  INVX1    g21631(.A(new_n24067_), .Y(new_n24068_));
  OAI21X1  g21632(.A0(new_n24068_), .A1(new_n24049_), .B0(new_n2954_), .Y(new_n24069_));
  INVX1    g21633(.A(new_n14594_), .Y(new_n24070_));
  AOI21X1  g21634(.A0(new_n24053_), .A1(new_n12182_), .B0(new_n24052_), .Y(new_n24071_));
  AOI21X1  g21635(.A0(new_n23670_), .A1(pi0642), .B0(new_n12060_), .Y(new_n24072_));
  AOI21X1  g21636(.A0(new_n24072_), .A1(new_n12144_), .B0(pi0681), .Y(new_n24073_));
  AOI21X1  g21637(.A0(new_n24073_), .A1(new_n11966_), .B0(new_n24071_), .Y(new_n24074_));
  INVX1    g21638(.A(new_n21936_), .Y(new_n24075_));
  OAI21X1  g21639(.A0(new_n24075_), .A1(new_n11968_), .B0(pi0681), .Y(new_n24076_));
  AND2X1   g21640(.A(new_n24076_), .B(new_n24074_), .Y(new_n24077_));
  OR2X1    g21641(.A(new_n24071_), .B(new_n5071_), .Y(new_n24078_));
  OAI21X1  g21642(.A0(new_n24078_), .A1(new_n24050_), .B0(new_n14590_), .Y(new_n24079_));
  AOI21X1  g21643(.A0(new_n24077_), .A1(new_n24070_), .B0(new_n24079_), .Y(new_n24080_));
  OAI21X1  g21644(.A0(new_n24077_), .A1(new_n14590_), .B0(new_n2964_), .Y(new_n24081_));
  AND2X1   g21645(.A(new_n12121_), .B(pi0642), .Y(new_n24082_));
  OAI21X1  g21646(.A0(new_n24082_), .A1(new_n23680_), .B0(new_n24031_), .Y(new_n24083_));
  INVX1    g21647(.A(new_n24083_), .Y(new_n24084_));
  NOR4X1   g21648(.A(new_n24030_), .B(new_n3003_), .C(new_n2740_), .D(new_n2555_), .Y(new_n24085_));
  INVX1    g21649(.A(new_n24085_), .Y(new_n24086_));
  NOR4X1   g21650(.A(new_n24086_), .B(new_n11971_), .C(new_n11970_), .D(new_n12060_), .Y(new_n24087_));
  NOR2X1   g21651(.A(new_n24087_), .B(pi0681), .Y(new_n24088_));
  OAI21X1  g21652(.A0(new_n24084_), .A1(new_n12059_), .B0(new_n24088_), .Y(new_n24089_));
  OAI21X1  g21653(.A0(new_n24083_), .A1(new_n11949_), .B0(new_n24089_), .Y(new_n24090_));
  NOR2X1   g21654(.A(new_n24090_), .B(new_n5071_), .Y(new_n24091_));
  MX2X1    g21655(.A(new_n12147_), .B(new_n11974_), .S0(new_n11968_), .Y(new_n24092_));
  INVX1    g21656(.A(new_n24092_), .Y(new_n24093_));
  OAI21X1  g21657(.A0(new_n24093_), .A1(new_n12059_), .B0(new_n24073_), .Y(new_n24094_));
  INVX1    g21658(.A(new_n24094_), .Y(new_n24095_));
  AOI21X1  g21659(.A0(new_n24093_), .A1(pi0681), .B0(new_n24095_), .Y(new_n24096_));
  AND2X1   g21660(.A(new_n24096_), .B(new_n5071_), .Y(new_n24097_));
  OR2X1    g21661(.A(new_n24097_), .B(new_n2964_), .Y(new_n24098_));
  OAI22X1  g21662(.A0(new_n24098_), .A1(new_n24091_), .B0(new_n24081_), .B1(new_n24080_), .Y(new_n24099_));
  AOI21X1  g21663(.A0(new_n24099_), .A1(pi0215), .B0(new_n2953_), .Y(new_n24100_));
  OAI21X1  g21664(.A0(new_n24069_), .A1(new_n24066_), .B0(new_n24100_), .Y(new_n24101_));
  AND2X1   g21665(.A(new_n24055_), .B(new_n5050_), .Y(new_n24102_));
  OAI21X1  g21666(.A0(new_n24060_), .A1(new_n5050_), .B0(new_n2971_), .Y(new_n24103_));
  AOI21X1  g21667(.A0(new_n24050_), .A1(new_n2970_), .B0(pi0223), .Y(new_n24104_));
  OAI21X1  g21668(.A0(new_n24103_), .A1(new_n24102_), .B0(new_n24104_), .Y(new_n24105_));
  AOI21X1  g21669(.A0(new_n24096_), .A1(new_n5051_), .B0(new_n2964_), .Y(new_n24106_));
  OAI21X1  g21670(.A0(new_n24090_), .A1(new_n5051_), .B0(new_n24106_), .Y(new_n24107_));
  NAND3X1  g21671(.A(new_n24107_), .B(new_n24105_), .C(new_n2953_), .Y(new_n24108_));
  AND2X1   g21672(.A(new_n24108_), .B(pi0039), .Y(new_n24109_));
  AND2X1   g21673(.A(pi0642), .B(new_n2964_), .Y(new_n24110_));
  AOI21X1  g21674(.A0(new_n24110_), .A1(new_n12165_), .B0(pi0299), .Y(new_n24111_));
  INVX1    g21675(.A(new_n12103_), .Y(new_n24112_));
  AOI21X1  g21676(.A0(new_n12165_), .A1(new_n11968_), .B0(new_n2964_), .Y(new_n24113_));
  NAND2X1  g21677(.A(new_n24113_), .B(new_n24112_), .Y(new_n24114_));
  AND2X1   g21678(.A(new_n24114_), .B(new_n24111_), .Y(new_n24115_));
  NAND3X1  g21679(.A(new_n24110_), .B(new_n12166_), .C(pi0603), .Y(new_n24116_));
  AND2X1   g21680(.A(new_n24116_), .B(pi0299), .Y(new_n24117_));
  INVX1    g21681(.A(new_n24117_), .Y(new_n24118_));
  AND2X1   g21682(.A(new_n12166_), .B(new_n11969_), .Y(new_n24119_));
  NOR3X1   g21683(.A(new_n24119_), .B(new_n12097_), .C(new_n2964_), .Y(new_n24120_));
  OAI21X1  g21684(.A0(new_n24120_), .A1(new_n24118_), .B0(new_n2959_), .Y(new_n24121_));
  OAI21X1  g21685(.A0(new_n24121_), .A1(new_n24115_), .B0(new_n2996_), .Y(new_n24122_));
  AOI21X1  g21686(.A0(new_n24109_), .A1(new_n24101_), .B0(new_n24122_), .Y(new_n24123_));
  AOI21X1  g21687(.A0(pi0223), .A1(pi0039), .B0(new_n2996_), .Y(new_n24124_));
  INVX1    g21688(.A(new_n24124_), .Y(new_n24125_));
  AOI21X1  g21689(.A0(new_n12416_), .A1(new_n2964_), .B0(pi0039), .Y(new_n24126_));
  AOI21X1  g21690(.A0(new_n24126_), .A1(new_n24086_), .B0(new_n24125_), .Y(new_n24127_));
  OR2X1    g21691(.A(new_n24127_), .B(new_n3810_), .Y(new_n24128_));
  OAI22X1  g21692(.A0(new_n24128_), .A1(new_n24123_), .B0(new_n3129_), .B1(new_n2964_), .Y(new_n24129_));
  MX2X1    g21693(.A(new_n24129_), .B(new_n24029_), .S0(new_n12601_), .Y(new_n24130_));
  AOI21X1  g21694(.A0(new_n24028_), .A1(new_n12590_), .B0(new_n12591_), .Y(new_n24131_));
  OAI21X1  g21695(.A0(new_n24130_), .A1(new_n12590_), .B0(new_n24131_), .Y(new_n24132_));
  AOI21X1  g21696(.A0(new_n24028_), .A1(pi0609), .B0(pi1155), .Y(new_n24133_));
  OAI21X1  g21697(.A0(new_n24130_), .A1(pi0609), .B0(new_n24133_), .Y(new_n24134_));
  AOI21X1  g21698(.A0(new_n24134_), .A1(new_n24132_), .B0(new_n11888_), .Y(new_n24135_));
  AOI21X1  g21699(.A0(new_n24130_), .A1(new_n11888_), .B0(new_n24135_), .Y(new_n24136_));
  NAND2X1  g21700(.A(new_n24136_), .B(pi0618), .Y(new_n24137_));
  AOI21X1  g21701(.A0(new_n24028_), .A1(new_n12614_), .B0(new_n12615_), .Y(new_n24138_));
  NAND2X1  g21702(.A(new_n24136_), .B(new_n12614_), .Y(new_n24139_));
  AOI21X1  g21703(.A0(new_n24028_), .A1(pi0618), .B0(pi1154), .Y(new_n24140_));
  AOI22X1  g21704(.A0(new_n24140_), .A1(new_n24139_), .B0(new_n24138_), .B1(new_n24137_), .Y(new_n24141_));
  MX2X1    g21705(.A(new_n24141_), .B(new_n24136_), .S0(new_n11887_), .Y(new_n24142_));
  OAI21X1  g21706(.A0(new_n24029_), .A1(pi0619), .B0(pi1159), .Y(new_n24143_));
  AOI21X1  g21707(.A0(new_n24142_), .A1(pi0619), .B0(new_n24143_), .Y(new_n24144_));
  OAI21X1  g21708(.A0(new_n24029_), .A1(new_n12637_), .B0(new_n12638_), .Y(new_n24145_));
  AOI21X1  g21709(.A0(new_n24142_), .A1(new_n12637_), .B0(new_n24145_), .Y(new_n24146_));
  OAI21X1  g21710(.A0(new_n24146_), .A1(new_n24144_), .B0(pi0789), .Y(new_n24147_));
  OAI21X1  g21711(.A0(new_n24142_), .A1(pi0789), .B0(new_n24147_), .Y(new_n24148_));
  MX2X1    g21712(.A(new_n24148_), .B(new_n24029_), .S0(new_n12841_), .Y(new_n24149_));
  MX2X1    g21713(.A(new_n24149_), .B(new_n24029_), .S0(new_n12711_), .Y(new_n24150_));
  AND2X1   g21714(.A(pi0681), .B(pi0680), .Y(new_n24151_));
  NOR2X1   g21715(.A(new_n24151_), .B(new_n12458_), .Y(new_n24152_));
  AND2X1   g21716(.A(new_n12458_), .B(new_n2964_), .Y(new_n24153_));
  OAI21X1  g21717(.A0(new_n12449_), .A1(new_n2964_), .B0(new_n2953_), .Y(new_n24154_));
  NOR3X1   g21718(.A(new_n24154_), .B(new_n24153_), .C(new_n24152_), .Y(new_n24155_));
  INVX1    g21719(.A(new_n24151_), .Y(new_n24156_));
  AND2X1   g21720(.A(new_n24156_), .B(new_n12463_), .Y(new_n24157_));
  NOR2X1   g21721(.A(new_n12463_), .B(pi0223), .Y(new_n24158_));
  OAI21X1  g21722(.A0(new_n12451_), .A1(new_n2964_), .B0(pi0299), .Y(new_n24159_));
  NOR3X1   g21723(.A(new_n24159_), .B(new_n24158_), .C(new_n24157_), .Y(new_n24160_));
  NOR3X1   g21724(.A(new_n24160_), .B(new_n24155_), .C(pi0039), .Y(new_n24161_));
  NOR4X1   g21725(.A(new_n12499_), .B(new_n11952_), .C(new_n2740_), .D(new_n11949_), .Y(new_n24162_));
  NOR2X1   g21726(.A(new_n24162_), .B(new_n24068_), .Y(new_n24163_));
  AND2X1   g21727(.A(new_n12072_), .B(new_n5070_), .Y(new_n24164_));
  OAI21X1  g21728(.A0(new_n12528_), .A1(new_n11949_), .B0(new_n24164_), .Y(new_n24165_));
  NOR2X1   g21729(.A(new_n23756_), .B(new_n11949_), .Y(new_n24166_));
  NOR3X1   g21730(.A(new_n24166_), .B(new_n12062_), .C(new_n5070_), .Y(new_n24167_));
  NOR2X1   g21731(.A(new_n24167_), .B(new_n2964_), .Y(new_n24168_));
  NAND3X1  g21732(.A(new_n12341_), .B(new_n12057_), .C(pi0681), .Y(new_n24169_));
  AND2X1   g21733(.A(new_n24169_), .B(new_n5071_), .Y(new_n24170_));
  NOR2X1   g21734(.A(new_n24156_), .B(new_n12502_), .Y(new_n24171_));
  OAI21X1  g21735(.A0(new_n24171_), .A1(new_n5071_), .B0(new_n2964_), .Y(new_n24172_));
  OAI21X1  g21736(.A0(new_n24172_), .A1(new_n24170_), .B0(new_n10137_), .Y(new_n24173_));
  AOI21X1  g21737(.A0(new_n24168_), .A1(new_n24165_), .B0(new_n24173_), .Y(new_n24174_));
  OAI21X1  g21738(.A0(new_n24174_), .A1(new_n24163_), .B0(new_n2954_), .Y(new_n24175_));
  AOI21X1  g21739(.A0(new_n12545_), .A1(pi0681), .B0(new_n11990_), .Y(new_n24176_));
  NAND2X1  g21740(.A(new_n24176_), .B(new_n5071_), .Y(new_n24177_));
  AOI21X1  g21741(.A0(new_n23767_), .A1(pi0681), .B0(new_n12008_), .Y(new_n24178_));
  AOI21X1  g21742(.A0(new_n24178_), .A1(new_n5070_), .B0(new_n2964_), .Y(new_n24179_));
  AND2X1   g21743(.A(pi0681), .B(new_n2964_), .Y(new_n24180_));
  AOI21X1  g21744(.A0(new_n24180_), .A1(new_n12518_), .B0(new_n2954_), .Y(new_n24181_));
  INVX1    g21745(.A(new_n24181_), .Y(new_n24182_));
  AOI21X1  g21746(.A0(new_n24179_), .A1(new_n24177_), .B0(new_n24182_), .Y(new_n24183_));
  NOR2X1   g21747(.A(new_n24183_), .B(new_n2953_), .Y(new_n24184_));
  NOR3X1   g21748(.A(new_n24156_), .B(new_n12502_), .C(new_n5051_), .Y(new_n24185_));
  OAI21X1  g21749(.A0(new_n24169_), .A1(new_n5050_), .B0(new_n2971_), .Y(new_n24186_));
  OAI22X1  g21750(.A0(new_n24186_), .A1(new_n24185_), .B0(new_n24162_), .B1(new_n2971_), .Y(new_n24187_));
  AND2X1   g21751(.A(new_n24187_), .B(new_n2964_), .Y(new_n24188_));
  NOR2X1   g21752(.A(new_n24176_), .B(new_n5050_), .Y(new_n24189_));
  OAI21X1  g21753(.A0(new_n24178_), .A1(new_n5051_), .B0(pi0223), .Y(new_n24190_));
  OAI21X1  g21754(.A0(new_n24190_), .A1(new_n24189_), .B0(new_n2953_), .Y(new_n24191_));
  OAI21X1  g21755(.A0(new_n24191_), .A1(new_n24188_), .B0(pi0039), .Y(new_n24192_));
  AOI21X1  g21756(.A0(new_n24184_), .A1(new_n24175_), .B0(new_n24192_), .Y(new_n24193_));
  OAI21X1  g21757(.A0(new_n24193_), .A1(new_n24161_), .B0(new_n2996_), .Y(new_n24194_));
  NOR4X1   g21758(.A(new_n13585_), .B(new_n3074_), .C(new_n11949_), .D(pi0039), .Y(new_n24195_));
  INVX1    g21759(.A(new_n24195_), .Y(new_n24196_));
  AOI21X1  g21760(.A0(new_n12901_), .A1(pi0223), .B0(new_n2996_), .Y(new_n24197_));
  AOI21X1  g21761(.A0(new_n24197_), .A1(new_n24196_), .B0(new_n3810_), .Y(new_n24198_));
  AOI22X1  g21762(.A0(new_n24198_), .A1(new_n24194_), .B0(new_n3810_), .B1(pi0223), .Y(new_n24199_));
  INVX1    g21763(.A(new_n24199_), .Y(new_n24200_));
  AOI21X1  g21764(.A0(new_n24028_), .A1(new_n12493_), .B0(new_n12494_), .Y(new_n24201_));
  OAI21X1  g21765(.A0(new_n24200_), .A1(new_n12493_), .B0(new_n24201_), .Y(new_n24202_));
  AOI21X1  g21766(.A0(new_n24028_), .A1(pi0625), .B0(pi1153), .Y(new_n24203_));
  OAI21X1  g21767(.A0(new_n24200_), .A1(pi0625), .B0(new_n24203_), .Y(new_n24204_));
  AND2X1   g21768(.A(new_n24204_), .B(new_n24202_), .Y(new_n24205_));
  MX2X1    g21769(.A(new_n24205_), .B(new_n24199_), .S0(new_n11889_), .Y(new_n24206_));
  MX2X1    g21770(.A(new_n24206_), .B(new_n24028_), .S0(new_n12618_), .Y(new_n24207_));
  MX2X1    g21771(.A(new_n24207_), .B(new_n24028_), .S0(new_n12641_), .Y(new_n24208_));
  AND2X1   g21772(.A(new_n24208_), .B(new_n22011_), .Y(new_n24209_));
  AOI22X1  g21773(.A0(new_n24209_), .A1(new_n17252_), .B0(new_n24028_), .B1(new_n22010_), .Y(new_n24210_));
  OAI22X1  g21774(.A0(new_n24210_), .A1(new_n13639_), .B0(new_n24029_), .B1(new_n22842_), .Y(new_n24211_));
  OAI21X1  g21775(.A0(new_n24029_), .A1(pi0647), .B0(pi1157), .Y(new_n24212_));
  AOI21X1  g21776(.A0(new_n24211_), .A1(pi0647), .B0(new_n24212_), .Y(new_n24213_));
  OAI21X1  g21777(.A0(new_n24029_), .A1(new_n12705_), .B0(new_n12706_), .Y(new_n24214_));
  AOI21X1  g21778(.A0(new_n24211_), .A1(new_n12705_), .B0(new_n24214_), .Y(new_n24215_));
  MX2X1    g21779(.A(new_n24215_), .B(new_n24213_), .S0(new_n12723_), .Y(new_n24216_));
  AOI21X1  g21780(.A0(new_n24150_), .A1(new_n14385_), .B0(new_n24216_), .Y(new_n24217_));
  NAND2X1  g21781(.A(new_n24149_), .B(new_n14394_), .Y(new_n24218_));
  AOI21X1  g21782(.A0(new_n24028_), .A1(pi0628), .B0(new_n12710_), .Y(new_n24219_));
  OAI21X1  g21783(.A0(new_n24210_), .A1(pi0628), .B0(new_n24219_), .Y(new_n24220_));
  AOI21X1  g21784(.A0(new_n24028_), .A1(new_n12683_), .B0(new_n12708_), .Y(new_n24221_));
  OAI21X1  g21785(.A0(new_n24210_), .A1(new_n12683_), .B0(new_n24221_), .Y(new_n24222_));
  NAND3X1  g21786(.A(new_n24222_), .B(new_n24220_), .C(new_n24218_), .Y(new_n24223_));
  OAI21X1  g21787(.A0(new_n24028_), .A1(pi0626), .B0(new_n16355_), .Y(new_n24224_));
  AOI21X1  g21788(.A0(new_n24148_), .A1(pi0626), .B0(new_n24224_), .Y(new_n24225_));
  AND2X1   g21789(.A(new_n24148_), .B(new_n12664_), .Y(new_n24226_));
  OAI21X1  g21790(.A0(new_n24028_), .A1(new_n12664_), .B0(new_n16351_), .Y(new_n24227_));
  AOI21X1  g21791(.A0(new_n24028_), .A1(new_n12659_), .B0(new_n24209_), .Y(new_n24228_));
  OAI22X1  g21792(.A0(new_n24228_), .A1(new_n12770_), .B0(new_n24227_), .B1(new_n24226_), .Y(new_n24229_));
  OAI21X1  g21793(.A0(new_n24229_), .A1(new_n24225_), .B0(pi0788), .Y(new_n24230_));
  INVX1    g21794(.A(new_n23390_), .Y(new_n24231_));
  OR2X1    g21795(.A(new_n12408_), .B(new_n11968_), .Y(new_n24232_));
  AOI21X1  g21796(.A0(new_n24232_), .A1(new_n12276_), .B0(new_n24231_), .Y(new_n24233_));
  NOR2X1   g21797(.A(new_n24233_), .B(new_n5029_), .Y(new_n24234_));
  INVX1    g21798(.A(new_n24234_), .Y(new_n24235_));
  OAI21X1  g21799(.A0(new_n12361_), .A1(new_n11968_), .B0(new_n12323_), .Y(new_n24236_));
  AOI21X1  g21800(.A0(new_n12314_), .A1(new_n11968_), .B0(new_n24236_), .Y(new_n24237_));
  OAI22X1  g21801(.A0(new_n24237_), .A1(new_n24235_), .B0(new_n24049_), .B1(pi0680), .Y(new_n24238_));
  AOI21X1  g21802(.A0(new_n24238_), .A1(pi0681), .B0(new_n24054_), .Y(new_n24239_));
  OAI21X1  g21803(.A0(new_n24057_), .A1(pi0680), .B0(pi0681), .Y(new_n24240_));
  NOR2X1   g21804(.A(new_n12323_), .B(pi0642), .Y(new_n24241_));
  AND2X1   g21805(.A(new_n24241_), .B(new_n12296_), .Y(new_n24242_));
  OAI21X1  g21806(.A0(new_n12354_), .A1(new_n11968_), .B0(pi0680), .Y(new_n24243_));
  NOR3X1   g21807(.A(new_n24243_), .B(new_n24242_), .C(new_n12300_), .Y(new_n24244_));
  OAI21X1  g21808(.A0(new_n24244_), .A1(new_n24240_), .B0(new_n24059_), .Y(new_n24245_));
  AOI21X1  g21809(.A0(new_n24245_), .A1(new_n5071_), .B0(pi0223), .Y(new_n24246_));
  OAI21X1  g21810(.A0(new_n24239_), .A1(new_n5071_), .B0(new_n24246_), .Y(new_n24247_));
  INVX1    g21811(.A(new_n24039_), .Y(new_n24248_));
  MX2X1    g21812(.A(new_n23825_), .B(new_n12211_), .S0(new_n11968_), .Y(new_n24249_));
  NOR4X1   g21813(.A(new_n24249_), .B(new_n3003_), .C(new_n2740_), .D(new_n2555_), .Y(new_n24250_));
  INVX1    g21814(.A(new_n24250_), .Y(new_n24251_));
  NOR2X1   g21815(.A(new_n24251_), .B(new_n12415_), .Y(new_n24252_));
  OAI21X1  g21816(.A0(new_n24252_), .A1(new_n12323_), .B0(pi0680), .Y(new_n24253_));
  AOI21X1  g21817(.A0(new_n24232_), .A1(new_n12247_), .B0(new_n12324_), .Y(new_n24254_));
  OAI22X1  g21818(.A0(new_n24254_), .A1(new_n24253_), .B0(new_n24151_), .B1(new_n24035_), .Y(new_n24255_));
  NAND2X1  g21819(.A(new_n24255_), .B(new_n24248_), .Y(new_n24256_));
  OAI21X1  g21820(.A0(new_n23826_), .A1(new_n11968_), .B0(pi0680), .Y(new_n24257_));
  AOI21X1  g21821(.A0(new_n24241_), .A1(new_n23821_), .B0(new_n24257_), .Y(new_n24258_));
  OAI21X1  g21822(.A0(new_n23819_), .A1(new_n12127_), .B0(new_n24258_), .Y(new_n24259_));
  OAI21X1  g21823(.A0(new_n24151_), .A1(new_n24042_), .B0(new_n24259_), .Y(new_n24260_));
  AOI21X1  g21824(.A0(new_n24260_), .A1(new_n24047_), .B0(new_n2964_), .Y(new_n24261_));
  AOI21X1  g21825(.A0(new_n24261_), .A1(new_n24256_), .B0(new_n10136_), .Y(new_n24262_));
  AOI21X1  g21826(.A0(new_n12276_), .A1(new_n11968_), .B0(new_n24156_), .Y(new_n24263_));
  AOI22X1  g21827(.A0(new_n24263_), .A1(new_n23942_), .B0(new_n24156_), .B1(new_n24030_), .Y(new_n24264_));
  NOR3X1   g21828(.A(new_n24264_), .B(new_n11953_), .C(pi0223), .Y(new_n24265_));
  OAI21X1  g21829(.A0(new_n24251_), .A1(new_n24156_), .B0(pi0223), .Y(new_n24266_));
  AOI21X1  g21830(.A0(new_n24156_), .A1(new_n24085_), .B0(new_n24266_), .Y(new_n24267_));
  NOR3X1   g21831(.A(new_n24267_), .B(new_n24265_), .C(new_n24068_), .Y(new_n24268_));
  OR2X1    g21832(.A(new_n24268_), .B(pi0215), .Y(new_n24269_));
  AOI21X1  g21833(.A0(new_n24262_), .A1(new_n24247_), .B0(new_n24269_), .Y(new_n24270_));
  OAI21X1  g21834(.A0(new_n24084_), .A1(pi0680), .B0(pi0681), .Y(new_n24271_));
  AOI22X1  g21835(.A0(new_n12409_), .A1(pi0642), .B0(new_n12225_), .B1(new_n12051_), .Y(new_n24272_));
  NOR2X1   g21836(.A(new_n24272_), .B(pi0616), .Y(new_n24273_));
  NOR2X1   g21837(.A(new_n24273_), .B(new_n24253_), .Y(new_n24274_));
  OAI21X1  g21838(.A0(new_n24274_), .A1(new_n24271_), .B0(new_n24089_), .Y(new_n24275_));
  NOR2X1   g21839(.A(new_n12238_), .B(new_n12323_), .Y(new_n24276_));
  NOR2X1   g21840(.A(new_n23871_), .B(new_n11968_), .Y(new_n24277_));
  OAI21X1  g21841(.A0(new_n12222_), .A1(new_n12127_), .B0(pi0680), .Y(new_n24278_));
  NOR3X1   g21842(.A(new_n24278_), .B(new_n24277_), .C(new_n24276_), .Y(new_n24279_));
  OR2X1    g21843(.A(new_n24279_), .B(new_n11949_), .Y(new_n24280_));
  AOI21X1  g21844(.A0(new_n24092_), .A1(new_n5029_), .B0(new_n24280_), .Y(new_n24281_));
  NOR2X1   g21845(.A(new_n24281_), .B(new_n24095_), .Y(new_n24282_));
  OAI21X1  g21846(.A0(new_n24282_), .A1(new_n5070_), .B0(pi0223), .Y(new_n24283_));
  AOI21X1  g21847(.A0(new_n24275_), .A1(new_n5070_), .B0(new_n24283_), .Y(new_n24284_));
  AOI21X1  g21848(.A0(new_n12327_), .A1(new_n11968_), .B0(new_n24236_), .Y(new_n24285_));
  OAI22X1  g21849(.A0(new_n24285_), .A1(new_n24235_), .B0(new_n24049_), .B1(pi0680), .Y(new_n24286_));
  AOI21X1  g21850(.A0(new_n24286_), .A1(pi0681), .B0(new_n24078_), .Y(new_n24287_));
  OAI21X1  g21851(.A0(new_n12385_), .A1(new_n12327_), .B0(new_n12125_), .Y(new_n24288_));
  OAI21X1  g21852(.A0(new_n23881_), .A1(new_n11968_), .B0(pi0680), .Y(new_n24289_));
  AOI21X1  g21853(.A0(new_n24241_), .A1(new_n12321_), .B0(new_n24289_), .Y(new_n24290_));
  AOI22X1  g21854(.A0(new_n24290_), .A1(new_n24288_), .B0(new_n24156_), .B1(new_n24076_), .Y(new_n24291_));
  NAND2X1  g21855(.A(new_n24074_), .B(new_n5071_), .Y(new_n24292_));
  OAI21X1  g21856(.A0(new_n24292_), .A1(new_n24291_), .B0(new_n2964_), .Y(new_n24293_));
  OAI21X1  g21857(.A0(new_n24293_), .A1(new_n24287_), .B0(pi0215), .Y(new_n24294_));
  OAI21X1  g21858(.A0(new_n24294_), .A1(new_n24284_), .B0(pi0299), .Y(new_n24295_));
  NOR2X1   g21859(.A(new_n24245_), .B(new_n5050_), .Y(new_n24296_));
  AND2X1   g21860(.A(new_n24239_), .B(new_n5050_), .Y(new_n24297_));
  OR2X1    g21861(.A(new_n24297_), .B(new_n2970_), .Y(new_n24298_));
  OAI21X1  g21862(.A0(new_n24264_), .A1(new_n11953_), .B0(new_n2970_), .Y(new_n24299_));
  AND2X1   g21863(.A(new_n24299_), .B(new_n2964_), .Y(new_n24300_));
  OAI21X1  g21864(.A0(new_n24298_), .A1(new_n24296_), .B0(new_n24300_), .Y(new_n24301_));
  AOI21X1  g21865(.A0(new_n24282_), .A1(new_n5051_), .B0(new_n2964_), .Y(new_n24302_));
  OAI21X1  g21866(.A0(new_n24275_), .A1(new_n5051_), .B0(new_n24302_), .Y(new_n24303_));
  NAND3X1  g21867(.A(new_n24303_), .B(new_n24301_), .C(new_n2953_), .Y(new_n24304_));
  AND2X1   g21868(.A(new_n24304_), .B(pi0039), .Y(new_n24305_));
  OAI21X1  g21869(.A0(new_n24295_), .A1(new_n24270_), .B0(new_n24305_), .Y(new_n24306_));
  INVX1    g21870(.A(new_n23922_), .Y(new_n24307_));
  NAND3X1  g21871(.A(new_n24156_), .B(new_n12461_), .C(new_n12459_), .Y(new_n24308_));
  NAND3X1  g21872(.A(new_n24308_), .B(new_n24113_), .C(new_n24307_), .Y(new_n24309_));
  NAND4X1  g21873(.A(new_n24180_), .B(new_n12461_), .C(new_n12459_), .D(pi0680), .Y(new_n24310_));
  NAND3X1  g21874(.A(new_n24310_), .B(new_n24309_), .C(new_n24111_), .Y(new_n24311_));
  NAND4X1  g21875(.A(new_n24180_), .B(new_n12465_), .C(new_n12464_), .D(pi0680), .Y(new_n24312_));
  AND2X1   g21876(.A(new_n24156_), .B(new_n23927_), .Y(new_n24313_));
  OR4X1    g21877(.A(new_n24313_), .B(new_n24119_), .C(new_n23932_), .D(new_n2964_), .Y(new_n24314_));
  NAND3X1  g21878(.A(new_n24314_), .B(new_n24312_), .C(new_n24117_), .Y(new_n24315_));
  NAND3X1  g21879(.A(new_n24315_), .B(new_n24311_), .C(new_n2959_), .Y(new_n24316_));
  NAND3X1  g21880(.A(new_n24316_), .B(new_n24306_), .C(new_n2996_), .Y(new_n24317_));
  INVX1    g21881(.A(new_n24264_), .Y(new_n24318_));
  OAI21X1  g21882(.A0(new_n24267_), .A1(new_n24318_), .B0(new_n24126_), .Y(new_n24319_));
  AOI21X1  g21883(.A0(new_n24319_), .A1(new_n24124_), .B0(new_n3810_), .Y(new_n24320_));
  AOI22X1  g21884(.A0(new_n24320_), .A1(new_n24317_), .B0(new_n3810_), .B1(pi0223), .Y(new_n24321_));
  INVX1    g21885(.A(new_n24202_), .Y(new_n24322_));
  INVX1    g21886(.A(new_n24204_), .Y(new_n24323_));
  AND2X1   g21887(.A(new_n24321_), .B(new_n12493_), .Y(new_n24324_));
  OAI21X1  g21888(.A0(new_n24129_), .A1(new_n12493_), .B0(new_n12494_), .Y(new_n24325_));
  OAI21X1  g21889(.A0(new_n24325_), .A1(new_n24324_), .B0(new_n12584_), .Y(new_n24326_));
  AND2X1   g21890(.A(new_n24321_), .B(pi0625), .Y(new_n24327_));
  OAI21X1  g21891(.A0(new_n24129_), .A1(pi0625), .B0(pi1153), .Y(new_n24328_));
  OAI21X1  g21892(.A0(new_n24328_), .A1(new_n24327_), .B0(pi0608), .Y(new_n24329_));
  OAI22X1  g21893(.A0(new_n24329_), .A1(new_n24323_), .B0(new_n24326_), .B1(new_n24322_), .Y(new_n24330_));
  MX2X1    g21894(.A(new_n24330_), .B(new_n24321_), .S0(new_n11889_), .Y(new_n24331_));
  NAND2X1  g21895(.A(new_n24331_), .B(new_n12590_), .Y(new_n24332_));
  AOI21X1  g21896(.A0(new_n24206_), .A1(pi0609), .B0(pi1155), .Y(new_n24333_));
  NAND2X1  g21897(.A(new_n24132_), .B(new_n12596_), .Y(new_n24334_));
  AOI21X1  g21898(.A0(new_n24333_), .A1(new_n24332_), .B0(new_n24334_), .Y(new_n24335_));
  NAND2X1  g21899(.A(new_n24331_), .B(pi0609), .Y(new_n24336_));
  AOI21X1  g21900(.A0(new_n24206_), .A1(new_n12590_), .B0(new_n12591_), .Y(new_n24337_));
  NAND2X1  g21901(.A(new_n24134_), .B(pi0660), .Y(new_n24338_));
  AOI21X1  g21902(.A0(new_n24337_), .A1(new_n24336_), .B0(new_n24338_), .Y(new_n24339_));
  OR2X1    g21903(.A(new_n24339_), .B(new_n24335_), .Y(new_n24340_));
  MX2X1    g21904(.A(new_n24340_), .B(new_n24331_), .S0(new_n11888_), .Y(new_n24341_));
  AND2X1   g21905(.A(new_n24341_), .B(new_n12614_), .Y(new_n24342_));
  INVX1    g21906(.A(new_n24207_), .Y(new_n24343_));
  OAI21X1  g21907(.A0(new_n24343_), .A1(new_n12614_), .B0(new_n12615_), .Y(new_n24344_));
  AOI21X1  g21908(.A0(new_n24138_), .A1(new_n24137_), .B0(pi0627), .Y(new_n24345_));
  OAI21X1  g21909(.A0(new_n24344_), .A1(new_n24342_), .B0(new_n24345_), .Y(new_n24346_));
  AND2X1   g21910(.A(new_n24341_), .B(pi0618), .Y(new_n24347_));
  OAI21X1  g21911(.A0(new_n24343_), .A1(pi0618), .B0(pi1154), .Y(new_n24348_));
  AOI21X1  g21912(.A0(new_n24140_), .A1(new_n24139_), .B0(new_n12622_), .Y(new_n24349_));
  OAI21X1  g21913(.A0(new_n24348_), .A1(new_n24347_), .B0(new_n24349_), .Y(new_n24350_));
  AOI21X1  g21914(.A0(new_n24350_), .A1(new_n24346_), .B0(new_n11887_), .Y(new_n24351_));
  AND2X1   g21915(.A(new_n24341_), .B(new_n11887_), .Y(new_n24352_));
  OAI21X1  g21916(.A0(new_n24352_), .A1(new_n24351_), .B0(new_n12637_), .Y(new_n24353_));
  AOI21X1  g21917(.A0(new_n24208_), .A1(pi0619), .B0(pi1159), .Y(new_n24354_));
  OR2X1    g21918(.A(new_n24144_), .B(pi0648), .Y(new_n24355_));
  AOI21X1  g21919(.A0(new_n24354_), .A1(new_n24353_), .B0(new_n24355_), .Y(new_n24356_));
  OAI21X1  g21920(.A0(new_n24352_), .A1(new_n24351_), .B0(pi0619), .Y(new_n24357_));
  AOI21X1  g21921(.A0(new_n24208_), .A1(new_n12637_), .B0(new_n12638_), .Y(new_n24358_));
  OR2X1    g21922(.A(new_n24146_), .B(new_n12645_), .Y(new_n24359_));
  AOI21X1  g21923(.A0(new_n24358_), .A1(new_n24357_), .B0(new_n24359_), .Y(new_n24360_));
  NOR3X1   g21924(.A(new_n24360_), .B(new_n24356_), .C(new_n11886_), .Y(new_n24361_));
  NOR3X1   g21925(.A(new_n24352_), .B(new_n24351_), .C(pi0789), .Y(new_n24362_));
  OR4X1    g21926(.A(new_n24362_), .B(new_n24361_), .C(new_n12841_), .D(new_n12691_), .Y(new_n24363_));
  AOI22X1  g21927(.A0(new_n24363_), .A1(new_n24230_), .B0(new_n24223_), .B1(pi0792), .Y(new_n24364_));
  OAI21X1  g21928(.A0(new_n24223_), .A1(new_n16350_), .B0(new_n14562_), .Y(new_n24365_));
  OAI22X1  g21929(.A0(new_n24365_), .A1(new_n24364_), .B0(new_n24217_), .B1(new_n11883_), .Y(new_n24366_));
  NOR2X1   g21930(.A(new_n24215_), .B(new_n24213_), .Y(new_n24367_));
  MX2X1    g21931(.A(new_n24367_), .B(new_n24211_), .S0(new_n11883_), .Y(new_n24368_));
  AOI21X1  g21932(.A0(new_n24368_), .A1(new_n12743_), .B0(new_n12739_), .Y(new_n24369_));
  OAI21X1  g21933(.A0(new_n24366_), .A1(new_n12743_), .B0(new_n24369_), .Y(new_n24370_));
  MX2X1    g21934(.A(new_n24150_), .B(new_n24029_), .S0(new_n12735_), .Y(new_n24371_));
  AOI21X1  g21935(.A0(new_n24028_), .A1(new_n12743_), .B0(pi0715), .Y(new_n24372_));
  OAI21X1  g21936(.A0(new_n24371_), .A1(new_n12743_), .B0(new_n24372_), .Y(new_n24373_));
  AND2X1   g21937(.A(new_n24373_), .B(pi1160), .Y(new_n24374_));
  AOI21X1  g21938(.A0(new_n24368_), .A1(pi0644), .B0(pi0715), .Y(new_n24375_));
  OAI21X1  g21939(.A0(new_n24366_), .A1(pi0644), .B0(new_n24375_), .Y(new_n24376_));
  AOI21X1  g21940(.A0(new_n24028_), .A1(pi0644), .B0(new_n12739_), .Y(new_n24377_));
  OAI21X1  g21941(.A0(new_n24371_), .A1(pi0644), .B0(new_n24377_), .Y(new_n24378_));
  AND2X1   g21942(.A(new_n24378_), .B(new_n11882_), .Y(new_n24379_));
  AOI22X1  g21943(.A0(new_n24379_), .A1(new_n24376_), .B0(new_n24374_), .B1(new_n24370_), .Y(new_n24380_));
  MX2X1    g21944(.A(new_n24380_), .B(new_n24366_), .S0(new_n12897_), .Y(new_n24381_));
  MX2X1    g21945(.A(new_n24381_), .B(pi0223), .S0(po1038), .Y(po0380));
  NOR2X1   g21946(.A(new_n23626_), .B(new_n2961_), .Y(new_n24383_));
  INVX1    g21947(.A(new_n24383_), .Y(new_n24384_));
  NOR3X1   g21948(.A(new_n12108_), .B(new_n12051_), .C(new_n5027_), .Y(new_n24385_));
  INVX1    g21949(.A(new_n24385_), .Y(new_n24386_));
  AOI21X1  g21950(.A0(new_n24386_), .A1(new_n12012_), .B0(new_n5028_), .Y(new_n24387_));
  AOI21X1  g21951(.A0(new_n12032_), .A1(new_n11950_), .B0(new_n24387_), .Y(new_n24388_));
  NOR2X1   g21952(.A(new_n24388_), .B(new_n11993_), .Y(new_n24389_));
  OAI21X1  g21953(.A0(new_n24385_), .A1(new_n12047_), .B0(pi0680), .Y(new_n24390_));
  OAI21X1  g21954(.A0(new_n24388_), .A1(pi0680), .B0(new_n24390_), .Y(new_n24391_));
  AOI21X1  g21955(.A0(new_n24391_), .A1(new_n11993_), .B0(new_n24389_), .Y(new_n24392_));
  NAND2X1  g21956(.A(new_n24392_), .B(new_n5070_), .Y(new_n24393_));
  AOI21X1  g21957(.A0(new_n12028_), .A1(new_n5033_), .B0(new_n12324_), .Y(new_n24394_));
  OAI21X1  g21958(.A0(new_n12031_), .A1(new_n5033_), .B0(new_n24394_), .Y(new_n24395_));
  AND2X1   g21959(.A(pi0616), .B(new_n12051_), .Y(new_n24396_));
  AOI22X1  g21960(.A0(new_n24396_), .A1(new_n12107_), .B0(new_n12291_), .B1(pi0614), .Y(new_n24397_));
  AOI21X1  g21961(.A0(new_n24397_), .A1(new_n24395_), .B0(new_n11993_), .Y(new_n24398_));
  AOI21X1  g21962(.A0(new_n24397_), .A1(new_n24395_), .B0(pi0680), .Y(new_n24399_));
  INVX1    g21963(.A(new_n24399_), .Y(new_n24400_));
  AOI21X1  g21964(.A0(new_n12352_), .A1(pi0614), .B0(new_n5029_), .Y(new_n24401_));
  AOI22X1  g21965(.A0(new_n24401_), .A1(new_n12046_), .B0(new_n24385_), .B1(pi0680), .Y(new_n24402_));
  AOI21X1  g21966(.A0(new_n24402_), .A1(new_n24400_), .B0(new_n12290_), .Y(new_n24403_));
  NOR3X1   g21967(.A(new_n24403_), .B(new_n24398_), .C(new_n5070_), .Y(new_n24404_));
  NOR2X1   g21968(.A(new_n24404_), .B(new_n2961_), .Y(new_n24405_));
  AND2X1   g21969(.A(new_n24385_), .B(new_n12056_), .Y(new_n24406_));
  AOI21X1  g21970(.A0(new_n24385_), .A1(new_n12056_), .B0(pi0680), .Y(new_n24407_));
  OAI21X1  g21971(.A0(new_n24407_), .A1(new_n24401_), .B0(new_n11993_), .Y(new_n24408_));
  OAI21X1  g21972(.A0(new_n24406_), .A1(new_n11993_), .B0(new_n24408_), .Y(new_n24409_));
  NOR2X1   g21973(.A(new_n23647_), .B(new_n12051_), .Y(new_n24410_));
  OAI21X1  g21974(.A0(new_n24410_), .A1(new_n5071_), .B0(new_n2961_), .Y(new_n24411_));
  AOI21X1  g21975(.A0(new_n24409_), .A1(new_n5071_), .B0(new_n24411_), .Y(new_n24412_));
  OR2X1    g21976(.A(new_n24412_), .B(new_n10136_), .Y(new_n24413_));
  AOI21X1  g21977(.A0(new_n24405_), .A1(new_n24393_), .B0(new_n24413_), .Y(new_n24414_));
  OAI21X1  g21978(.A0(new_n12012_), .A1(new_n2961_), .B0(new_n10136_), .Y(new_n24415_));
  NOR4X1   g21979(.A(new_n12171_), .B(new_n11952_), .C(new_n2740_), .D(new_n12051_), .Y(new_n24416_));
  OAI21X1  g21980(.A0(new_n24416_), .A1(new_n24415_), .B0(new_n2954_), .Y(new_n24417_));
  OAI21X1  g21981(.A0(new_n23667_), .A1(new_n12182_), .B0(pi0614), .Y(new_n24418_));
  OR2X1    g21982(.A(new_n24418_), .B(pi0224), .Y(new_n24419_));
  INVX1    g21983(.A(new_n24387_), .Y(new_n24420_));
  AOI21X1  g21984(.A0(new_n24420_), .A1(new_n11981_), .B0(new_n11993_), .Y(new_n24421_));
  AND2X1   g21985(.A(new_n24420_), .B(new_n11981_), .Y(new_n24422_));
  AOI21X1  g21986(.A0(new_n24385_), .A1(pi0680), .B0(new_n12003_), .Y(new_n24423_));
  OAI21X1  g21987(.A0(new_n24422_), .A1(pi0680), .B0(new_n24423_), .Y(new_n24424_));
  AOI21X1  g21988(.A0(new_n24424_), .A1(new_n11993_), .B0(new_n24421_), .Y(new_n24425_));
  AND2X1   g21989(.A(new_n24425_), .B(new_n5070_), .Y(new_n24426_));
  INVX1    g21990(.A(new_n23469_), .Y(new_n24427_));
  OAI21X1  g21991(.A0(new_n12147_), .A1(new_n12051_), .B0(new_n23468_), .Y(new_n24428_));
  AND2X1   g21992(.A(new_n12149_), .B(pi0680), .Y(new_n24429_));
  AOI22X1  g21993(.A0(new_n24429_), .A1(new_n24427_), .B0(new_n24428_), .B1(new_n5029_), .Y(new_n24430_));
  NAND2X1  g21994(.A(new_n24428_), .B(new_n12290_), .Y(new_n24431_));
  OAI21X1  g21995(.A0(new_n24430_), .A1(new_n12290_), .B0(new_n24431_), .Y(new_n24432_));
  OAI21X1  g21996(.A0(new_n24432_), .A1(new_n5070_), .B0(pi0224), .Y(new_n24433_));
  OAI22X1  g21997(.A0(new_n24433_), .A1(new_n24426_), .B0(new_n24419_), .B1(new_n12186_), .Y(new_n24434_));
  AOI21X1  g21998(.A0(new_n24434_), .A1(pi0215), .B0(new_n2953_), .Y(new_n24435_));
  OAI21X1  g21999(.A0(new_n24417_), .A1(new_n24414_), .B0(new_n24435_), .Y(new_n24436_));
  OAI21X1  g22000(.A0(new_n24432_), .A1(new_n5050_), .B0(pi0224), .Y(new_n24437_));
  AOI21X1  g22001(.A0(new_n24425_), .A1(new_n5050_), .B0(new_n24437_), .Y(new_n24438_));
  OAI21X1  g22002(.A0(new_n24419_), .A1(new_n12194_), .B0(pi0223), .Y(new_n24439_));
  AND2X1   g22003(.A(new_n24392_), .B(new_n5050_), .Y(new_n24440_));
  NOR3X1   g22004(.A(new_n24403_), .B(new_n24398_), .C(new_n5050_), .Y(new_n24441_));
  NOR3X1   g22005(.A(new_n24441_), .B(new_n24440_), .C(new_n2961_), .Y(new_n24442_));
  AND2X1   g22006(.A(new_n24409_), .B(new_n5051_), .Y(new_n24443_));
  OAI21X1  g22007(.A0(new_n24410_), .A1(new_n5051_), .B0(new_n6400_), .Y(new_n24444_));
  AOI21X1  g22008(.A0(new_n12190_), .A1(pi0614), .B0(pi0223), .Y(new_n24445_));
  OAI21X1  g22009(.A0(new_n24444_), .A1(new_n24443_), .B0(new_n24445_), .Y(new_n24446_));
  OAI22X1  g22010(.A0(new_n24446_), .A1(new_n24442_), .B0(new_n24439_), .B1(new_n24438_), .Y(new_n24447_));
  AOI21X1  g22011(.A0(new_n24447_), .A1(new_n2953_), .B0(new_n2959_), .Y(new_n24448_));
  AOI21X1  g22012(.A0(new_n12165_), .A1(new_n12051_), .B0(new_n2961_), .Y(new_n24449_));
  NOR4X1   g22013(.A(new_n12102_), .B(new_n12051_), .C(new_n5027_), .D(pi0224), .Y(new_n24450_));
  OR2X1    g22014(.A(new_n24450_), .B(pi0299), .Y(new_n24451_));
  AOI21X1  g22015(.A0(new_n24449_), .A1(new_n24112_), .B0(new_n24451_), .Y(new_n24452_));
  NAND3X1  g22016(.A(new_n12166_), .B(pi0614), .C(pi0603), .Y(new_n24453_));
  NOR2X1   g22017(.A(new_n12096_), .B(new_n2961_), .Y(new_n24454_));
  OAI22X1  g22018(.A0(new_n24454_), .A1(new_n24453_), .B0(new_n11943_), .B1(new_n2961_), .Y(new_n24455_));
  OAI21X1  g22019(.A0(new_n24455_), .A1(new_n2953_), .B0(new_n2959_), .Y(new_n24456_));
  OAI21X1  g22020(.A0(new_n24456_), .A1(new_n24452_), .B0(new_n2996_), .Y(new_n24457_));
  AOI21X1  g22021(.A0(new_n24448_), .A1(new_n24436_), .B0(new_n24457_), .Y(new_n24458_));
  OAI21X1  g22022(.A0(new_n12202_), .A1(new_n2961_), .B0(pi0038), .Y(new_n24459_));
  AOI21X1  g22023(.A0(new_n12205_), .A1(pi0614), .B0(new_n24459_), .Y(new_n24460_));
  OR2X1    g22024(.A(new_n24460_), .B(new_n3810_), .Y(new_n24461_));
  OAI22X1  g22025(.A0(new_n24461_), .A1(new_n24458_), .B0(new_n3129_), .B1(new_n2961_), .Y(new_n24462_));
  MX2X1    g22026(.A(new_n24462_), .B(new_n24383_), .S0(new_n12601_), .Y(new_n24463_));
  NAND2X1  g22027(.A(new_n24463_), .B(new_n11888_), .Y(new_n24464_));
  OR2X1    g22028(.A(new_n24463_), .B(new_n12590_), .Y(new_n24465_));
  AOI21X1  g22029(.A0(new_n24384_), .A1(new_n12590_), .B0(new_n12591_), .Y(new_n24466_));
  OR2X1    g22030(.A(new_n24463_), .B(pi0609), .Y(new_n24467_));
  AOI21X1  g22031(.A0(new_n24384_), .A1(pi0609), .B0(pi1155), .Y(new_n24468_));
  AOI22X1  g22032(.A0(new_n24468_), .A1(new_n24467_), .B0(new_n24466_), .B1(new_n24465_), .Y(new_n24469_));
  OAI21X1  g22033(.A0(new_n24469_), .A1(new_n11888_), .B0(new_n24464_), .Y(new_n24470_));
  AND2X1   g22034(.A(new_n24470_), .B(new_n11887_), .Y(new_n24471_));
  AOI21X1  g22035(.A0(new_n24384_), .A1(new_n12614_), .B0(new_n12615_), .Y(new_n24472_));
  OAI21X1  g22036(.A0(new_n24470_), .A1(new_n12614_), .B0(new_n24472_), .Y(new_n24473_));
  AOI21X1  g22037(.A0(new_n24384_), .A1(pi0618), .B0(pi1154), .Y(new_n24474_));
  OAI21X1  g22038(.A0(new_n24470_), .A1(pi0618), .B0(new_n24474_), .Y(new_n24475_));
  AOI21X1  g22039(.A0(new_n24475_), .A1(new_n24473_), .B0(new_n11887_), .Y(new_n24476_));
  OAI21X1  g22040(.A0(new_n24476_), .A1(new_n24471_), .B0(new_n11886_), .Y(new_n24477_));
  NOR3X1   g22041(.A(new_n24476_), .B(new_n24471_), .C(new_n12637_), .Y(new_n24478_));
  OAI21X1  g22042(.A0(new_n24383_), .A1(pi0619), .B0(pi1159), .Y(new_n24479_));
  NOR2X1   g22043(.A(new_n24479_), .B(new_n24478_), .Y(new_n24480_));
  NOR3X1   g22044(.A(new_n24476_), .B(new_n24471_), .C(pi0619), .Y(new_n24481_));
  OAI21X1  g22045(.A0(new_n24383_), .A1(new_n12637_), .B0(new_n12638_), .Y(new_n24482_));
  NOR2X1   g22046(.A(new_n24482_), .B(new_n24481_), .Y(new_n24483_));
  OAI21X1  g22047(.A0(new_n24483_), .A1(new_n24480_), .B0(pi0789), .Y(new_n24484_));
  AND2X1   g22048(.A(new_n24484_), .B(new_n24477_), .Y(new_n24485_));
  MX2X1    g22049(.A(new_n24485_), .B(new_n24384_), .S0(new_n12841_), .Y(new_n24486_));
  NOR2X1   g22050(.A(new_n3129_), .B(new_n2961_), .Y(new_n24487_));
  AND2X1   g22051(.A(pi0680), .B(pi0662), .Y(new_n24488_));
  NOR2X1   g22052(.A(new_n24488_), .B(new_n12458_), .Y(new_n24489_));
  AND2X1   g22053(.A(new_n12458_), .B(new_n2961_), .Y(new_n24490_));
  OAI21X1  g22054(.A0(new_n12449_), .A1(new_n2961_), .B0(new_n2953_), .Y(new_n24491_));
  NOR3X1   g22055(.A(new_n24491_), .B(new_n24490_), .C(new_n24489_), .Y(new_n24492_));
  INVX1    g22056(.A(new_n24488_), .Y(new_n24493_));
  AND2X1   g22057(.A(new_n24493_), .B(new_n12463_), .Y(new_n24494_));
  AOI21X1  g22058(.A0(new_n13240_), .A1(pi0224), .B0(new_n2953_), .Y(new_n24495_));
  OAI21X1  g22059(.A0(new_n12463_), .A1(pi0224), .B0(new_n24495_), .Y(new_n24496_));
  OAI21X1  g22060(.A0(new_n24496_), .A1(new_n24494_), .B0(new_n2959_), .Y(new_n24497_));
  NOR4X1   g22061(.A(new_n24493_), .B(new_n12210_), .C(new_n11952_), .D(new_n2740_), .Y(new_n24498_));
  MX2X1    g22062(.A(new_n12528_), .B(new_n12055_), .S0(new_n11977_), .Y(new_n24499_));
  OAI21X1  g22063(.A0(new_n23756_), .A1(new_n11978_), .B0(new_n12063_), .Y(new_n24500_));
  OAI21X1  g22064(.A0(new_n24500_), .A1(new_n5070_), .B0(pi0224), .Y(new_n24501_));
  AOI21X1  g22065(.A0(new_n24499_), .A1(new_n5070_), .B0(new_n24501_), .Y(new_n24502_));
  AND2X1   g22066(.A(new_n12341_), .B(new_n12057_), .Y(new_n24503_));
  AOI21X1  g22067(.A0(new_n24503_), .A1(pi0662), .B0(new_n5070_), .Y(new_n24504_));
  INVX1    g22068(.A(new_n12502_), .Y(new_n24505_));
  AOI21X1  g22069(.A0(new_n24488_), .A1(new_n24505_), .B0(new_n5071_), .Y(new_n24506_));
  NOR3X1   g22070(.A(new_n24506_), .B(new_n24504_), .C(pi0224), .Y(new_n24507_));
  OR2X1    g22071(.A(new_n24507_), .B(new_n10136_), .Y(new_n24508_));
  OAI22X1  g22072(.A0(new_n24508_), .A1(new_n24502_), .B0(new_n24498_), .B1(new_n24415_), .Y(new_n24509_));
  INVX1    g22073(.A(new_n12545_), .Y(new_n24510_));
  MX2X1    g22074(.A(new_n24510_), .B(new_n12082_), .S0(new_n11977_), .Y(new_n24511_));
  MX2X1    g22075(.A(new_n23767_), .B(new_n12009_), .S0(new_n11977_), .Y(new_n24512_));
  OAI21X1  g22076(.A0(new_n24512_), .A1(new_n5071_), .B0(pi0224), .Y(new_n24513_));
  AOI21X1  g22077(.A0(new_n24511_), .A1(new_n5071_), .B0(new_n24513_), .Y(new_n24514_));
  OR2X1    g22078(.A(new_n11977_), .B(pi0224), .Y(new_n24515_));
  NOR4X1   g22079(.A(new_n24515_), .B(new_n12378_), .C(new_n12186_), .D(new_n5029_), .Y(new_n24516_));
  OR2X1    g22080(.A(new_n24516_), .B(new_n2954_), .Y(new_n24517_));
  OAI21X1  g22081(.A0(new_n24517_), .A1(new_n24514_), .B0(pi0299), .Y(new_n24518_));
  AOI21X1  g22082(.A0(new_n24509_), .A1(new_n2954_), .B0(new_n24518_), .Y(new_n24519_));
  OAI21X1  g22083(.A0(new_n24500_), .A1(new_n5050_), .B0(pi0224), .Y(new_n24520_));
  AOI21X1  g22084(.A0(new_n24499_), .A1(new_n5050_), .B0(new_n24520_), .Y(new_n24521_));
  AOI21X1  g22085(.A0(new_n24503_), .A1(pi0662), .B0(new_n5050_), .Y(new_n24522_));
  AOI21X1  g22086(.A0(new_n24488_), .A1(new_n24505_), .B0(new_n5051_), .Y(new_n24523_));
  NOR3X1   g22087(.A(new_n24523_), .B(new_n24522_), .C(new_n6401_), .Y(new_n24524_));
  OAI21X1  g22088(.A0(new_n12500_), .A1(new_n11977_), .B0(new_n2964_), .Y(new_n24525_));
  NOR3X1   g22089(.A(new_n24525_), .B(new_n24524_), .C(new_n24521_), .Y(new_n24526_));
  OAI21X1  g22090(.A0(new_n24512_), .A1(new_n5051_), .B0(pi0224), .Y(new_n24527_));
  AOI21X1  g22091(.A0(new_n24511_), .A1(new_n5051_), .B0(new_n24527_), .Y(new_n24528_));
  NOR4X1   g22092(.A(new_n24515_), .B(new_n12378_), .C(new_n12194_), .D(new_n5029_), .Y(new_n24529_));
  OR2X1    g22093(.A(new_n24529_), .B(new_n2964_), .Y(new_n24530_));
  OAI21X1  g22094(.A0(new_n24530_), .A1(new_n24528_), .B0(new_n2953_), .Y(new_n24531_));
  OAI21X1  g22095(.A0(new_n24531_), .A1(new_n24526_), .B0(pi0039), .Y(new_n24532_));
  OAI22X1  g22096(.A0(new_n24532_), .A1(new_n24519_), .B0(new_n24497_), .B1(new_n24492_), .Y(new_n24533_));
  NOR4X1   g22097(.A(new_n13585_), .B(new_n3074_), .C(new_n11977_), .D(pi0039), .Y(new_n24534_));
  OAI21X1  g22098(.A0(new_n24534_), .A1(new_n24459_), .B0(new_n3129_), .Y(new_n24535_));
  AOI21X1  g22099(.A0(new_n24533_), .A1(new_n2996_), .B0(new_n24535_), .Y(new_n24536_));
  NOR2X1   g22100(.A(new_n24536_), .B(new_n24487_), .Y(new_n24537_));
  NAND2X1  g22101(.A(new_n24537_), .B(pi0625), .Y(new_n24538_));
  AOI21X1  g22102(.A0(new_n24384_), .A1(new_n12493_), .B0(new_n12494_), .Y(new_n24539_));
  NAND2X1  g22103(.A(new_n24537_), .B(new_n12493_), .Y(new_n24540_));
  AOI21X1  g22104(.A0(new_n24384_), .A1(pi0625), .B0(pi1153), .Y(new_n24541_));
  AOI22X1  g22105(.A0(new_n24541_), .A1(new_n24540_), .B0(new_n24539_), .B1(new_n24538_), .Y(new_n24542_));
  MX2X1    g22106(.A(new_n24542_), .B(new_n24537_), .S0(new_n11889_), .Y(new_n24543_));
  MX2X1    g22107(.A(new_n24543_), .B(new_n24384_), .S0(new_n12618_), .Y(new_n24544_));
  MX2X1    g22108(.A(new_n24544_), .B(new_n24384_), .S0(new_n12641_), .Y(new_n24545_));
  AND2X1   g22109(.A(new_n24545_), .B(new_n22011_), .Y(new_n24546_));
  AOI22X1  g22110(.A0(new_n24546_), .A1(new_n17252_), .B0(new_n24384_), .B1(new_n22010_), .Y(new_n24547_));
  AOI21X1  g22111(.A0(new_n24384_), .A1(pi0628), .B0(new_n12710_), .Y(new_n24548_));
  OAI21X1  g22112(.A0(new_n24547_), .A1(pi0628), .B0(new_n24548_), .Y(new_n24549_));
  AOI21X1  g22113(.A0(new_n24384_), .A1(new_n12683_), .B0(new_n12708_), .Y(new_n24550_));
  OAI21X1  g22114(.A0(new_n24547_), .A1(new_n12683_), .B0(new_n24550_), .Y(new_n24551_));
  AND2X1   g22115(.A(new_n24551_), .B(new_n24549_), .Y(new_n24552_));
  OAI21X1  g22116(.A0(new_n24486_), .A1(new_n14395_), .B0(new_n24552_), .Y(new_n24553_));
  NOR2X1   g22117(.A(new_n24388_), .B(pi0680), .Y(new_n24554_));
  MX2X1    g22118(.A(new_n23941_), .B(new_n16526_), .S0(new_n12051_), .Y(new_n24555_));
  OAI21X1  g22119(.A0(new_n11959_), .A1(pi0120), .B0(new_n24555_), .Y(new_n24556_));
  AND2X1   g22120(.A(new_n24556_), .B(pi0616), .Y(new_n24557_));
  INVX1    g22121(.A(new_n24557_), .Y(new_n24558_));
  NOR2X1   g22122(.A(new_n12408_), .B(new_n12051_), .Y(new_n24559_));
  OAI21X1  g22123(.A0(new_n24559_), .A1(new_n12248_), .B0(new_n11950_), .Y(new_n24560_));
  AOI21X1  g22124(.A0(new_n24560_), .A1(new_n24558_), .B0(new_n5029_), .Y(new_n24561_));
  OAI21X1  g22125(.A0(new_n24561_), .A1(new_n24554_), .B0(pi0662), .Y(new_n24562_));
  NOR2X1   g22126(.A(new_n23382_), .B(pi0662), .Y(new_n24563_));
  INVX1    g22127(.A(new_n24563_), .Y(new_n24564_));
  NOR2X1   g22128(.A(new_n24564_), .B(new_n24388_), .Y(new_n24565_));
  AOI21X1  g22129(.A0(new_n24391_), .A1(new_n11993_), .B0(new_n24565_), .Y(new_n24566_));
  NAND2X1  g22130(.A(new_n24566_), .B(new_n24562_), .Y(new_n24567_));
  INVX1    g22131(.A(new_n24410_), .Y(new_n24568_));
  INVX1    g22132(.A(new_n24396_), .Y(new_n24569_));
  OAI22X1  g22133(.A0(new_n24569_), .A1(new_n12308_), .B0(new_n12361_), .B1(new_n11950_), .Y(new_n24570_));
  NAND2X1  g22134(.A(new_n24570_), .B(pi0680), .Y(new_n24571_));
  OAI21X1  g22135(.A0(new_n24416_), .A1(new_n23849_), .B0(new_n24571_), .Y(new_n24572_));
  MX2X1    g22136(.A(new_n24572_), .B(new_n24568_), .S0(new_n11977_), .Y(new_n24573_));
  AOI21X1  g22137(.A0(new_n24573_), .A1(new_n2961_), .B0(new_n5071_), .Y(new_n24574_));
  OAI21X1  g22138(.A0(new_n24567_), .A1(new_n2961_), .B0(new_n24574_), .Y(new_n24575_));
  AOI21X1  g22139(.A0(new_n12354_), .A1(pi0614), .B0(new_n5029_), .Y(new_n24576_));
  OAI21X1  g22140(.A0(new_n12305_), .A1(pi0614), .B0(new_n24576_), .Y(new_n24577_));
  OAI21X1  g22141(.A0(new_n24406_), .A1(pi0680), .B0(new_n24577_), .Y(new_n24578_));
  OAI21X1  g22142(.A0(new_n24564_), .A1(new_n24406_), .B0(new_n24408_), .Y(new_n24579_));
  AOI21X1  g22143(.A0(new_n24578_), .A1(pi0662), .B0(new_n24579_), .Y(new_n24580_));
  OAI22X1  g22144(.A0(new_n24569_), .A1(new_n23820_), .B0(new_n23826_), .B1(new_n12051_), .Y(new_n24581_));
  OAI21X1  g22145(.A0(new_n24581_), .A1(new_n23823_), .B0(pi0680), .Y(new_n24582_));
  AOI21X1  g22146(.A0(new_n24582_), .A1(new_n24400_), .B0(new_n11977_), .Y(new_n24583_));
  AOI21X1  g22147(.A0(new_n24397_), .A1(new_n24395_), .B0(new_n24564_), .Y(new_n24584_));
  NOR3X1   g22148(.A(new_n24584_), .B(new_n24583_), .C(new_n24403_), .Y(new_n24585_));
  AOI21X1  g22149(.A0(new_n24585_), .A1(pi0224), .B0(new_n5070_), .Y(new_n24586_));
  OAI21X1  g22150(.A0(new_n24580_), .A1(pi0224), .B0(new_n24586_), .Y(new_n24587_));
  NAND3X1  g22151(.A(new_n24587_), .B(new_n24575_), .C(new_n10137_), .Y(new_n24588_));
  AOI21X1  g22152(.A0(new_n24488_), .A1(new_n12308_), .B0(new_n24416_), .Y(new_n24589_));
  OR2X1    g22153(.A(new_n24589_), .B(pi0224), .Y(new_n24590_));
  OR2X1    g22154(.A(new_n24488_), .B(new_n24385_), .Y(new_n24591_));
  OAI21X1  g22155(.A0(new_n24591_), .A1(new_n12416_), .B0(pi0224), .Y(new_n24592_));
  AOI21X1  g22156(.A0(new_n24555_), .A1(new_n24488_), .B0(new_n24592_), .Y(new_n24593_));
  NOR2X1   g22157(.A(new_n24593_), .B(new_n24415_), .Y(new_n24594_));
  AOI21X1  g22158(.A0(new_n24594_), .A1(new_n24590_), .B0(pi0215), .Y(new_n24595_));
  OAI21X1  g22159(.A0(new_n12408_), .A1(new_n12051_), .B0(new_n12226_), .Y(new_n24596_));
  AOI21X1  g22160(.A0(new_n24596_), .A1(new_n11950_), .B0(new_n24557_), .Y(new_n24597_));
  MX2X1    g22161(.A(new_n24597_), .B(new_n24422_), .S0(new_n5029_), .Y(new_n24598_));
  AOI21X1  g22162(.A0(new_n24420_), .A1(new_n11981_), .B0(new_n24564_), .Y(new_n24599_));
  AOI21X1  g22163(.A0(new_n24424_), .A1(new_n11993_), .B0(new_n24599_), .Y(new_n24600_));
  OAI21X1  g22164(.A0(new_n24598_), .A1(new_n11977_), .B0(new_n24600_), .Y(new_n24601_));
  OAI21X1  g22165(.A0(new_n23871_), .A1(new_n12051_), .B0(new_n12239_), .Y(new_n24602_));
  MX2X1    g22166(.A(new_n24602_), .B(new_n24428_), .S0(new_n5029_), .Y(new_n24603_));
  NAND2X1  g22167(.A(new_n24563_), .B(new_n24428_), .Y(new_n24604_));
  OAI21X1  g22168(.A0(new_n24430_), .A1(new_n12290_), .B0(new_n24604_), .Y(new_n24605_));
  AOI21X1  g22169(.A0(new_n24603_), .A1(pi0662), .B0(new_n24605_), .Y(new_n24606_));
  OAI21X1  g22170(.A0(new_n24606_), .A1(new_n5070_), .B0(pi0224), .Y(new_n24607_));
  AOI21X1  g22171(.A0(new_n24601_), .A1(new_n5070_), .B0(new_n24607_), .Y(new_n24608_));
  AND2X1   g22172(.A(new_n12334_), .B(pi0680), .Y(new_n24609_));
  OAI21X1  g22173(.A0(new_n24609_), .A1(new_n24416_), .B0(new_n24571_), .Y(new_n24610_));
  MX2X1    g22174(.A(new_n24610_), .B(new_n24418_), .S0(new_n11977_), .Y(new_n24611_));
  NOR2X1   g22175(.A(new_n24611_), .B(new_n5071_), .Y(new_n24612_));
  OAI21X1  g22176(.A0(new_n24418_), .A1(new_n11966_), .B0(new_n11977_), .Y(new_n24613_));
  OR2X1    g22177(.A(new_n12328_), .B(new_n12324_), .Y(new_n24614_));
  OAI21X1  g22178(.A0(new_n23881_), .A1(new_n12051_), .B0(pi0680), .Y(new_n24615_));
  AOI21X1  g22179(.A0(new_n12322_), .A1(new_n12051_), .B0(new_n24615_), .Y(new_n24616_));
  AND2X1   g22180(.A(new_n24616_), .B(new_n24614_), .Y(new_n24617_));
  OR2X1    g22181(.A(pi0680), .B(new_n12051_), .Y(new_n24618_));
  OAI21X1  g22182(.A0(new_n24618_), .A1(new_n24075_), .B0(pi0662), .Y(new_n24619_));
  OAI21X1  g22183(.A0(new_n24619_), .A1(new_n24617_), .B0(new_n24613_), .Y(new_n24620_));
  OAI21X1  g22184(.A0(new_n24620_), .A1(new_n5070_), .B0(new_n2961_), .Y(new_n24621_));
  OAI21X1  g22185(.A0(new_n24621_), .A1(new_n24612_), .B0(pi0215), .Y(new_n24622_));
  OAI21X1  g22186(.A0(new_n24622_), .A1(new_n24608_), .B0(pi0299), .Y(new_n24623_));
  AOI21X1  g22187(.A0(new_n24595_), .A1(new_n24588_), .B0(new_n24623_), .Y(new_n24624_));
  AOI21X1  g22188(.A0(new_n24585_), .A1(new_n5051_), .B0(new_n2961_), .Y(new_n24625_));
  OAI21X1  g22189(.A0(new_n24567_), .A1(new_n5051_), .B0(new_n24625_), .Y(new_n24626_));
  OR2X1    g22190(.A(new_n24580_), .B(new_n5050_), .Y(new_n24627_));
  AOI21X1  g22191(.A0(new_n24573_), .A1(new_n5050_), .B0(new_n6401_), .Y(new_n24628_));
  OAI21X1  g22192(.A0(new_n24590_), .A1(pi0222), .B0(new_n2964_), .Y(new_n24629_));
  AOI21X1  g22193(.A0(new_n24628_), .A1(new_n24627_), .B0(new_n24629_), .Y(new_n24630_));
  AOI21X1  g22194(.A0(new_n24611_), .A1(new_n2961_), .B0(new_n5051_), .Y(new_n24631_));
  OAI21X1  g22195(.A0(new_n24601_), .A1(new_n2961_), .B0(new_n24631_), .Y(new_n24632_));
  NAND2X1  g22196(.A(new_n24606_), .B(pi0224), .Y(new_n24633_));
  AOI21X1  g22197(.A0(new_n24620_), .A1(new_n2961_), .B0(new_n5050_), .Y(new_n24634_));
  AOI21X1  g22198(.A0(new_n24634_), .A1(new_n24633_), .B0(new_n2964_), .Y(new_n24635_));
  AOI22X1  g22199(.A0(new_n24635_), .A1(new_n24632_), .B0(new_n24630_), .B1(new_n24626_), .Y(new_n24636_));
  OAI21X1  g22200(.A0(new_n24636_), .A1(pi0299), .B0(pi0039), .Y(new_n24637_));
  OAI22X1  g22201(.A0(new_n24493_), .A1(new_n23918_), .B0(new_n13222_), .B1(new_n12051_), .Y(new_n24638_));
  NAND3X1  g22202(.A(new_n24493_), .B(new_n12461_), .C(new_n12459_), .Y(new_n24639_));
  AND2X1   g22203(.A(new_n24449_), .B(new_n24307_), .Y(new_n24640_));
  AOI22X1  g22204(.A0(new_n24640_), .A1(new_n24639_), .B0(new_n24638_), .B1(new_n2961_), .Y(new_n24641_));
  OAI22X1  g22205(.A0(new_n23931_), .A1(new_n23929_), .B0(new_n13239_), .B1(pi0614), .Y(new_n24642_));
  NAND2X1  g22206(.A(new_n24642_), .B(pi0224), .Y(new_n24643_));
  NAND3X1  g22207(.A(new_n24453_), .B(new_n23928_), .C(new_n2961_), .Y(new_n24644_));
  AOI21X1  g22208(.A0(new_n24644_), .A1(new_n24643_), .B0(new_n24493_), .Y(new_n24645_));
  OAI21X1  g22209(.A0(new_n24488_), .A1(new_n24455_), .B0(pi0299), .Y(new_n24646_));
  OAI22X1  g22210(.A0(new_n24646_), .A1(new_n24645_), .B0(new_n24641_), .B1(pi0299), .Y(new_n24647_));
  AOI21X1  g22211(.A0(new_n24647_), .A1(new_n2959_), .B0(pi0038), .Y(new_n24648_));
  OAI21X1  g22212(.A0(new_n24637_), .A1(new_n24624_), .B0(new_n24648_), .Y(new_n24649_));
  NAND3X1  g22213(.A(new_n12269_), .B(new_n12202_), .C(pi0662), .Y(new_n24650_));
  AOI21X1  g22214(.A0(new_n24650_), .A1(new_n24460_), .B0(new_n3810_), .Y(new_n24651_));
  AOI21X1  g22215(.A0(new_n24651_), .A1(new_n24649_), .B0(new_n24487_), .Y(new_n24652_));
  AND2X1   g22216(.A(new_n24652_), .B(new_n12493_), .Y(new_n24653_));
  OAI21X1  g22217(.A0(new_n24462_), .A1(new_n12493_), .B0(new_n12494_), .Y(new_n24654_));
  AOI21X1  g22218(.A0(new_n24539_), .A1(new_n24538_), .B0(pi0608), .Y(new_n24655_));
  OAI21X1  g22219(.A0(new_n24654_), .A1(new_n24653_), .B0(new_n24655_), .Y(new_n24656_));
  AND2X1   g22220(.A(new_n24652_), .B(pi0625), .Y(new_n24657_));
  OAI21X1  g22221(.A0(new_n24462_), .A1(pi0625), .B0(pi1153), .Y(new_n24658_));
  AOI21X1  g22222(.A0(new_n24541_), .A1(new_n24540_), .B0(new_n12584_), .Y(new_n24659_));
  OAI21X1  g22223(.A0(new_n24658_), .A1(new_n24657_), .B0(new_n24659_), .Y(new_n24660_));
  AOI21X1  g22224(.A0(new_n24660_), .A1(new_n24656_), .B0(new_n11889_), .Y(new_n24661_));
  AOI21X1  g22225(.A0(new_n24652_), .A1(new_n11889_), .B0(new_n24661_), .Y(new_n24662_));
  AOI21X1  g22226(.A0(new_n24543_), .A1(pi0609), .B0(pi1155), .Y(new_n24663_));
  OAI21X1  g22227(.A0(new_n24662_), .A1(pi0609), .B0(new_n24663_), .Y(new_n24664_));
  AOI21X1  g22228(.A0(new_n24466_), .A1(new_n24465_), .B0(pi0660), .Y(new_n24665_));
  AOI21X1  g22229(.A0(new_n24543_), .A1(new_n12590_), .B0(new_n12591_), .Y(new_n24666_));
  OAI21X1  g22230(.A0(new_n24662_), .A1(new_n12590_), .B0(new_n24666_), .Y(new_n24667_));
  AOI21X1  g22231(.A0(new_n24468_), .A1(new_n24467_), .B0(new_n12596_), .Y(new_n24668_));
  AOI22X1  g22232(.A0(new_n24668_), .A1(new_n24667_), .B0(new_n24665_), .B1(new_n24664_), .Y(new_n24669_));
  MX2X1    g22233(.A(new_n24669_), .B(new_n24662_), .S0(new_n11888_), .Y(new_n24670_));
  AOI21X1  g22234(.A0(new_n24544_), .A1(pi0618), .B0(pi1154), .Y(new_n24671_));
  OAI21X1  g22235(.A0(new_n24670_), .A1(pi0618), .B0(new_n24671_), .Y(new_n24672_));
  AND2X1   g22236(.A(new_n24473_), .B(new_n12622_), .Y(new_n24673_));
  AOI21X1  g22237(.A0(new_n24544_), .A1(new_n12614_), .B0(new_n12615_), .Y(new_n24674_));
  OAI21X1  g22238(.A0(new_n24670_), .A1(new_n12614_), .B0(new_n24674_), .Y(new_n24675_));
  AND2X1   g22239(.A(new_n24475_), .B(pi0627), .Y(new_n24676_));
  AOI22X1  g22240(.A0(new_n24676_), .A1(new_n24675_), .B0(new_n24673_), .B1(new_n24672_), .Y(new_n24677_));
  MX2X1    g22241(.A(new_n24677_), .B(new_n24670_), .S0(new_n11887_), .Y(new_n24678_));
  AOI21X1  g22242(.A0(new_n24545_), .A1(pi0619), .B0(pi1159), .Y(new_n24679_));
  OAI21X1  g22243(.A0(new_n24678_), .A1(pi0619), .B0(new_n24679_), .Y(new_n24680_));
  NOR2X1   g22244(.A(new_n24480_), .B(pi0648), .Y(new_n24681_));
  AND2X1   g22245(.A(new_n24681_), .B(new_n24680_), .Y(new_n24682_));
  OR2X1    g22246(.A(new_n24678_), .B(new_n12637_), .Y(new_n24683_));
  AOI21X1  g22247(.A0(new_n24545_), .A1(new_n12637_), .B0(new_n12638_), .Y(new_n24684_));
  OAI21X1  g22248(.A0(new_n24482_), .A1(new_n24481_), .B0(pi0648), .Y(new_n24685_));
  AOI21X1  g22249(.A0(new_n24684_), .A1(new_n24683_), .B0(new_n24685_), .Y(new_n24686_));
  OR2X1    g22250(.A(new_n24686_), .B(new_n11886_), .Y(new_n24687_));
  AOI21X1  g22251(.A0(new_n24678_), .A1(new_n11886_), .B0(new_n14264_), .Y(new_n24688_));
  OAI21X1  g22252(.A0(new_n24687_), .A1(new_n24682_), .B0(new_n24688_), .Y(new_n24689_));
  AOI21X1  g22253(.A0(new_n24383_), .A1(new_n12664_), .B0(new_n16356_), .Y(new_n24690_));
  OAI21X1  g22254(.A0(new_n24485_), .A1(new_n12664_), .B0(new_n24690_), .Y(new_n24691_));
  AOI21X1  g22255(.A0(new_n24383_), .A1(pi0626), .B0(new_n16352_), .Y(new_n24692_));
  OAI21X1  g22256(.A0(new_n24485_), .A1(pi0626), .B0(new_n24692_), .Y(new_n24693_));
  MX2X1    g22257(.A(new_n24545_), .B(new_n24384_), .S0(new_n12659_), .Y(new_n24694_));
  NAND2X1  g22258(.A(new_n24694_), .B(new_n12769_), .Y(new_n24695_));
  NAND3X1  g22259(.A(new_n24695_), .B(new_n24693_), .C(new_n24691_), .Y(new_n24696_));
  AOI21X1  g22260(.A0(new_n24696_), .A1(pi0788), .B0(new_n14273_), .Y(new_n24697_));
  AOI22X1  g22261(.A0(new_n24697_), .A1(new_n24689_), .B0(new_n24553_), .B1(pi0792), .Y(new_n24698_));
  NAND2X1  g22262(.A(new_n24383_), .B(new_n12711_), .Y(new_n24699_));
  OAI21X1  g22263(.A0(new_n24486_), .A1(new_n12711_), .B0(new_n24699_), .Y(new_n24700_));
  OAI22X1  g22264(.A0(new_n24547_), .A1(new_n13639_), .B0(new_n24383_), .B1(new_n22842_), .Y(new_n24701_));
  OAI21X1  g22265(.A0(new_n24383_), .A1(pi0647), .B0(pi1157), .Y(new_n24702_));
  AOI21X1  g22266(.A0(new_n24701_), .A1(pi0647), .B0(new_n24702_), .Y(new_n24703_));
  OAI21X1  g22267(.A0(new_n24383_), .A1(new_n12705_), .B0(new_n12706_), .Y(new_n24704_));
  AOI21X1  g22268(.A0(new_n24701_), .A1(new_n12705_), .B0(new_n24704_), .Y(new_n24705_));
  MX2X1    g22269(.A(new_n24705_), .B(new_n24703_), .S0(new_n12723_), .Y(new_n24706_));
  AOI21X1  g22270(.A0(new_n24700_), .A1(new_n14385_), .B0(new_n24706_), .Y(new_n24707_));
  OAI22X1  g22271(.A0(new_n24707_), .A1(new_n11883_), .B0(new_n24698_), .B1(new_n14269_), .Y(new_n24708_));
  NOR2X1   g22272(.A(new_n24705_), .B(new_n24703_), .Y(new_n24709_));
  MX2X1    g22273(.A(new_n24709_), .B(new_n24701_), .S0(new_n11883_), .Y(new_n24710_));
  AOI21X1  g22274(.A0(new_n24710_), .A1(new_n12743_), .B0(new_n12739_), .Y(new_n24711_));
  OAI21X1  g22275(.A0(new_n24708_), .A1(new_n12743_), .B0(new_n24711_), .Y(new_n24712_));
  MX2X1    g22276(.A(new_n24700_), .B(new_n24383_), .S0(new_n12735_), .Y(new_n24713_));
  AOI21X1  g22277(.A0(new_n24384_), .A1(new_n12743_), .B0(pi0715), .Y(new_n24714_));
  OAI21X1  g22278(.A0(new_n24713_), .A1(new_n12743_), .B0(new_n24714_), .Y(new_n24715_));
  AND2X1   g22279(.A(new_n24715_), .B(pi1160), .Y(new_n24716_));
  AOI21X1  g22280(.A0(new_n24710_), .A1(pi0644), .B0(pi0715), .Y(new_n24717_));
  OAI21X1  g22281(.A0(new_n24708_), .A1(pi0644), .B0(new_n24717_), .Y(new_n24718_));
  AOI21X1  g22282(.A0(new_n24384_), .A1(pi0644), .B0(new_n12739_), .Y(new_n24719_));
  OAI21X1  g22283(.A0(new_n24713_), .A1(pi0644), .B0(new_n24719_), .Y(new_n24720_));
  AND2X1   g22284(.A(new_n24720_), .B(new_n11882_), .Y(new_n24721_));
  AOI22X1  g22285(.A0(new_n24721_), .A1(new_n24718_), .B0(new_n24716_), .B1(new_n24712_), .Y(new_n24722_));
  MX2X1    g22286(.A(new_n24722_), .B(new_n24708_), .S0(new_n12897_), .Y(new_n24723_));
  MX2X1    g22287(.A(new_n24723_), .B(pi0224), .S0(po1038), .Y(po0381));
  OR2X1    g22288(.A(new_n5822_), .B(pi0056), .Y(new_n24725_));
  AOI21X1  g22289(.A0(new_n5083_), .A1(new_n7169_), .B0(pi0137), .Y(new_n24726_));
  NOR4X1   g22290(.A(new_n24726_), .B(new_n5086_), .C(new_n3074_), .D(pi0039), .Y(new_n24727_));
  NAND3X1  g22291(.A(new_n8529_), .B(new_n2873_), .C(new_n2706_), .Y(new_n24728_));
  AOI21X1  g22292(.A0(new_n24728_), .A1(new_n2553_), .B0(new_n2547_), .Y(new_n24729_));
  OAI21X1  g22293(.A0(new_n24729_), .A1(new_n2730_), .B0(new_n2540_), .Y(new_n24730_));
  AOI21X1  g22294(.A0(new_n24730_), .A1(new_n2815_), .B0(new_n2453_), .Y(new_n24731_));
  OR2X1    g22295(.A(new_n2723_), .B(pi0137), .Y(new_n24732_));
  NOR2X1   g22296(.A(new_n2769_), .B(pi0032), .Y(new_n24733_));
  OAI21X1  g22297(.A0(new_n8529_), .A1(new_n2458_), .B0(new_n24733_), .Y(new_n24734_));
  AND2X1   g22298(.A(new_n24734_), .B(new_n2776_), .Y(new_n24735_));
  NOR3X1   g22299(.A(new_n2785_), .B(new_n2730_), .C(pi0095), .Y(new_n24736_));
  OR2X1    g22300(.A(new_n5916_), .B(new_n2458_), .Y(new_n24737_));
  NOR4X1   g22301(.A(new_n24737_), .B(new_n2709_), .C(new_n5134_), .D(pi0051), .Y(new_n24738_));
  AOI22X1  g22302(.A0(new_n24738_), .A1(new_n24736_), .B0(new_n24735_), .B1(new_n2785_), .Y(new_n24739_));
  INVX1    g22303(.A(new_n24739_), .Y(new_n24740_));
  INVX1    g22304(.A(new_n24735_), .Y(new_n24741_));
  OAI21X1  g22305(.A0(new_n24737_), .A1(new_n2525_), .B0(new_n2456_), .Y(new_n24742_));
  AOI21X1  g22306(.A0(new_n24742_), .A1(new_n24736_), .B0(pi1093), .Y(new_n24743_));
  AOI22X1  g22307(.A0(new_n24739_), .A1(new_n24743_), .B0(new_n24741_), .B1(pi1093), .Y(new_n24744_));
  OR2X1    g22308(.A(new_n2805_), .B(new_n2784_), .Y(new_n24745_));
  AND2X1   g22309(.A(new_n24745_), .B(new_n24743_), .Y(new_n24746_));
  OAI21X1  g22310(.A0(new_n24737_), .A1(new_n2752_), .B0(new_n2456_), .Y(new_n24747_));
  OAI21X1  g22311(.A0(new_n2805_), .A1(new_n2784_), .B0(pi1093), .Y(new_n24748_));
  AOI21X1  g22312(.A0(new_n24747_), .A1(new_n24736_), .B0(new_n24748_), .Y(new_n24749_));
  OAI21X1  g22313(.A0(new_n24749_), .A1(new_n24746_), .B0(new_n8598_), .Y(new_n24750_));
  OAI22X1  g22314(.A0(new_n24750_), .A1(new_n24740_), .B0(new_n24744_), .B1(new_n24732_), .Y(new_n24751_));
  OAI21X1  g22315(.A0(new_n24751_), .A1(new_n24731_), .B0(pi0332), .Y(new_n24752_));
  AOI21X1  g22316(.A0(new_n2731_), .A1(new_n2815_), .B0(new_n2453_), .Y(new_n24753_));
  AOI22X1  g22317(.A0(new_n24745_), .A1(new_n24743_), .B0(new_n2805_), .B1(pi1093), .Y(new_n24754_));
  OAI21X1  g22318(.A0(new_n24754_), .A1(new_n24732_), .B0(new_n24750_), .Y(new_n24755_));
  OAI21X1  g22319(.A0(new_n24755_), .A1(new_n24753_), .B0(new_n2445_), .Y(new_n24756_));
  NAND3X1  g22320(.A(new_n24756_), .B(new_n24752_), .C(new_n3056_), .Y(new_n24757_));
  AOI21X1  g22321(.A0(new_n24741_), .A1(new_n2453_), .B0(new_n24731_), .Y(new_n24758_));
  NOR2X1   g22322(.A(new_n24753_), .B(new_n2806_), .Y(new_n24759_));
  MX2X1    g22323(.A(new_n24759_), .B(new_n24758_), .S0(pi0332), .Y(new_n24760_));
  AOI21X1  g22324(.A0(new_n24760_), .A1(new_n2830_), .B0(pi0210), .Y(new_n24761_));
  AOI21X1  g22325(.A0(new_n2815_), .A1(new_n2714_), .B0(new_n2453_), .Y(new_n24762_));
  OR2X1    g22326(.A(new_n24762_), .B(new_n2771_), .Y(new_n24763_));
  OAI21X1  g22327(.A0(new_n24729_), .A1(new_n2489_), .B0(new_n2540_), .Y(new_n24764_));
  NAND2X1  g22328(.A(new_n24764_), .B(new_n2848_), .Y(new_n24765_));
  NOR3X1   g22329(.A(new_n2489_), .B(pi0137), .C(pi0095), .Y(new_n24766_));
  AOI21X1  g22330(.A0(new_n24766_), .A1(new_n24734_), .B0(new_n2445_), .Y(new_n24767_));
  AOI22X1  g22331(.A0(new_n24767_), .A1(new_n24765_), .B0(new_n24763_), .B1(new_n2445_), .Y(new_n24768_));
  OAI21X1  g22332(.A0(new_n24768_), .A1(new_n2766_), .B0(pi0299), .Y(new_n24769_));
  AOI21X1  g22333(.A0(new_n24761_), .A1(new_n24757_), .B0(new_n24769_), .Y(new_n24770_));
  NAND2X1  g22334(.A(new_n24760_), .B(new_n5081_), .Y(new_n24771_));
  NAND3X1  g22335(.A(new_n24756_), .B(new_n24752_), .C(new_n5082_), .Y(new_n24772_));
  AND2X1   g22336(.A(new_n24772_), .B(new_n2973_), .Y(new_n24773_));
  OAI21X1  g22337(.A0(new_n24768_), .A1(new_n2973_), .B0(new_n2953_), .Y(new_n24774_));
  AOI21X1  g22338(.A0(new_n24773_), .A1(new_n24771_), .B0(new_n24774_), .Y(new_n24775_));
  OAI21X1  g22339(.A0(new_n24775_), .A1(new_n24770_), .B0(new_n2959_), .Y(new_n24776_));
  AOI21X1  g22340(.A0(new_n3017_), .A1(pi0039), .B0(pi0038), .Y(new_n24777_));
  OAI21X1  g22341(.A0(pi0137), .A1(new_n2996_), .B0(new_n4997_), .Y(new_n24778_));
  AOI21X1  g22342(.A0(new_n24777_), .A1(new_n24776_), .B0(new_n24778_), .Y(new_n24779_));
  OAI21X1  g22343(.A0(new_n24779_), .A1(new_n24727_), .B0(new_n3156_), .Y(new_n24780_));
  NOR4X1   g22344(.A(new_n3157_), .B(new_n3003_), .C(new_n2555_), .D(new_n2453_), .Y(new_n24781_));
  AOI21X1  g22345(.A0(new_n24781_), .A1(pi0087), .B0(pi0075), .Y(new_n24782_));
  NOR4X1   g22346(.A(new_n24726_), .B(new_n5788_), .C(new_n3074_), .D(pi0039), .Y(new_n24783_));
  OAI21X1  g22347(.A0(new_n24783_), .A1(new_n3095_), .B0(new_n3100_), .Y(new_n24784_));
  AOI21X1  g22348(.A0(new_n24782_), .A1(new_n24780_), .B0(new_n24784_), .Y(new_n24785_));
  NAND3X1  g22349(.A(new_n24781_), .B(new_n3098_), .C(pi0092), .Y(new_n24786_));
  NAND2X1  g22350(.A(new_n24786_), .B(new_n3112_), .Y(new_n24787_));
  NAND3X1  g22351(.A(new_n24781_), .B(new_n3098_), .C(new_n3100_), .Y(new_n24788_));
  AOI21X1  g22352(.A0(new_n24788_), .A1(pi0054), .B0(pi0074), .Y(new_n24789_));
  OAI21X1  g22353(.A0(new_n24787_), .A1(new_n24785_), .B0(new_n24789_), .Y(new_n24790_));
  AND2X1   g22354(.A(new_n4992_), .B(pi0074), .Y(new_n24791_));
  AOI21X1  g22355(.A0(new_n24791_), .A1(new_n24781_), .B0(pi0055), .Y(new_n24792_));
  AOI21X1  g22356(.A0(new_n24792_), .A1(new_n24790_), .B0(new_n24725_), .Y(new_n24793_));
  NOR4X1   g22357(.A(new_n3139_), .B(new_n3136_), .C(new_n3143_), .D(pi0055), .Y(new_n24794_));
  AND2X1   g22358(.A(new_n24794_), .B(new_n24781_), .Y(new_n24795_));
  OAI21X1  g22359(.A0(new_n24795_), .A1(new_n24793_), .B0(new_n3245_), .Y(new_n24796_));
  NAND3X1  g22360(.A(new_n24781_), .B(new_n3247_), .C(pi0062), .Y(new_n24797_));
  AND2X1   g22361(.A(new_n24797_), .B(new_n3246_), .Y(new_n24798_));
  NAND2X1  g22362(.A(new_n24781_), .B(new_n3247_), .Y(new_n24799_));
  OAI21X1  g22363(.A0(new_n24799_), .A1(pi0062), .B0(new_n3393_), .Y(new_n24800_));
  NAND2X1  g22364(.A(new_n24800_), .B(new_n4983_), .Y(new_n24801_));
  AOI21X1  g22365(.A0(new_n24798_), .A1(new_n24796_), .B0(new_n24801_), .Y(po0382));
  AND2X1   g22366(.A(pi0231), .B(pi0228), .Y(new_n24803_));
  OAI21X1  g22367(.A0(new_n2868_), .A1(new_n2521_), .B0(new_n5134_), .Y(new_n24804_));
  AOI21X1  g22368(.A0(new_n24804_), .A1(new_n2516_), .B0(new_n2557_), .Y(new_n24805_));
  OAI21X1  g22369(.A0(new_n24805_), .A1(new_n3194_), .B0(new_n2553_), .Y(new_n24806_));
  AOI21X1  g22370(.A0(new_n24806_), .A1(new_n2546_), .B0(new_n5023_), .Y(new_n24807_));
  OAI21X1  g22371(.A0(new_n24807_), .A1(pi0095), .B0(new_n2772_), .Y(new_n24808_));
  AND2X1   g22372(.A(new_n24808_), .B(new_n2959_), .Y(new_n24809_));
  NOR3X1   g22373(.A(new_n24809_), .B(new_n3193_), .C(pi0038), .Y(new_n24810_));
  MX2X1    g22374(.A(new_n24810_), .B(pi0231), .S0(pi0228), .Y(new_n24811_));
  AOI21X1  g22375(.A0(new_n3631_), .A1(new_n3065_), .B0(new_n24803_), .Y(new_n24812_));
  OAI21X1  g22376(.A0(new_n24812_), .A1(new_n3026_), .B0(new_n3156_), .Y(new_n24813_));
  AOI21X1  g22377(.A0(new_n24811_), .A1(new_n3026_), .B0(new_n24813_), .Y(new_n24814_));
  NOR3X1   g22378(.A(new_n24803_), .B(new_n5827_), .C(new_n3156_), .Y(new_n24815_));
  NOR3X1   g22379(.A(new_n24815_), .B(new_n24814_), .C(pi0075), .Y(new_n24816_));
  AOI21X1  g22380(.A0(new_n10121_), .A1(new_n5836_), .B0(new_n24803_), .Y(new_n24817_));
  OAI21X1  g22381(.A0(new_n24817_), .A1(new_n3095_), .B0(new_n3100_), .Y(new_n24818_));
  OR2X1    g22382(.A(new_n24803_), .B(new_n3100_), .Y(new_n24819_));
  OAI22X1  g22383(.A0(new_n24819_), .A1(new_n5844_), .B0(new_n24818_), .B1(new_n24816_), .Y(new_n24820_));
  OAI21X1  g22384(.A0(new_n24803_), .A1(new_n3112_), .B0(new_n4991_), .Y(new_n24821_));
  AOI21X1  g22385(.A0(new_n24820_), .A1(new_n3112_), .B0(new_n24821_), .Y(new_n24822_));
  OAI21X1  g22386(.A0(new_n24803_), .A1(new_n5851_), .B0(pi0074), .Y(new_n24823_));
  NAND2X1  g22387(.A(new_n24823_), .B(new_n3128_), .Y(new_n24824_));
  OR2X1    g22388(.A(new_n24803_), .B(new_n3128_), .Y(new_n24825_));
  AND2X1   g22389(.A(new_n24825_), .B(new_n3143_), .Y(new_n24826_));
  OAI21X1  g22390(.A0(new_n24824_), .A1(new_n24822_), .B0(new_n24826_), .Y(new_n24827_));
  OAI21X1  g22391(.A0(new_n24803_), .A1(new_n5855_), .B0(pi0056), .Y(new_n24828_));
  AND2X1   g22392(.A(new_n24828_), .B(new_n3245_), .Y(new_n24829_));
  NOR3X1   g22393(.A(new_n24803_), .B(new_n5828_), .C(new_n3245_), .Y(new_n24830_));
  AOI21X1  g22394(.A0(new_n24829_), .A1(new_n24827_), .B0(new_n24830_), .Y(new_n24831_));
  MX2X1    g22395(.A(new_n24831_), .B(new_n24803_), .S0(new_n3393_), .Y(po0383));
  AND2X1   g22396(.A(new_n5172_), .B(new_n2486_), .Y(new_n24833_));
  NAND4X1  g22397(.A(new_n8268_), .B(new_n8260_), .C(new_n5252_), .D(new_n2528_), .Y(new_n24834_));
  NOR4X1   g22398(.A(new_n12015_), .B(new_n2511_), .C(new_n2478_), .D(pi0047), .Y(new_n24835_));
  OR4X1    g22399(.A(new_n2473_), .B(new_n2461_), .C(pi0081), .D(new_n2567_), .Y(new_n24836_));
  OAI21X1  g22400(.A0(new_n24836_), .A1(new_n11909_), .B0(new_n2530_), .Y(new_n24837_));
  AOI21X1  g22401(.A0(new_n24835_), .A1(new_n8276_), .B0(new_n24837_), .Y(new_n24838_));
  NAND2X1  g22402(.A(new_n24838_), .B(new_n24834_), .Y(new_n24839_));
  AOI21X1  g22403(.A0(new_n24839_), .A1(new_n24833_), .B0(pi0072), .Y(new_n24840_));
  OR2X1    g22404(.A(new_n24840_), .B(new_n5191_), .Y(new_n24841_));
  AOI21X1  g22405(.A0(new_n2724_), .A1(pi1093), .B0(new_n5258_), .Y(new_n24842_));
  INVX1    g22406(.A(new_n5260_), .Y(new_n24843_));
  NAND4X1  g22407(.A(new_n9582_), .B(new_n9565_), .C(new_n5189_), .D(new_n2552_), .Y(new_n24844_));
  AOI21X1  g22408(.A0(new_n24844_), .A1(new_n24843_), .B0(new_n2756_), .Y(new_n24845_));
  AOI21X1  g22409(.A0(new_n24837_), .A1(new_n24833_), .B0(pi0072), .Y(new_n24846_));
  NOR2X1   g22410(.A(new_n8269_), .B(new_n8261_), .Y(new_n24847_));
  AND2X1   g22411(.A(new_n24833_), .B(new_n24847_), .Y(new_n24848_));
  AOI22X1  g22412(.A0(new_n24848_), .A1(new_n5939_), .B0(new_n2756_), .B1(pi0829), .Y(new_n24849_));
  AOI21X1  g22413(.A0(new_n24849_), .A1(new_n24846_), .B0(new_n5191_), .Y(new_n24850_));
  INVX1    g22414(.A(new_n24848_), .Y(new_n24851_));
  AOI21X1  g22415(.A0(new_n24851_), .A1(new_n24846_), .B0(new_n5191_), .Y(new_n24852_));
  OAI22X1  g22416(.A0(new_n24852_), .A1(new_n9767_), .B0(new_n24850_), .B1(new_n24845_), .Y(new_n24853_));
  AOI21X1  g22417(.A0(new_n24842_), .A1(new_n24841_), .B0(new_n24853_), .Y(new_n24854_));
  OAI21X1  g22418(.A0(new_n24854_), .A1(pi0039), .B0(new_n8569_), .Y(po0384));
  OR2X1    g22419(.A(new_n8535_), .B(new_n8532_), .Y(new_n24856_));
  AND2X1   g22420(.A(new_n24856_), .B(pi0039), .Y(new_n24857_));
  NOR2X1   g22421(.A(new_n6772_), .B(new_n2781_), .Y(new_n24858_));
  NAND2X1  g22422(.A(new_n7718_), .B(new_n2456_), .Y(new_n24859_));
  NOR4X1   g22423(.A(new_n24859_), .B(new_n24858_), .C(new_n8583_), .D(new_n2537_), .Y(new_n24860_));
  AOI21X1  g22424(.A0(new_n24857_), .A1(new_n5256_), .B0(new_n24860_), .Y(new_n24861_));
  OAI22X1  g22425(.A0(new_n24861_), .A1(new_n7690_), .B0(new_n3013_), .B1(pi0039), .Y(po0385));
  OAI21X1  g22426(.A0(new_n4995_), .A1(new_n2996_), .B0(new_n7686_), .Y(new_n24863_));
  NOR3X1   g22427(.A(new_n5041_), .B(new_n2829_), .C(new_n2756_), .Y(new_n24864_));
  AND2X1   g22428(.A(new_n24864_), .B(new_n12023_), .Y(new_n24865_));
  OAI21X1  g22429(.A0(new_n24864_), .A1(new_n11951_), .B0(pi1091), .Y(new_n24866_));
  OR2X1    g22430(.A(new_n24866_), .B(new_n24865_), .Y(new_n24867_));
  AOI21X1  g22431(.A0(new_n11959_), .A1(new_n6881_), .B0(pi1091), .Y(new_n24868_));
  OAI21X1  g22432(.A0(new_n12016_), .A1(new_n6881_), .B0(new_n24868_), .Y(new_n24869_));
  AND2X1   g22433(.A(new_n24869_), .B(new_n24867_), .Y(new_n24870_));
  MX2X1    g22434(.A(new_n24870_), .B(new_n3630_), .S0(pi0120), .Y(new_n24871_));
  MX2X1    g22435(.A(new_n24871_), .B(new_n13365_), .S0(new_n5052_), .Y(new_n24872_));
  NOR2X1   g22436(.A(new_n11952_), .B(new_n6269_), .Y(new_n24873_));
  AOI21X1  g22437(.A0(new_n24871_), .A1(new_n6269_), .B0(new_n24873_), .Y(new_n24874_));
  AOI21X1  g22438(.A0(new_n24874_), .A1(new_n5050_), .B0(new_n2970_), .Y(new_n24875_));
  OAI21X1  g22439(.A0(new_n24872_), .A1(new_n5050_), .B0(new_n24875_), .Y(new_n24876_));
  AOI21X1  g22440(.A0(new_n13365_), .A1(new_n2970_), .B0(pi0223), .Y(new_n24877_));
  OR2X1    g22441(.A(new_n11952_), .B(new_n5053_), .Y(new_n24878_));
  AND2X1   g22442(.A(new_n5044_), .B(pi0120), .Y(new_n24879_));
  NOR2X1   g22443(.A(new_n24879_), .B(new_n11952_), .Y(new_n24880_));
  INVX1    g22444(.A(new_n24880_), .Y(new_n24881_));
  AOI21X1  g22445(.A0(new_n24881_), .A1(new_n24878_), .B0(new_n5050_), .Y(new_n24882_));
  NOR2X1   g22446(.A(new_n24880_), .B(new_n24873_), .Y(new_n24883_));
  OAI21X1  g22447(.A0(new_n24883_), .A1(new_n5051_), .B0(pi0223), .Y(new_n24884_));
  OAI21X1  g22448(.A0(new_n24884_), .A1(new_n24882_), .B0(new_n2953_), .Y(new_n24885_));
  AOI21X1  g22449(.A0(new_n24877_), .A1(new_n24876_), .B0(new_n24885_), .Y(new_n24886_));
  AOI21X1  g22450(.A0(new_n24874_), .A1(new_n5070_), .B0(new_n10136_), .Y(new_n24887_));
  OAI21X1  g22451(.A0(new_n24872_), .A1(new_n5070_), .B0(new_n24887_), .Y(new_n24888_));
  NOR2X1   g22452(.A(new_n12179_), .B(pi0215), .Y(new_n24889_));
  AOI21X1  g22453(.A0(new_n24881_), .A1(new_n24878_), .B0(new_n5070_), .Y(new_n24890_));
  OAI21X1  g22454(.A0(new_n24883_), .A1(new_n5071_), .B0(pi0215), .Y(new_n24891_));
  OAI21X1  g22455(.A0(new_n24891_), .A1(new_n24890_), .B0(pi0299), .Y(new_n24892_));
  AOI21X1  g22456(.A0(new_n24889_), .A1(new_n24888_), .B0(new_n24892_), .Y(new_n24893_));
  OAI21X1  g22457(.A0(new_n24893_), .A1(new_n24886_), .B0(pi0039), .Y(new_n24894_));
  INVX1    g22458(.A(new_n11922_), .Y(new_n24895_));
  AND2X1   g22459(.A(pi1091), .B(pi0829), .Y(new_n24896_));
  AOI21X1  g22460(.A0(new_n24896_), .A1(new_n11938_), .B0(pi0824), .Y(new_n24897_));
  NOR2X1   g22461(.A(new_n11935_), .B(new_n5251_), .Y(new_n24898_));
  NOR3X1   g22462(.A(new_n24898_), .B(new_n24897_), .C(new_n5253_), .Y(new_n24899_));
  NOR2X1   g22463(.A(new_n24899_), .B(new_n24895_), .Y(new_n24900_));
  AOI21X1  g22464(.A0(new_n24897_), .A1(new_n24896_), .B0(new_n24898_), .Y(new_n24901_));
  OR2X1    g22465(.A(new_n5253_), .B(new_n5252_), .Y(new_n24902_));
  OAI22X1  g22466(.A0(new_n24902_), .A1(new_n24901_), .B0(new_n5253_), .B1(new_n5019_), .Y(new_n24903_));
  NOR2X1   g22467(.A(new_n5253_), .B(new_n5019_), .Y(new_n24904_));
  OAI21X1  g22468(.A0(new_n11922_), .A1(new_n5938_), .B0(new_n11920_), .Y(new_n24905_));
  AOI21X1  g22469(.A0(new_n24905_), .A1(new_n24904_), .B0(new_n2756_), .Y(new_n24906_));
  OAI21X1  g22470(.A0(new_n24903_), .A1(new_n24900_), .B0(new_n24906_), .Y(new_n24907_));
  OR4X1    g22471(.A(new_n11907_), .B(new_n5894_), .C(pi0095), .D(pi0032), .Y(new_n24908_));
  NOR4X1   g22472(.A(new_n6998_), .B(new_n2570_), .C(new_n2744_), .D(pi0091), .Y(new_n24909_));
  AOI21X1  g22473(.A0(new_n24909_), .A1(new_n11901_), .B0(pi0040), .Y(new_n24910_));
  OAI21X1  g22474(.A0(new_n24910_), .A1(new_n7750_), .B0(pi0252), .Y(new_n24911_));
  NAND3X1  g22475(.A(new_n24911_), .B(new_n11897_), .C(new_n5894_), .Y(new_n24912_));
  AND2X1   g22476(.A(new_n24912_), .B(new_n2756_), .Y(new_n24913_));
  AOI21X1  g22477(.A0(new_n24913_), .A1(new_n24908_), .B0(pi0039), .Y(new_n24914_));
  AOI21X1  g22478(.A0(new_n24914_), .A1(new_n24907_), .B0(pi0038), .Y(new_n24915_));
  AOI21X1  g22479(.A0(new_n24915_), .A1(new_n24894_), .B0(new_n24863_), .Y(po0387));
  INVX1    g22480(.A(new_n5795_), .Y(new_n24917_));
  INVX1    g22481(.A(new_n2709_), .Y(new_n24918_));
  INVX1    g22482(.A(new_n2685_), .Y(new_n24919_));
  NOR2X1   g22483(.A(new_n2678_), .B(pi0081), .Y(new_n24920_));
  NOR2X1   g22484(.A(new_n24920_), .B(new_n5162_), .Y(new_n24921_));
  OAI21X1  g22485(.A0(new_n24921_), .A1(new_n2577_), .B0(new_n24919_), .Y(new_n24922_));
  AOI21X1  g22486(.A0(new_n24922_), .A1(new_n2601_), .B0(new_n5139_), .Y(new_n24923_));
  OAI21X1  g22487(.A0(new_n24923_), .A1(new_n2745_), .B0(new_n5138_), .Y(new_n24924_));
  AOI21X1  g22488(.A0(new_n24924_), .A1(new_n2474_), .B0(new_n2598_), .Y(new_n24925_));
  OAI21X1  g22489(.A0(new_n24925_), .A1(new_n2596_), .B0(new_n2589_), .Y(new_n24926_));
  AOI21X1  g22490(.A0(new_n24926_), .A1(new_n2576_), .B0(new_n2585_), .Y(new_n24927_));
  OAI21X1  g22491(.A0(new_n24927_), .A1(new_n2697_), .B0(new_n2575_), .Y(new_n24928_));
  AOI21X1  g22492(.A0(new_n24928_), .A1(new_n2573_), .B0(new_n2572_), .Y(new_n24929_));
  OAI21X1  g22493(.A0(new_n24929_), .A1(new_n2565_), .B0(new_n2857_), .Y(new_n24930_));
  AOI21X1  g22494(.A0(new_n24930_), .A1(new_n2541_), .B0(new_n11228_), .Y(new_n24931_));
  MX2X1    g22495(.A(new_n24931_), .B(new_n24918_), .S0(pi0070), .Y(new_n24932_));
  OAI21X1  g22496(.A0(new_n24932_), .A1(pi0051), .B0(new_n2556_), .Y(new_n24933_));
  AOI21X1  g22497(.A0(new_n24933_), .A1(new_n2873_), .B0(new_n2554_), .Y(new_n24934_));
  OAI21X1  g22498(.A0(new_n7639_), .A1(pi1082), .B0(new_n2456_), .Y(new_n24935_));
  OAI22X1  g22499(.A0(new_n24935_), .A1(new_n24934_), .B0(new_n2488_), .B1(new_n2456_), .Y(new_n24936_));
  AOI21X1  g22500(.A0(new_n24936_), .A1(new_n2540_), .B0(new_n2716_), .Y(new_n24937_));
  MX2X1    g22501(.A(new_n5074_), .B(new_n5058_), .S0(new_n2953_), .Y(new_n24938_));
  OR4X1    g22502(.A(new_n5043_), .B(new_n5041_), .C(new_n2755_), .D(new_n5096_), .Y(po0950));
  NOR3X1   g22503(.A(po0950), .B(new_n24938_), .C(new_n5245_), .Y(new_n24940_));
  NOR4X1   g22504(.A(new_n24940_), .B(new_n8500_), .C(new_n7692_), .D(pi0287), .Y(new_n24941_));
  AOI21X1  g22505(.A0(new_n3074_), .A1(pi0039), .B0(new_n24941_), .Y(new_n24942_));
  OAI21X1  g22506(.A0(new_n24937_), .A1(pi0039), .B0(new_n24942_), .Y(new_n24943_));
  AOI21X1  g22507(.A0(new_n24943_), .A1(new_n2996_), .B0(new_n4998_), .Y(new_n24944_));
  NOR2X1   g22508(.A(new_n5087_), .B(pi0087), .Y(new_n24945_));
  INVX1    g22509(.A(new_n24945_), .Y(new_n24946_));
  OAI21X1  g22510(.A0(new_n24946_), .A1(new_n24944_), .B0(new_n5104_), .Y(new_n24947_));
  AOI21X1  g22511(.A0(new_n24947_), .A1(new_n3105_), .B0(new_n24917_), .Y(new_n24948_));
  MX2X1    g22512(.A(new_n24948_), .B(new_n5817_), .S0(pi0054), .Y(new_n24949_));
  OAI21X1  g22513(.A0(new_n24949_), .A1(new_n6755_), .B0(new_n11283_), .Y(new_n24950_));
  AOI21X1  g22514(.A0(new_n24950_), .A1(new_n3143_), .B0(new_n4989_), .Y(new_n24951_));
  OAI21X1  g22515(.A0(new_n24951_), .A1(pi0062), .B0(new_n11282_), .Y(new_n24952_));
  AOI21X1  g22516(.A0(new_n24952_), .A1(new_n3246_), .B0(new_n4985_), .Y(po0389));
  INVX1    g22517(.A(pi0230), .Y(new_n24954_));
  NOR2X1   g22518(.A(pi0214), .B(pi0212), .Y(new_n24955_));
  NOR2X1   g22519(.A(new_n24955_), .B(pi0211), .Y(new_n24956_));
  NOR2X1   g22520(.A(new_n24956_), .B(new_n23539_), .Y(new_n24957_));
  NOR2X1   g22521(.A(new_n24957_), .B(new_n6520_), .Y(new_n24958_));
  MX2X1    g22522(.A(new_n2439_), .B(new_n3495_), .S0(pi0211), .Y(new_n24959_));
  INVX1    g22523(.A(new_n24959_), .Y(new_n24960_));
  INVX1    g22524(.A(pi0212), .Y(new_n24961_));
  XOR2X1   g22525(.A(pi0214), .B(new_n24961_), .Y(new_n24962_));
  INVX1    g22526(.A(new_n24962_), .Y(new_n24963_));
  AND2X1   g22527(.A(pi1143), .B(new_n8548_), .Y(new_n24964_));
  AOI22X1  g22528(.A0(new_n24964_), .A1(new_n8074_), .B0(new_n24963_), .B1(new_n24960_), .Y(new_n24965_));
  OAI22X1  g22529(.A0(new_n24965_), .A1(pi0219), .B0(new_n8034_), .B1(new_n3706_), .Y(new_n24966_));
  AND2X1   g22530(.A(new_n24966_), .B(new_n24958_), .Y(new_n24967_));
  NOR2X1   g22531(.A(new_n24959_), .B(new_n2953_), .Y(new_n24968_));
  AOI21X1  g22532(.A0(pi1142), .A1(pi0199), .B0(pi0200), .Y(new_n24969_));
  OAI21X1  g22533(.A0(new_n2439_), .A1(pi0199), .B0(new_n24969_), .Y(new_n24970_));
  AOI21X1  g22534(.A0(pi1143), .A1(new_n7941_), .B0(new_n8009_), .Y(new_n24971_));
  INVX1    g22535(.A(new_n24971_), .Y(new_n24972_));
  AND2X1   g22536(.A(new_n24972_), .B(new_n24970_), .Y(new_n24973_));
  AOI21X1  g22537(.A0(new_n24972_), .A1(new_n24970_), .B0(pi0299), .Y(new_n24974_));
  OAI21X1  g22538(.A0(new_n3495_), .A1(pi0199), .B0(new_n24969_), .Y(new_n24975_));
  AOI21X1  g22539(.A0(pi1142), .A1(new_n7941_), .B0(new_n8009_), .Y(new_n24976_));
  NOR3X1   g22540(.A(new_n24976_), .B(pi0299), .C(new_n22803_), .Y(new_n24977_));
  NAND2X1  g22541(.A(new_n24977_), .B(new_n24975_), .Y(new_n24978_));
  OAI21X1  g22542(.A0(new_n24974_), .A1(pi0207), .B0(new_n24978_), .Y(new_n24979_));
  AND2X1   g22543(.A(new_n23109_), .B(pi0207), .Y(new_n24980_));
  AOI22X1  g22544(.A0(new_n24980_), .A1(new_n24973_), .B0(new_n24979_), .B1(pi0208), .Y(new_n24981_));
  NOR2X1   g22545(.A(new_n24981_), .B(pi0299), .Y(new_n24982_));
  NOR3X1   g22546(.A(new_n24982_), .B(new_n24968_), .C(pi0214), .Y(new_n24983_));
  INVX1    g22547(.A(pi0214), .Y(new_n24984_));
  MX2X1    g22548(.A(pi1143), .B(pi1142), .S0(pi0211), .Y(new_n24985_));
  AND2X1   g22549(.A(new_n24985_), .B(pi0299), .Y(new_n24986_));
  OR2X1    g22550(.A(new_n24986_), .B(new_n24984_), .Y(new_n24987_));
  OAI21X1  g22551(.A0(new_n24987_), .A1(new_n24982_), .B0(pi0212), .Y(new_n24988_));
  NOR2X1   g22552(.A(new_n24988_), .B(new_n24983_), .Y(new_n24989_));
  NOR2X1   g22553(.A(new_n24982_), .B(pi0214), .Y(new_n24990_));
  OAI21X1  g22554(.A0(new_n24982_), .A1(new_n24968_), .B0(new_n24961_), .Y(new_n24991_));
  OAI21X1  g22555(.A0(new_n24991_), .A1(new_n24990_), .B0(new_n23539_), .Y(new_n24992_));
  OR2X1    g22556(.A(new_n24992_), .B(new_n24989_), .Y(new_n24993_));
  INVX1    g22557(.A(new_n24956_), .Y(new_n24994_));
  NAND2X1  g22558(.A(new_n24982_), .B(new_n24994_), .Y(new_n24995_));
  AND2X1   g22559(.A(new_n24981_), .B(new_n2953_), .Y(new_n24996_));
  AND2X1   g22560(.A(new_n3706_), .B(pi0299), .Y(new_n24997_));
  OR4X1    g22561(.A(new_n24997_), .B(new_n24996_), .C(new_n24955_), .D(pi0211), .Y(new_n24998_));
  NAND3X1  g22562(.A(new_n24998_), .B(new_n24995_), .C(pi0219), .Y(new_n24999_));
  AND2X1   g22563(.A(new_n24999_), .B(new_n6520_), .Y(new_n25000_));
  AOI21X1  g22564(.A0(new_n25000_), .A1(new_n24993_), .B0(new_n24967_), .Y(new_n25001_));
  NAND2X1  g22565(.A(new_n25001_), .B(pi0213), .Y(new_n25002_));
  INVX1    g22566(.A(pi0213), .Y(new_n25003_));
  MX2X1    g22567(.A(pi1157), .B(pi1156), .S0(pi0211), .Y(new_n25004_));
  AOI21X1  g22568(.A0(new_n25004_), .A1(pi0214), .B0(pi0212), .Y(new_n25005_));
  MX2X1    g22569(.A(new_n12684_), .B(new_n12591_), .S0(pi0211), .Y(new_n25006_));
  MX2X1    g22570(.A(new_n12591_), .B(new_n12615_), .S0(pi0211), .Y(new_n25007_));
  MX2X1    g22571(.A(new_n25007_), .B(new_n25006_), .S0(new_n24984_), .Y(new_n25008_));
  AOI21X1  g22572(.A0(new_n25008_), .A1(pi0212), .B0(new_n25005_), .Y(new_n25009_));
  NOR2X1   g22573(.A(new_n25009_), .B(pi0219), .Y(new_n25010_));
  AND2X1   g22574(.A(pi0214), .B(new_n8548_), .Y(new_n25011_));
  AOI21X1  g22575(.A0(new_n25011_), .A1(pi1155), .B0(pi0212), .Y(new_n25012_));
  AOI21X1  g22576(.A0(pi1154), .A1(new_n8548_), .B0(pi0214), .Y(new_n25013_));
  INVX1    g22577(.A(new_n8074_), .Y(new_n25014_));
  AND2X1   g22578(.A(pi1153), .B(new_n8548_), .Y(new_n25015_));
  NOR2X1   g22579(.A(new_n25015_), .B(new_n25014_), .Y(new_n25016_));
  NOR3X1   g22580(.A(new_n25016_), .B(new_n25013_), .C(new_n25012_), .Y(new_n25017_));
  OAI21X1  g22581(.A0(new_n25017_), .A1(new_n23539_), .B0(po1038), .Y(new_n25018_));
  OAI21X1  g22582(.A0(new_n25018_), .A1(new_n25010_), .B0(new_n25003_), .Y(new_n25019_));
  INVX1    g22583(.A(new_n25019_), .Y(new_n25020_));
  AND2X1   g22584(.A(pi0299), .B(new_n23539_), .Y(new_n25021_));
  NAND2X1  g22585(.A(new_n25021_), .B(new_n25009_), .Y(new_n25022_));
  AND2X1   g22586(.A(pi0214), .B(new_n24961_), .Y(new_n25023_));
  AND2X1   g22587(.A(pi1155), .B(pi0299), .Y(new_n25024_));
  OAI21X1  g22588(.A0(new_n12494_), .A1(new_n2953_), .B0(pi0214), .Y(new_n25025_));
  AND2X1   g22589(.A(pi1154), .B(pi0299), .Y(new_n25026_));
  INVX1    g22590(.A(new_n25026_), .Y(new_n25027_));
  AOI21X1  g22591(.A0(new_n25027_), .A1(new_n24984_), .B0(new_n24961_), .Y(new_n25028_));
  AOI22X1  g22592(.A0(new_n25028_), .A1(new_n25025_), .B0(new_n25024_), .B1(new_n25023_), .Y(new_n25029_));
  AND2X1   g22593(.A(pi0219), .B(new_n8548_), .Y(new_n25030_));
  INVX1    g22594(.A(new_n25030_), .Y(new_n25031_));
  OAI21X1  g22595(.A0(new_n25031_), .A1(new_n25029_), .B0(new_n25022_), .Y(new_n25032_));
  OAI21X1  g22596(.A0(new_n25032_), .A1(new_n24982_), .B0(new_n6520_), .Y(new_n25033_));
  AOI21X1  g22597(.A0(new_n25033_), .A1(new_n25020_), .B0(new_n23244_), .Y(new_n25034_));
  NAND2X1  g22598(.A(new_n25034_), .B(new_n25002_), .Y(new_n25035_));
  NOR4X1   g22599(.A(new_n12591_), .B(pi0299), .C(pi0200), .D(new_n7941_), .Y(new_n25036_));
  NOR2X1   g22600(.A(new_n25036_), .B(pi1156), .Y(new_n25037_));
  NOR2X1   g22601(.A(pi1155), .B(pi0200), .Y(new_n25038_));
  XOR2X1   g22602(.A(pi0200), .B(pi0199), .Y(new_n25039_));
  AND2X1   g22603(.A(new_n25039_), .B(new_n2953_), .Y(new_n25040_));
  INVX1    g22604(.A(new_n25040_), .Y(new_n25041_));
  NOR4X1   g22605(.A(new_n25041_), .B(new_n25038_), .C(new_n25037_), .D(new_n22803_), .Y(new_n25042_));
  INVX1    g22606(.A(new_n25042_), .Y(new_n25043_));
  AOI21X1  g22607(.A0(pi0200), .A1(pi0199), .B0(pi0299), .Y(new_n25044_));
  NOR2X1   g22608(.A(new_n25044_), .B(new_n12494_), .Y(new_n25045_));
  NOR2X1   g22609(.A(new_n25045_), .B(new_n12615_), .Y(new_n25046_));
  NOR4X1   g22610(.A(new_n12591_), .B(pi0299), .C(pi0200), .D(pi0199), .Y(new_n25047_));
  INVX1    g22611(.A(new_n25039_), .Y(new_n25048_));
  NOR2X1   g22612(.A(new_n8502_), .B(pi1153), .Y(new_n25049_));
  NOR3X1   g22613(.A(new_n25049_), .B(new_n25048_), .C(new_n12615_), .Y(new_n25050_));
  NOR2X1   g22614(.A(new_n25050_), .B(new_n25047_), .Y(new_n25051_));
  INVX1    g22615(.A(new_n25051_), .Y(new_n25052_));
  NOR2X1   g22616(.A(pi0299), .B(pi0200), .Y(new_n25053_));
  INVX1    g22617(.A(new_n25053_), .Y(new_n25054_));
  AND2X1   g22618(.A(new_n12494_), .B(pi0199), .Y(new_n25055_));
  OAI21X1  g22619(.A0(pi1155), .A1(pi0199), .B0(new_n12615_), .Y(new_n25056_));
  NOR3X1   g22620(.A(new_n25056_), .B(new_n25055_), .C(new_n25054_), .Y(new_n25057_));
  AOI21X1  g22621(.A0(new_n25052_), .A1(new_n25046_), .B0(new_n25057_), .Y(new_n25058_));
  NOR4X1   g22622(.A(new_n12591_), .B(pi0299), .C(new_n8009_), .D(pi0199), .Y(new_n25059_));
  NOR2X1   g22623(.A(new_n25059_), .B(pi1154), .Y(new_n25060_));
  INVX1    g22624(.A(new_n25060_), .Y(new_n25061_));
  AOI21X1  g22625(.A0(pi1155), .A1(new_n7941_), .B0(new_n8009_), .Y(new_n25062_));
  NOR3X1   g22626(.A(new_n25062_), .B(new_n8130_), .C(pi0299), .Y(new_n25063_));
  AND2X1   g22627(.A(new_n12591_), .B(pi0200), .Y(new_n25064_));
  NOR3X1   g22628(.A(new_n25064_), .B(new_n8503_), .C(new_n12684_), .Y(new_n25065_));
  AOI21X1  g22629(.A0(new_n25063_), .A1(new_n25061_), .B0(new_n25065_), .Y(new_n25066_));
  MX2X1    g22630(.A(new_n25066_), .B(new_n25058_), .S0(pi0207), .Y(new_n25067_));
  MX2X1    g22631(.A(new_n25067_), .B(new_n25043_), .S0(new_n23109_), .Y(new_n25068_));
  INVX1    g22632(.A(new_n25044_), .Y(new_n25069_));
  AND2X1   g22633(.A(new_n12591_), .B(pi0199), .Y(new_n25070_));
  NOR3X1   g22634(.A(new_n25070_), .B(new_n25069_), .C(new_n12684_), .Y(new_n25071_));
  NOR3X1   g22635(.A(new_n25070_), .B(new_n25054_), .C(pi1156), .Y(new_n25072_));
  OR2X1    g22636(.A(new_n25072_), .B(new_n25071_), .Y(new_n25073_));
  AND2X1   g22637(.A(new_n25073_), .B(pi0207), .Y(new_n25074_));
  INVX1    g22638(.A(new_n25074_), .Y(new_n25075_));
  MX2X1    g22639(.A(new_n25075_), .B(new_n25067_), .S0(pi0208), .Y(new_n25076_));
  MX2X1    g22640(.A(new_n25076_), .B(new_n25068_), .S0(new_n12706_), .Y(new_n25077_));
  AND2X1   g22641(.A(new_n25077_), .B(pi0211), .Y(new_n25078_));
  AOI21X1  g22642(.A0(new_n25077_), .A1(new_n24984_), .B0(pi0212), .Y(new_n25079_));
  INVX1    g22643(.A(new_n25011_), .Y(new_n25080_));
  NOR4X1   g22644(.A(pi1155), .B(pi0299), .C(pi0200), .D(new_n7941_), .Y(new_n25081_));
  AND2X1   g22645(.A(new_n2953_), .B(pi0200), .Y(new_n25082_));
  MX2X1    g22646(.A(new_n25082_), .B(new_n8131_), .S0(new_n12494_), .Y(new_n25083_));
  INVX1    g22647(.A(new_n25083_), .Y(new_n25084_));
  AOI22X1  g22648(.A0(new_n25084_), .A1(pi1155), .B0(new_n25081_), .B1(pi1153), .Y(new_n25085_));
  AND2X1   g22649(.A(new_n2953_), .B(pi0199), .Y(new_n25086_));
  INVX1    g22650(.A(new_n25086_), .Y(new_n25087_));
  NOR3X1   g22651(.A(new_n25055_), .B(new_n25048_), .C(pi0299), .Y(new_n25088_));
  AOI21X1  g22652(.A0(new_n25087_), .A1(pi1155), .B0(new_n25088_), .Y(new_n25089_));
  MX2X1    g22653(.A(new_n25089_), .B(new_n25085_), .S0(new_n12615_), .Y(new_n25090_));
  AND2X1   g22654(.A(new_n25090_), .B(pi0207), .Y(new_n25091_));
  INVX1    g22655(.A(new_n25066_), .Y(new_n25092_));
  NOR3X1   g22656(.A(new_n25092_), .B(new_n25024_), .C(pi0207), .Y(new_n25093_));
  NOR3X1   g22657(.A(new_n25093_), .B(new_n25091_), .C(new_n23109_), .Y(new_n25094_));
  OAI21X1  g22658(.A0(new_n25082_), .A1(new_n12591_), .B0(new_n8503_), .Y(new_n25095_));
  AOI21X1  g22659(.A0(new_n8009_), .A1(pi0199), .B0(pi0299), .Y(new_n25096_));
  OR2X1    g22660(.A(new_n25096_), .B(pi1155), .Y(new_n25097_));
  AOI21X1  g22661(.A0(new_n2953_), .A1(pi0200), .B0(pi1156), .Y(new_n25098_));
  AOI22X1  g22662(.A0(new_n25098_), .A1(new_n25097_), .B0(new_n25095_), .B1(pi1156), .Y(new_n25099_));
  INVX1    g22663(.A(new_n25024_), .Y(new_n25100_));
  AOI21X1  g22664(.A0(new_n25100_), .A1(new_n22803_), .B0(pi0208), .Y(new_n25101_));
  NAND2X1  g22665(.A(new_n25101_), .B(pi1157), .Y(new_n25102_));
  AOI21X1  g22666(.A0(new_n25099_), .A1(pi0207), .B0(new_n25102_), .Y(new_n25103_));
  INVX1    g22667(.A(new_n25101_), .Y(new_n25104_));
  NOR3X1   g22668(.A(new_n12591_), .B(pi0200), .C(new_n7941_), .Y(new_n25105_));
  NOR3X1   g22669(.A(new_n25105_), .B(pi1156), .C(pi0299), .Y(new_n25106_));
  NOR2X1   g22670(.A(new_n25039_), .B(pi0299), .Y(new_n25107_));
  NOR2X1   g22671(.A(new_n8502_), .B(pi1155), .Y(new_n25108_));
  NOR4X1   g22672(.A(new_n25108_), .B(new_n25107_), .C(new_n25106_), .D(new_n25104_), .Y(new_n25109_));
  OR4X1    g22673(.A(new_n25109_), .B(new_n25103_), .C(new_n25094_), .D(new_n25080_), .Y(new_n25110_));
  MX2X1    g22674(.A(new_n25107_), .B(new_n25096_), .S0(new_n12591_), .Y(new_n25111_));
  OAI21X1  g22675(.A0(new_n25111_), .A1(new_n12615_), .B0(new_n25066_), .Y(new_n25112_));
  AOI21X1  g22676(.A0(new_n25089_), .A1(new_n2953_), .B0(new_n12615_), .Y(new_n25113_));
  OR2X1    g22677(.A(new_n25113_), .B(new_n25057_), .Y(new_n25114_));
  MX2X1    g22678(.A(new_n25114_), .B(new_n25112_), .S0(new_n22803_), .Y(new_n25115_));
  AND2X1   g22679(.A(new_n25115_), .B(pi0208), .Y(new_n25116_));
  MX2X1    g22680(.A(new_n25082_), .B(new_n8131_), .S0(new_n12591_), .Y(new_n25117_));
  AOI21X1  g22681(.A0(pi1155), .A1(new_n8009_), .B0(new_n25087_), .Y(new_n25118_));
  MX2X1    g22682(.A(new_n25118_), .B(new_n25117_), .S0(new_n12684_), .Y(new_n25119_));
  NOR2X1   g22683(.A(pi0299), .B(pi0207), .Y(new_n25120_));
  NOR2X1   g22684(.A(new_n25120_), .B(pi0208), .Y(new_n25121_));
  INVX1    g22685(.A(new_n25121_), .Y(new_n25122_));
  AOI21X1  g22686(.A0(new_n25119_), .A1(pi0207), .B0(new_n25122_), .Y(new_n25123_));
  INVX1    g22687(.A(new_n25123_), .Y(new_n25124_));
  OAI21X1  g22688(.A0(pi1154), .A1(new_n2953_), .B0(pi1157), .Y(new_n25125_));
  AOI21X1  g22689(.A0(new_n25043_), .A1(new_n25027_), .B0(pi0208), .Y(new_n25126_));
  NAND2X1  g22690(.A(new_n25126_), .B(new_n12706_), .Y(new_n25127_));
  OAI21X1  g22691(.A0(new_n25125_), .A1(new_n25124_), .B0(new_n25127_), .Y(new_n25128_));
  OR4X1    g22692(.A(new_n25128_), .B(new_n25116_), .C(pi0214), .D(pi0211), .Y(new_n25129_));
  INVX1    g22693(.A(new_n25096_), .Y(new_n25130_));
  AOI21X1  g22694(.A0(new_n25130_), .A1(pi1153), .B0(new_n25052_), .Y(new_n25131_));
  NOR2X1   g22695(.A(new_n25131_), .B(new_n22803_), .Y(new_n25132_));
  MX2X1    g22696(.A(new_n25086_), .B(new_n8131_), .S0(new_n12591_), .Y(new_n25133_));
  OAI22X1  g22697(.A0(new_n25133_), .A1(new_n12684_), .B0(new_n25111_), .B1(new_n12615_), .Y(new_n25134_));
  AOI21X1  g22698(.A0(pi0200), .A1(new_n7941_), .B0(pi0299), .Y(new_n25135_));
  MX2X1    g22699(.A(new_n25135_), .B(new_n2953_), .S0(new_n12591_), .Y(new_n25136_));
  INVX1    g22700(.A(new_n25136_), .Y(new_n25137_));
  NOR2X1   g22701(.A(new_n25137_), .B(new_n25134_), .Y(new_n25138_));
  AND2X1   g22702(.A(new_n12494_), .B(pi0299), .Y(new_n25139_));
  NOR3X1   g22703(.A(new_n25139_), .B(new_n25138_), .C(pi0207), .Y(new_n25140_));
  OAI21X1  g22704(.A0(new_n25140_), .A1(new_n25132_), .B0(pi0208), .Y(new_n25141_));
  INVX1    g22705(.A(new_n25037_), .Y(new_n25142_));
  AND2X1   g22706(.A(pi0200), .B(new_n7941_), .Y(new_n25143_));
  OR4X1    g22707(.A(new_n25105_), .B(new_n25143_), .C(new_n12684_), .D(pi0299), .Y(new_n25144_));
  AND2X1   g22708(.A(new_n25144_), .B(new_n25142_), .Y(new_n25145_));
  AOI21X1  g22709(.A0(new_n25145_), .A1(pi0207), .B0(pi0299), .Y(new_n25146_));
  OR2X1    g22710(.A(new_n25146_), .B(pi0208), .Y(new_n25147_));
  AND2X1   g22711(.A(new_n25147_), .B(new_n12706_), .Y(new_n25148_));
  NOR2X1   g22712(.A(new_n25123_), .B(new_n12706_), .Y(new_n25149_));
  NOR3X1   g22713(.A(new_n25149_), .B(new_n25148_), .C(new_n25139_), .Y(new_n25150_));
  NOR2X1   g22714(.A(new_n25150_), .B(new_n25080_), .Y(new_n25151_));
  AOI21X1  g22715(.A0(new_n25151_), .A1(new_n25141_), .B0(new_n24961_), .Y(new_n25152_));
  AOI22X1  g22716(.A0(new_n25152_), .A1(new_n25129_), .B0(new_n25110_), .B1(new_n25079_), .Y(new_n25153_));
  OAI21X1  g22717(.A0(new_n25153_), .A1(new_n25078_), .B0(pi0219), .Y(new_n25154_));
  NAND2X1  g22718(.A(new_n25068_), .B(new_n12706_), .Y(new_n25155_));
  AND2X1   g22719(.A(new_n12591_), .B(pi0299), .Y(new_n25156_));
  NOR2X1   g22720(.A(new_n25135_), .B(new_n12591_), .Y(new_n25157_));
  OR4X1    g22721(.A(new_n25157_), .B(new_n25156_), .C(new_n25134_), .D(pi0207), .Y(new_n25158_));
  AND2X1   g22722(.A(new_n2953_), .B(pi0207), .Y(new_n25159_));
  AOI21X1  g22723(.A0(new_n25131_), .A1(new_n25159_), .B0(new_n23109_), .Y(new_n25160_));
  NAND2X1  g22724(.A(new_n25160_), .B(new_n25158_), .Y(new_n25161_));
  AOI21X1  g22725(.A0(new_n25161_), .A1(new_n25149_), .B0(pi0211), .Y(new_n25162_));
  AND2X1   g22726(.A(new_n25162_), .B(new_n25155_), .Y(new_n25163_));
  NOR2X1   g22727(.A(new_n25133_), .B(new_n12684_), .Y(new_n25164_));
  AOI21X1  g22728(.A0(new_n25063_), .A1(new_n25061_), .B0(new_n25164_), .Y(new_n25165_));
  AND2X1   g22729(.A(pi1156), .B(pi0299), .Y(new_n25166_));
  INVX1    g22730(.A(new_n25166_), .Y(new_n25167_));
  MX2X1    g22731(.A(new_n25167_), .B(new_n25165_), .S0(new_n22803_), .Y(new_n25168_));
  OAI21X1  g22732(.A0(new_n25058_), .A1(new_n22803_), .B0(new_n25168_), .Y(new_n25169_));
  AND2X1   g22733(.A(new_n25169_), .B(pi0208), .Y(new_n25170_));
  NOR3X1   g22734(.A(new_n25146_), .B(new_n25037_), .C(pi0208), .Y(new_n25171_));
  AND2X1   g22735(.A(pi1157), .B(new_n23109_), .Y(new_n25172_));
  INVX1    g22736(.A(new_n25172_), .Y(new_n25173_));
  AOI21X1  g22737(.A0(new_n25167_), .A1(new_n25075_), .B0(new_n25173_), .Y(new_n25174_));
  NOR3X1   g22738(.A(new_n25174_), .B(new_n25171_), .C(new_n25170_), .Y(new_n25175_));
  OAI21X1  g22739(.A0(new_n25175_), .A1(new_n8548_), .B0(pi0214), .Y(new_n25176_));
  OAI21X1  g22740(.A0(new_n25176_), .A1(new_n25163_), .B0(new_n25079_), .Y(new_n25177_));
  OAI21X1  g22741(.A0(new_n25128_), .A1(new_n25116_), .B0(new_n8033_), .Y(new_n25178_));
  OR2X1    g22742(.A(new_n25109_), .B(new_n25103_), .Y(new_n25179_));
  XOR2X1   g22743(.A(pi0214), .B(pi0211), .Y(new_n25180_));
  OAI21X1  g22744(.A0(new_n25179_), .A1(new_n25094_), .B0(new_n25180_), .Y(new_n25181_));
  NOR2X1   g22745(.A(pi0214), .B(pi0211), .Y(new_n25182_));
  INVX1    g22746(.A(new_n25182_), .Y(new_n25183_));
  OR2X1    g22747(.A(new_n25175_), .B(new_n25183_), .Y(new_n25184_));
  NAND3X1  g22748(.A(new_n25184_), .B(new_n25181_), .C(new_n25178_), .Y(new_n25185_));
  AOI21X1  g22749(.A0(new_n25185_), .A1(pi0212), .B0(pi0219), .Y(new_n25186_));
  AOI21X1  g22750(.A0(new_n25186_), .A1(new_n25177_), .B0(po1038), .Y(new_n25187_));
  AOI21X1  g22751(.A0(new_n25187_), .A1(new_n25154_), .B0(new_n25019_), .Y(new_n25188_));
  AND2X1   g22752(.A(pi1143), .B(pi0299), .Y(new_n25189_));
  INVX1    g22753(.A(new_n25189_), .Y(new_n25190_));
  NAND3X1  g22754(.A(new_n25190_), .B(new_n25058_), .C(pi0207), .Y(new_n25191_));
  OAI21X1  g22755(.A0(new_n25039_), .A1(pi0299), .B0(pi1155), .Y(new_n25192_));
  AND2X1   g22756(.A(new_n3495_), .B(pi0299), .Y(new_n25193_));
  NOR2X1   g22757(.A(new_n25193_), .B(new_n25192_), .Y(new_n25194_));
  AND2X1   g22758(.A(new_n25189_), .B(new_n12591_), .Y(new_n25195_));
  NOR4X1   g22759(.A(new_n25195_), .B(new_n25194_), .C(new_n25081_), .D(new_n12615_), .Y(new_n25196_));
  INVX1    g22760(.A(new_n25196_), .Y(new_n25197_));
  AOI21X1  g22761(.A0(new_n25190_), .A1(new_n25060_), .B0(pi1156), .Y(new_n25198_));
  OAI21X1  g22762(.A0(new_n25193_), .A1(new_n25133_), .B0(new_n12615_), .Y(new_n25199_));
  OAI21X1  g22763(.A0(new_n25062_), .A1(pi0299), .B0(pi1154), .Y(new_n25200_));
  INVX1    g22764(.A(new_n25200_), .Y(new_n25201_));
  AOI21X1  g22765(.A0(new_n25201_), .A1(new_n25190_), .B0(new_n12684_), .Y(new_n25202_));
  AOI22X1  g22766(.A0(new_n25202_), .A1(new_n25199_), .B0(new_n25198_), .B1(new_n25197_), .Y(new_n25203_));
  AOI21X1  g22767(.A0(new_n25203_), .A1(new_n22803_), .B0(new_n23109_), .Y(new_n25204_));
  AND2X1   g22768(.A(new_n25204_), .B(new_n25191_), .Y(new_n25205_));
  OR2X1    g22769(.A(new_n25147_), .B(pi1157), .Y(new_n25206_));
  OAI21X1  g22770(.A0(pi1155), .A1(new_n7941_), .B0(pi1156), .Y(new_n25207_));
  OAI21X1  g22771(.A0(new_n25207_), .A1(new_n25069_), .B0(new_n25117_), .Y(new_n25208_));
  AOI21X1  g22772(.A0(new_n3495_), .A1(pi0299), .B0(new_n22803_), .Y(new_n25209_));
  AOI21X1  g22773(.A0(new_n25209_), .A1(new_n25208_), .B0(new_n25189_), .Y(new_n25210_));
  OAI22X1  g22774(.A0(new_n25210_), .A1(new_n25173_), .B0(new_n25206_), .B1(new_n25193_), .Y(new_n25211_));
  OR4X1    g22775(.A(new_n25211_), .B(new_n25205_), .C(new_n25014_), .D(pi0211), .Y(new_n25212_));
  OAI21X1  g22776(.A0(new_n25211_), .A1(new_n25205_), .B0(pi0211), .Y(new_n25213_));
  AND2X1   g22777(.A(new_n25058_), .B(pi0207), .Y(new_n25214_));
  AND2X1   g22778(.A(pi1144), .B(pi0299), .Y(new_n25215_));
  INVX1    g22779(.A(new_n25215_), .Y(new_n25216_));
  AND2X1   g22780(.A(new_n2439_), .B(pi0299), .Y(new_n25217_));
  NOR2X1   g22781(.A(new_n25217_), .B(new_n25192_), .Y(new_n25218_));
  AND2X1   g22782(.A(new_n25215_), .B(new_n12591_), .Y(new_n25219_));
  NOR4X1   g22783(.A(new_n25219_), .B(new_n25218_), .C(new_n25081_), .D(new_n12615_), .Y(new_n25220_));
  OAI21X1  g22784(.A0(new_n25215_), .A1(new_n25061_), .B0(new_n12684_), .Y(new_n25221_));
  OR2X1    g22785(.A(new_n25217_), .B(new_n25133_), .Y(new_n25222_));
  AND2X1   g22786(.A(new_n25222_), .B(new_n12615_), .Y(new_n25223_));
  OAI21X1  g22787(.A0(new_n25215_), .A1(new_n25200_), .B0(pi1156), .Y(new_n25224_));
  OAI22X1  g22788(.A0(new_n25224_), .A1(new_n25223_), .B0(new_n25221_), .B1(new_n25220_), .Y(new_n25225_));
  OAI21X1  g22789(.A0(new_n25225_), .A1(pi0207), .B0(pi0208), .Y(new_n25226_));
  AOI21X1  g22790(.A0(new_n25216_), .A1(new_n25214_), .B0(new_n25226_), .Y(new_n25227_));
  AOI21X1  g22791(.A0(new_n2439_), .A1(pi0299), .B0(new_n22803_), .Y(new_n25228_));
  AOI21X1  g22792(.A0(new_n25228_), .A1(new_n25208_), .B0(new_n25215_), .Y(new_n25229_));
  OAI22X1  g22793(.A0(new_n25229_), .A1(new_n25173_), .B0(new_n25217_), .B1(new_n25206_), .Y(new_n25230_));
  OAI21X1  g22794(.A0(new_n25230_), .A1(new_n25227_), .B0(new_n8548_), .Y(new_n25231_));
  XOR2X1   g22795(.A(pi0214), .B(pi0212), .Y(new_n25232_));
  NAND3X1  g22796(.A(new_n25232_), .B(new_n25231_), .C(new_n25213_), .Y(new_n25233_));
  AOI21X1  g22797(.A0(new_n25233_), .A1(new_n25212_), .B0(pi0219), .Y(new_n25234_));
  OAI22X1  g22798(.A0(new_n23539_), .A1(new_n8548_), .B0(pi0214), .B1(pi0212), .Y(new_n25235_));
  AND2X1   g22799(.A(new_n25235_), .B(new_n25077_), .Y(new_n25236_));
  NOR3X1   g22800(.A(new_n25149_), .B(new_n25148_), .C(new_n24997_), .Y(new_n25237_));
  INVX1    g22801(.A(new_n25090_), .Y(new_n25238_));
  OAI21X1  g22802(.A0(new_n3706_), .A1(new_n2953_), .B0(pi0207), .Y(new_n25239_));
  AOI21X1  g22803(.A0(new_n25238_), .A1(new_n2953_), .B0(new_n25239_), .Y(new_n25240_));
  INVX1    g22804(.A(new_n24997_), .Y(new_n25241_));
  AOI21X1  g22805(.A0(pi1142), .A1(pi0299), .B0(new_n25059_), .Y(new_n25242_));
  OR2X1    g22806(.A(pi1156), .B(pi1154), .Y(new_n25243_));
  OAI21X1  g22807(.A0(new_n25243_), .A1(new_n25242_), .B0(new_n22803_), .Y(new_n25244_));
  AOI21X1  g22808(.A0(new_n25134_), .A1(new_n25241_), .B0(new_n25244_), .Y(new_n25245_));
  NOR3X1   g22809(.A(new_n25245_), .B(new_n25240_), .C(new_n23109_), .Y(new_n25246_));
  NOR4X1   g22810(.A(new_n25246_), .B(new_n25237_), .C(new_n25235_), .D(new_n8034_), .Y(new_n25247_));
  NOR4X1   g22811(.A(new_n25247_), .B(new_n25236_), .C(new_n25234_), .D(po1038), .Y(new_n25248_));
  OR2X1    g22812(.A(new_n24967_), .B(new_n25003_), .Y(new_n25249_));
  OAI21X1  g22813(.A0(new_n25249_), .A1(new_n25248_), .B0(new_n23244_), .Y(new_n25250_));
  OAI21X1  g22814(.A0(new_n25250_), .A1(new_n25188_), .B0(new_n25035_), .Y(new_n25251_));
  MX2X1    g22815(.A(new_n25251_), .B(new_n22718_), .S0(new_n24954_), .Y(po0390));
  NOR2X1   g22816(.A(new_n24955_), .B(pi0219), .Y(new_n25253_));
  MX2X1    g22817(.A(new_n12615_), .B(new_n12494_), .S0(pi0211), .Y(new_n25254_));
  INVX1    g22818(.A(new_n25254_), .Y(new_n25255_));
  OAI21X1  g22819(.A0(new_n25255_), .A1(new_n8074_), .B0(new_n25253_), .Y(new_n25256_));
  NOR2X1   g22820(.A(new_n25256_), .B(new_n25016_), .Y(new_n25257_));
  AOI21X1  g22821(.A0(new_n25257_), .A1(po1038), .B0(pi1152), .Y(new_n25258_));
  XOR2X1   g22822(.A(pi0208), .B(pi0207), .Y(new_n25259_));
  AOI21X1  g22823(.A0(new_n25038_), .A1(new_n7941_), .B0(new_n25069_), .Y(new_n25260_));
  OAI21X1  g22824(.A0(new_n25047_), .A1(pi1154), .B0(new_n25260_), .Y(new_n25261_));
  NOR2X1   g22825(.A(new_n25261_), .B(new_n22803_), .Y(new_n25262_));
  OAI22X1  g22826(.A0(new_n25262_), .A1(new_n25259_), .B0(new_n25092_), .B1(new_n7896_), .Y(new_n25263_));
  INVX1    g22827(.A(new_n25263_), .Y(new_n25264_));
  OAI21X1  g22828(.A0(new_n25264_), .A1(pi0214), .B0(new_n24961_), .Y(new_n25265_));
  MX2X1    g22829(.A(new_n25112_), .B(new_n25026_), .S0(new_n22803_), .Y(new_n25266_));
  AND2X1   g22830(.A(new_n25266_), .B(new_n23109_), .Y(new_n25267_));
  AND2X1   g22831(.A(pi0200), .B(pi0199), .Y(new_n25268_));
  AOI21X1  g22832(.A0(new_n8130_), .A1(new_n12591_), .B0(new_n25268_), .Y(new_n25269_));
  OAI22X1  g22833(.A0(new_n25269_), .A1(pi0299), .B0(new_n25047_), .B1(pi1154), .Y(new_n25270_));
  INVX1    g22834(.A(new_n25270_), .Y(new_n25271_));
  MX2X1    g22835(.A(new_n25271_), .B(new_n25112_), .S0(new_n22803_), .Y(new_n25272_));
  AOI21X1  g22836(.A0(new_n25272_), .A1(pi0208), .B0(new_n25267_), .Y(new_n25273_));
  NOR3X1   g22837(.A(new_n25137_), .B(new_n25134_), .C(new_n22803_), .Y(new_n25274_));
  INVX1    g22838(.A(new_n25274_), .Y(new_n25275_));
  AOI21X1  g22839(.A0(new_n25270_), .A1(new_n25159_), .B0(new_n23109_), .Y(new_n25276_));
  AOI22X1  g22840(.A0(new_n25276_), .A1(new_n25158_), .B0(new_n25275_), .B1(new_n25121_), .Y(new_n25277_));
  OR2X1    g22841(.A(new_n25277_), .B(new_n25139_), .Y(new_n25278_));
  MX2X1    g22842(.A(new_n25278_), .B(new_n25273_), .S0(new_n8548_), .Y(new_n25279_));
  AOI21X1  g22843(.A0(new_n25279_), .A1(pi0214), .B0(new_n25265_), .Y(new_n25280_));
  OR2X1    g22844(.A(new_n25280_), .B(pi0219), .Y(new_n25281_));
  OAI21X1  g22845(.A0(new_n25277_), .A1(new_n25139_), .B0(new_n8548_), .Y(new_n25282_));
  NAND2X1  g22846(.A(new_n25282_), .B(pi0214), .Y(new_n25283_));
  AND2X1   g22847(.A(new_n25263_), .B(pi0211), .Y(new_n25284_));
  OAI22X1  g22848(.A0(new_n25284_), .A1(new_n25283_), .B0(new_n25279_), .B1(pi0214), .Y(new_n25285_));
  AOI21X1  g22849(.A0(new_n25285_), .A1(pi0212), .B0(new_n25281_), .Y(new_n25286_));
  OAI21X1  g22850(.A0(new_n25264_), .A1(new_n23539_), .B0(new_n6520_), .Y(new_n25287_));
  OAI21X1  g22851(.A0(new_n25287_), .A1(new_n25286_), .B0(new_n25258_), .Y(new_n25288_));
  INVX1    g22852(.A(pi1152), .Y(new_n25289_));
  NOR2X1   g22853(.A(new_n25013_), .B(new_n25011_), .Y(new_n25290_));
  AOI21X1  g22854(.A0(new_n25183_), .A1(pi1153), .B0(new_n25290_), .Y(new_n25291_));
  AOI21X1  g22855(.A0(new_n25255_), .A1(new_n25023_), .B0(pi0219), .Y(new_n25292_));
  OAI21X1  g22856(.A0(new_n25291_), .A1(new_n24961_), .B0(new_n25292_), .Y(new_n25293_));
  AOI21X1  g22857(.A0(new_n25293_), .A1(new_n24958_), .B0(new_n25289_), .Y(new_n25294_));
  OAI22X1  g22858(.A0(new_n25283_), .A1(new_n25277_), .B0(new_n25279_), .B1(pi0214), .Y(new_n25295_));
  AND2X1   g22859(.A(new_n25295_), .B(pi0212), .Y(new_n25296_));
  AOI21X1  g22860(.A0(new_n25264_), .A1(new_n24994_), .B0(new_n23539_), .Y(new_n25297_));
  OR2X1    g22861(.A(new_n25277_), .B(new_n24994_), .Y(new_n25298_));
  AOI21X1  g22862(.A0(new_n25298_), .A1(new_n25297_), .B0(po1038), .Y(new_n25299_));
  OAI21X1  g22863(.A0(new_n25296_), .A1(new_n25281_), .B0(new_n25299_), .Y(new_n25300_));
  AOI21X1  g22864(.A0(new_n25300_), .A1(new_n25294_), .B0(pi0213), .Y(new_n25301_));
  OAI21X1  g22865(.A0(new_n25165_), .A1(new_n22803_), .B0(new_n25167_), .Y(new_n25302_));
  AND2X1   g22866(.A(new_n25302_), .B(new_n23109_), .Y(new_n25303_));
  OAI21X1  g22867(.A0(new_n25261_), .A1(new_n22803_), .B0(new_n25168_), .Y(new_n25304_));
  AOI21X1  g22868(.A0(new_n25304_), .A1(pi0208), .B0(new_n25303_), .Y(new_n25305_));
  INVX1    g22869(.A(new_n25093_), .Y(new_n25306_));
  AOI21X1  g22870(.A0(new_n25066_), .A1(new_n25100_), .B0(new_n25104_), .Y(new_n25307_));
  NOR2X1   g22871(.A(new_n25024_), .B(new_n22803_), .Y(new_n25308_));
  AOI21X1  g22872(.A0(new_n25308_), .A1(new_n25261_), .B0(new_n23109_), .Y(new_n25309_));
  AOI21X1  g22873(.A0(new_n25309_), .A1(new_n25306_), .B0(new_n25307_), .Y(new_n25310_));
  MX2X1    g22874(.A(new_n25310_), .B(new_n25305_), .S0(new_n8548_), .Y(new_n25311_));
  AOI21X1  g22875(.A0(new_n25311_), .A1(pi0214), .B0(new_n25265_), .Y(new_n25312_));
  NOR2X1   g22876(.A(new_n25273_), .B(new_n8548_), .Y(new_n25313_));
  OAI21X1  g22877(.A0(new_n25310_), .A1(pi0211), .B0(pi0214), .Y(new_n25314_));
  OAI21X1  g22878(.A0(new_n25314_), .A1(new_n25313_), .B0(pi0212), .Y(new_n25315_));
  AOI21X1  g22879(.A0(new_n25311_), .A1(new_n24984_), .B0(new_n25315_), .Y(new_n25316_));
  NOR3X1   g22880(.A(new_n25316_), .B(new_n25312_), .C(pi0219), .Y(new_n25317_));
  INVX1    g22881(.A(new_n25297_), .Y(new_n25318_));
  NOR3X1   g22882(.A(new_n25273_), .B(new_n24955_), .C(pi0211), .Y(new_n25319_));
  OAI21X1  g22883(.A0(new_n25319_), .A1(new_n25318_), .B0(new_n23355_), .Y(new_n25320_));
  OAI21X1  g22884(.A0(new_n25320_), .A1(new_n25317_), .B0(pi0209), .Y(new_n25321_));
  AOI21X1  g22885(.A0(new_n25301_), .A1(new_n25288_), .B0(new_n25321_), .Y(new_n25322_));
  INVX1    g22886(.A(new_n24955_), .Y(new_n25323_));
  NOR4X1   g22887(.A(new_n12494_), .B(pi0299), .C(new_n8009_), .D(pi0199), .Y(new_n25324_));
  NOR2X1   g22888(.A(new_n25324_), .B(pi1154), .Y(new_n25325_));
  INVX1    g22889(.A(new_n25325_), .Y(new_n25326_));
  AND2X1   g22890(.A(pi1153), .B(new_n7941_), .Y(new_n25327_));
  NOR4X1   g22891(.A(new_n25327_), .B(new_n12615_), .C(pi0299), .D(new_n8009_), .Y(new_n25328_));
  INVX1    g22892(.A(new_n25328_), .Y(new_n25329_));
  AOI21X1  g22893(.A0(new_n25329_), .A1(new_n25326_), .B0(new_n25130_), .Y(new_n25330_));
  INVX1    g22894(.A(new_n25330_), .Y(new_n25331_));
  AND2X1   g22895(.A(new_n8009_), .B(pi0199), .Y(new_n25332_));
  INVX1    g22896(.A(new_n25332_), .Y(new_n25333_));
  NOR2X1   g22897(.A(pi1153), .B(pi0200), .Y(new_n25334_));
  OR2X1    g22898(.A(new_n25334_), .B(pi0199), .Y(new_n25335_));
  AND2X1   g22899(.A(new_n25335_), .B(new_n2953_), .Y(new_n25336_));
  AND2X1   g22900(.A(new_n25336_), .B(new_n25333_), .Y(new_n25337_));
  AOI21X1  g22901(.A0(new_n25337_), .A1(pi0207), .B0(new_n23109_), .Y(new_n25338_));
  OAI21X1  g22902(.A0(new_n25331_), .A1(pi0207), .B0(new_n25338_), .Y(new_n25339_));
  INVX1    g22903(.A(new_n25339_), .Y(new_n25340_));
  AOI21X1  g22904(.A0(new_n25331_), .A1(new_n25121_), .B0(new_n25340_), .Y(new_n25341_));
  NOR3X1   g22905(.A(pi0299), .B(pi0200), .C(pi0199), .Y(new_n25342_));
  OAI21X1  g22906(.A0(new_n25342_), .A1(pi1153), .B0(new_n25046_), .Y(new_n25343_));
  NOR2X1   g22907(.A(pi1153), .B(pi0199), .Y(new_n25344_));
  NOR4X1   g22908(.A(new_n25344_), .B(new_n25268_), .C(new_n8130_), .D(pi0299), .Y(new_n25345_));
  INVX1    g22909(.A(new_n25345_), .Y(new_n25346_));
  AND2X1   g22910(.A(new_n25346_), .B(new_n25343_), .Y(new_n25347_));
  INVX1    g22911(.A(new_n25347_), .Y(new_n25348_));
  NOR2X1   g22912(.A(pi0208), .B(pi0207), .Y(new_n25349_));
  NOR3X1   g22913(.A(pi1153), .B(pi0200), .C(pi0199), .Y(new_n25350_));
  NOR3X1   g22914(.A(new_n25350_), .B(new_n25268_), .C(pi0299), .Y(new_n25351_));
  INVX1    g22915(.A(new_n25351_), .Y(new_n25352_));
  AOI21X1  g22916(.A0(new_n25352_), .A1(new_n7896_), .B0(new_n25349_), .Y(new_n25353_));
  OAI21X1  g22917(.A0(new_n25348_), .A1(new_n7896_), .B0(new_n25353_), .Y(new_n25354_));
  AND2X1   g22918(.A(new_n25354_), .B(pi0211), .Y(new_n25355_));
  AOI21X1  g22919(.A0(new_n25341_), .A1(new_n8548_), .B0(new_n25355_), .Y(new_n25356_));
  OAI21X1  g22920(.A0(new_n25354_), .A1(new_n25323_), .B0(pi0219), .Y(new_n25357_));
  AOI21X1  g22921(.A0(new_n25356_), .A1(new_n25323_), .B0(new_n25357_), .Y(new_n25358_));
  NOR2X1   g22922(.A(new_n25358_), .B(po1038), .Y(new_n25359_));
  OAI21X1  g22923(.A0(new_n25347_), .A1(new_n22803_), .B0(new_n25027_), .Y(new_n25360_));
  AND2X1   g22924(.A(new_n12615_), .B(pi0299), .Y(new_n25361_));
  INVX1    g22925(.A(new_n25361_), .Y(new_n25362_));
  AOI21X1  g22926(.A0(new_n25336_), .A1(new_n25333_), .B0(new_n22803_), .Y(new_n25363_));
  AND2X1   g22927(.A(new_n25363_), .B(new_n25362_), .Y(new_n25364_));
  INVX1    g22928(.A(new_n25343_), .Y(new_n25365_));
  AOI21X1  g22929(.A0(new_n8132_), .A1(pi1154), .B0(new_n25365_), .Y(new_n25366_));
  AOI21X1  g22930(.A0(new_n25366_), .A1(new_n25346_), .B0(pi0207), .Y(new_n25367_));
  OR2X1    g22931(.A(new_n25367_), .B(new_n25364_), .Y(new_n25368_));
  MX2X1    g22932(.A(new_n25368_), .B(new_n25360_), .S0(new_n23109_), .Y(new_n25369_));
  AND2X1   g22933(.A(new_n25369_), .B(new_n8548_), .Y(new_n25370_));
  NOR3X1   g22934(.A(new_n12494_), .B(new_n2953_), .C(pi0207), .Y(new_n25371_));
  NOR2X1   g22935(.A(new_n25053_), .B(pi1153), .Y(new_n25372_));
  OAI21X1  g22936(.A0(pi0299), .A1(new_n7941_), .B0(pi1154), .Y(new_n25373_));
  AOI21X1  g22937(.A0(new_n25373_), .A1(new_n25107_), .B0(new_n25372_), .Y(new_n25374_));
  AOI21X1  g22938(.A0(new_n25374_), .A1(pi0207), .B0(new_n25371_), .Y(new_n25375_));
  NOR2X1   g22939(.A(new_n8131_), .B(pi1153), .Y(new_n25376_));
  AND2X1   g22940(.A(new_n25268_), .B(new_n2953_), .Y(new_n25377_));
  NOR3X1   g22941(.A(new_n25377_), .B(new_n25376_), .C(new_n22803_), .Y(new_n25378_));
  AOI21X1  g22942(.A0(new_n25374_), .A1(new_n22803_), .B0(new_n25378_), .Y(new_n25379_));
  MX2X1    g22943(.A(new_n25379_), .B(new_n25375_), .S0(new_n23109_), .Y(new_n25380_));
  NOR2X1   g22944(.A(new_n25380_), .B(new_n8548_), .Y(new_n25381_));
  OR2X1    g22945(.A(new_n25381_), .B(new_n25370_), .Y(new_n25382_));
  OR2X1    g22946(.A(new_n25380_), .B(pi0211), .Y(new_n25383_));
  OR2X1    g22947(.A(new_n25341_), .B(new_n8548_), .Y(new_n25384_));
  NAND3X1  g22948(.A(new_n25384_), .B(new_n25383_), .C(pi0214), .Y(new_n25385_));
  AND2X1   g22949(.A(new_n25385_), .B(pi0212), .Y(new_n25386_));
  OAI21X1  g22950(.A0(new_n25382_), .A1(pi0214), .B0(new_n25386_), .Y(new_n25387_));
  AOI21X1  g22951(.A0(new_n25354_), .A1(new_n24984_), .B0(pi0212), .Y(new_n25388_));
  OAI21X1  g22952(.A0(new_n25382_), .A1(new_n24984_), .B0(new_n25388_), .Y(new_n25389_));
  NAND3X1  g22953(.A(new_n25389_), .B(new_n25387_), .C(new_n23539_), .Y(new_n25390_));
  NAND2X1  g22954(.A(new_n25390_), .B(new_n25359_), .Y(new_n25391_));
  AND2X1   g22955(.A(new_n8074_), .B(new_n8548_), .Y(new_n25392_));
  OR2X1    g22956(.A(pi1154), .B(new_n12494_), .Y(new_n25393_));
  OAI22X1  g22957(.A0(new_n25393_), .A1(new_n25135_), .B0(new_n25373_), .B1(new_n25372_), .Y(new_n25394_));
  AOI21X1  g22958(.A0(new_n25394_), .A1(pi0207), .B0(new_n25371_), .Y(new_n25395_));
  NOR2X1   g22959(.A(new_n8131_), .B(new_n22803_), .Y(new_n25396_));
  AOI22X1  g22960(.A0(new_n25396_), .A1(pi1153), .B0(new_n25394_), .B1(new_n22803_), .Y(new_n25397_));
  MX2X1    g22961(.A(new_n25397_), .B(new_n25395_), .S0(new_n23109_), .Y(new_n25398_));
  INVX1    g22962(.A(new_n25376_), .Y(new_n25399_));
  AOI21X1  g22963(.A0(new_n2953_), .A1(pi0199), .B0(new_n12494_), .Y(new_n25400_));
  INVX1    g22964(.A(new_n25400_), .Y(new_n25401_));
  AOI21X1  g22965(.A0(new_n25401_), .A1(new_n25399_), .B0(new_n12615_), .Y(new_n25402_));
  OR2X1    g22966(.A(new_n25402_), .B(new_n25324_), .Y(new_n25403_));
  MX2X1    g22967(.A(new_n25403_), .B(new_n25026_), .S0(new_n22803_), .Y(new_n25404_));
  OR2X1    g22968(.A(new_n25403_), .B(pi0207), .Y(new_n25405_));
  OAI21X1  g22969(.A0(new_n8135_), .A1(new_n12494_), .B0(new_n2953_), .Y(new_n25406_));
  AOI21X1  g22970(.A0(new_n25406_), .A1(new_n25362_), .B0(new_n22803_), .Y(new_n25407_));
  NOR2X1   g22971(.A(new_n25407_), .B(new_n23109_), .Y(new_n25408_));
  AOI22X1  g22972(.A0(new_n25408_), .A1(new_n25405_), .B0(new_n25404_), .B1(new_n23109_), .Y(new_n25409_));
  MX2X1    g22973(.A(new_n25409_), .B(new_n25398_), .S0(pi0211), .Y(new_n25410_));
  AOI22X1  g22974(.A0(new_n25410_), .A1(new_n25232_), .B0(new_n25398_), .B1(new_n25392_), .Y(new_n25411_));
  AOI21X1  g22975(.A0(new_n12494_), .A1(pi0200), .B0(new_n8503_), .Y(new_n25412_));
  MX2X1    g22976(.A(new_n25412_), .B(new_n25324_), .S0(new_n12615_), .Y(new_n25413_));
  NOR3X1   g22977(.A(pi0299), .B(new_n23109_), .C(new_n22803_), .Y(new_n25414_));
  NOR2X1   g22978(.A(new_n8131_), .B(new_n12494_), .Y(new_n25415_));
  AOI22X1  g22979(.A0(new_n25415_), .A1(new_n25414_), .B0(new_n25413_), .B1(new_n25259_), .Y(new_n25416_));
  INVX1    g22980(.A(new_n25416_), .Y(new_n25417_));
  OAI21X1  g22981(.A0(new_n25417_), .A1(new_n23539_), .B0(new_n6520_), .Y(new_n25418_));
  AOI21X1  g22982(.A0(pi0214), .A1(new_n8548_), .B0(new_n25232_), .Y(new_n25419_));
  AOI21X1  g22983(.A0(new_n25419_), .A1(new_n25416_), .B0(new_n25418_), .Y(new_n25420_));
  OAI21X1  g22984(.A0(new_n25411_), .A1(pi0219), .B0(new_n25420_), .Y(new_n25421_));
  AOI22X1  g22985(.A0(new_n25421_), .A1(new_n25258_), .B0(new_n25391_), .B1(new_n25294_), .Y(new_n25422_));
  AND2X1   g22986(.A(new_n6520_), .B(new_n25289_), .Y(new_n25423_));
  NOR3X1   g22987(.A(new_n12494_), .B(new_n8009_), .C(pi0199), .Y(new_n25424_));
  OAI21X1  g22988(.A0(new_n25424_), .A1(pi0299), .B0(new_n12615_), .Y(new_n25425_));
  OAI21X1  g22989(.A0(new_n8502_), .A1(pi1155), .B0(new_n25402_), .Y(new_n25426_));
  OAI21X1  g22990(.A0(new_n25425_), .A1(new_n25156_), .B0(new_n25426_), .Y(new_n25427_));
  NOR2X1   g22991(.A(new_n25427_), .B(new_n22803_), .Y(new_n25428_));
  INVX1    g22992(.A(new_n25156_), .Y(new_n25429_));
  AOI21X1  g22993(.A0(new_n25406_), .A1(new_n25429_), .B0(new_n22803_), .Y(new_n25430_));
  NOR2X1   g22994(.A(new_n25430_), .B(new_n23109_), .Y(new_n25431_));
  OAI21X1  g22995(.A0(new_n25427_), .A1(pi0207), .B0(new_n25431_), .Y(new_n25432_));
  OAI21X1  g22996(.A0(new_n25428_), .A1(new_n25104_), .B0(new_n25432_), .Y(new_n25433_));
  AOI21X1  g22997(.A0(new_n25409_), .A1(pi0211), .B0(new_n25014_), .Y(new_n25434_));
  OAI21X1  g22998(.A0(new_n25433_), .A1(pi0211), .B0(new_n25434_), .Y(new_n25435_));
  AOI21X1  g22999(.A0(pi1156), .A1(pi0299), .B0(pi0211), .Y(new_n25436_));
  AOI21X1  g23000(.A0(new_n25436_), .A1(new_n25416_), .B0(new_n24962_), .Y(new_n25437_));
  OAI21X1  g23001(.A0(new_n25433_), .A1(new_n8548_), .B0(new_n25437_), .Y(new_n25438_));
  AND2X1   g23002(.A(new_n25438_), .B(new_n25435_), .Y(new_n25439_));
  NAND2X1  g23003(.A(new_n25409_), .B(new_n8548_), .Y(new_n25440_));
  NOR2X1   g23004(.A(new_n24955_), .B(new_n23539_), .Y(new_n25441_));
  INVX1    g23005(.A(new_n25441_), .Y(new_n25442_));
  AOI21X1  g23006(.A0(new_n25416_), .A1(pi0211), .B0(new_n25442_), .Y(new_n25443_));
  AOI22X1  g23007(.A0(new_n25443_), .A1(new_n25440_), .B0(new_n25417_), .B1(new_n24955_), .Y(new_n25444_));
  OAI21X1  g23008(.A0(new_n25439_), .A1(pi0219), .B0(new_n25444_), .Y(new_n25445_));
  INVX1    g23009(.A(new_n25354_), .Y(new_n25446_));
  AOI22X1  g23010(.A0(new_n25370_), .A1(new_n25323_), .B0(new_n25446_), .B1(new_n24994_), .Y(new_n25447_));
  AND2X1   g23011(.A(new_n25369_), .B(pi0211), .Y(new_n25448_));
  OAI21X1  g23012(.A0(new_n25330_), .A1(new_n25104_), .B0(new_n25339_), .Y(new_n25449_));
  NOR3X1   g23013(.A(pi1154), .B(pi0200), .C(pi0199), .Y(new_n25450_));
  AOI22X1  g23014(.A0(new_n25450_), .A1(new_n25120_), .B0(new_n12591_), .B1(pi0299), .Y(new_n25451_));
  NAND3X1  g23015(.A(new_n25451_), .B(new_n25449_), .C(new_n8548_), .Y(new_n25452_));
  NAND2X1  g23016(.A(new_n25452_), .B(new_n8074_), .Y(new_n25453_));
  NAND3X1  g23017(.A(new_n25451_), .B(new_n25449_), .C(pi0211), .Y(new_n25454_));
  OAI21X1  g23018(.A0(new_n25348_), .A1(new_n25166_), .B0(new_n22803_), .Y(new_n25455_));
  OAI21X1  g23019(.A0(pi1156), .A1(new_n2953_), .B0(new_n25363_), .Y(new_n25456_));
  NAND3X1  g23020(.A(new_n25456_), .B(new_n25455_), .C(pi0208), .Y(new_n25457_));
  AOI21X1  g23021(.A0(pi1156), .A1(pi0299), .B0(pi0208), .Y(new_n25458_));
  OAI21X1  g23022(.A0(new_n25347_), .A1(new_n22803_), .B0(new_n25458_), .Y(new_n25459_));
  AND2X1   g23023(.A(new_n25459_), .B(new_n8548_), .Y(new_n25460_));
  AOI21X1  g23024(.A0(new_n25460_), .A1(new_n25457_), .B0(new_n24962_), .Y(new_n25461_));
  NAND3X1  g23025(.A(new_n25354_), .B(new_n24984_), .C(new_n24961_), .Y(new_n25462_));
  NAND2X1  g23026(.A(new_n25462_), .B(new_n23539_), .Y(new_n25463_));
  AOI21X1  g23027(.A0(new_n25461_), .A1(new_n25454_), .B0(new_n25463_), .Y(new_n25464_));
  OAI21X1  g23028(.A0(new_n25453_), .A1(new_n25448_), .B0(new_n25464_), .Y(new_n25465_));
  OAI21X1  g23029(.A0(new_n25447_), .A1(new_n23539_), .B0(new_n25465_), .Y(new_n25466_));
  AND2X1   g23030(.A(new_n6520_), .B(pi1152), .Y(new_n25467_));
  AOI22X1  g23031(.A0(new_n25467_), .A1(new_n25466_), .B0(new_n25445_), .B1(new_n25423_), .Y(new_n25468_));
  OAI21X1  g23032(.A0(new_n25468_), .A1(new_n25003_), .B0(new_n23244_), .Y(new_n25469_));
  AOI21X1  g23033(.A0(new_n25422_), .A1(new_n25003_), .B0(new_n25469_), .Y(new_n25470_));
  NOR2X1   g23034(.A(new_n25008_), .B(new_n24961_), .Y(new_n25471_));
  NOR3X1   g23035(.A(new_n25006_), .B(new_n24984_), .C(pi0212), .Y(new_n25472_));
  NOR3X1   g23036(.A(new_n25472_), .B(new_n25471_), .C(pi0219), .Y(new_n25473_));
  AOI21X1  g23037(.A0(pi1154), .A1(new_n8548_), .B0(new_n23539_), .Y(new_n25474_));
  OR4X1    g23038(.A(new_n25474_), .B(new_n24957_), .C(new_n6520_), .D(new_n25003_), .Y(new_n25475_));
  OAI22X1  g23039(.A0(new_n25475_), .A1(new_n25473_), .B0(new_n25470_), .B1(new_n25322_), .Y(new_n25476_));
  MX2X1    g23040(.A(new_n25476_), .B(pi0234), .S0(new_n24954_), .Y(po0391));
  INVX1    g23041(.A(new_n25109_), .Y(new_n25478_));
  OAI21X1  g23042(.A0(new_n25157_), .A1(new_n25065_), .B0(pi0207), .Y(new_n25479_));
  INVX1    g23043(.A(new_n25479_), .Y(new_n25480_));
  NOR4X1   g23044(.A(new_n25108_), .B(new_n25107_), .C(new_n25106_), .D(pi0207), .Y(new_n25481_));
  OAI21X1  g23045(.A0(new_n25481_), .A1(new_n25480_), .B0(pi0208), .Y(new_n25482_));
  AOI21X1  g23046(.A0(new_n25482_), .A1(new_n25478_), .B0(pi1157), .Y(new_n25483_));
  AND2X1   g23047(.A(pi1157), .B(pi0208), .Y(new_n25484_));
  INVX1    g23048(.A(new_n25484_), .Y(new_n25485_));
  OR2X1    g23049(.A(new_n25099_), .B(pi0207), .Y(new_n25486_));
  AOI21X1  g23050(.A0(new_n25486_), .A1(new_n25479_), .B0(new_n25485_), .Y(new_n25487_));
  NOR3X1   g23051(.A(new_n25487_), .B(new_n25483_), .C(new_n25103_), .Y(new_n25488_));
  AND2X1   g23052(.A(new_n25059_), .B(new_n12684_), .Y(new_n25489_));
  OAI21X1  g23053(.A0(new_n25489_), .A1(new_n25164_), .B0(pi0207), .Y(new_n25490_));
  NAND3X1  g23054(.A(new_n25144_), .B(new_n25142_), .C(new_n22803_), .Y(new_n25491_));
  AOI21X1  g23055(.A0(new_n25491_), .A1(new_n25490_), .B0(new_n23109_), .Y(new_n25492_));
  NOR2X1   g23056(.A(new_n25492_), .B(new_n25171_), .Y(new_n25493_));
  NOR2X1   g23057(.A(new_n25493_), .B(pi1157), .Y(new_n25494_));
  INVX1    g23058(.A(new_n25174_), .Y(new_n25495_));
  NOR2X1   g23059(.A(new_n25118_), .B(new_n12684_), .Y(new_n25496_));
  OAI21X1  g23060(.A0(new_n25496_), .A1(new_n25072_), .B0(new_n22803_), .Y(new_n25497_));
  AND2X1   g23061(.A(new_n25497_), .B(new_n25490_), .Y(new_n25498_));
  OR2X1    g23062(.A(new_n25498_), .B(new_n25485_), .Y(new_n25499_));
  NAND2X1  g23063(.A(new_n25499_), .B(new_n25495_), .Y(new_n25500_));
  OR2X1    g23064(.A(new_n25500_), .B(new_n25494_), .Y(new_n25501_));
  AOI21X1  g23065(.A0(new_n25501_), .A1(new_n8548_), .B0(new_n25014_), .Y(new_n25502_));
  OAI21X1  g23066(.A0(new_n25488_), .A1(new_n8548_), .B0(new_n25502_), .Y(new_n25503_));
  NOR2X1   g23067(.A(new_n25042_), .B(pi0208), .Y(new_n25504_));
  NOR3X1   g23068(.A(new_n25489_), .B(new_n25065_), .C(new_n7897_), .Y(new_n25505_));
  NOR3X1   g23069(.A(new_n25041_), .B(new_n25038_), .C(new_n25037_), .Y(new_n25506_));
  NOR2X1   g23070(.A(new_n25506_), .B(pi0207), .Y(new_n25507_));
  NOR3X1   g23071(.A(new_n25507_), .B(new_n25505_), .C(new_n25504_), .Y(new_n25508_));
  OR2X1    g23072(.A(new_n25508_), .B(pi1157), .Y(new_n25509_));
  AOI21X1  g23073(.A0(new_n25073_), .A1(pi0207), .B0(pi0208), .Y(new_n25510_));
  NOR3X1   g23074(.A(new_n25072_), .B(new_n25071_), .C(pi0207), .Y(new_n25511_));
  NOR3X1   g23075(.A(new_n25511_), .B(new_n25505_), .C(new_n25510_), .Y(new_n25512_));
  OAI21X1  g23076(.A0(new_n25512_), .A1(new_n12706_), .B0(new_n25509_), .Y(new_n25513_));
  AND2X1   g23077(.A(new_n25513_), .B(new_n24955_), .Y(new_n25514_));
  OAI21X1  g23078(.A0(new_n25500_), .A1(new_n25494_), .B0(pi0211), .Y(new_n25515_));
  INVX1    g23079(.A(new_n25232_), .Y(new_n25516_));
  AOI21X1  g23080(.A0(new_n25119_), .A1(new_n22803_), .B0(new_n23109_), .Y(new_n25517_));
  OR4X1    g23081(.A(new_n25157_), .B(new_n25156_), .C(new_n25164_), .D(new_n22803_), .Y(new_n25518_));
  AOI21X1  g23082(.A0(new_n25518_), .A1(new_n25517_), .B0(new_n25123_), .Y(new_n25519_));
  OAI21X1  g23083(.A0(new_n25508_), .A1(pi1157), .B0(new_n8548_), .Y(new_n25520_));
  AOI21X1  g23084(.A0(new_n25519_), .A1(pi1157), .B0(new_n25520_), .Y(new_n25521_));
  NOR2X1   g23085(.A(new_n25521_), .B(new_n25516_), .Y(new_n25522_));
  AOI21X1  g23086(.A0(new_n25522_), .A1(new_n25515_), .B0(new_n25514_), .Y(new_n25523_));
  AOI21X1  g23087(.A0(new_n25523_), .A1(new_n25503_), .B0(pi0219), .Y(new_n25524_));
  OR4X1    g23088(.A(new_n25487_), .B(new_n25483_), .C(new_n25103_), .D(pi0211), .Y(new_n25525_));
  AOI21X1  g23089(.A0(new_n25513_), .A1(pi0211), .B0(new_n24962_), .Y(new_n25526_));
  OAI21X1  g23090(.A0(new_n25513_), .A1(new_n24963_), .B0(pi0219), .Y(new_n25527_));
  AOI21X1  g23091(.A0(new_n25526_), .A1(new_n25525_), .B0(new_n25527_), .Y(new_n25528_));
  NOR3X1   g23092(.A(new_n25528_), .B(new_n25524_), .C(new_n23244_), .Y(new_n25529_));
  AOI21X1  g23093(.A0(new_n25131_), .A1(new_n25159_), .B0(new_n25122_), .Y(new_n25530_));
  AND2X1   g23094(.A(new_n25131_), .B(new_n25120_), .Y(new_n25531_));
  INVX1    g23095(.A(new_n25425_), .Y(new_n25532_));
  NOR3X1   g23096(.A(new_n25532_), .B(new_n25402_), .C(new_n22803_), .Y(new_n25533_));
  NOR3X1   g23097(.A(new_n25533_), .B(new_n25531_), .C(new_n23109_), .Y(new_n25534_));
  OAI21X1  g23098(.A0(new_n25534_), .A1(new_n25530_), .B0(pi1157), .Y(new_n25535_));
  OAI21X1  g23099(.A0(new_n25349_), .A1(new_n25058_), .B0(new_n7897_), .Y(new_n25536_));
  OAI21X1  g23100(.A0(new_n25413_), .A1(new_n7897_), .B0(new_n25536_), .Y(new_n25537_));
  INVX1    g23101(.A(new_n25537_), .Y(new_n25538_));
  AOI21X1  g23102(.A0(new_n25538_), .A1(new_n12706_), .B0(pi0211), .Y(new_n25539_));
  AND2X1   g23103(.A(new_n25537_), .B(new_n25167_), .Y(new_n25540_));
  AOI22X1  g23104(.A0(new_n25540_), .A1(pi0211), .B0(new_n25539_), .B1(new_n25535_), .Y(new_n25541_));
  NAND2X1  g23105(.A(new_n25090_), .B(new_n22803_), .Y(new_n25542_));
  NOR2X1   g23106(.A(new_n25428_), .B(new_n23109_), .Y(new_n25543_));
  AOI22X1  g23107(.A0(new_n25543_), .A1(new_n25542_), .B0(new_n25101_), .B1(new_n25238_), .Y(new_n25544_));
  OR2X1    g23108(.A(new_n25544_), .B(new_n8548_), .Y(new_n25545_));
  AOI21X1  g23109(.A0(new_n25537_), .A1(new_n25167_), .B0(pi0211), .Y(new_n25546_));
  NOR2X1   g23110(.A(new_n25546_), .B(new_n25014_), .Y(new_n25547_));
  AOI22X1  g23111(.A0(new_n25547_), .A1(new_n25545_), .B0(new_n25537_), .B1(new_n24955_), .Y(new_n25548_));
  OAI21X1  g23112(.A0(new_n25541_), .A1(new_n25516_), .B0(new_n25548_), .Y(new_n25549_));
  AOI21X1  g23113(.A0(new_n25537_), .A1(pi0211), .B0(new_n24962_), .Y(new_n25550_));
  INVX1    g23114(.A(new_n25550_), .Y(new_n25551_));
  AOI21X1  g23115(.A0(new_n25544_), .A1(new_n8548_), .B0(new_n25551_), .Y(new_n25552_));
  AOI21X1  g23116(.A0(new_n25538_), .A1(new_n24962_), .B0(new_n23539_), .Y(new_n25553_));
  INVX1    g23117(.A(new_n25553_), .Y(new_n25554_));
  OAI21X1  g23118(.A0(new_n25554_), .A1(new_n25552_), .B0(new_n23244_), .Y(new_n25555_));
  AOI21X1  g23119(.A0(new_n25549_), .A1(new_n23539_), .B0(new_n25555_), .Y(new_n25556_));
  OAI21X1  g23120(.A0(new_n25556_), .A1(new_n25529_), .B0(new_n6520_), .Y(new_n25557_));
  NAND3X1  g23121(.A(new_n25004_), .B(pi0214), .C(new_n24961_), .Y(new_n25558_));
  NAND2X1  g23122(.A(new_n25004_), .B(new_n24984_), .Y(new_n25559_));
  OAI21X1  g23123(.A0(new_n25006_), .A1(new_n24984_), .B0(new_n25559_), .Y(new_n25560_));
  AOI21X1  g23124(.A0(new_n25560_), .A1(pi0212), .B0(pi0219), .Y(new_n25561_));
  NAND2X1  g23125(.A(new_n25561_), .B(new_n25558_), .Y(new_n25562_));
  AOI21X1  g23126(.A0(pi1155), .A1(new_n8548_), .B0(new_n23539_), .Y(new_n25563_));
  NOR2X1   g23127(.A(new_n25232_), .B(new_n23539_), .Y(new_n25564_));
  NOR3X1   g23128(.A(new_n25564_), .B(new_n25563_), .C(new_n6520_), .Y(new_n25565_));
  AOI21X1  g23129(.A0(new_n25565_), .A1(new_n25562_), .B0(new_n25003_), .Y(new_n25566_));
  NOR2X1   g23130(.A(new_n25519_), .B(new_n12706_), .Y(new_n25567_));
  INVX1    g23131(.A(new_n25567_), .Y(new_n25568_));
  AOI21X1  g23132(.A0(new_n12706_), .A1(pi0299), .B0(new_n25494_), .Y(new_n25569_));
  AOI21X1  g23133(.A0(new_n25569_), .A1(new_n25568_), .B0(new_n25139_), .Y(new_n25570_));
  OR2X1    g23134(.A(new_n25570_), .B(pi0211), .Y(new_n25571_));
  AOI21X1  g23135(.A0(new_n25571_), .A1(new_n25526_), .B0(new_n25527_), .Y(new_n25572_));
  NAND2X1  g23136(.A(new_n25570_), .B(pi0211), .Y(new_n25573_));
  AOI21X1  g23137(.A0(new_n25137_), .A1(new_n25061_), .B0(new_n25065_), .Y(new_n25574_));
  NOR4X1   g23138(.A(new_n25268_), .B(new_n25038_), .C(new_n8130_), .D(pi0299), .Y(new_n25575_));
  AOI21X1  g23139(.A0(new_n25144_), .A1(pi1154), .B0(new_n25575_), .Y(new_n25576_));
  OR2X1    g23140(.A(new_n25106_), .B(pi0207), .Y(new_n25577_));
  OAI22X1  g23141(.A0(new_n25577_), .A1(new_n25576_), .B0(new_n25574_), .B1(new_n22803_), .Y(new_n25578_));
  AOI21X1  g23142(.A0(new_n25578_), .A1(pi0208), .B0(new_n25126_), .Y(new_n25579_));
  OAI22X1  g23143(.A0(new_n25579_), .A1(pi1157), .B0(new_n25519_), .B1(new_n25125_), .Y(new_n25580_));
  AOI21X1  g23144(.A0(new_n25580_), .A1(new_n8548_), .B0(new_n25014_), .Y(new_n25581_));
  NAND2X1  g23145(.A(new_n25581_), .B(new_n25573_), .Y(new_n25582_));
  OAI21X1  g23146(.A0(new_n25580_), .A1(new_n8548_), .B0(new_n25525_), .Y(new_n25583_));
  AOI21X1  g23147(.A0(new_n25583_), .A1(new_n25232_), .B0(new_n25514_), .Y(new_n25584_));
  AOI21X1  g23148(.A0(new_n25584_), .A1(new_n25582_), .B0(pi0219), .Y(new_n25585_));
  OAI21X1  g23149(.A0(new_n25585_), .A1(new_n25572_), .B0(pi0209), .Y(new_n25586_));
  INVX1    g23150(.A(new_n25371_), .Y(new_n25587_));
  OAI21X1  g23151(.A0(new_n25131_), .A1(new_n22803_), .B0(new_n25587_), .Y(new_n25588_));
  AND2X1   g23152(.A(new_n25588_), .B(new_n23109_), .Y(new_n25589_));
  INVX1    g23153(.A(new_n25131_), .Y(new_n25590_));
  MX2X1    g23154(.A(new_n25394_), .B(new_n25590_), .S0(new_n22803_), .Y(new_n25591_));
  AOI21X1  g23155(.A0(new_n25591_), .A1(pi0208), .B0(new_n25589_), .Y(new_n25592_));
  AND2X1   g23156(.A(new_n25592_), .B(new_n8548_), .Y(new_n25593_));
  OAI21X1  g23157(.A0(new_n25593_), .A1(new_n25551_), .B0(new_n25553_), .Y(new_n25594_));
  NAND2X1  g23158(.A(new_n25544_), .B(new_n8548_), .Y(new_n25595_));
  MX2X1    g23159(.A(new_n25114_), .B(new_n25026_), .S0(new_n22803_), .Y(new_n25596_));
  MX2X1    g23160(.A(new_n25403_), .B(new_n25114_), .S0(new_n22803_), .Y(new_n25597_));
  MX2X1    g23161(.A(new_n25597_), .B(new_n25596_), .S0(new_n23109_), .Y(new_n25598_));
  OAI21X1  g23162(.A0(new_n25598_), .A1(new_n8548_), .B0(new_n25595_), .Y(new_n25599_));
  AND2X1   g23163(.A(new_n25598_), .B(new_n8548_), .Y(new_n25600_));
  OAI21X1  g23164(.A0(new_n25592_), .A1(new_n8548_), .B0(new_n8074_), .Y(new_n25601_));
  OAI22X1  g23165(.A0(new_n25601_), .A1(new_n25600_), .B0(new_n25538_), .B1(new_n25323_), .Y(new_n25602_));
  AOI21X1  g23166(.A0(new_n25599_), .A1(new_n24963_), .B0(new_n25602_), .Y(new_n25603_));
  OAI21X1  g23167(.A0(new_n25603_), .A1(pi0219), .B0(new_n25594_), .Y(new_n25604_));
  AOI21X1  g23168(.A0(new_n25604_), .A1(new_n23244_), .B0(po1038), .Y(new_n25605_));
  AOI21X1  g23169(.A0(pi1153), .A1(new_n8548_), .B0(new_n23539_), .Y(new_n25606_));
  OR2X1    g23170(.A(new_n25606_), .B(new_n6520_), .Y(new_n25607_));
  AOI21X1  g23171(.A0(new_n25255_), .A1(new_n8074_), .B0(pi0219), .Y(new_n25608_));
  OAI21X1  g23172(.A0(new_n25516_), .A1(new_n25007_), .B0(new_n25608_), .Y(new_n25609_));
  OAI21X1  g23173(.A0(new_n25232_), .A1(new_n23539_), .B0(new_n25609_), .Y(new_n25610_));
  OAI21X1  g23174(.A0(new_n25610_), .A1(new_n25607_), .B0(new_n25003_), .Y(new_n25611_));
  AOI21X1  g23175(.A0(new_n25605_), .A1(new_n25586_), .B0(new_n25611_), .Y(new_n25612_));
  AOI21X1  g23176(.A0(new_n25566_), .A1(new_n25557_), .B0(new_n25612_), .Y(new_n25613_));
  MX2X1    g23177(.A(new_n25613_), .B(pi0235), .S0(new_n24954_), .Y(po0392));
  NOR4X1   g23178(.A(new_n24809_), .B(new_n3193_), .C(pi0100), .D(pi0038), .Y(new_n25615_));
  OAI21X1  g23179(.A0(new_n25615_), .A1(new_n24946_), .B0(new_n5104_), .Y(new_n25616_));
  AOI21X1  g23180(.A0(new_n25616_), .A1(new_n3095_), .B0(new_n5790_), .Y(new_n25617_));
  OAI21X1  g23181(.A0(new_n25617_), .A1(pi0092), .B0(new_n9927_), .Y(new_n25618_));
  AOI21X1  g23182(.A0(new_n25618_), .A1(new_n4991_), .B0(new_n4994_), .Y(new_n25619_));
  OAI21X1  g23183(.A0(new_n25619_), .A1(pi0056), .B0(new_n4990_), .Y(new_n25620_));
  AOI21X1  g23184(.A0(new_n25620_), .A1(new_n3245_), .B0(new_n9931_), .Y(po0393));
  MX2X1    g23185(.A(pi1158), .B(pi1157), .S0(pi0211), .Y(new_n25622_));
  NAND3X1  g23186(.A(new_n25622_), .B(pi0214), .C(new_n24961_), .Y(new_n25623_));
  AND2X1   g23187(.A(new_n25623_), .B(new_n25561_), .Y(new_n25624_));
  NOR4X1   g23188(.A(new_n12684_), .B(new_n24984_), .C(pi0212), .D(pi0211), .Y(new_n25625_));
  OAI22X1  g23189(.A0(new_n25625_), .A1(new_n23539_), .B0(new_n5118_), .B1(pi0057), .Y(new_n25626_));
  INVX1    g23190(.A(new_n25626_), .Y(new_n25627_));
  AND2X1   g23191(.A(pi1154), .B(new_n8548_), .Y(new_n25628_));
  AOI22X1  g23192(.A0(new_n25182_), .A1(pi1155), .B0(new_n25628_), .B1(pi0214), .Y(new_n25629_));
  NOR3X1   g23193(.A(new_n25629_), .B(new_n6520_), .C(new_n24961_), .Y(new_n25630_));
  NOR2X1   g23194(.A(new_n25630_), .B(new_n25627_), .Y(new_n25631_));
  OAI21X1  g23195(.A0(new_n25631_), .A1(new_n25624_), .B0(new_n25003_), .Y(new_n25632_));
  INVX1    g23196(.A(new_n25021_), .Y(new_n25633_));
  AOI21X1  g23197(.A0(pi1143), .A1(pi0199), .B0(pi0200), .Y(new_n25634_));
  OAI21X1  g23198(.A0(new_n2439_), .A1(pi0199), .B0(new_n25634_), .Y(new_n25635_));
  NAND3X1  g23199(.A(new_n25635_), .B(new_n25414_), .C(new_n24972_), .Y(new_n25636_));
  OAI21X1  g23200(.A0(new_n3346_), .A1(pi0199), .B0(new_n25634_), .Y(new_n25637_));
  OAI21X1  g23201(.A0(new_n2439_), .A1(pi0199), .B0(pi0200), .Y(new_n25638_));
  NAND3X1  g23202(.A(new_n25638_), .B(new_n25637_), .C(new_n25259_), .Y(new_n25639_));
  AOI21X1  g23203(.A0(new_n25639_), .A1(new_n25636_), .B0(pi0299), .Y(new_n25640_));
  INVX1    g23204(.A(new_n25023_), .Y(new_n25641_));
  NOR2X1   g23205(.A(new_n25026_), .B(new_n24984_), .Y(new_n25642_));
  OAI21X1  g23206(.A0(new_n25024_), .A1(pi0214), .B0(pi0212), .Y(new_n25643_));
  OAI22X1  g23207(.A0(new_n25643_), .A1(new_n25642_), .B0(new_n25167_), .B1(new_n25641_), .Y(new_n25644_));
  AOI21X1  g23208(.A0(new_n25644_), .A1(new_n25030_), .B0(new_n25640_), .Y(new_n25645_));
  OAI21X1  g23209(.A0(new_n25624_), .A1(new_n25633_), .B0(new_n25645_), .Y(new_n25646_));
  AOI21X1  g23210(.A0(new_n25646_), .A1(new_n6520_), .B0(new_n25632_), .Y(new_n25647_));
  MX2X1    g23211(.A(new_n3346_), .B(new_n2439_), .S0(pi0211), .Y(new_n25648_));
  AOI21X1  g23212(.A0(new_n25648_), .A1(new_n25014_), .B0(new_n24955_), .Y(new_n25649_));
  OAI21X1  g23213(.A0(new_n24960_), .A1(new_n25014_), .B0(new_n25649_), .Y(new_n25650_));
  NAND2X1  g23214(.A(new_n25650_), .B(new_n23539_), .Y(new_n25651_));
  OAI21X1  g23215(.A0(new_n3495_), .A1(pi0211), .B0(pi0219), .Y(new_n25652_));
  NAND3X1  g23216(.A(new_n25652_), .B(new_n25651_), .C(new_n24958_), .Y(new_n25653_));
  NAND3X1  g23217(.A(new_n25441_), .B(new_n24964_), .C(pi0299), .Y(new_n25654_));
  OAI21X1  g23218(.A0(new_n25650_), .A1(new_n25633_), .B0(new_n25654_), .Y(new_n25655_));
  OAI21X1  g23219(.A0(new_n25655_), .A1(new_n25640_), .B0(new_n6520_), .Y(new_n25656_));
  NAND2X1  g23220(.A(new_n25656_), .B(new_n25653_), .Y(new_n25657_));
  OAI21X1  g23221(.A0(new_n25657_), .A1(new_n25003_), .B0(pi0209), .Y(new_n25658_));
  NAND3X1  g23222(.A(new_n25053_), .B(new_n23109_), .C(pi0207), .Y(new_n25659_));
  OR2X1    g23223(.A(pi1158), .B(pi0199), .Y(new_n25660_));
  AOI22X1  g23224(.A0(new_n25660_), .A1(pi1156), .B0(new_n25342_), .B1(pi1158), .Y(new_n25661_));
  NOR2X1   g23225(.A(new_n25661_), .B(new_n25659_), .Y(new_n25662_));
  AND2X1   g23226(.A(new_n25066_), .B(pi0207), .Y(new_n25663_));
  NOR3X1   g23227(.A(new_n25663_), .B(new_n25507_), .C(new_n23109_), .Y(new_n25664_));
  OAI21X1  g23228(.A0(new_n25664_), .A1(new_n25662_), .B0(new_n12706_), .Y(new_n25665_));
  INVX1    g23229(.A(new_n25159_), .Y(new_n25666_));
  NOR3X1   g23230(.A(new_n12684_), .B(pi0200), .C(new_n7941_), .Y(new_n25667_));
  AOI21X1  g23231(.A0(new_n12676_), .A1(new_n8009_), .B0(pi0199), .Y(new_n25668_));
  NOR2X1   g23232(.A(new_n25668_), .B(new_n25667_), .Y(new_n25669_));
  NOR2X1   g23233(.A(new_n25669_), .B(new_n25666_), .Y(new_n25670_));
  NOR3X1   g23234(.A(new_n25663_), .B(new_n25511_), .C(new_n23109_), .Y(new_n25671_));
  AOI21X1  g23235(.A0(new_n25670_), .A1(new_n23109_), .B0(new_n25671_), .Y(new_n25672_));
  OAI21X1  g23236(.A0(new_n25672_), .A1(new_n12706_), .B0(new_n25665_), .Y(new_n25673_));
  NOR2X1   g23237(.A(new_n25673_), .B(new_n24956_), .Y(new_n25674_));
  OAI21X1  g23238(.A0(new_n25165_), .A1(new_n22803_), .B0(new_n25497_), .Y(new_n25675_));
  AND2X1   g23239(.A(new_n25675_), .B(new_n25484_), .Y(new_n25676_));
  AND2X1   g23240(.A(new_n25491_), .B(pi0208), .Y(new_n25677_));
  OAI21X1  g23241(.A0(new_n25165_), .A1(new_n22803_), .B0(new_n25677_), .Y(new_n25678_));
  NOR3X1   g23242(.A(new_n25661_), .B(new_n22803_), .C(pi0200), .Y(new_n25679_));
  INVX1    g23243(.A(new_n25679_), .Y(new_n25680_));
  AOI21X1  g23244(.A0(new_n25680_), .A1(new_n25458_), .B0(pi1157), .Y(new_n25681_));
  AND2X1   g23245(.A(new_n25681_), .B(new_n25678_), .Y(new_n25682_));
  OAI21X1  g23246(.A0(new_n25670_), .A1(new_n25166_), .B0(new_n25172_), .Y(new_n25683_));
  INVX1    g23247(.A(new_n25683_), .Y(new_n25684_));
  OR4X1    g23248(.A(new_n25684_), .B(new_n25682_), .C(new_n25676_), .D(new_n25641_), .Y(new_n25685_));
  AOI21X1  g23249(.A0(new_n25066_), .A1(new_n25100_), .B0(new_n22803_), .Y(new_n25686_));
  OAI21X1  g23250(.A0(new_n25686_), .A1(new_n25481_), .B0(pi0208), .Y(new_n25687_));
  AOI21X1  g23251(.A0(new_n25024_), .A1(new_n23109_), .B0(new_n25662_), .Y(new_n25688_));
  AOI21X1  g23252(.A0(new_n25688_), .A1(new_n25687_), .B0(pi1157), .Y(new_n25689_));
  INVX1    g23253(.A(new_n25686_), .Y(new_n25690_));
  AOI21X1  g23254(.A0(new_n25690_), .A1(new_n25486_), .B0(new_n25485_), .Y(new_n25691_));
  AOI21X1  g23255(.A0(new_n25039_), .A1(new_n2953_), .B0(pi1158), .Y(new_n25692_));
  NOR3X1   g23256(.A(new_n25692_), .B(new_n25377_), .C(new_n12684_), .Y(new_n25693_));
  OAI21X1  g23257(.A0(new_n25693_), .A1(new_n25668_), .B0(new_n25159_), .Y(new_n25694_));
  AOI21X1  g23258(.A0(new_n25694_), .A1(new_n25100_), .B0(new_n25173_), .Y(new_n25695_));
  NOR3X1   g23259(.A(new_n25695_), .B(new_n25691_), .C(new_n25689_), .Y(new_n25696_));
  NOR3X1   g23260(.A(new_n25361_), .B(new_n25119_), .C(pi0207), .Y(new_n25697_));
  NOR2X1   g23261(.A(new_n25662_), .B(pi1157), .Y(new_n25698_));
  OAI21X1  g23262(.A0(new_n25577_), .A1(new_n25576_), .B0(new_n25698_), .Y(new_n25699_));
  OAI21X1  g23263(.A0(new_n25697_), .A1(new_n12706_), .B0(new_n25699_), .Y(new_n25700_));
  AOI21X1  g23264(.A0(new_n25112_), .A1(pi0207), .B0(new_n23109_), .Y(new_n25701_));
  AOI21X1  g23265(.A0(pi1154), .A1(pi0299), .B0(pi0208), .Y(new_n25702_));
  OAI21X1  g23266(.A0(new_n25698_), .A1(new_n25694_), .B0(new_n25702_), .Y(new_n25703_));
  NAND2X1  g23267(.A(new_n25703_), .B(pi0214), .Y(new_n25704_));
  AOI21X1  g23268(.A0(new_n25701_), .A1(new_n25700_), .B0(new_n25704_), .Y(new_n25705_));
  NOR2X1   g23269(.A(new_n25705_), .B(new_n24961_), .Y(new_n25706_));
  OAI21X1  g23270(.A0(new_n25696_), .A1(pi0214), .B0(new_n25706_), .Y(new_n25707_));
  AOI21X1  g23271(.A0(new_n25707_), .A1(new_n25685_), .B0(pi0211), .Y(new_n25708_));
  OAI21X1  g23272(.A0(new_n25708_), .A1(new_n25674_), .B0(pi0219), .Y(new_n25709_));
  OR2X1    g23273(.A(new_n25673_), .B(pi0214), .Y(new_n25710_));
  AND2X1   g23274(.A(new_n25710_), .B(new_n24961_), .Y(new_n25711_));
  NOR3X1   g23275(.A(new_n25668_), .B(new_n25667_), .C(pi0299), .Y(new_n25712_));
  NOR2X1   g23276(.A(new_n25712_), .B(new_n25122_), .Y(new_n25713_));
  AOI21X1  g23277(.A0(new_n25517_), .A1(new_n25275_), .B0(new_n25713_), .Y(new_n25714_));
  OAI21X1  g23278(.A0(new_n25714_), .A1(new_n12706_), .B0(new_n25665_), .Y(new_n25715_));
  NOR2X1   g23279(.A(new_n25715_), .B(new_n8548_), .Y(new_n25716_));
  OR4X1    g23280(.A(new_n25157_), .B(new_n25156_), .C(new_n25134_), .D(new_n12676_), .Y(new_n25717_));
  AOI21X1  g23281(.A0(new_n25066_), .A1(new_n12676_), .B0(new_n22803_), .Y(new_n25718_));
  AND2X1   g23282(.A(new_n25718_), .B(new_n25717_), .Y(new_n25719_));
  AOI21X1  g23283(.A0(new_n25144_), .A1(new_n25142_), .B0(pi0299), .Y(new_n25720_));
  OAI21X1  g23284(.A0(pi1158), .A1(new_n2953_), .B0(new_n22803_), .Y(new_n25721_));
  OAI21X1  g23285(.A0(new_n25721_), .A1(new_n25720_), .B0(pi0208), .Y(new_n25722_));
  OAI21X1  g23286(.A0(new_n25396_), .A1(pi0299), .B0(pi1158), .Y(new_n25723_));
  AOI21X1  g23287(.A0(new_n25667_), .A1(new_n25159_), .B0(pi0208), .Y(new_n25724_));
  AOI21X1  g23288(.A0(new_n25724_), .A1(new_n25723_), .B0(pi1157), .Y(new_n25725_));
  OAI21X1  g23289(.A0(new_n25722_), .A1(new_n25719_), .B0(new_n25725_), .Y(new_n25726_));
  AND2X1   g23290(.A(new_n12676_), .B(pi0299), .Y(new_n25727_));
  NOR3X1   g23291(.A(new_n25727_), .B(new_n25119_), .C(pi0207), .Y(new_n25728_));
  OR2X1    g23292(.A(new_n25728_), .B(new_n25719_), .Y(new_n25729_));
  NOR3X1   g23293(.A(new_n25098_), .B(new_n25048_), .C(pi0299), .Y(new_n25730_));
  INVX1    g23294(.A(new_n25730_), .Y(new_n25731_));
  AOI21X1  g23295(.A0(new_n25342_), .A1(pi1158), .B0(new_n12706_), .Y(new_n25732_));
  AOI21X1  g23296(.A0(new_n25732_), .A1(new_n25731_), .B0(new_n22803_), .Y(new_n25733_));
  INVX1    g23297(.A(new_n25733_), .Y(new_n25734_));
  AOI21X1  g23298(.A0(new_n25734_), .A1(new_n25723_), .B0(new_n25173_), .Y(new_n25735_));
  OR2X1    g23299(.A(new_n25735_), .B(pi0211), .Y(new_n25736_));
  AOI21X1  g23300(.A0(new_n25729_), .A1(new_n25484_), .B0(new_n25736_), .Y(new_n25737_));
  AOI21X1  g23301(.A0(new_n25737_), .A1(new_n25726_), .B0(new_n25716_), .Y(new_n25738_));
  OAI21X1  g23302(.A0(new_n25738_), .A1(new_n24984_), .B0(new_n25711_), .Y(new_n25739_));
  INVX1    g23303(.A(new_n8033_), .Y(new_n25740_));
  INVX1    g23304(.A(new_n25180_), .Y(new_n25741_));
  NOR3X1   g23305(.A(new_n25684_), .B(new_n25682_), .C(new_n25676_), .Y(new_n25742_));
  NOR2X1   g23306(.A(new_n25742_), .B(new_n25741_), .Y(new_n25743_));
  AOI21X1  g23307(.A0(new_n25715_), .A1(new_n25182_), .B0(new_n25743_), .Y(new_n25744_));
  OAI21X1  g23308(.A0(new_n25696_), .A1(new_n25740_), .B0(new_n25744_), .Y(new_n25745_));
  AOI21X1  g23309(.A0(new_n25745_), .A1(pi0212), .B0(pi0219), .Y(new_n25746_));
  AOI21X1  g23310(.A0(new_n25746_), .A1(new_n25739_), .B0(po1038), .Y(new_n25747_));
  AOI21X1  g23311(.A0(new_n25747_), .A1(new_n25709_), .B0(new_n25632_), .Y(new_n25748_));
  AND2X1   g23312(.A(new_n3346_), .B(pi0299), .Y(new_n25749_));
  OAI21X1  g23313(.A0(new_n25749_), .A1(new_n25111_), .B0(pi1154), .Y(new_n25750_));
  AND2X1   g23314(.A(pi1145), .B(pi0299), .Y(new_n25751_));
  INVX1    g23315(.A(new_n25751_), .Y(new_n25752_));
  AOI21X1  g23316(.A0(new_n25752_), .A1(new_n25060_), .B0(pi1156), .Y(new_n25753_));
  OAI21X1  g23317(.A0(new_n25749_), .A1(new_n25133_), .B0(new_n12615_), .Y(new_n25754_));
  AOI21X1  g23318(.A0(new_n25752_), .A1(new_n25201_), .B0(new_n12684_), .Y(new_n25755_));
  AOI22X1  g23319(.A0(new_n25755_), .A1(new_n25754_), .B0(new_n25753_), .B1(new_n25750_), .Y(new_n25756_));
  NOR2X1   g23320(.A(new_n25756_), .B(new_n22803_), .Y(new_n25757_));
  INVX1    g23321(.A(new_n25757_), .Y(new_n25758_));
  AND2X1   g23322(.A(pi1157), .B(new_n8009_), .Y(new_n25759_));
  INVX1    g23323(.A(new_n25759_), .Y(new_n25760_));
  OAI21X1  g23324(.A0(new_n25760_), .A1(pi0199), .B0(new_n25720_), .Y(new_n25761_));
  AOI21X1  g23325(.A0(new_n3346_), .A1(pi0299), .B0(pi0207), .Y(new_n25762_));
  AOI21X1  g23326(.A0(new_n25762_), .A1(new_n25761_), .B0(new_n23109_), .Y(new_n25763_));
  OR4X1    g23327(.A(new_n12684_), .B(pi0299), .C(pi0200), .D(new_n7941_), .Y(new_n25764_));
  AOI21X1  g23328(.A0(new_n25342_), .A1(pi1158), .B0(pi1157), .Y(new_n25765_));
  NAND2X1  g23329(.A(new_n25765_), .B(new_n25764_), .Y(new_n25766_));
  OR2X1    g23330(.A(new_n25751_), .B(pi0208), .Y(new_n25767_));
  AOI21X1  g23331(.A0(new_n25766_), .A1(new_n25733_), .B0(new_n25767_), .Y(new_n25768_));
  AOI21X1  g23332(.A0(new_n25763_), .A1(new_n25758_), .B0(new_n25768_), .Y(new_n25769_));
  OAI21X1  g23333(.A0(new_n25679_), .A1(pi1157), .B0(new_n23109_), .Y(new_n25770_));
  NOR2X1   g23334(.A(new_n25770_), .B(new_n25694_), .Y(new_n25771_));
  NOR2X1   g23335(.A(new_n25771_), .B(pi0208), .Y(new_n25772_));
  AND2X1   g23336(.A(new_n25225_), .B(pi0207), .Y(new_n25773_));
  INVX1    g23337(.A(new_n25773_), .Y(new_n25774_));
  AOI21X1  g23338(.A0(new_n2439_), .A1(pi0299), .B0(pi0207), .Y(new_n25775_));
  AOI21X1  g23339(.A0(new_n25775_), .A1(new_n25761_), .B0(new_n23109_), .Y(new_n25776_));
  AOI22X1  g23340(.A0(new_n25776_), .A1(new_n25774_), .B0(new_n25772_), .B1(new_n25216_), .Y(new_n25777_));
  MX2X1    g23341(.A(new_n25777_), .B(new_n25769_), .S0(new_n8548_), .Y(new_n25778_));
  OAI21X1  g23342(.A0(new_n25778_), .A1(new_n24984_), .B0(new_n25711_), .Y(new_n25779_));
  OR2X1    g23343(.A(new_n25778_), .B(pi0214), .Y(new_n25780_));
  NAND2X1  g23344(.A(new_n25777_), .B(new_n8548_), .Y(new_n25781_));
  OR2X1    g23345(.A(new_n25203_), .B(new_n22803_), .Y(new_n25782_));
  AOI21X1  g23346(.A0(new_n3495_), .A1(pi0299), .B0(pi0207), .Y(new_n25783_));
  AOI21X1  g23347(.A0(new_n25783_), .A1(new_n25761_), .B0(new_n23109_), .Y(new_n25784_));
  AOI22X1  g23348(.A0(new_n25784_), .A1(new_n25782_), .B0(new_n25772_), .B1(new_n25190_), .Y(new_n25785_));
  AOI21X1  g23349(.A0(new_n25785_), .A1(pi0211), .B0(new_n24984_), .Y(new_n25786_));
  AOI21X1  g23350(.A0(new_n25786_), .A1(new_n25781_), .B0(new_n24961_), .Y(new_n25787_));
  AOI21X1  g23351(.A0(new_n25787_), .A1(new_n25780_), .B0(pi0219), .Y(new_n25788_));
  MX2X1    g23352(.A(new_n25785_), .B(new_n25673_), .S0(new_n24994_), .Y(new_n25789_));
  OAI21X1  g23353(.A0(new_n25789_), .A1(new_n23539_), .B0(new_n6520_), .Y(new_n25790_));
  AOI21X1  g23354(.A0(new_n25788_), .A1(new_n25779_), .B0(new_n25790_), .Y(new_n25791_));
  NAND2X1  g23355(.A(new_n25653_), .B(pi0213), .Y(new_n25792_));
  OAI21X1  g23356(.A0(new_n25792_), .A1(new_n25791_), .B0(new_n23244_), .Y(new_n25793_));
  OAI22X1  g23357(.A0(new_n25793_), .A1(new_n25748_), .B0(new_n25658_), .B1(new_n25647_), .Y(new_n25794_));
  MX2X1    g23358(.A(new_n25794_), .B(new_n22797_), .S0(new_n24954_), .Y(po0394));
  NOR2X1   g23359(.A(pi1153), .B(pi0211), .Y(new_n25796_));
  NAND2X1  g23360(.A(new_n25796_), .B(pi0219), .Y(new_n25797_));
  NAND3X1  g23361(.A(new_n25797_), .B(new_n25609_), .C(new_n24958_), .Y(new_n25798_));
  NOR4X1   g23362(.A(new_n25349_), .B(new_n7896_), .C(pi0299), .D(pi0200), .Y(new_n25799_));
  AOI21X1  g23363(.A0(new_n25414_), .A1(new_n25039_), .B0(new_n25799_), .Y(new_n25800_));
  OAI21X1  g23364(.A0(new_n25800_), .A1(new_n25350_), .B0(new_n24984_), .Y(new_n25801_));
  AND2X1   g23365(.A(new_n25801_), .B(new_n24961_), .Y(new_n25802_));
  MX2X1    g23366(.A(new_n25096_), .B(new_n25082_), .S0(pi1153), .Y(new_n25803_));
  OAI22X1  g23367(.A0(new_n25803_), .A1(new_n12591_), .B0(new_n25344_), .B1(new_n25054_), .Y(new_n25804_));
  AOI21X1  g23368(.A0(new_n25048_), .A1(new_n25159_), .B0(new_n23109_), .Y(new_n25805_));
  OR2X1    g23369(.A(new_n25805_), .B(new_n25101_), .Y(new_n25806_));
  AOI22X1  g23370(.A0(new_n25806_), .A1(new_n25804_), .B0(new_n25414_), .B1(new_n25039_), .Y(new_n25807_));
  NOR2X1   g23371(.A(new_n25007_), .B(new_n2953_), .Y(new_n25808_));
  NOR2X1   g23372(.A(new_n25808_), .B(new_n24984_), .Y(new_n25809_));
  OAI21X1  g23373(.A0(new_n25807_), .A1(pi0299), .B0(new_n25809_), .Y(new_n25810_));
  AND2X1   g23374(.A(new_n25807_), .B(new_n25182_), .Y(new_n25811_));
  OAI21X1  g23375(.A0(new_n22803_), .A1(pi0200), .B0(new_n2953_), .Y(new_n25812_));
  AND2X1   g23376(.A(new_n25812_), .B(new_n23109_), .Y(new_n25813_));
  NAND2X1  g23377(.A(new_n25120_), .B(pi0200), .Y(new_n25814_));
  AOI21X1  g23378(.A0(new_n25814_), .A1(new_n25805_), .B0(new_n25813_), .Y(new_n25815_));
  OAI21X1  g23379(.A0(new_n25815_), .A1(new_n25376_), .B0(new_n8033_), .Y(new_n25816_));
  NOR2X1   g23380(.A(new_n25800_), .B(new_n25350_), .Y(new_n25817_));
  OR4X1    g23381(.A(new_n25817_), .B(new_n25182_), .C(new_n25026_), .D(new_n8033_), .Y(new_n25818_));
  NAND3X1  g23382(.A(new_n25818_), .B(new_n25816_), .C(pi0212), .Y(new_n25819_));
  OAI21X1  g23383(.A0(new_n25819_), .A1(new_n25811_), .B0(new_n23539_), .Y(new_n25820_));
  AOI21X1  g23384(.A0(new_n25810_), .A1(new_n25802_), .B0(new_n25820_), .Y(new_n25821_));
  AND2X1   g23385(.A(new_n6520_), .B(pi1151), .Y(new_n25822_));
  MX2X1    g23386(.A(new_n25815_), .B(new_n25800_), .S0(pi0211), .Y(new_n25823_));
  NOR2X1   g23387(.A(new_n25817_), .B(new_n25323_), .Y(new_n25824_));
  NOR3X1   g23388(.A(new_n25824_), .B(new_n25823_), .C(new_n25376_), .Y(new_n25825_));
  OAI21X1  g23389(.A0(new_n25825_), .A1(new_n23539_), .B0(new_n25822_), .Y(new_n25826_));
  AND2X1   g23390(.A(new_n25342_), .B(new_n25259_), .Y(new_n25827_));
  AND2X1   g23391(.A(new_n25827_), .B(pi1153), .Y(new_n25828_));
  OAI21X1  g23392(.A0(new_n25828_), .A1(new_n25026_), .B0(new_n8548_), .Y(new_n25829_));
  AND2X1   g23393(.A(pi1153), .B(pi0211), .Y(new_n25830_));
  AOI21X1  g23394(.A0(new_n25259_), .A1(new_n8130_), .B0(pi0299), .Y(new_n25831_));
  INVX1    g23395(.A(new_n25831_), .Y(new_n25832_));
  AOI21X1  g23396(.A0(new_n25832_), .A1(new_n25830_), .B0(new_n25014_), .Y(new_n25833_));
  NOR3X1   g23397(.A(new_n25828_), .B(new_n25808_), .C(new_n24962_), .Y(new_n25834_));
  AOI21X1  g23398(.A0(new_n25833_), .A1(new_n25829_), .B0(new_n25834_), .Y(new_n25835_));
  OR2X1    g23399(.A(new_n25835_), .B(pi0219), .Y(new_n25836_));
  INVX1    g23400(.A(pi1151), .Y(new_n25837_));
  NAND3X1  g23401(.A(new_n5117_), .B(new_n25837_), .C(new_n2436_), .Y(new_n25838_));
  NOR2X1   g23402(.A(new_n25831_), .B(new_n9544_), .Y(new_n25839_));
  AOI21X1  g23403(.A0(new_n25342_), .A1(new_n25259_), .B0(pi0214), .Y(new_n25840_));
  NAND2X1  g23404(.A(new_n25840_), .B(new_n24961_), .Y(new_n25841_));
  NAND2X1  g23405(.A(new_n25841_), .B(new_n25839_), .Y(new_n25842_));
  NOR2X1   g23406(.A(new_n25842_), .B(new_n12494_), .Y(new_n25843_));
  NOR2X1   g23407(.A(new_n25843_), .B(new_n25253_), .Y(new_n25844_));
  NOR2X1   g23408(.A(new_n25844_), .B(new_n25838_), .Y(new_n25845_));
  AOI21X1  g23409(.A0(new_n25845_), .A1(new_n25836_), .B0(pi1152), .Y(new_n25846_));
  OAI21X1  g23410(.A0(new_n25826_), .A1(new_n25821_), .B0(new_n25846_), .Y(new_n25847_));
  INVX1    g23411(.A(new_n25253_), .Y(new_n25848_));
  OAI21X1  g23412(.A0(new_n25400_), .A1(new_n8547_), .B0(pi0207), .Y(new_n25849_));
  NAND2X1  g23413(.A(new_n25849_), .B(new_n25587_), .Y(new_n25850_));
  AOI21X1  g23414(.A0(pi0207), .A1(pi0200), .B0(pi0199), .Y(new_n25851_));
  OAI21X1  g23415(.A0(new_n25851_), .A1(pi0299), .B0(pi0208), .Y(new_n25852_));
  NOR3X1   g23416(.A(pi0207), .B(pi0200), .C(pi0199), .Y(new_n25853_));
  OR2X1    g23417(.A(new_n25853_), .B(pi0299), .Y(new_n25854_));
  AOI21X1  g23418(.A0(new_n25854_), .A1(new_n12494_), .B0(new_n25852_), .Y(new_n25855_));
  AOI21X1  g23419(.A0(new_n25850_), .A1(new_n23109_), .B0(new_n25855_), .Y(new_n25856_));
  OR2X1    g23420(.A(new_n25856_), .B(new_n8548_), .Y(new_n25857_));
  MX2X1    g23421(.A(new_n25336_), .B(new_n8131_), .S0(pi0207), .Y(new_n25858_));
  OAI22X1  g23422(.A0(new_n25858_), .A1(new_n23109_), .B0(new_n25336_), .B1(new_n25122_), .Y(new_n25859_));
  NAND3X1  g23423(.A(new_n25859_), .B(new_n25362_), .C(new_n8548_), .Y(new_n25860_));
  AND2X1   g23424(.A(new_n25860_), .B(new_n25857_), .Y(new_n25861_));
  AND2X1   g23425(.A(new_n25007_), .B(pi0299), .Y(new_n25862_));
  AND2X1   g23426(.A(new_n25859_), .B(new_n24963_), .Y(new_n25863_));
  INVX1    g23427(.A(new_n25863_), .Y(new_n25864_));
  OAI22X1  g23428(.A0(new_n25864_), .A1(new_n25862_), .B0(new_n25861_), .B1(new_n25014_), .Y(new_n25865_));
  AOI21X1  g23429(.A0(pi0207), .A1(new_n8009_), .B0(new_n25259_), .Y(new_n25866_));
  NOR2X1   g23430(.A(new_n25866_), .B(new_n8503_), .Y(new_n25867_));
  INVX1    g23431(.A(new_n25867_), .Y(new_n25868_));
  AOI21X1  g23432(.A0(new_n25334_), .A1(new_n7897_), .B0(new_n25868_), .Y(new_n25869_));
  INVX1    g23433(.A(new_n25869_), .Y(new_n25870_));
  NOR3X1   g23434(.A(new_n12494_), .B(new_n2953_), .C(pi0211), .Y(new_n25871_));
  INVX1    g23435(.A(new_n25871_), .Y(new_n25872_));
  OAI21X1  g23436(.A0(new_n25872_), .A1(new_n24955_), .B0(new_n25870_), .Y(new_n25873_));
  AOI22X1  g23437(.A0(new_n25873_), .A1(new_n25848_), .B0(new_n25865_), .B1(new_n23539_), .Y(new_n25874_));
  OAI21X1  g23438(.A0(new_n25377_), .A1(new_n22803_), .B0(new_n25337_), .Y(new_n25875_));
  AOI21X1  g23439(.A0(new_n25337_), .A1(pi0207), .B0(new_n25122_), .Y(new_n25876_));
  AOI21X1  g23440(.A0(new_n25875_), .A1(pi0208), .B0(new_n25876_), .Y(new_n25877_));
  INVX1    g23441(.A(new_n25877_), .Y(new_n25878_));
  NAND3X1  g23442(.A(new_n25878_), .B(new_n25429_), .C(new_n8548_), .Y(new_n25879_));
  NAND3X1  g23443(.A(new_n25878_), .B(new_n25362_), .C(pi0211), .Y(new_n25880_));
  AOI21X1  g23444(.A0(new_n25880_), .A1(new_n25879_), .B0(new_n24962_), .Y(new_n25881_));
  NOR4X1   g23445(.A(new_n25853_), .B(new_n25268_), .C(pi0299), .D(new_n23109_), .Y(new_n25882_));
  AOI21X1  g23446(.A0(new_n25039_), .A1(new_n25159_), .B0(new_n25882_), .Y(new_n25883_));
  INVX1    g23447(.A(new_n25883_), .Y(new_n25884_));
  AOI21X1  g23448(.A0(new_n25832_), .A1(new_n25830_), .B0(new_n25884_), .Y(new_n25885_));
  AOI21X1  g23449(.A0(new_n25885_), .A1(new_n25860_), .B0(new_n25014_), .Y(new_n25886_));
  INVX1    g23450(.A(new_n25828_), .Y(new_n25887_));
  AND2X1   g23451(.A(new_n25883_), .B(new_n24984_), .Y(new_n25888_));
  AOI21X1  g23452(.A0(new_n25888_), .A1(new_n25887_), .B0(pi0212), .Y(new_n25889_));
  AND2X1   g23453(.A(new_n25889_), .B(new_n24984_), .Y(new_n25890_));
  OR4X1    g23454(.A(new_n25890_), .B(new_n25886_), .C(new_n25881_), .D(pi0219), .Y(new_n25891_));
  NOR3X1   g23455(.A(new_n25884_), .B(new_n25843_), .C(new_n23539_), .Y(new_n25892_));
  NOR3X1   g23456(.A(new_n25892_), .B(po1038), .C(new_n25837_), .Y(new_n25893_));
  AOI21X1  g23457(.A0(new_n25893_), .A1(new_n25891_), .B0(new_n25289_), .Y(new_n25894_));
  OAI21X1  g23458(.A0(new_n25874_), .A1(new_n25838_), .B0(new_n25894_), .Y(new_n25895_));
  AOI21X1  g23459(.A0(new_n25895_), .A1(new_n25847_), .B0(pi0209), .Y(new_n25896_));
  NOR3X1   g23460(.A(new_n25393_), .B(new_n25048_), .C(pi0299), .Y(new_n25897_));
  INVX1    g23461(.A(new_n25897_), .Y(new_n25898_));
  NAND2X1  g23462(.A(new_n25898_), .B(new_n25366_), .Y(new_n25899_));
  MX2X1    g23463(.A(new_n25899_), .B(new_n25114_), .S0(new_n22803_), .Y(new_n25900_));
  MX2X1    g23464(.A(new_n25900_), .B(new_n25596_), .S0(new_n23109_), .Y(new_n25901_));
  INVX1    g23465(.A(new_n25366_), .Y(new_n25902_));
  OAI21X1  g23466(.A0(pi1153), .A1(pi0299), .B0(new_n12615_), .Y(new_n25903_));
  OAI21X1  g23467(.A0(new_n25903_), .A1(new_n25107_), .B0(pi0207), .Y(new_n25904_));
  OAI21X1  g23468(.A0(new_n25904_), .A1(new_n25902_), .B0(pi0208), .Y(new_n25905_));
  AOI21X1  g23469(.A0(new_n25430_), .A1(new_n25069_), .B0(new_n25905_), .Y(new_n25906_));
  AOI22X1  g23470(.A0(new_n25906_), .A1(new_n25542_), .B0(new_n25101_), .B1(new_n25238_), .Y(new_n25907_));
  OAI21X1  g23471(.A0(new_n25907_), .A1(pi0211), .B0(new_n25023_), .Y(new_n25908_));
  AOI21X1  g23472(.A0(new_n25901_), .A1(pi0211), .B0(new_n25908_), .Y(new_n25909_));
  AND2X1   g23473(.A(new_n25901_), .B(new_n25180_), .Y(new_n25910_));
  NOR2X1   g23474(.A(new_n25907_), .B(new_n25183_), .Y(new_n25911_));
  OAI21X1  g23475(.A0(new_n25107_), .A1(new_n12494_), .B0(new_n25343_), .Y(new_n25912_));
  MX2X1    g23476(.A(new_n25912_), .B(new_n25590_), .S0(new_n22803_), .Y(new_n25913_));
  AOI21X1  g23477(.A0(new_n25913_), .A1(pi0208), .B0(new_n25589_), .Y(new_n25914_));
  OAI21X1  g23478(.A0(new_n25914_), .A1(new_n25740_), .B0(pi0212), .Y(new_n25915_));
  NOR3X1   g23479(.A(new_n25915_), .B(new_n25911_), .C(new_n25910_), .Y(new_n25916_));
  OAI21X1  g23480(.A0(new_n25916_), .A1(new_n25909_), .B0(new_n23539_), .Y(new_n25917_));
  INVX1    g23481(.A(new_n25536_), .Y(new_n25918_));
  NOR3X1   g23482(.A(new_n25897_), .B(new_n25365_), .C(new_n7897_), .Y(new_n25919_));
  NOR2X1   g23483(.A(new_n25919_), .B(new_n25918_), .Y(new_n25920_));
  NOR2X1   g23484(.A(new_n25914_), .B(pi0211), .Y(new_n25921_));
  AOI21X1  g23485(.A0(new_n25920_), .A1(pi0211), .B0(new_n25921_), .Y(new_n25922_));
  OAI21X1  g23486(.A0(new_n25919_), .A1(new_n25918_), .B0(new_n24984_), .Y(new_n25923_));
  OAI21X1  g23487(.A0(new_n25923_), .A1(pi0212), .B0(new_n6520_), .Y(new_n25924_));
  AOI21X1  g23488(.A0(new_n25922_), .A1(new_n25441_), .B0(new_n25924_), .Y(new_n25925_));
  AOI21X1  g23489(.A0(new_n25925_), .A1(new_n25917_), .B0(new_n23244_), .Y(new_n25926_));
  OAI21X1  g23490(.A0(new_n25926_), .A1(new_n25896_), .B0(new_n25798_), .Y(new_n25927_));
  NAND2X1  g23491(.A(new_n25927_), .B(pi0213), .Y(new_n25928_));
  INVX1    g23492(.A(new_n24958_), .Y(new_n25929_));
  AND2X1   g23493(.A(new_n8033_), .B(pi0212), .Y(new_n25930_));
  NOR4X1   g23494(.A(new_n24955_), .B(new_n8074_), .C(new_n12494_), .D(pi0211), .Y(new_n25931_));
  NOR3X1   g23495(.A(new_n25931_), .B(new_n25930_), .C(pi0219), .Y(new_n25932_));
  OAI21X1  g23496(.A0(new_n25932_), .A1(new_n25929_), .B0(pi1151), .Y(new_n25933_));
  INVX1    g23497(.A(new_n25933_), .Y(new_n25934_));
  AND2X1   g23498(.A(new_n25131_), .B(new_n25159_), .Y(new_n25935_));
  OAI22X1  g23499(.A0(new_n25905_), .A1(new_n25531_), .B0(new_n25935_), .B1(new_n25122_), .Y(new_n25936_));
  MX2X1    g23500(.A(new_n25936_), .B(new_n25920_), .S0(pi0211), .Y(new_n25937_));
  OAI22X1  g23501(.A0(new_n25937_), .A1(new_n24955_), .B0(new_n25923_), .B1(pi0212), .Y(new_n25938_));
  AOI21X1  g23502(.A0(new_n25938_), .A1(pi0219), .B0(po1038), .Y(new_n25939_));
  INVX1    g23503(.A(new_n25920_), .Y(new_n25940_));
  MX2X1    g23504(.A(new_n25922_), .B(new_n25940_), .S0(new_n24984_), .Y(new_n25941_));
  OR2X1    g23505(.A(new_n25922_), .B(pi0214), .Y(new_n25942_));
  MX2X1    g23506(.A(new_n25936_), .B(new_n25920_), .S0(new_n8548_), .Y(new_n25943_));
  AOI21X1  g23507(.A0(new_n25943_), .A1(pi0214), .B0(new_n24961_), .Y(new_n25944_));
  AOI22X1  g23508(.A0(new_n25944_), .A1(new_n25942_), .B0(new_n25941_), .B1(new_n24961_), .Y(new_n25945_));
  OAI21X1  g23509(.A0(new_n25945_), .A1(pi0219), .B0(new_n25939_), .Y(new_n25946_));
  AOI21X1  g23510(.A0(new_n5117_), .A1(new_n2436_), .B0(pi0219), .Y(new_n25947_));
  AOI21X1  g23511(.A0(new_n25931_), .A1(new_n25947_), .B0(pi1151), .Y(new_n25948_));
  INVX1    g23512(.A(new_n25948_), .Y(new_n25949_));
  AND2X1   g23513(.A(new_n25232_), .B(new_n23539_), .Y(new_n25950_));
  OAI21X1  g23514(.A0(new_n25950_), .A1(new_n25920_), .B0(new_n6520_), .Y(new_n25951_));
  AOI21X1  g23515(.A0(new_n25950_), .A1(new_n25922_), .B0(new_n25951_), .Y(new_n25952_));
  OAI21X1  g23516(.A0(new_n25952_), .A1(new_n25949_), .B0(new_n25289_), .Y(new_n25953_));
  AOI21X1  g23517(.A0(new_n25946_), .A1(new_n25934_), .B0(new_n25953_), .Y(new_n25954_));
  NOR4X1   g23518(.A(new_n24955_), .B(new_n25930_), .C(new_n6520_), .D(pi0219), .Y(new_n25955_));
  MX2X1    g23519(.A(new_n25796_), .B(pi0211), .S0(new_n8074_), .Y(new_n25956_));
  INVX1    g23520(.A(new_n25956_), .Y(new_n25957_));
  AOI21X1  g23521(.A0(new_n25957_), .A1(new_n25955_), .B0(pi1151), .Y(new_n25958_));
  INVX1    g23522(.A(new_n25958_), .Y(new_n25959_));
  AOI21X1  g23523(.A0(new_n25936_), .A1(pi0211), .B0(new_n25921_), .Y(new_n25960_));
  NAND2X1  g23524(.A(new_n25960_), .B(pi0214), .Y(new_n25961_));
  AND2X1   g23525(.A(new_n25923_), .B(new_n24961_), .Y(new_n25962_));
  AOI21X1  g23526(.A0(new_n25962_), .A1(new_n25961_), .B0(pi0219), .Y(new_n25963_));
  NOR2X1   g23527(.A(new_n25960_), .B(pi0214), .Y(new_n25964_));
  AOI21X1  g23528(.A0(new_n25937_), .A1(pi0214), .B0(new_n25964_), .Y(new_n25965_));
  OAI21X1  g23529(.A0(new_n25965_), .A1(new_n24961_), .B0(new_n25963_), .Y(new_n25966_));
  AOI21X1  g23530(.A0(new_n25940_), .A1(pi0219), .B0(po1038), .Y(new_n25967_));
  AOI21X1  g23531(.A0(new_n25967_), .A1(new_n25966_), .B0(new_n25959_), .Y(new_n25968_));
  INVX1    g23532(.A(new_n25955_), .Y(new_n25969_));
  NOR3X1   g23533(.A(new_n24957_), .B(new_n8034_), .C(new_n6520_), .Y(new_n25970_));
  NOR2X1   g23534(.A(new_n25970_), .B(new_n25837_), .Y(new_n25971_));
  OAI21X1  g23535(.A0(new_n25956_), .A1(new_n25969_), .B0(new_n25971_), .Y(new_n25972_));
  AOI21X1  g23536(.A0(new_n25936_), .A1(pi0214), .B0(new_n25964_), .Y(new_n25973_));
  OAI21X1  g23537(.A0(new_n25973_), .A1(new_n24961_), .B0(new_n25963_), .Y(new_n25974_));
  AOI21X1  g23538(.A0(new_n25974_), .A1(new_n25939_), .B0(new_n25972_), .Y(new_n25975_));
  NOR3X1   g23539(.A(new_n25975_), .B(new_n25968_), .C(new_n25289_), .Y(new_n25976_));
  NOR3X1   g23540(.A(new_n25976_), .B(new_n25954_), .C(new_n23244_), .Y(new_n25977_));
  NOR3X1   g23541(.A(new_n25823_), .B(new_n25376_), .C(pi0214), .Y(new_n25978_));
  AOI21X1  g23542(.A0(new_n25827_), .A1(pi1153), .B0(new_n9544_), .Y(new_n25979_));
  INVX1    g23543(.A(new_n25979_), .Y(new_n25980_));
  OAI21X1  g23544(.A0(new_n25980_), .A1(new_n25817_), .B0(pi0214), .Y(new_n25981_));
  NAND2X1  g23545(.A(new_n25981_), .B(pi0212), .Y(new_n25982_));
  OAI22X1  g23546(.A0(new_n25982_), .A1(new_n25978_), .B0(new_n25825_), .B1(pi0212), .Y(new_n25983_));
  AND2X1   g23547(.A(pi0299), .B(new_n8548_), .Y(new_n25984_));
  NOR3X1   g23548(.A(new_n25984_), .B(new_n25828_), .C(new_n25817_), .Y(new_n25985_));
  NOR2X1   g23549(.A(new_n25985_), .B(new_n25824_), .Y(new_n25986_));
  OAI21X1  g23550(.A0(new_n25986_), .A1(new_n23539_), .B0(new_n6520_), .Y(new_n25987_));
  AOI21X1  g23551(.A0(new_n25983_), .A1(new_n23539_), .B0(new_n25987_), .Y(new_n25988_));
  OR2X1    g23552(.A(new_n25988_), .B(new_n25933_), .Y(new_n25989_));
  NAND4X1  g23553(.A(new_n25840_), .B(new_n25839_), .C(pi1153), .D(pi0212), .Y(new_n25990_));
  NOR3X1   g23554(.A(new_n25979_), .B(new_n25840_), .C(new_n24961_), .Y(new_n25991_));
  NOR2X1   g23555(.A(new_n25991_), .B(pi0219), .Y(new_n25992_));
  AOI21X1  g23556(.A0(new_n25871_), .A1(new_n25023_), .B0(new_n25827_), .Y(new_n25993_));
  NAND3X1  g23557(.A(new_n25993_), .B(new_n25992_), .C(new_n25990_), .Y(new_n25994_));
  INVX1    g23558(.A(new_n25827_), .Y(new_n25995_));
  AOI21X1  g23559(.A0(new_n25995_), .A1(pi0219), .B0(po1038), .Y(new_n25996_));
  NAND3X1  g23560(.A(new_n25996_), .B(new_n25994_), .C(new_n25843_), .Y(new_n25997_));
  AOI21X1  g23561(.A0(new_n25997_), .A1(new_n25948_), .B0(pi1152), .Y(new_n25998_));
  INVX1    g23562(.A(new_n25972_), .Y(new_n25999_));
  AND2X1   g23563(.A(new_n25883_), .B(new_n25887_), .Y(new_n26000_));
  OAI21X1  g23564(.A0(new_n25877_), .A1(pi0211), .B0(new_n26000_), .Y(new_n26001_));
  NAND2X1  g23565(.A(new_n25888_), .B(new_n25887_), .Y(new_n26002_));
  OAI21X1  g23566(.A0(new_n26001_), .A1(new_n24984_), .B0(new_n26002_), .Y(new_n26003_));
  NAND2X1  g23567(.A(new_n26003_), .B(new_n24961_), .Y(new_n26004_));
  AOI21X1  g23568(.A0(new_n26004_), .A1(new_n26001_), .B0(new_n23539_), .Y(new_n26005_));
  NOR2X1   g23569(.A(new_n26005_), .B(po1038), .Y(new_n26006_));
  INVX1    g23570(.A(new_n26006_), .Y(new_n26007_));
  INVX1    g23571(.A(new_n25889_), .Y(new_n26008_));
  AOI22X1  g23572(.A0(new_n25878_), .A1(pi0211), .B0(new_n25832_), .B1(pi1153), .Y(new_n26009_));
  AND2X1   g23573(.A(new_n25883_), .B(pi0214), .Y(new_n26010_));
  AOI21X1  g23574(.A0(new_n26010_), .A1(new_n26009_), .B0(new_n26008_), .Y(new_n26011_));
  AND2X1   g23575(.A(new_n26009_), .B(new_n25888_), .Y(new_n26012_));
  AND2X1   g23576(.A(new_n25877_), .B(pi0214), .Y(new_n26013_));
  NOR3X1   g23577(.A(new_n26013_), .B(new_n26012_), .C(new_n24961_), .Y(new_n26014_));
  NOR3X1   g23578(.A(new_n26014_), .B(new_n26011_), .C(pi0219), .Y(new_n26015_));
  OAI21X1  g23579(.A0(new_n26015_), .A1(new_n26007_), .B0(new_n25999_), .Y(new_n26016_));
  AOI21X1  g23580(.A0(new_n25870_), .A1(pi0219), .B0(po1038), .Y(new_n26017_));
  AOI21X1  g23581(.A0(new_n25856_), .A1(new_n8548_), .B0(new_n25864_), .Y(new_n26018_));
  AOI21X1  g23582(.A0(new_n25392_), .A1(pi0299), .B0(pi0219), .Y(new_n26019_));
  OAI21X1  g23583(.A0(new_n25870_), .A1(new_n25232_), .B0(new_n26019_), .Y(new_n26020_));
  OAI21X1  g23584(.A0(new_n26020_), .A1(new_n26018_), .B0(new_n26017_), .Y(new_n26021_));
  AOI21X1  g23585(.A0(new_n26021_), .A1(new_n25958_), .B0(new_n25289_), .Y(new_n26022_));
  AOI22X1  g23586(.A0(new_n26022_), .A1(new_n26016_), .B0(new_n25998_), .B1(new_n25989_), .Y(new_n26023_));
  AND2X1   g23587(.A(new_n26023_), .B(new_n23244_), .Y(new_n26024_));
  OR2X1    g23588(.A(new_n26024_), .B(pi0213), .Y(new_n26025_));
  OAI21X1  g23589(.A0(new_n26025_), .A1(new_n25977_), .B0(new_n25928_), .Y(new_n26026_));
  MX2X1    g23590(.A(new_n26026_), .B(pi0238), .S0(new_n24954_), .Y(po0395));
  INVX1    g23591(.A(new_n24980_), .Y(new_n26028_));
  NOR2X1   g23592(.A(new_n25066_), .B(new_n26028_), .Y(new_n26029_));
  AOI21X1  g23593(.A0(new_n26029_), .A1(new_n24984_), .B0(pi0212), .Y(new_n26030_));
  AND2X1   g23594(.A(new_n26030_), .B(new_n23539_), .Y(new_n26031_));
  INVX1    g23595(.A(new_n26031_), .Y(new_n26032_));
  AND2X1   g23596(.A(pi1158), .B(pi0299), .Y(new_n26033_));
  AOI22X1  g23597(.A0(new_n26033_), .A1(new_n26028_), .B0(new_n25719_), .B1(new_n23109_), .Y(new_n26034_));
  OR2X1    g23598(.A(new_n25274_), .B(new_n25122_), .Y(new_n26035_));
  AOI21X1  g23599(.A0(pi0299), .A1(pi0208), .B0(new_n12706_), .Y(new_n26036_));
  AND2X1   g23600(.A(new_n26036_), .B(new_n26035_), .Y(new_n26037_));
  OAI21X1  g23601(.A0(new_n26029_), .A1(pi1157), .B0(pi0211), .Y(new_n26038_));
  OAI22X1  g23602(.A0(new_n26038_), .A1(new_n26037_), .B0(new_n26034_), .B1(pi0211), .Y(new_n26039_));
  AOI21X1  g23603(.A0(new_n26039_), .A1(pi0214), .B0(new_n26032_), .Y(new_n26040_));
  AND2X1   g23604(.A(new_n26030_), .B(pi0219), .Y(new_n26041_));
  INVX1    g23605(.A(new_n26029_), .Y(new_n26042_));
  AOI21X1  g23606(.A0(new_n26042_), .A1(pi0211), .B0(new_n24984_), .Y(new_n26043_));
  INVX1    g23607(.A(new_n26043_), .Y(new_n26044_));
  NOR3X1   g23608(.A(new_n25303_), .B(new_n25166_), .C(pi0211), .Y(new_n26045_));
  OAI21X1  g23609(.A0(new_n26045_), .A1(new_n26044_), .B0(new_n26041_), .Y(new_n26046_));
  AOI21X1  g23610(.A0(new_n26042_), .A1(pi0212), .B0(po1038), .Y(new_n26047_));
  NAND3X1  g23611(.A(new_n26047_), .B(new_n26046_), .C(new_n23244_), .Y(new_n26048_));
  NOR4X1   g23612(.A(new_n25698_), .B(new_n25669_), .C(new_n25666_), .D(pi0208), .Y(new_n26049_));
  INVX1    g23613(.A(new_n26049_), .Y(new_n26050_));
  OAI21X1  g23614(.A0(new_n26050_), .A1(pi0214), .B0(new_n24961_), .Y(new_n26051_));
  NOR2X1   g23615(.A(new_n26051_), .B(pi0219), .Y(new_n26052_));
  NAND2X1  g23616(.A(new_n25724_), .B(new_n25723_), .Y(new_n26053_));
  MX2X1    g23617(.A(new_n26033_), .B(new_n12706_), .S0(new_n23109_), .Y(new_n26054_));
  AOI21X1  g23618(.A0(new_n26054_), .A1(new_n26053_), .B0(new_n25736_), .Y(new_n26055_));
  INVX1    g23619(.A(new_n25713_), .Y(new_n26056_));
  AOI21X1  g23620(.A0(new_n26036_), .A1(new_n26056_), .B0(new_n25698_), .Y(new_n26057_));
  OAI21X1  g23621(.A0(new_n26057_), .A1(new_n8548_), .B0(pi0214), .Y(new_n26058_));
  OAI21X1  g23622(.A0(new_n26058_), .A1(new_n26055_), .B0(new_n26052_), .Y(new_n26059_));
  NOR2X1   g23623(.A(new_n26051_), .B(new_n23539_), .Y(new_n26060_));
  AOI21X1  g23624(.A0(new_n26050_), .A1(new_n25436_), .B0(new_n24984_), .Y(new_n26061_));
  OAI21X1  g23625(.A0(new_n26049_), .A1(new_n8548_), .B0(new_n26061_), .Y(new_n26062_));
  AOI21X1  g23626(.A0(new_n26050_), .A1(pi0212), .B0(po1038), .Y(new_n26063_));
  NAND2X1  g23627(.A(new_n26063_), .B(pi0209), .Y(new_n26064_));
  AOI21X1  g23628(.A0(new_n26062_), .A1(new_n26060_), .B0(new_n26064_), .Y(new_n26065_));
  AND2X1   g23629(.A(new_n25623_), .B(new_n23539_), .Y(new_n26066_));
  OAI21X1  g23630(.A0(new_n26066_), .A1(new_n25626_), .B0(pi0213), .Y(new_n26067_));
  AOI21X1  g23631(.A0(new_n26065_), .A1(new_n26059_), .B0(new_n26067_), .Y(new_n26068_));
  OAI21X1  g23632(.A0(new_n26048_), .A1(new_n26040_), .B0(new_n26068_), .Y(new_n26069_));
  OR2X1    g23633(.A(new_n25024_), .B(new_n8548_), .Y(new_n26070_));
  OAI21X1  g23634(.A0(new_n26070_), .A1(new_n25771_), .B0(new_n26061_), .Y(new_n26071_));
  NAND2X1  g23635(.A(new_n26071_), .B(new_n26052_), .Y(new_n26072_));
  INVX1    g23636(.A(new_n26063_), .Y(new_n26073_));
  OR2X1    g23637(.A(new_n25026_), .B(pi0211), .Y(new_n26074_));
  AOI21X1  g23638(.A0(new_n26050_), .A1(pi0211), .B0(new_n24984_), .Y(new_n26075_));
  OAI21X1  g23639(.A0(new_n26074_), .A1(new_n25771_), .B0(new_n26075_), .Y(new_n26076_));
  AOI21X1  g23640(.A0(new_n26076_), .A1(new_n26060_), .B0(new_n26073_), .Y(new_n26077_));
  AOI21X1  g23641(.A0(new_n26077_), .A1(new_n26072_), .B0(new_n23244_), .Y(new_n26078_));
  OAI21X1  g23642(.A0(new_n25267_), .A1(new_n25026_), .B0(new_n26043_), .Y(new_n26079_));
  NAND2X1  g23643(.A(new_n26079_), .B(new_n26041_), .Y(new_n26080_));
  OAI21X1  g23644(.A0(new_n26070_), .A1(new_n25307_), .B0(pi0214), .Y(new_n26081_));
  OAI21X1  g23645(.A0(new_n26081_), .A1(new_n26045_), .B0(new_n26031_), .Y(new_n26082_));
  NAND3X1  g23646(.A(new_n26082_), .B(new_n26080_), .C(new_n26047_), .Y(new_n26083_));
  AOI21X1  g23647(.A0(new_n26083_), .A1(new_n23244_), .B0(new_n26078_), .Y(new_n26084_));
  OR2X1    g23648(.A(new_n25474_), .B(new_n6520_), .Y(new_n26085_));
  OAI21X1  g23649(.A0(new_n25472_), .A1(pi0219), .B0(new_n25023_), .Y(new_n26086_));
  OAI21X1  g23650(.A0(new_n26086_), .A1(new_n26085_), .B0(new_n25003_), .Y(new_n26087_));
  OAI21X1  g23651(.A0(new_n26087_), .A1(new_n26084_), .B0(new_n26069_), .Y(new_n26088_));
  NOR2X1   g23652(.A(pi0239), .B(pi0230), .Y(new_n26089_));
  AOI21X1  g23653(.A0(new_n26088_), .A1(pi0230), .B0(new_n26089_), .Y(po0396));
  INVX1    g23654(.A(pi1147), .Y(new_n26091_));
  INVX1    g23655(.A(new_n25996_), .Y(new_n26092_));
  NOR4X1   g23656(.A(new_n25866_), .B(new_n8503_), .C(new_n5118_), .D(pi0057), .Y(new_n26093_));
  INVX1    g23657(.A(new_n26093_), .Y(new_n26094_));
  NOR2X1   g23658(.A(new_n25867_), .B(pi0214), .Y(new_n26095_));
  NOR2X1   g23659(.A(new_n26095_), .B(pi0212), .Y(new_n26096_));
  NOR4X1   g23660(.A(pi0299), .B(pi0208), .C(new_n22803_), .D(pi0199), .Y(new_n26097_));
  INVX1    g23661(.A(new_n26097_), .Y(new_n26098_));
  NAND4X1  g23662(.A(new_n26098_), .B(new_n25852_), .C(new_n2953_), .D(pi0214), .Y(new_n26099_));
  AOI21X1  g23663(.A0(new_n26099_), .A1(new_n26096_), .B0(pi0219), .Y(new_n26100_));
  NAND3X1  g23664(.A(new_n26098_), .B(new_n25852_), .C(new_n2953_), .Y(new_n26101_));
  AND2X1   g23665(.A(new_n26101_), .B(new_n8548_), .Y(new_n26102_));
  NOR3X1   g23666(.A(new_n25866_), .B(new_n8503_), .C(new_n8548_), .Y(new_n26103_));
  NOR3X1   g23667(.A(new_n26103_), .B(new_n26102_), .C(new_n24984_), .Y(new_n26104_));
  NOR2X1   g23668(.A(new_n26104_), .B(new_n24961_), .Y(new_n26105_));
  NAND2X1  g23669(.A(new_n26105_), .B(new_n26101_), .Y(new_n26106_));
  AOI22X1  g23670(.A0(new_n26106_), .A1(new_n26100_), .B0(new_n26094_), .B1(new_n26092_), .Y(new_n26107_));
  NOR2X1   g23671(.A(new_n26107_), .B(new_n25955_), .Y(new_n26108_));
  NAND2X1  g23672(.A(new_n26108_), .B(new_n26091_), .Y(new_n26109_));
  AOI22X1  g23673(.A0(new_n5117_), .A1(new_n2436_), .B0(pi0219), .B1(pi0211), .Y(new_n26110_));
  AND2X1   g23674(.A(new_n26110_), .B(new_n25323_), .Y(new_n26111_));
  NOR2X1   g23675(.A(new_n24955_), .B(new_n2953_), .Y(new_n26112_));
  INVX1    g23676(.A(new_n26112_), .Y(new_n26113_));
  NOR3X1   g23677(.A(new_n26113_), .B(new_n24957_), .C(po1038), .Y(new_n26114_));
  NOR3X1   g23678(.A(new_n25349_), .B(new_n25268_), .C(pi0299), .Y(new_n26115_));
  AND2X1   g23679(.A(new_n26115_), .B(new_n6520_), .Y(new_n26116_));
  OR4X1    g23680(.A(new_n26116_), .B(new_n26114_), .C(new_n26111_), .D(new_n26091_), .Y(new_n26117_));
  NAND3X1  g23681(.A(new_n26117_), .B(new_n26109_), .C(pi1149), .Y(new_n26118_));
  NOR3X1   g23682(.A(new_n24984_), .B(pi0212), .C(new_n8548_), .Y(new_n26119_));
  AOI21X1  g23683(.A0(new_n25180_), .A1(pi0212), .B0(new_n26119_), .Y(new_n26120_));
  NOR3X1   g23684(.A(new_n26120_), .B(new_n6520_), .C(pi0219), .Y(new_n26121_));
  INVX1    g23685(.A(new_n25135_), .Y(new_n26122_));
  OAI22X1  g23686(.A0(new_n25396_), .A1(new_n25259_), .B0(new_n26122_), .B1(new_n7896_), .Y(new_n26123_));
  NOR2X1   g23687(.A(new_n26123_), .B(new_n25854_), .Y(new_n26124_));
  AND2X1   g23688(.A(new_n8033_), .B(pi0299), .Y(new_n26125_));
  OAI21X1  g23689(.A0(new_n26125_), .A1(new_n26124_), .B0(new_n24961_), .Y(new_n26126_));
  NAND2X1  g23690(.A(new_n26126_), .B(new_n23539_), .Y(new_n26127_));
  AOI21X1  g23691(.A0(new_n26123_), .A1(new_n2953_), .B0(new_n24984_), .Y(new_n26128_));
  AOI21X1  g23692(.A0(new_n26124_), .A1(new_n24984_), .B0(pi0212), .Y(new_n26129_));
  INVX1    g23693(.A(new_n26129_), .Y(new_n26130_));
  AND2X1   g23694(.A(new_n26123_), .B(new_n2953_), .Y(new_n26131_));
  INVX1    g23695(.A(new_n26131_), .Y(new_n26132_));
  AOI21X1  g23696(.A0(new_n26132_), .A1(new_n8548_), .B0(new_n26124_), .Y(new_n26133_));
  OR2X1    g23697(.A(new_n26133_), .B(new_n24984_), .Y(new_n26134_));
  AND2X1   g23698(.A(new_n26134_), .B(pi0212), .Y(new_n26135_));
  OAI21X1  g23699(.A0(new_n26131_), .A1(pi0214), .B0(new_n26135_), .Y(new_n26136_));
  OAI21X1  g23700(.A0(new_n26130_), .A1(new_n26128_), .B0(new_n26136_), .Y(new_n26137_));
  INVX1    g23701(.A(new_n26137_), .Y(new_n26138_));
  NOR3X1   g23702(.A(new_n26128_), .B(new_n26124_), .C(new_n9544_), .Y(new_n26139_));
  NOR2X1   g23703(.A(new_n26139_), .B(new_n24961_), .Y(new_n26140_));
  AOI21X1  g23704(.A0(new_n26140_), .A1(new_n26138_), .B0(new_n26127_), .Y(new_n26141_));
  OAI21X1  g23705(.A0(new_n26123_), .A1(new_n25854_), .B0(pi0219), .Y(new_n26142_));
  AND2X1   g23706(.A(new_n26142_), .B(new_n6520_), .Y(new_n26143_));
  INVX1    g23707(.A(new_n26143_), .Y(new_n26144_));
  NOR2X1   g23708(.A(new_n26144_), .B(new_n26141_), .Y(new_n26145_));
  NOR3X1   g23709(.A(new_n26145_), .B(new_n26121_), .C(pi1147), .Y(new_n26146_));
  INVX1    g23710(.A(pi1149), .Y(new_n26147_));
  NOR2X1   g23711(.A(new_n25182_), .B(new_n24961_), .Y(new_n26148_));
  NOR3X1   g23712(.A(new_n26148_), .B(new_n26119_), .C(pi0219), .Y(new_n26149_));
  NOR4X1   g23713(.A(new_n26149_), .B(new_n26113_), .C(new_n24957_), .D(po1038), .Y(new_n26150_));
  NOR2X1   g23714(.A(new_n25883_), .B(po1038), .Y(new_n26151_));
  NOR3X1   g23715(.A(new_n26149_), .B(new_n24957_), .C(new_n6520_), .Y(new_n26152_));
  NOR3X1   g23716(.A(new_n26152_), .B(new_n26151_), .C(new_n26150_), .Y(new_n26153_));
  INVX1    g23717(.A(new_n26153_), .Y(new_n26154_));
  OAI21X1  g23718(.A0(new_n26154_), .A1(new_n26091_), .B0(new_n26147_), .Y(new_n26155_));
  OAI21X1  g23719(.A0(new_n26155_), .A1(new_n26146_), .B0(new_n26118_), .Y(new_n26156_));
  AND2X1   g23720(.A(new_n25232_), .B(new_n8548_), .Y(new_n26157_));
  NOR3X1   g23721(.A(new_n26157_), .B(new_n25930_), .C(pi0219), .Y(new_n26158_));
  NOR3X1   g23722(.A(new_n26158_), .B(new_n24957_), .C(new_n6520_), .Y(new_n26159_));
  INVX1    g23723(.A(new_n25815_), .Y(new_n26160_));
  AOI21X1  g23724(.A0(new_n26160_), .A1(pi0211), .B0(new_n24984_), .Y(new_n26161_));
  OAI21X1  g23725(.A0(new_n25800_), .A1(pi0211), .B0(new_n26161_), .Y(new_n26162_));
  AND2X1   g23726(.A(new_n26162_), .B(new_n8074_), .Y(new_n26163_));
  AOI21X1  g23727(.A0(new_n25800_), .A1(new_n24984_), .B0(pi0212), .Y(new_n26164_));
  INVX1    g23728(.A(new_n26164_), .Y(new_n26165_));
  AOI21X1  g23729(.A0(new_n25823_), .A1(pi0214), .B0(new_n26165_), .Y(new_n26166_));
  NOR2X1   g23730(.A(new_n26166_), .B(pi0219), .Y(new_n26167_));
  NAND2X1  g23731(.A(new_n26162_), .B(pi0212), .Y(new_n26168_));
  OAI21X1  g23732(.A0(new_n26168_), .A1(new_n25823_), .B0(new_n26167_), .Y(new_n26169_));
  NOR2X1   g23733(.A(new_n26169_), .B(new_n26163_), .Y(new_n26170_));
  INVX1    g23734(.A(new_n26166_), .Y(new_n26171_));
  INVX1    g23735(.A(new_n25823_), .Y(new_n26172_));
  AOI21X1  g23736(.A0(new_n26172_), .A1(pi0212), .B0(new_n23539_), .Y(new_n26173_));
  AOI21X1  g23737(.A0(new_n26173_), .A1(new_n26171_), .B0(po1038), .Y(new_n26174_));
  INVX1    g23738(.A(new_n26174_), .Y(new_n26175_));
  NOR2X1   g23739(.A(new_n26175_), .B(new_n26170_), .Y(new_n26176_));
  NOR3X1   g23740(.A(new_n26176_), .B(new_n26159_), .C(new_n26091_), .Y(new_n26177_));
  INVX1    g23741(.A(new_n25259_), .Y(new_n26178_));
  NOR4X1   g23742(.A(new_n26178_), .B(new_n8135_), .C(po1038), .D(pi0299), .Y(new_n26179_));
  AOI21X1  g23743(.A0(new_n6520_), .A1(new_n2953_), .B0(pi0219), .Y(new_n26180_));
  AND2X1   g23744(.A(new_n26180_), .B(new_n26157_), .Y(new_n26181_));
  NOR2X1   g23745(.A(new_n26181_), .B(new_n26179_), .Y(new_n26182_));
  INVX1    g23746(.A(new_n26182_), .Y(new_n26183_));
  OAI21X1  g23747(.A0(new_n26183_), .A1(pi1147), .B0(pi1149), .Y(new_n26184_));
  AOI21X1  g23748(.A0(new_n8033_), .A1(pi0299), .B0(pi0212), .Y(new_n26185_));
  INVX1    g23749(.A(new_n25984_), .Y(new_n26186_));
  OAI21X1  g23750(.A0(new_n26186_), .A1(new_n24984_), .B0(new_n25883_), .Y(new_n26187_));
  INVX1    g23751(.A(new_n26187_), .Y(new_n26188_));
  AOI21X1  g23752(.A0(new_n9544_), .A1(new_n24984_), .B0(new_n24961_), .Y(new_n26189_));
  AOI22X1  g23753(.A0(new_n26189_), .A1(new_n26188_), .B0(new_n26185_), .B1(new_n25883_), .Y(new_n26190_));
  OR2X1    g23754(.A(new_n26190_), .B(pi0219), .Y(new_n26191_));
  AND2X1   g23755(.A(pi0207), .B(pi0200), .Y(new_n26192_));
  OAI21X1  g23756(.A0(new_n26192_), .A1(new_n25130_), .B0(pi0208), .Y(new_n26193_));
  AOI21X1  g23757(.A0(new_n26193_), .A1(new_n7941_), .B0(new_n25883_), .Y(new_n26194_));
  NOR2X1   g23758(.A(new_n26194_), .B(pi0299), .Y(new_n26195_));
  INVX1    g23759(.A(new_n26195_), .Y(new_n26196_));
  OAI21X1  g23760(.A0(new_n26196_), .A1(pi0219), .B0(new_n26191_), .Y(new_n26197_));
  NAND2X1  g23761(.A(new_n26197_), .B(new_n8548_), .Y(new_n26198_));
  INVX1    g23762(.A(new_n9544_), .Y(new_n26199_));
  NAND3X1  g23763(.A(new_n25883_), .B(new_n26199_), .C(pi0214), .Y(new_n26200_));
  AND2X1   g23764(.A(new_n26186_), .B(new_n25883_), .Y(new_n26201_));
  AOI21X1  g23765(.A0(new_n26201_), .A1(new_n24984_), .B0(new_n24961_), .Y(new_n26202_));
  AND2X1   g23766(.A(new_n26202_), .B(new_n26200_), .Y(new_n26203_));
  AOI21X1  g23767(.A0(new_n26187_), .A1(new_n24961_), .B0(pi0219), .Y(new_n26204_));
  INVX1    g23768(.A(new_n26204_), .Y(new_n26205_));
  NOR2X1   g23769(.A(new_n26205_), .B(new_n26203_), .Y(new_n26206_));
  NOR2X1   g23770(.A(new_n24957_), .B(po1038), .Y(new_n26207_));
  INVX1    g23771(.A(new_n26207_), .Y(new_n26208_));
  AOI21X1  g23772(.A0(new_n26186_), .A1(pi0219), .B0(new_n26208_), .Y(new_n26209_));
  NOR2X1   g23773(.A(new_n26209_), .B(new_n26151_), .Y(new_n26210_));
  NOR3X1   g23774(.A(new_n26210_), .B(new_n26206_), .C(new_n26195_), .Y(new_n26211_));
  AOI21X1  g23775(.A0(new_n26211_), .A1(new_n26198_), .B0(new_n25970_), .Y(new_n26212_));
  OR2X1    g23776(.A(pi1149), .B(new_n26091_), .Y(new_n26213_));
  OAI22X1  g23777(.A0(new_n26213_), .A1(new_n26212_), .B0(new_n26184_), .B1(new_n26177_), .Y(new_n26214_));
  MX2X1    g23778(.A(new_n26214_), .B(new_n26156_), .S0(pi1148), .Y(new_n26215_));
  AND2X1   g23779(.A(pi1146), .B(pi0211), .Y(new_n26216_));
  MX2X1    g23780(.A(new_n3165_), .B(new_n3346_), .S0(pi0211), .Y(new_n26217_));
  INVX1    g23781(.A(new_n26216_), .Y(new_n26218_));
  MX2X1    g23782(.A(new_n26218_), .B(new_n26217_), .S0(pi0214), .Y(new_n26219_));
  NOR2X1   g23783(.A(new_n26219_), .B(new_n24961_), .Y(new_n26220_));
  AOI21X1  g23784(.A0(new_n26216_), .A1(new_n25023_), .B0(new_n26220_), .Y(new_n26221_));
  AND2X1   g23785(.A(pi1145), .B(new_n8548_), .Y(new_n26222_));
  OAI22X1  g23786(.A0(new_n26222_), .A1(new_n23539_), .B0(new_n5118_), .B1(pi0057), .Y(new_n26223_));
  AOI21X1  g23787(.A0(new_n26221_), .A1(new_n25442_), .B0(new_n26223_), .Y(new_n26224_));
  NOR4X1   g23788(.A(new_n24955_), .B(new_n8328_), .C(new_n6520_), .D(pi0219), .Y(new_n26225_));
  OR2X1    g23789(.A(new_n26225_), .B(new_n26091_), .Y(new_n26226_));
  NOR2X1   g23790(.A(new_n26226_), .B(new_n26224_), .Y(new_n26227_));
  INVX1    g23791(.A(new_n26227_), .Y(new_n26228_));
  AND2X1   g23792(.A(new_n25751_), .B(new_n8548_), .Y(new_n26229_));
  INVX1    g23793(.A(new_n26229_), .Y(new_n26230_));
  AOI21X1  g23794(.A0(new_n26230_), .A1(pi0219), .B0(new_n26208_), .Y(new_n26231_));
  OR2X1    g23795(.A(new_n26231_), .B(new_n26151_), .Y(new_n26232_));
  NOR2X1   g23796(.A(new_n26217_), .B(new_n2953_), .Y(new_n26233_));
  INVX1    g23797(.A(new_n26233_), .Y(new_n26234_));
  AOI21X1  g23798(.A0(new_n26234_), .A1(new_n25883_), .B0(new_n25014_), .Y(new_n26235_));
  OAI21X1  g23799(.A0(pi1146), .A1(new_n8548_), .B0(pi0299), .Y(new_n26236_));
  AOI21X1  g23800(.A0(new_n26236_), .A1(new_n25883_), .B0(new_n25516_), .Y(new_n26237_));
  NOR2X1   g23801(.A(new_n25883_), .B(new_n25323_), .Y(new_n26238_));
  OR4X1    g23802(.A(new_n26238_), .B(new_n26237_), .C(new_n26235_), .D(pi0219), .Y(new_n26239_));
  AND2X1   g23803(.A(new_n26239_), .B(new_n26232_), .Y(new_n26240_));
  NOR3X1   g23804(.A(new_n26123_), .B(new_n25854_), .C(po1038), .Y(new_n26241_));
  INVX1    g23805(.A(new_n26241_), .Y(new_n26242_));
  NOR2X1   g23806(.A(new_n26224_), .B(pi1147), .Y(new_n26243_));
  NOR3X1   g23807(.A(new_n26221_), .B(new_n23540_), .C(new_n2953_), .Y(new_n26244_));
  AOI21X1  g23808(.A0(new_n26231_), .A1(pi0219), .B0(new_n26244_), .Y(new_n26245_));
  NAND3X1  g23809(.A(new_n26245_), .B(new_n26243_), .C(new_n26242_), .Y(new_n26246_));
  AND2X1   g23810(.A(new_n26246_), .B(pi1148), .Y(new_n26247_));
  OAI21X1  g23811(.A0(new_n26240_), .A1(new_n26228_), .B0(new_n26247_), .Y(new_n26248_));
  AOI21X1  g23812(.A0(new_n9544_), .A1(new_n3165_), .B0(new_n25516_), .Y(new_n26249_));
  NOR2X1   g23813(.A(new_n26195_), .B(pi0219), .Y(new_n26250_));
  OAI21X1  g23814(.A0(new_n26249_), .A1(new_n26235_), .B0(new_n26250_), .Y(new_n26251_));
  INVX1    g23815(.A(new_n26222_), .Y(new_n26252_));
  NOR3X1   g23816(.A(new_n26252_), .B(new_n25442_), .C(new_n2953_), .Y(new_n26253_));
  AOI21X1  g23817(.A0(new_n26194_), .A1(new_n25848_), .B0(new_n26253_), .Y(new_n26254_));
  AOI21X1  g23818(.A0(new_n26254_), .A1(new_n26251_), .B0(po1038), .Y(new_n26255_));
  AOI21X1  g23819(.A0(new_n26245_), .A1(new_n26243_), .B0(pi1148), .Y(new_n26256_));
  OAI21X1  g23820(.A0(new_n26255_), .A1(new_n26228_), .B0(new_n26256_), .Y(new_n26257_));
  AOI21X1  g23821(.A0(new_n26257_), .A1(new_n26248_), .B0(pi1149), .Y(new_n26258_));
  AOI21X1  g23822(.A0(new_n25800_), .A1(pi0219), .B0(po1038), .Y(new_n26259_));
  OR2X1    g23823(.A(new_n26259_), .B(new_n26231_), .Y(new_n26260_));
  AND2X1   g23824(.A(pi1146), .B(pi0299), .Y(new_n26261_));
  INVX1    g23825(.A(new_n26261_), .Y(new_n26262_));
  NAND3X1  g23826(.A(new_n25814_), .B(new_n25805_), .C(new_n2953_), .Y(new_n26263_));
  NAND3X1  g23827(.A(new_n26263_), .B(new_n26262_), .C(new_n25659_), .Y(new_n26264_));
  MX2X1    g23828(.A(new_n26264_), .B(new_n26160_), .S0(new_n8548_), .Y(new_n26265_));
  OAI21X1  g23829(.A0(new_n26265_), .A1(new_n24984_), .B0(new_n26164_), .Y(new_n26266_));
  NOR2X1   g23830(.A(new_n26233_), .B(new_n24984_), .Y(new_n26267_));
  NAND3X1  g23831(.A(new_n26267_), .B(new_n26263_), .C(new_n25659_), .Y(new_n26268_));
  AND2X1   g23832(.A(new_n26268_), .B(pi0212), .Y(new_n26269_));
  OAI21X1  g23833(.A0(new_n26265_), .A1(pi0214), .B0(new_n26269_), .Y(new_n26270_));
  NAND3X1  g23834(.A(new_n26270_), .B(new_n26266_), .C(new_n23539_), .Y(new_n26271_));
  AOI21X1  g23835(.A0(new_n26271_), .A1(new_n26260_), .B0(new_n26228_), .Y(new_n26272_));
  INVX1    g23836(.A(pi1148), .Y(new_n26273_));
  INVX1    g23837(.A(new_n26179_), .Y(new_n26274_));
  NAND3X1  g23838(.A(new_n26245_), .B(new_n26243_), .C(new_n26274_), .Y(new_n26275_));
  NAND2X1  g23839(.A(new_n26275_), .B(new_n26273_), .Y(new_n26276_));
  OAI21X1  g23840(.A0(new_n25868_), .A1(new_n24956_), .B0(pi0219), .Y(new_n26277_));
  AOI21X1  g23841(.A0(new_n26102_), .A1(new_n25323_), .B0(new_n26277_), .Y(new_n26278_));
  NOR2X1   g23842(.A(new_n26278_), .B(po1038), .Y(new_n26279_));
  AOI21X1  g23843(.A0(new_n26279_), .A1(new_n8502_), .B0(new_n26231_), .Y(new_n26280_));
  INVX1    g23844(.A(new_n26096_), .Y(new_n26281_));
  NAND3X1  g23845(.A(pi1146), .B(pi0299), .C(pi0211), .Y(new_n26282_));
  AOI21X1  g23846(.A0(new_n26282_), .A1(new_n25868_), .B0(new_n26281_), .Y(new_n26283_));
  NAND2X1  g23847(.A(new_n26101_), .B(pi0212), .Y(new_n26284_));
  AOI21X1  g23848(.A0(new_n26219_), .A1(new_n25868_), .B0(new_n26284_), .Y(new_n26285_));
  NOR3X1   g23849(.A(new_n26285_), .B(new_n26283_), .C(pi0219), .Y(new_n26286_));
  OAI21X1  g23850(.A0(new_n26286_), .A1(new_n26280_), .B0(new_n26243_), .Y(new_n26287_));
  INVX1    g23851(.A(new_n26115_), .Y(new_n26288_));
  AOI21X1  g23852(.A0(new_n26288_), .A1(pi0219), .B0(po1038), .Y(new_n26289_));
  INVX1    g23853(.A(new_n26289_), .Y(new_n26290_));
  NOR2X1   g23854(.A(new_n26115_), .B(new_n8548_), .Y(new_n26291_));
  INVX1    g23855(.A(new_n26291_), .Y(new_n26292_));
  AND2X1   g23856(.A(pi0299), .B(pi0214), .Y(new_n26293_));
  INVX1    g23857(.A(new_n26293_), .Y(new_n26294_));
  AOI21X1  g23858(.A0(new_n26294_), .A1(new_n26288_), .B0(pi0212), .Y(new_n26295_));
  AND2X1   g23859(.A(new_n26295_), .B(new_n26292_), .Y(new_n26296_));
  INVX1    g23860(.A(new_n26296_), .Y(new_n26297_));
  AOI21X1  g23861(.A0(new_n26288_), .A1(new_n2953_), .B0(new_n24961_), .Y(new_n26298_));
  NOR3X1   g23862(.A(new_n25182_), .B(new_n2953_), .C(new_n24961_), .Y(new_n26299_));
  INVX1    g23863(.A(new_n26299_), .Y(new_n26300_));
  AOI21X1  g23864(.A0(new_n26300_), .A1(new_n26298_), .B0(pi0219), .Y(new_n26301_));
  AOI21X1  g23865(.A0(new_n26301_), .A1(new_n26297_), .B0(new_n26290_), .Y(new_n26302_));
  INVX1    g23866(.A(new_n26302_), .Y(new_n26303_));
  NAND3X1  g23867(.A(new_n26303_), .B(new_n26245_), .C(new_n26227_), .Y(new_n26304_));
  NAND3X1  g23868(.A(new_n26304_), .B(new_n26287_), .C(pi1148), .Y(new_n26305_));
  OAI21X1  g23869(.A0(new_n26276_), .A1(new_n26272_), .B0(new_n26305_), .Y(new_n26306_));
  AOI21X1  g23870(.A0(new_n26306_), .A1(pi1149), .B0(new_n26258_), .Y(new_n26307_));
  OAI21X1  g23871(.A0(new_n26307_), .A1(pi0213), .B0(pi0209), .Y(new_n26308_));
  AOI21X1  g23872(.A0(new_n26215_), .A1(pi0213), .B0(new_n26308_), .Y(new_n26309_));
  AOI21X1  g23873(.A0(pi1146), .A1(new_n7941_), .B0(new_n8009_), .Y(new_n26310_));
  NOR3X1   g23874(.A(pi1145), .B(pi0200), .C(new_n7941_), .Y(new_n26311_));
  OR4X1    g23875(.A(new_n26311_), .B(new_n26310_), .C(pi0299), .D(pi0207), .Y(new_n26312_));
  AOI21X1  g23876(.A0(pi1145), .A1(pi0199), .B0(pi0200), .Y(new_n26313_));
  OAI21X1  g23877(.A0(new_n3165_), .A1(pi0199), .B0(new_n26313_), .Y(new_n26314_));
  OAI21X1  g23878(.A0(new_n3346_), .A1(pi0199), .B0(pi0200), .Y(new_n26315_));
  NAND3X1  g23879(.A(new_n26315_), .B(new_n26314_), .C(new_n25159_), .Y(new_n26316_));
  NAND3X1  g23880(.A(new_n26316_), .B(new_n26312_), .C(new_n26262_), .Y(new_n26317_));
  NOR3X1   g23881(.A(new_n26311_), .B(new_n26310_), .C(pi0299), .Y(new_n26318_));
  AND2X1   g23882(.A(new_n26318_), .B(new_n24980_), .Y(new_n26319_));
  AOI21X1  g23883(.A0(new_n26317_), .A1(pi0208), .B0(new_n26319_), .Y(new_n26320_));
  AOI21X1  g23884(.A0(new_n26320_), .A1(new_n2953_), .B0(new_n8548_), .Y(new_n26321_));
  INVX1    g23885(.A(new_n26313_), .Y(new_n26322_));
  OR2X1    g23886(.A(new_n26322_), .B(new_n26312_), .Y(new_n26323_));
  NAND3X1  g23887(.A(new_n26323_), .B(new_n26317_), .C(pi0208), .Y(new_n26324_));
  NOR3X1   g23888(.A(new_n26313_), .B(new_n26310_), .C(pi0299), .Y(new_n26325_));
  INVX1    g23889(.A(new_n26325_), .Y(new_n26326_));
  OAI21X1  g23890(.A0(new_n26326_), .A1(new_n26028_), .B0(new_n26324_), .Y(new_n26327_));
  NOR2X1   g23891(.A(new_n26327_), .B(pi0299), .Y(new_n26328_));
  NOR2X1   g23892(.A(new_n26328_), .B(new_n24984_), .Y(new_n26329_));
  OAI21X1  g23893(.A0(new_n26329_), .A1(new_n26321_), .B0(pi0212), .Y(new_n26330_));
  AND2X1   g23894(.A(new_n26320_), .B(new_n2953_), .Y(new_n26331_));
  OR2X1    g23895(.A(new_n26331_), .B(new_n25740_), .Y(new_n26332_));
  NAND2X1  g23896(.A(new_n26316_), .B(new_n26178_), .Y(new_n26333_));
  OAI21X1  g23897(.A0(new_n26318_), .A1(new_n7896_), .B0(new_n26333_), .Y(new_n26334_));
  AND2X1   g23898(.A(new_n26334_), .B(new_n23539_), .Y(new_n26335_));
  NAND3X1  g23899(.A(new_n26335_), .B(new_n26332_), .C(new_n26330_), .Y(new_n26336_));
  AOI22X1  g23900(.A0(new_n26326_), .A1(new_n7897_), .B0(new_n26316_), .B1(new_n26178_), .Y(new_n26337_));
  AND2X1   g23901(.A(new_n26337_), .B(new_n24955_), .Y(new_n26338_));
  INVX1    g23902(.A(new_n26334_), .Y(new_n26339_));
  AOI21X1  g23903(.A0(new_n26320_), .A1(new_n2953_), .B0(pi0211), .Y(new_n26340_));
  NOR2X1   g23904(.A(new_n26340_), .B(new_n26339_), .Y(new_n26341_));
  AOI21X1  g23905(.A0(new_n26341_), .A1(pi0214), .B0(new_n26328_), .Y(new_n26342_));
  INVX1    g23906(.A(new_n26337_), .Y(new_n26343_));
  OAI21X1  g23907(.A0(new_n26343_), .A1(pi0214), .B0(new_n24961_), .Y(new_n26344_));
  OAI22X1  g23908(.A0(new_n26344_), .A1(new_n26329_), .B0(new_n26342_), .B1(new_n24961_), .Y(new_n26345_));
  OAI21X1  g23909(.A0(new_n26337_), .A1(new_n23539_), .B0(new_n6520_), .Y(new_n26346_));
  AOI21X1  g23910(.A0(new_n26345_), .A1(new_n23539_), .B0(new_n26346_), .Y(new_n26347_));
  OAI21X1  g23911(.A0(new_n26338_), .A1(new_n26336_), .B0(new_n26347_), .Y(new_n26348_));
  NOR2X1   g23912(.A(new_n26121_), .B(pi1147), .Y(new_n26349_));
  AOI21X1  g23913(.A0(new_n26339_), .A1(new_n24994_), .B0(new_n23539_), .Y(new_n26350_));
  NAND2X1  g23914(.A(new_n26340_), .B(new_n25323_), .Y(new_n26351_));
  AOI21X1  g23915(.A0(new_n26351_), .A1(new_n26350_), .B0(po1038), .Y(new_n26352_));
  OR2X1    g23916(.A(new_n26152_), .B(new_n26091_), .Y(new_n26353_));
  AOI21X1  g23917(.A0(new_n26352_), .A1(new_n26336_), .B0(new_n26353_), .Y(new_n26354_));
  OR2X1    g23918(.A(new_n26354_), .B(pi1149), .Y(new_n26355_));
  AOI21X1  g23919(.A0(new_n26349_), .A1(new_n26348_), .B0(new_n26355_), .Y(new_n26356_));
  NOR3X1   g23920(.A(new_n26347_), .B(new_n25955_), .C(pi1147), .Y(new_n26357_));
  INVX1    g23921(.A(new_n26352_), .Y(new_n26358_));
  AOI21X1  g23922(.A0(new_n26335_), .A1(new_n26113_), .B0(new_n26358_), .Y(new_n26359_));
  OR2X1    g23923(.A(new_n26111_), .B(new_n26091_), .Y(new_n26360_));
  OAI21X1  g23924(.A0(new_n26360_), .A1(new_n26359_), .B0(pi1149), .Y(new_n26361_));
  OAI21X1  g23925(.A0(new_n26361_), .A1(new_n26357_), .B0(pi1148), .Y(new_n26362_));
  AND2X1   g23926(.A(new_n6520_), .B(new_n26091_), .Y(new_n26363_));
  AND2X1   g23927(.A(new_n26363_), .B(new_n26337_), .Y(new_n26364_));
  INVX1    g23928(.A(new_n25970_), .Y(new_n26365_));
  NOR3X1   g23929(.A(new_n26339_), .B(new_n26321_), .C(new_n24984_), .Y(new_n26366_));
  NAND2X1  g23930(.A(new_n26334_), .B(new_n24984_), .Y(new_n26367_));
  OAI21X1  g23931(.A0(new_n26367_), .A1(new_n26340_), .B0(pi0212), .Y(new_n26368_));
  NOR2X1   g23932(.A(new_n26368_), .B(new_n26366_), .Y(new_n26369_));
  AOI21X1  g23933(.A0(new_n26334_), .A1(new_n24984_), .B0(pi0212), .Y(new_n26370_));
  INVX1    g23934(.A(new_n26370_), .Y(new_n26371_));
  OAI21X1  g23935(.A0(new_n26371_), .A1(new_n26341_), .B0(new_n23539_), .Y(new_n26372_));
  NOR2X1   g23936(.A(new_n26372_), .B(new_n26369_), .Y(new_n26373_));
  INVX1    g23937(.A(new_n26373_), .Y(new_n26374_));
  NAND3X1  g23938(.A(new_n26374_), .B(new_n26352_), .C(new_n26336_), .Y(new_n26375_));
  AOI21X1  g23939(.A0(new_n26375_), .A1(new_n26365_), .B0(new_n26091_), .Y(new_n26376_));
  OAI21X1  g23940(.A0(new_n26376_), .A1(new_n26364_), .B0(new_n26147_), .Y(new_n26377_));
  AOI21X1  g23941(.A0(new_n26374_), .A1(new_n26352_), .B0(new_n26159_), .Y(new_n26378_));
  NOR4X1   g23942(.A(new_n24955_), .B(new_n8074_), .C(pi0219), .D(pi0211), .Y(new_n26379_));
  AOI22X1  g23943(.A0(new_n26363_), .A1(new_n26337_), .B0(new_n26379_), .B1(new_n26091_), .Y(new_n26380_));
  INVX1    g23944(.A(new_n26379_), .Y(new_n26381_));
  NOR3X1   g23945(.A(new_n26327_), .B(new_n26381_), .C(new_n11777_), .Y(new_n26382_));
  OAI22X1  g23946(.A0(new_n26382_), .A1(new_n26380_), .B0(new_n26378_), .B1(new_n26091_), .Y(new_n26383_));
  AOI21X1  g23947(.A0(new_n26383_), .A1(pi1149), .B0(pi1148), .Y(new_n26384_));
  AOI21X1  g23948(.A0(new_n26384_), .A1(new_n26377_), .B0(new_n25003_), .Y(new_n26385_));
  OAI21X1  g23949(.A0(new_n26362_), .A1(new_n26356_), .B0(new_n26385_), .Y(new_n26386_));
  OR2X1    g23950(.A(new_n26338_), .B(new_n23539_), .Y(new_n26387_));
  AOI21X1  g23951(.A0(new_n26337_), .A1(new_n25323_), .B0(new_n24956_), .Y(new_n26388_));
  AND2X1   g23952(.A(new_n26327_), .B(new_n2953_), .Y(new_n26389_));
  NOR3X1   g23953(.A(new_n26389_), .B(new_n25751_), .C(pi0211), .Y(new_n26390_));
  NOR2X1   g23954(.A(new_n26390_), .B(new_n26388_), .Y(new_n26391_));
  AOI21X1  g23955(.A0(new_n26261_), .A1(pi0211), .B0(new_n26337_), .Y(new_n26392_));
  INVX1    g23956(.A(new_n26392_), .Y(new_n26393_));
  AOI21X1  g23957(.A0(new_n26343_), .A1(new_n24984_), .B0(pi0212), .Y(new_n26394_));
  AOI21X1  g23958(.A0(new_n26394_), .A1(new_n26393_), .B0(pi0219), .Y(new_n26395_));
  INVX1    g23959(.A(new_n26267_), .Y(new_n26396_));
  AOI21X1  g23960(.A0(new_n26392_), .A1(new_n24984_), .B0(new_n24961_), .Y(new_n26397_));
  OAI21X1  g23961(.A0(new_n26389_), .A1(new_n26396_), .B0(new_n26397_), .Y(new_n26398_));
  AOI21X1  g23962(.A0(new_n26398_), .A1(new_n26395_), .B0(po1038), .Y(new_n26399_));
  OAI21X1  g23963(.A0(new_n26391_), .A1(new_n26387_), .B0(new_n26399_), .Y(new_n26400_));
  INVX1    g23964(.A(new_n25749_), .Y(new_n26401_));
  NAND2X1  g23965(.A(new_n26321_), .B(new_n26401_), .Y(new_n26402_));
  NAND2X1  g23966(.A(new_n26320_), .B(new_n26267_), .Y(new_n26403_));
  OAI21X1  g23967(.A0(new_n26331_), .A1(new_n25740_), .B0(new_n26403_), .Y(new_n26404_));
  NAND3X1  g23968(.A(new_n26320_), .B(new_n26236_), .C(new_n24984_), .Y(new_n26405_));
  NAND2X1  g23969(.A(new_n26405_), .B(pi0212), .Y(new_n26406_));
  AOI21X1  g23970(.A0(new_n26404_), .A1(new_n26402_), .B0(new_n26406_), .Y(new_n26407_));
  OAI21X1  g23971(.A0(new_n26371_), .A1(new_n26341_), .B0(new_n26395_), .Y(new_n26408_));
  NAND3X1  g23972(.A(new_n26340_), .B(new_n26401_), .C(new_n25323_), .Y(new_n26409_));
  AOI21X1  g23973(.A0(new_n26409_), .A1(new_n26350_), .B0(po1038), .Y(new_n26410_));
  OAI21X1  g23974(.A0(new_n26408_), .A1(new_n26407_), .B0(new_n26410_), .Y(new_n26411_));
  AOI22X1  g23975(.A0(new_n26411_), .A1(new_n26227_), .B0(new_n26400_), .B1(new_n26243_), .Y(new_n26412_));
  AOI21X1  g23976(.A0(new_n26412_), .A1(new_n25003_), .B0(pi0209), .Y(new_n26413_));
  AOI21X1  g23977(.A0(new_n26413_), .A1(new_n26386_), .B0(new_n26309_), .Y(new_n26414_));
  MX2X1    g23978(.A(new_n26414_), .B(pi0240), .S0(new_n24954_), .Y(po0397));
  OR2X1    g23979(.A(new_n26379_), .B(new_n6520_), .Y(new_n26416_));
  AND2X1   g23980(.A(new_n26416_), .B(pi1151), .Y(new_n26417_));
  OAI21X1  g23981(.A0(new_n26381_), .A1(new_n25877_), .B0(new_n26000_), .Y(new_n26418_));
  AND2X1   g23982(.A(new_n26418_), .B(pi1152), .Y(new_n26419_));
  OAI21X1  g23983(.A0(new_n26419_), .A1(po1038), .B0(new_n26417_), .Y(new_n26420_));
  AND2X1   g23984(.A(new_n26157_), .B(new_n25021_), .Y(new_n26421_));
  OAI21X1  g23985(.A0(new_n26421_), .A1(new_n25817_), .B0(new_n26417_), .Y(new_n26422_));
  OAI21X1  g23986(.A0(new_n25838_), .A1(new_n25887_), .B0(new_n26422_), .Y(new_n26423_));
  NOR2X1   g23987(.A(new_n25838_), .B(new_n25289_), .Y(new_n26424_));
  AOI22X1  g23988(.A0(new_n26424_), .A1(new_n25869_), .B0(new_n26423_), .B1(new_n25289_), .Y(new_n26425_));
  AOI21X1  g23989(.A0(new_n26425_), .A1(new_n26420_), .B0(pi1150), .Y(new_n26426_));
  NOR2X1   g23990(.A(new_n25955_), .B(new_n25837_), .Y(new_n26427_));
  AOI21X1  g23991(.A0(new_n25887_), .A1(pi0219), .B0(po1038), .Y(new_n26428_));
  OAI21X1  g23992(.A0(new_n26013_), .A1(new_n26008_), .B0(new_n23539_), .Y(new_n26429_));
  INVX1    g23993(.A(new_n26429_), .Y(new_n26430_));
  AOI21X1  g23994(.A0(new_n25877_), .A1(new_n24984_), .B0(new_n24961_), .Y(new_n26431_));
  OAI21X1  g23995(.A0(new_n26001_), .A1(new_n24984_), .B0(new_n26431_), .Y(new_n26432_));
  AOI21X1  g23996(.A0(new_n26432_), .A1(new_n26430_), .B0(new_n25289_), .Y(new_n26433_));
  NOR2X1   g23997(.A(new_n25815_), .B(new_n25376_), .Y(new_n26434_));
  NAND2X1  g23998(.A(new_n25823_), .B(pi0214), .Y(new_n26435_));
  AOI21X1  g23999(.A0(new_n25815_), .A1(new_n24984_), .B0(new_n24961_), .Y(new_n26436_));
  AND2X1   g24000(.A(new_n26436_), .B(new_n26435_), .Y(new_n26437_));
  OAI22X1  g24001(.A0(new_n26437_), .A1(new_n25802_), .B0(new_n26434_), .B1(pi0299), .Y(new_n26438_));
  INVX1    g24002(.A(new_n25800_), .Y(new_n26439_));
  OAI21X1  g24003(.A0(new_n26439_), .A1(new_n23539_), .B0(new_n25289_), .Y(new_n26440_));
  AOI21X1  g24004(.A0(new_n26438_), .A1(new_n23539_), .B0(new_n26440_), .Y(new_n26441_));
  OAI22X1  g24005(.A0(new_n26441_), .A1(new_n26433_), .B0(new_n26428_), .B1(new_n26151_), .Y(new_n26442_));
  NOR2X1   g24006(.A(new_n26121_), .B(pi1151), .Y(new_n26443_));
  INVX1    g24007(.A(new_n26443_), .Y(new_n26444_));
  NOR3X1   g24008(.A(new_n25840_), .B(new_n25831_), .C(pi0212), .Y(new_n26445_));
  AOI21X1  g24009(.A0(new_n26445_), .A1(new_n26186_), .B0(pi0219), .Y(new_n26446_));
  NOR2X1   g24010(.A(new_n25839_), .B(new_n24984_), .Y(new_n26447_));
  AND2X1   g24011(.A(new_n25840_), .B(new_n8548_), .Y(new_n26448_));
  NOR3X1   g24012(.A(new_n26448_), .B(new_n25831_), .C(new_n24961_), .Y(new_n26449_));
  INVX1    g24013(.A(new_n26449_), .Y(new_n26450_));
  OAI21X1  g24014(.A0(new_n26450_), .A1(new_n26447_), .B0(new_n26446_), .Y(new_n26451_));
  OR4X1    g24015(.A(new_n25991_), .B(new_n25828_), .C(pi0299), .D(pi0219), .Y(new_n26452_));
  NAND3X1  g24016(.A(new_n26452_), .B(new_n26451_), .C(new_n26428_), .Y(new_n26453_));
  AND2X1   g24017(.A(new_n26453_), .B(new_n25289_), .Y(new_n26454_));
  AND2X1   g24018(.A(new_n26452_), .B(new_n26451_), .Y(new_n26455_));
  OAI21X1  g24019(.A0(new_n26455_), .A1(new_n25869_), .B0(new_n26017_), .Y(new_n26456_));
  AOI21X1  g24020(.A0(new_n26456_), .A1(pi1152), .B0(new_n26454_), .Y(new_n26457_));
  OAI21X1  g24021(.A0(new_n26457_), .A1(new_n26444_), .B0(pi1150), .Y(new_n26458_));
  AOI21X1  g24022(.A0(new_n26442_), .A1(new_n26427_), .B0(new_n26458_), .Y(new_n26459_));
  OAI21X1  g24023(.A0(new_n26459_), .A1(new_n26426_), .B0(new_n26147_), .Y(new_n26460_));
  NOR3X1   g24024(.A(new_n25884_), .B(new_n25828_), .C(new_n24961_), .Y(new_n26461_));
  OAI21X1  g24025(.A0(new_n25877_), .A1(new_n25180_), .B0(new_n26461_), .Y(new_n26462_));
  AOI21X1  g24026(.A0(new_n26462_), .A1(new_n26004_), .B0(pi0219), .Y(new_n26463_));
  OR4X1    g24027(.A(new_n26463_), .B(new_n26005_), .C(po1038), .D(new_n25289_), .Y(new_n26464_));
  OR2X1    g24028(.A(new_n26159_), .B(new_n25837_), .Y(new_n26465_));
  NOR2X1   g24029(.A(new_n25985_), .B(pi0214), .Y(new_n26466_));
  OAI22X1  g24030(.A0(new_n26466_), .A1(new_n25982_), .B0(new_n25986_), .B1(pi0212), .Y(new_n26467_));
  NAND2X1  g24031(.A(new_n26467_), .B(new_n23539_), .Y(new_n26468_));
  NOR2X1   g24032(.A(new_n25987_), .B(pi1152), .Y(new_n26469_));
  AOI21X1  g24033(.A0(new_n26469_), .A1(new_n26468_), .B0(new_n26465_), .Y(new_n26470_));
  INVX1    g24034(.A(pi1150), .Y(new_n26471_));
  NOR2X1   g24035(.A(new_n26428_), .B(new_n26209_), .Y(new_n26472_));
  AOI21X1  g24036(.A0(new_n25992_), .A1(new_n25887_), .B0(new_n26472_), .Y(new_n26473_));
  AND2X1   g24037(.A(new_n26473_), .B(new_n25289_), .Y(new_n26474_));
  NOR3X1   g24038(.A(new_n26428_), .B(new_n26209_), .C(new_n26017_), .Y(new_n26475_));
  NOR3X1   g24039(.A(new_n25991_), .B(new_n25869_), .C(pi0219), .Y(new_n26476_));
  OR2X1    g24040(.A(new_n26476_), .B(new_n25289_), .Y(new_n26477_));
  NOR2X1   g24041(.A(new_n25970_), .B(pi1151), .Y(new_n26478_));
  OAI21X1  g24042(.A0(new_n26477_), .A1(new_n26475_), .B0(new_n26478_), .Y(new_n26479_));
  OAI21X1  g24043(.A0(new_n26479_), .A1(new_n26474_), .B0(new_n26471_), .Y(new_n26480_));
  AOI21X1  g24044(.A0(new_n26470_), .A1(new_n26464_), .B0(new_n26480_), .Y(new_n26481_));
  NOR2X1   g24045(.A(new_n25877_), .B(new_n24961_), .Y(new_n26482_));
  OAI21X1  g24046(.A0(new_n26482_), .A1(new_n26429_), .B0(pi1152), .Y(new_n26483_));
  AOI21X1  g24047(.A0(new_n26110_), .A1(new_n25323_), .B0(new_n25837_), .Y(new_n26484_));
  INVX1    g24048(.A(new_n26484_), .Y(new_n26485_));
  OAI22X1  g24049(.A0(new_n26434_), .A1(pi0299), .B0(new_n25817_), .B1(new_n25323_), .Y(new_n26486_));
  NAND2X1  g24050(.A(new_n26486_), .B(new_n23539_), .Y(new_n26487_));
  AOI21X1  g24051(.A0(new_n26487_), .A1(new_n26469_), .B0(new_n26485_), .Y(new_n26488_));
  OAI21X1  g24052(.A0(new_n26483_), .A1(new_n26007_), .B0(new_n26488_), .Y(new_n26489_));
  NOR2X1   g24053(.A(new_n26152_), .B(pi1151), .Y(new_n26490_));
  INVX1    g24054(.A(new_n26454_), .Y(new_n26491_));
  AOI21X1  g24055(.A0(new_n25840_), .A1(new_n24961_), .B0(new_n25979_), .Y(new_n26492_));
  OR2X1    g24056(.A(new_n25869_), .B(new_n8074_), .Y(new_n26493_));
  OAI22X1  g24057(.A0(new_n26493_), .A1(new_n26492_), .B0(new_n25859_), .B1(new_n25014_), .Y(new_n26494_));
  AOI21X1  g24058(.A0(new_n26494_), .A1(new_n23539_), .B0(new_n26475_), .Y(new_n26495_));
  OAI22X1  g24059(.A0(new_n26495_), .A1(new_n25289_), .B0(new_n26473_), .B1(new_n26491_), .Y(new_n26496_));
  AOI21X1  g24060(.A0(new_n26496_), .A1(new_n26490_), .B0(new_n26471_), .Y(new_n26497_));
  AOI21X1  g24061(.A0(new_n26497_), .A1(new_n26489_), .B0(new_n26481_), .Y(new_n26498_));
  OAI21X1  g24062(.A0(new_n26498_), .A1(new_n26147_), .B0(new_n26460_), .Y(new_n26499_));
  OAI21X1  g24063(.A0(new_n26023_), .A1(new_n25003_), .B0(pi0209), .Y(new_n26500_));
  AOI21X1  g24064(.A0(new_n26499_), .A1(new_n25003_), .B0(new_n26500_), .Y(new_n26501_));
  OAI21X1  g24065(.A0(new_n26144_), .A1(new_n26141_), .B0(new_n26443_), .Y(new_n26502_));
  INVX1    g24066(.A(new_n26427_), .Y(new_n26503_));
  NOR2X1   g24067(.A(new_n26503_), .B(new_n26107_), .Y(new_n26504_));
  NOR2X1   g24068(.A(new_n26504_), .B(new_n26471_), .Y(new_n26505_));
  NAND2X1  g24069(.A(new_n26505_), .B(new_n26502_), .Y(new_n26506_));
  AND2X1   g24070(.A(pi1151), .B(new_n26471_), .Y(new_n26507_));
  AOI21X1  g24071(.A0(new_n26507_), .A1(new_n26183_), .B0(pi1149), .Y(new_n26508_));
  INVX1    g24072(.A(new_n26478_), .Y(new_n26509_));
  AOI21X1  g24073(.A0(new_n26211_), .A1(new_n26198_), .B0(new_n26509_), .Y(new_n26510_));
  NOR2X1   g24074(.A(new_n26510_), .B(pi1150), .Y(new_n26511_));
  OAI21X1  g24075(.A0(new_n26465_), .A1(new_n26176_), .B0(new_n26511_), .Y(new_n26512_));
  NOR3X1   g24076(.A(new_n26485_), .B(new_n26116_), .C(new_n26114_), .Y(new_n26513_));
  INVX1    g24077(.A(new_n26513_), .Y(new_n26514_));
  AOI21X1  g24078(.A0(new_n26153_), .A1(new_n25837_), .B0(new_n26471_), .Y(new_n26515_));
  AOI21X1  g24079(.A0(new_n26515_), .A1(new_n26514_), .B0(new_n26147_), .Y(new_n26516_));
  AOI22X1  g24080(.A0(new_n26516_), .A1(new_n26512_), .B0(new_n26508_), .B1(new_n26506_), .Y(new_n26517_));
  INVX1    g24081(.A(new_n26163_), .Y(new_n26518_));
  INVX1    g24082(.A(new_n25139_), .Y(new_n26519_));
  NOR2X1   g24083(.A(new_n25815_), .B(pi0211), .Y(new_n26520_));
  AOI22X1  g24084(.A0(new_n26520_), .A1(new_n26519_), .B0(new_n26439_), .B1(pi0211), .Y(new_n26521_));
  AOI22X1  g24085(.A0(new_n26521_), .A1(new_n26518_), .B0(new_n26168_), .B1(new_n26165_), .Y(new_n26522_));
  OAI21X1  g24086(.A0(new_n26522_), .A1(pi0219), .B0(new_n26174_), .Y(new_n26523_));
  AND2X1   g24087(.A(new_n25796_), .B(pi0299), .Y(new_n26524_));
  OAI21X1  g24088(.A0(new_n26421_), .A1(new_n26194_), .B0(new_n6520_), .Y(new_n26525_));
  OAI21X1  g24089(.A0(new_n26525_), .A1(new_n26524_), .B0(new_n25948_), .Y(new_n26526_));
  NAND2X1  g24090(.A(new_n26526_), .B(new_n25289_), .Y(new_n26527_));
  AOI21X1  g24091(.A0(new_n26523_), .A1(new_n25934_), .B0(new_n26527_), .Y(new_n26528_));
  OAI21X1  g24092(.A0(new_n26439_), .A1(pi0214), .B0(new_n26162_), .Y(new_n26529_));
  NOR3X1   g24093(.A(new_n26299_), .B(new_n25825_), .C(pi0219), .Y(new_n26530_));
  NAND2X1  g24094(.A(new_n26530_), .B(new_n26529_), .Y(new_n26531_));
  AOI21X1  g24095(.A0(new_n26531_), .A1(new_n26174_), .B0(new_n25972_), .Y(new_n26532_));
  OAI22X1  g24096(.A0(new_n26194_), .A1(new_n26112_), .B0(new_n25957_), .B1(new_n25040_), .Y(new_n26533_));
  NOR2X1   g24097(.A(new_n26194_), .B(new_n23539_), .Y(new_n26534_));
  NOR2X1   g24098(.A(new_n26534_), .B(po1038), .Y(new_n26535_));
  INVX1    g24099(.A(new_n26535_), .Y(new_n26536_));
  AOI21X1  g24100(.A0(new_n26533_), .A1(new_n23539_), .B0(new_n26536_), .Y(new_n26537_));
  OAI21X1  g24101(.A0(new_n26537_), .A1(new_n25959_), .B0(pi1152), .Y(new_n26538_));
  OAI21X1  g24102(.A0(new_n26538_), .A1(new_n26532_), .B0(new_n26471_), .Y(new_n26539_));
  OR2X1    g24103(.A(new_n26539_), .B(new_n26528_), .Y(new_n26540_));
  NOR4X1   g24104(.A(new_n26299_), .B(new_n26115_), .C(pi1153), .D(pi0219), .Y(new_n26541_));
  NOR4X1   g24105(.A(new_n2953_), .B(new_n24984_), .C(new_n24961_), .D(new_n8548_), .Y(new_n26542_));
  NOR2X1   g24106(.A(new_n26542_), .B(pi0219), .Y(new_n26543_));
  INVX1    g24107(.A(new_n26543_), .Y(new_n26544_));
  AND2X1   g24108(.A(new_n26544_), .B(new_n26209_), .Y(new_n26545_));
  NOR2X1   g24109(.A(new_n26545_), .B(new_n26302_), .Y(new_n26546_));
  OAI21X1  g24110(.A0(new_n26546_), .A1(new_n26541_), .B0(new_n25934_), .Y(new_n26547_));
  NAND3X1  g24111(.A(new_n26157_), .B(new_n25021_), .C(pi1153), .Y(new_n26548_));
  AOI21X1  g24112(.A0(new_n26548_), .A1(new_n25948_), .B0(pi1152), .Y(new_n26549_));
  OAI21X1  g24113(.A0(new_n25883_), .A1(po1038), .B0(new_n25837_), .Y(new_n26550_));
  AND2X1   g24114(.A(new_n26550_), .B(new_n25289_), .Y(new_n26551_));
  OAI21X1  g24115(.A0(new_n26551_), .A1(new_n26549_), .B0(new_n26547_), .Y(new_n26552_));
  NOR2X1   g24116(.A(new_n26116_), .B(new_n26114_), .Y(new_n26553_));
  NOR4X1   g24117(.A(new_n26299_), .B(new_n26115_), .C(pi0219), .D(pi0211), .Y(new_n26554_));
  NOR2X1   g24118(.A(new_n26554_), .B(new_n26553_), .Y(new_n26555_));
  NOR2X1   g24119(.A(new_n26555_), .B(new_n25972_), .Y(new_n26556_));
  OAI21X1  g24120(.A0(new_n26546_), .A1(new_n26541_), .B0(new_n26556_), .Y(new_n26557_));
  AOI21X1  g24121(.A0(new_n25883_), .A1(pi0219), .B0(po1038), .Y(new_n26558_));
  AOI21X1  g24122(.A0(new_n26186_), .A1(new_n25883_), .B0(new_n25014_), .Y(new_n26559_));
  OR2X1    g24123(.A(new_n26524_), .B(new_n24962_), .Y(new_n26560_));
  AOI21X1  g24124(.A0(new_n25883_), .A1(new_n2953_), .B0(new_n26560_), .Y(new_n26561_));
  OR4X1    g24125(.A(new_n26561_), .B(new_n26559_), .C(new_n26238_), .D(pi0219), .Y(new_n26562_));
  AOI21X1  g24126(.A0(new_n26562_), .A1(new_n26558_), .B0(new_n25959_), .Y(new_n26563_));
  NOR2X1   g24127(.A(new_n26563_), .B(new_n25289_), .Y(new_n26564_));
  AOI21X1  g24128(.A0(new_n26564_), .A1(new_n26557_), .B0(new_n26471_), .Y(new_n26565_));
  AOI21X1  g24129(.A0(new_n26565_), .A1(new_n26552_), .B0(new_n26147_), .Y(new_n26566_));
  INVX1    g24130(.A(new_n26135_), .Y(new_n26567_));
  NOR3X1   g24131(.A(new_n26524_), .B(new_n26131_), .C(new_n24984_), .Y(new_n26568_));
  NOR3X1   g24132(.A(new_n26524_), .B(new_n26131_), .C(pi0214), .Y(new_n26569_));
  OAI22X1  g24133(.A0(new_n26569_), .A1(new_n26567_), .B0(new_n26568_), .B1(new_n26130_), .Y(new_n26570_));
  AOI21X1  g24134(.A0(new_n26570_), .A1(new_n23539_), .B0(new_n26144_), .Y(new_n26571_));
  INVX1    g24135(.A(new_n26279_), .Y(new_n26572_));
  OAI21X1  g24136(.A0(new_n25122_), .A1(new_n25086_), .B0(new_n25852_), .Y(new_n26573_));
  AOI21X1  g24137(.A0(new_n12494_), .A1(pi0299), .B0(pi0211), .Y(new_n26574_));
  AOI22X1  g24138(.A0(new_n26574_), .A1(new_n26573_), .B0(new_n26101_), .B1(pi0211), .Y(new_n26575_));
  AOI21X1  g24139(.A0(new_n26575_), .A1(pi0214), .B0(new_n26281_), .Y(new_n26576_));
  AOI21X1  g24140(.A0(new_n26575_), .A1(new_n24984_), .B0(new_n26284_), .Y(new_n26577_));
  NOR3X1   g24141(.A(new_n26577_), .B(new_n26576_), .C(pi0219), .Y(new_n26578_));
  OAI21X1  g24142(.A0(new_n26578_), .A1(new_n26572_), .B0(new_n25999_), .Y(new_n26579_));
  AND2X1   g24143(.A(new_n26579_), .B(pi1152), .Y(new_n26580_));
  OAI21X1  g24144(.A0(new_n26571_), .A1(new_n25959_), .B0(new_n26580_), .Y(new_n26581_));
  INVX1    g24145(.A(new_n25950_), .Y(new_n26582_));
  OAI21X1  g24146(.A0(new_n26131_), .A1(new_n25139_), .B0(new_n8548_), .Y(new_n26583_));
  NOR2X1   g24147(.A(new_n26133_), .B(new_n26582_), .Y(new_n26584_));
  AOI22X1  g24148(.A0(new_n26584_), .A1(new_n26583_), .B0(new_n26124_), .B1(new_n26582_), .Y(new_n26585_));
  OAI21X1  g24149(.A0(new_n26585_), .A1(po1038), .B0(new_n25948_), .Y(new_n26586_));
  INVX1    g24150(.A(new_n26575_), .Y(new_n26587_));
  AOI21X1  g24151(.A0(new_n26101_), .A1(pi0211), .B0(new_n25867_), .Y(new_n26588_));
  INVX1    g24152(.A(new_n26095_), .Y(new_n26589_));
  OAI21X1  g24153(.A0(new_n26102_), .A1(new_n26589_), .B0(pi0212), .Y(new_n26590_));
  AOI21X1  g24154(.A0(new_n26588_), .A1(pi0214), .B0(new_n26590_), .Y(new_n26591_));
  AOI21X1  g24155(.A0(new_n26574_), .A1(new_n26573_), .B0(new_n26103_), .Y(new_n26592_));
  OAI21X1  g24156(.A0(new_n26592_), .A1(new_n26281_), .B0(new_n23539_), .Y(new_n26593_));
  AOI21X1  g24157(.A0(new_n26591_), .A1(new_n26587_), .B0(new_n26593_), .Y(new_n26594_));
  OAI21X1  g24158(.A0(new_n26594_), .A1(new_n26572_), .B0(new_n25934_), .Y(new_n26595_));
  NAND3X1  g24159(.A(new_n26595_), .B(new_n26586_), .C(new_n25289_), .Y(new_n26596_));
  NAND3X1  g24160(.A(new_n26596_), .B(new_n26581_), .C(pi1150), .Y(new_n26597_));
  AOI21X1  g24161(.A0(new_n25842_), .A1(pi0219), .B0(po1038), .Y(new_n26598_));
  AND2X1   g24162(.A(new_n26598_), .B(new_n25994_), .Y(new_n26599_));
  INVX1    g24163(.A(new_n26598_), .Y(new_n26600_));
  AOI21X1  g24164(.A0(new_n26450_), .A1(new_n26446_), .B0(new_n26600_), .Y(new_n26601_));
  OR2X1    g24165(.A(new_n26601_), .B(new_n25972_), .Y(new_n26602_));
  NOR3X1   g24166(.A(new_n24955_), .B(new_n25930_), .C(pi0219), .Y(new_n26603_));
  NAND3X1  g24167(.A(new_n25957_), .B(new_n26603_), .C(pi0299), .Y(new_n26604_));
  AOI21X1  g24168(.A0(new_n26604_), .A1(new_n25958_), .B0(new_n25289_), .Y(new_n26605_));
  OAI21X1  g24169(.A0(new_n26602_), .A1(new_n26599_), .B0(new_n26605_), .Y(new_n26606_));
  OAI21X1  g24170(.A0(new_n26599_), .A1(new_n25933_), .B0(new_n26549_), .Y(new_n26607_));
  AND2X1   g24171(.A(new_n26607_), .B(new_n26471_), .Y(new_n26608_));
  AOI21X1  g24172(.A0(new_n26608_), .A1(new_n26606_), .B0(pi1149), .Y(new_n26609_));
  AOI22X1  g24173(.A0(new_n26609_), .A1(new_n26597_), .B0(new_n26566_), .B1(new_n26540_), .Y(new_n26610_));
  OAI21X1  g24174(.A0(new_n26610_), .A1(new_n25003_), .B0(new_n23244_), .Y(new_n26611_));
  AOI21X1  g24175(.A0(new_n26517_), .A1(new_n25003_), .B0(new_n26611_), .Y(new_n26612_));
  NOR2X1   g24176(.A(new_n26612_), .B(new_n26501_), .Y(new_n26613_));
  MX2X1    g24177(.A(new_n26613_), .B(pi0241), .S0(new_n24954_), .Y(po0398));
  NOR2X1   g24178(.A(pi0242), .B(pi0230), .Y(new_n26615_));
  MX2X1    g24179(.A(new_n26217_), .B(new_n25648_), .S0(pi0214), .Y(new_n26616_));
  NOR3X1   g24180(.A(new_n26217_), .B(new_n24984_), .C(pi0212), .Y(new_n26617_));
  NOR2X1   g24181(.A(new_n26617_), .B(pi0219), .Y(new_n26618_));
  OAI21X1  g24182(.A0(new_n26616_), .A1(new_n24961_), .B0(new_n26618_), .Y(new_n26619_));
  INVX1    g24183(.A(new_n26619_), .Y(new_n26620_));
  AOI21X1  g24184(.A0(pi1144), .A1(new_n8548_), .B0(new_n23539_), .Y(new_n26621_));
  NOR3X1   g24185(.A(new_n26621_), .B(new_n26620_), .C(new_n25929_), .Y(new_n26622_));
  INVX1    g24186(.A(new_n26622_), .Y(new_n26623_));
  AOI21X1  g24187(.A0(pi1144), .A1(pi0199), .B0(pi0200), .Y(new_n26624_));
  OAI21X1  g24188(.A0(new_n3165_), .A1(pi0199), .B0(new_n26624_), .Y(new_n26625_));
  NAND3X1  g24189(.A(new_n26625_), .B(new_n26315_), .C(new_n2953_), .Y(new_n26626_));
  NAND2X1  g24190(.A(new_n26626_), .B(new_n22803_), .Y(new_n26627_));
  OAI21X1  g24191(.A0(new_n3346_), .A1(pi0199), .B0(new_n26624_), .Y(new_n26628_));
  NAND3X1  g24192(.A(new_n26628_), .B(new_n25638_), .C(new_n2953_), .Y(new_n26629_));
  AOI21X1  g24193(.A0(new_n26629_), .A1(pi0207), .B0(new_n23109_), .Y(new_n26630_));
  AND2X1   g24194(.A(new_n26630_), .B(new_n26627_), .Y(new_n26631_));
  NOR2X1   g24195(.A(new_n26626_), .B(new_n26028_), .Y(new_n26632_));
  NOR3X1   g24196(.A(new_n26632_), .B(new_n26631_), .C(new_n25751_), .Y(new_n26633_));
  NOR2X1   g24197(.A(new_n26633_), .B(pi0211), .Y(new_n26634_));
  NOR3X1   g24198(.A(new_n26632_), .B(new_n26631_), .C(new_n25215_), .Y(new_n26635_));
  OAI21X1  g24199(.A0(new_n26635_), .A1(new_n8548_), .B0(pi0214), .Y(new_n26636_));
  NOR2X1   g24200(.A(new_n26636_), .B(new_n26634_), .Y(new_n26637_));
  OAI21X1  g24201(.A0(new_n26626_), .A1(new_n26028_), .B0(new_n26262_), .Y(new_n26638_));
  AOI21X1  g24202(.A0(new_n26630_), .A1(new_n26627_), .B0(new_n26638_), .Y(new_n26639_));
  MX2X1    g24203(.A(new_n26639_), .B(new_n26633_), .S0(pi0211), .Y(new_n26640_));
  AND2X1   g24204(.A(new_n26640_), .B(new_n24984_), .Y(new_n26641_));
  NOR3X1   g24205(.A(new_n26641_), .B(new_n26637_), .C(new_n24961_), .Y(new_n26642_));
  NOR2X1   g24206(.A(new_n26626_), .B(new_n26178_), .Y(new_n26643_));
  AOI21X1  g24207(.A0(new_n26630_), .A1(new_n26627_), .B0(new_n26643_), .Y(new_n26644_));
  AOI21X1  g24208(.A0(new_n26644_), .A1(new_n24984_), .B0(pi0212), .Y(new_n26645_));
  INVX1    g24209(.A(new_n26645_), .Y(new_n26646_));
  AOI21X1  g24210(.A0(new_n26640_), .A1(pi0214), .B0(new_n26646_), .Y(new_n26647_));
  OR2X1    g24211(.A(new_n26647_), .B(pi0219), .Y(new_n26648_));
  INVX1    g24212(.A(new_n26644_), .Y(new_n26649_));
  AOI21X1  g24213(.A0(new_n26649_), .A1(new_n24994_), .B0(new_n23539_), .Y(new_n26650_));
  OR2X1    g24214(.A(new_n26635_), .B(new_n24994_), .Y(new_n26651_));
  AOI21X1  g24215(.A0(new_n26651_), .A1(new_n26650_), .B0(po1038), .Y(new_n26652_));
  OAI21X1  g24216(.A0(new_n26648_), .A1(new_n26642_), .B0(new_n26652_), .Y(new_n26653_));
  AND2X1   g24217(.A(new_n26653_), .B(new_n26623_), .Y(new_n26654_));
  OAI21X1  g24218(.A0(new_n3706_), .A1(new_n2953_), .B0(new_n24956_), .Y(new_n26655_));
  OAI22X1  g24219(.A0(new_n26655_), .A1(new_n26632_), .B0(new_n26643_), .B1(new_n8548_), .Y(new_n26656_));
  OAI22X1  g24220(.A0(new_n25516_), .A1(new_n24968_), .B0(new_n24986_), .B1(new_n25014_), .Y(new_n26657_));
  NOR2X1   g24221(.A(new_n26632_), .B(pi0219), .Y(new_n26658_));
  NAND2X1  g24222(.A(new_n26658_), .B(new_n26657_), .Y(new_n26659_));
  OAI21X1  g24223(.A0(new_n26643_), .A1(new_n25323_), .B0(new_n26659_), .Y(new_n26660_));
  AOI21X1  g24224(.A0(new_n26656_), .A1(pi0219), .B0(new_n26660_), .Y(new_n26661_));
  OAI21X1  g24225(.A0(new_n26661_), .A1(new_n26631_), .B0(new_n6520_), .Y(new_n26662_));
  AOI21X1  g24226(.A0(new_n24966_), .A1(new_n24958_), .B0(pi0213), .Y(new_n26663_));
  AOI22X1  g24227(.A0(new_n26663_), .A1(new_n26662_), .B0(new_n26654_), .B1(pi0213), .Y(new_n26664_));
  AND2X1   g24228(.A(new_n24955_), .B(pi0219), .Y(new_n26665_));
  NOR3X1   g24229(.A(new_n26665_), .B(new_n26621_), .C(new_n26620_), .Y(new_n26666_));
  OAI21X1  g24230(.A0(new_n26666_), .A1(new_n2953_), .B0(new_n6520_), .Y(new_n26667_));
  OAI21X1  g24231(.A0(new_n26667_), .A1(new_n24996_), .B0(new_n26623_), .Y(new_n26668_));
  AOI21X1  g24232(.A0(new_n26668_), .A1(pi0213), .B0(pi0209), .Y(new_n26669_));
  OAI21X1  g24233(.A0(new_n25001_), .A1(pi0213), .B0(new_n26669_), .Y(new_n26670_));
  OAI21X1  g24234(.A0(new_n26664_), .A1(new_n23244_), .B0(new_n26670_), .Y(new_n26671_));
  AOI21X1  g24235(.A0(new_n26671_), .A1(pi0230), .B0(new_n26615_), .Y(po0399));
  INVX1    g24236(.A(pi0243), .Y(new_n26673_));
  INVX1    g24237(.A(pi0273), .Y(new_n26674_));
  AOI21X1  g24238(.A0(new_n5145_), .A1(new_n2614_), .B0(new_n7734_), .Y(new_n26675_));
  NAND2X1  g24239(.A(new_n26675_), .B(pi0802), .Y(new_n26676_));
  NOR2X1   g24240(.A(new_n26676_), .B(new_n3175_), .Y(new_n26677_));
  AOI21X1  g24241(.A0(new_n26677_), .A1(pi0271), .B0(pi1091), .Y(new_n26678_));
  NOR2X1   g24242(.A(new_n26678_), .B(new_n26674_), .Y(new_n26679_));
  NOR2X1   g24243(.A(new_n26679_), .B(pi1091), .Y(new_n26680_));
  INVX1    g24244(.A(new_n26680_), .Y(new_n26681_));
  OAI21X1  g24245(.A0(new_n26679_), .A1(pi1091), .B0(pi0199), .Y(new_n26682_));
  INVX1    g24246(.A(pi0802), .Y(new_n26683_));
  NOR3X1   g24247(.A(pi0085), .B(pi0083), .C(pi0081), .Y(new_n26684_));
  OR4X1    g24248(.A(new_n26684_), .B(new_n26683_), .C(new_n7734_), .D(new_n3175_), .Y(new_n26685_));
  NOR2X1   g24249(.A(new_n26685_), .B(pi1091), .Y(new_n26686_));
  INVX1    g24250(.A(new_n26686_), .Y(new_n26687_));
  INVX1    g24251(.A(pi0271), .Y(new_n26688_));
  NOR4X1   g24252(.A(new_n26685_), .B(pi1091), .C(new_n26674_), .D(new_n26688_), .Y(new_n26689_));
  NOR2X1   g24253(.A(new_n26689_), .B(new_n26679_), .Y(new_n26690_));
  AOI21X1  g24254(.A0(new_n26690_), .A1(new_n2722_), .B0(pi0199), .Y(new_n26691_));
  INVX1    g24255(.A(new_n26691_), .Y(new_n26692_));
  AOI21X1  g24256(.A0(new_n26692_), .A1(new_n26682_), .B0(new_n26687_), .Y(new_n26693_));
  NOR2X1   g24257(.A(new_n26693_), .B(pi0299), .Y(new_n26694_));
  AND2X1   g24258(.A(new_n26694_), .B(new_n26682_), .Y(new_n26695_));
  INVX1    g24259(.A(new_n26695_), .Y(new_n26696_));
  AOI21X1  g24260(.A0(new_n26681_), .A1(new_n8009_), .B0(new_n26696_), .Y(new_n26697_));
  NOR2X1   g24261(.A(new_n26689_), .B(new_n2953_), .Y(new_n26698_));
  OAI22X1  g24262(.A0(new_n26698_), .A1(new_n26697_), .B0(pi1091), .B1(new_n26673_), .Y(new_n26699_));
  AOI22X1  g24263(.A0(new_n26692_), .A1(new_n26682_), .B0(new_n26687_), .B1(new_n8009_), .Y(new_n26700_));
  NOR2X1   g24264(.A(new_n26700_), .B(pi0299), .Y(new_n26701_));
  AND2X1   g24265(.A(new_n26701_), .B(new_n26682_), .Y(new_n26702_));
  NOR4X1   g24266(.A(new_n26676_), .B(pi1091), .C(new_n3175_), .D(new_n26688_), .Y(new_n26703_));
  AOI21X1  g24267(.A0(new_n26703_), .A1(pi0273), .B0(new_n2953_), .Y(new_n26704_));
  INVX1    g24268(.A(new_n26694_), .Y(new_n26705_));
  AOI21X1  g24269(.A0(new_n26681_), .A1(new_n8009_), .B0(new_n26705_), .Y(new_n26706_));
  AOI21X1  g24270(.A0(new_n26706_), .A1(new_n26692_), .B0(new_n26704_), .Y(new_n26707_));
  INVX1    g24271(.A(new_n26707_), .Y(new_n26708_));
  INVX1    g24272(.A(new_n26706_), .Y(new_n26709_));
  NOR3X1   g24273(.A(new_n26679_), .B(pi1091), .C(new_n2953_), .Y(new_n26710_));
  INVX1    g24274(.A(new_n26710_), .Y(new_n26711_));
  AOI21X1  g24275(.A0(new_n26711_), .A1(new_n26709_), .B0(new_n26673_), .Y(new_n26712_));
  OAI21X1  g24276(.A0(new_n26708_), .A1(new_n26702_), .B0(new_n26712_), .Y(new_n26713_));
  AND2X1   g24277(.A(new_n26713_), .B(pi1155), .Y(new_n26714_));
  AND2X1   g24278(.A(new_n26706_), .B(new_n26692_), .Y(new_n26715_));
  NOR4X1   g24279(.A(new_n26689_), .B(new_n26679_), .C(pi1091), .D(new_n2953_), .Y(new_n26716_));
  NOR3X1   g24280(.A(new_n26716_), .B(new_n26715_), .C(new_n12591_), .Y(new_n26717_));
  OR2X1    g24281(.A(new_n26717_), .B(new_n26714_), .Y(new_n26718_));
  OR4X1    g24282(.A(new_n26701_), .B(new_n26698_), .C(new_n26697_), .D(pi0243), .Y(new_n26719_));
  NOR3X1   g24283(.A(new_n26700_), .B(new_n26691_), .C(pi0299), .Y(new_n26720_));
  NOR3X1   g24284(.A(new_n26720_), .B(new_n26716_), .C(new_n26697_), .Y(new_n26721_));
  OR4X1    g24285(.A(new_n26715_), .B(new_n26702_), .C(new_n26698_), .D(new_n26673_), .Y(new_n26722_));
  OAI21X1  g24286(.A0(new_n26721_), .A1(pi0243), .B0(new_n26722_), .Y(new_n26723_));
  AOI22X1  g24287(.A0(new_n26723_), .A1(new_n12591_), .B0(new_n26719_), .B1(new_n26718_), .Y(new_n26724_));
  AOI21X1  g24288(.A0(new_n26724_), .A1(new_n26699_), .B0(new_n12684_), .Y(new_n26725_));
  NOR2X1   g24289(.A(new_n26720_), .B(new_n26710_), .Y(new_n26726_));
  NOR2X1   g24290(.A(new_n26726_), .B(pi0243), .Y(new_n26727_));
  MX2X1    g24291(.A(new_n26693_), .B(new_n26689_), .S0(pi0299), .Y(new_n26728_));
  INVX1    g24292(.A(new_n26728_), .Y(new_n26729_));
  AOI21X1  g24293(.A0(new_n26729_), .A1(new_n26727_), .B0(pi1155), .Y(new_n26730_));
  NOR4X1   g24294(.A(new_n26706_), .B(new_n26698_), .C(new_n26695_), .D(new_n26673_), .Y(new_n26731_));
  INVX1    g24295(.A(new_n26731_), .Y(new_n26732_));
  AOI21X1  g24296(.A0(new_n26732_), .A1(new_n26730_), .B0(pi1156), .Y(new_n26733_));
  INVX1    g24297(.A(new_n26733_), .Y(new_n26734_));
  NOR2X1   g24298(.A(new_n26706_), .B(new_n26698_), .Y(new_n26735_));
  NOR2X1   g24299(.A(new_n26716_), .B(new_n26701_), .Y(new_n26736_));
  NOR2X1   g24300(.A(new_n26736_), .B(pi0243), .Y(new_n26737_));
  NOR2X1   g24301(.A(new_n26737_), .B(new_n12591_), .Y(new_n26738_));
  INVX1    g24302(.A(new_n26738_), .Y(new_n26739_));
  AOI21X1  g24303(.A0(new_n26735_), .A1(pi0243), .B0(new_n26739_), .Y(new_n26740_));
  OAI21X1  g24304(.A0(new_n26740_), .A1(new_n26734_), .B0(pi1157), .Y(new_n26741_));
  AND2X1   g24305(.A(new_n26728_), .B(new_n12591_), .Y(new_n26742_));
  NOR2X1   g24306(.A(pi1091), .B(pi0243), .Y(new_n26743_));
  AND2X1   g24307(.A(new_n26703_), .B(pi0273), .Y(new_n26744_));
  MX2X1    g24308(.A(new_n26744_), .B(new_n26693_), .S0(new_n2953_), .Y(new_n26745_));
  INVX1    g24309(.A(new_n26745_), .Y(new_n26746_));
  AOI21X1  g24310(.A0(new_n26746_), .A1(new_n26743_), .B0(pi1155), .Y(new_n26747_));
  OAI22X1  g24311(.A0(new_n26747_), .A1(new_n26742_), .B0(new_n26729_), .B1(new_n26673_), .Y(new_n26748_));
  INVX1    g24312(.A(new_n26748_), .Y(new_n26749_));
  AND2X1   g24313(.A(new_n2722_), .B(pi0243), .Y(new_n26750_));
  NOR3X1   g24314(.A(new_n26682_), .B(new_n26750_), .C(new_n12591_), .Y(new_n26751_));
  OR4X1    g24315(.A(new_n26751_), .B(new_n26749_), .C(new_n26740_), .D(pi1156), .Y(new_n26752_));
  NOR4X1   g24316(.A(new_n26706_), .B(new_n26698_), .C(new_n26686_), .D(pi1155), .Y(new_n26753_));
  NOR3X1   g24317(.A(new_n26693_), .B(new_n26691_), .C(pi0299), .Y(new_n26754_));
  NOR2X1   g24318(.A(new_n26754_), .B(new_n26716_), .Y(new_n26755_));
  AOI21X1  g24319(.A0(new_n26694_), .A1(new_n26682_), .B0(new_n26698_), .Y(new_n26756_));
  INVX1    g24320(.A(new_n26756_), .Y(new_n26757_));
  MX2X1    g24321(.A(new_n26757_), .B(new_n26755_), .S0(pi0243), .Y(new_n26758_));
  INVX1    g24322(.A(new_n26758_), .Y(new_n26759_));
  NOR3X1   g24323(.A(new_n26759_), .B(new_n26753_), .C(new_n12684_), .Y(new_n26760_));
  NOR2X1   g24324(.A(new_n26760_), .B(pi1157), .Y(new_n26761_));
  AOI21X1  g24325(.A0(new_n26761_), .A1(new_n26752_), .B0(new_n8548_), .Y(new_n26762_));
  OAI21X1  g24326(.A0(new_n26741_), .A1(new_n26725_), .B0(new_n26762_), .Y(new_n26763_));
  MX2X1    g24327(.A(new_n26700_), .B(new_n26689_), .S0(pi0299), .Y(new_n26764_));
  NOR2X1   g24328(.A(new_n26716_), .B(new_n26706_), .Y(new_n26765_));
  INVX1    g24329(.A(new_n26765_), .Y(new_n26766_));
  MX2X1    g24330(.A(new_n26766_), .B(new_n26764_), .S0(new_n26673_), .Y(new_n26767_));
  INVX1    g24331(.A(new_n26767_), .Y(new_n26768_));
  AOI21X1  g24332(.A0(new_n26768_), .A1(new_n26733_), .B0(new_n12706_), .Y(new_n26769_));
  OAI21X1  g24333(.A0(new_n26724_), .A1(new_n12684_), .B0(new_n26769_), .Y(new_n26770_));
  NOR4X1   g24334(.A(new_n26764_), .B(new_n26716_), .C(new_n26706_), .D(pi1155), .Y(new_n26771_));
  OR4X1    g24335(.A(new_n26771_), .B(new_n26759_), .C(new_n26753_), .D(new_n12684_), .Y(new_n26772_));
  AND2X1   g24336(.A(new_n26748_), .B(new_n12684_), .Y(new_n26773_));
  OAI21X1  g24337(.A0(new_n26767_), .A1(new_n26759_), .B0(pi1155), .Y(new_n26774_));
  AOI21X1  g24338(.A0(new_n26774_), .A1(new_n26773_), .B0(pi1157), .Y(new_n26775_));
  AOI21X1  g24339(.A0(new_n26775_), .A1(new_n26772_), .B0(pi0211), .Y(new_n26776_));
  AOI21X1  g24340(.A0(new_n26776_), .A1(new_n26770_), .B0(pi0219), .Y(new_n26777_));
  INVX1    g24341(.A(pi0253), .Y(new_n26778_));
  INVX1    g24342(.A(pi0254), .Y(new_n26779_));
  INVX1    g24343(.A(pi0267), .Y(new_n26780_));
  NOR4X1   g24344(.A(new_n26780_), .B(pi0263), .C(new_n26779_), .D(new_n26778_), .Y(new_n26781_));
  MX2X1    g24345(.A(new_n26744_), .B(new_n26700_), .S0(new_n2953_), .Y(new_n26782_));
  INVX1    g24346(.A(new_n26782_), .Y(new_n26783_));
  OR4X1    g24347(.A(new_n26783_), .B(new_n26710_), .C(new_n26697_), .D(pi0243), .Y(new_n26784_));
  NAND3X1  g24348(.A(new_n26784_), .B(new_n26713_), .C(pi1155), .Y(new_n26785_));
  INVX1    g24349(.A(new_n26702_), .Y(new_n26786_));
  AND2X1   g24350(.A(new_n26707_), .B(new_n26786_), .Y(new_n26787_));
  NOR2X1   g24351(.A(new_n26710_), .B(new_n26697_), .Y(new_n26788_));
  INVX1    g24352(.A(new_n26788_), .Y(new_n26789_));
  MX2X1    g24353(.A(new_n26789_), .B(new_n26787_), .S0(pi0243), .Y(new_n26790_));
  OAI21X1  g24354(.A0(new_n26726_), .A1(pi0243), .B0(new_n26699_), .Y(new_n26791_));
  OAI21X1  g24355(.A0(new_n26791_), .A1(new_n26790_), .B0(new_n12591_), .Y(new_n26792_));
  AOI21X1  g24356(.A0(new_n26792_), .A1(new_n26785_), .B0(new_n12684_), .Y(new_n26793_));
  NOR2X1   g24357(.A(new_n26720_), .B(new_n26704_), .Y(new_n26794_));
  NOR2X1   g24358(.A(new_n26794_), .B(pi0243), .Y(new_n26795_));
  OAI21X1  g24359(.A0(new_n26695_), .A1(new_n26673_), .B0(new_n12591_), .Y(new_n26796_));
  NOR2X1   g24360(.A(new_n26796_), .B(new_n26795_), .Y(new_n26797_));
  NOR4X1   g24361(.A(new_n26704_), .B(new_n26701_), .C(new_n12591_), .D(pi0243), .Y(new_n26798_));
  NOR4X1   g24362(.A(new_n26798_), .B(new_n26797_), .C(new_n26712_), .D(pi1156), .Y(new_n26799_));
  NOR4X1   g24363(.A(new_n26799_), .B(new_n26793_), .C(new_n12706_), .D(pi0211), .Y(new_n26800_));
  INVX1    g24364(.A(new_n26790_), .Y(new_n26801_));
  AND2X1   g24365(.A(new_n26707_), .B(pi0243), .Y(new_n26802_));
  OAI22X1  g24366(.A0(new_n26802_), .A1(new_n26739_), .B0(new_n26727_), .B1(pi1155), .Y(new_n26803_));
  AOI21X1  g24367(.A0(new_n26803_), .A1(new_n26801_), .B0(new_n12684_), .Y(new_n26804_));
  NOR3X1   g24368(.A(new_n26706_), .B(new_n26704_), .C(new_n26673_), .Y(new_n26805_));
  OAI21X1  g24369(.A0(new_n26805_), .A1(new_n26737_), .B0(pi1155), .Y(new_n26806_));
  NOR2X1   g24370(.A(new_n26706_), .B(new_n26704_), .Y(new_n26807_));
  NAND2X1  g24371(.A(new_n26807_), .B(new_n26696_), .Y(new_n26808_));
  MX2X1    g24372(.A(new_n26808_), .B(new_n26726_), .S0(new_n26673_), .Y(new_n26809_));
  AOI21X1  g24373(.A0(new_n26809_), .A1(new_n26806_), .B0(pi1156), .Y(new_n26810_));
  NOR4X1   g24374(.A(new_n26810_), .B(new_n26804_), .C(new_n12706_), .D(new_n8548_), .Y(new_n26811_));
  NOR3X1   g24375(.A(new_n26754_), .B(new_n26704_), .C(new_n12591_), .Y(new_n26812_));
  NOR3X1   g24376(.A(new_n26754_), .B(new_n26704_), .C(new_n26701_), .Y(new_n26813_));
  OAI21X1  g24377(.A0(new_n26813_), .A1(new_n26812_), .B0(pi0243), .Y(new_n26814_));
  AOI21X1  g24378(.A0(new_n26694_), .A1(new_n26682_), .B0(new_n26710_), .Y(new_n26815_));
  OR2X1    g24379(.A(new_n26815_), .B(pi0243), .Y(new_n26816_));
  OAI21X1  g24380(.A0(new_n26816_), .A1(new_n26753_), .B0(new_n26814_), .Y(new_n26817_));
  AND2X1   g24381(.A(new_n26817_), .B(pi1156), .Y(new_n26818_));
  OR4X1    g24382(.A(new_n26754_), .B(new_n26706_), .C(new_n26704_), .D(new_n26673_), .Y(new_n26819_));
  AOI21X1  g24383(.A0(new_n26701_), .A1(new_n26682_), .B0(new_n26710_), .Y(new_n26820_));
  INVX1    g24384(.A(new_n26820_), .Y(new_n26821_));
  AOI21X1  g24385(.A0(new_n26821_), .A1(new_n26673_), .B0(new_n12591_), .Y(new_n26822_));
  OAI21X1  g24386(.A0(new_n26746_), .A1(new_n26673_), .B0(new_n26747_), .Y(new_n26823_));
  NAND2X1  g24387(.A(new_n26823_), .B(new_n12684_), .Y(new_n26824_));
  AOI21X1  g24388(.A0(new_n26822_), .A1(new_n26819_), .B0(new_n26824_), .Y(new_n26825_));
  NOR3X1   g24389(.A(new_n26825_), .B(new_n26818_), .C(pi1157), .Y(new_n26826_));
  NOR3X1   g24390(.A(new_n26826_), .B(new_n26811_), .C(new_n26800_), .Y(new_n26827_));
  OAI21X1  g24391(.A0(new_n26827_), .A1(new_n23539_), .B0(new_n26781_), .Y(new_n26828_));
  AOI21X1  g24392(.A0(new_n26777_), .A1(new_n26763_), .B0(new_n26828_), .Y(new_n26829_));
  AOI21X1  g24393(.A0(new_n25268_), .A1(new_n2953_), .B0(new_n12684_), .Y(new_n26830_));
  AND2X1   g24394(.A(pi1091), .B(new_n2953_), .Y(new_n26831_));
  AOI21X1  g24395(.A0(new_n26831_), .A1(new_n25269_), .B0(new_n26743_), .Y(new_n26832_));
  NOR2X1   g24396(.A(new_n26832_), .B(new_n12684_), .Y(new_n26833_));
  NOR2X1   g24397(.A(new_n25342_), .B(new_n2722_), .Y(new_n26834_));
  AOI21X1  g24398(.A0(new_n26834_), .A1(new_n26830_), .B0(new_n26833_), .Y(new_n26835_));
  NOR3X1   g24399(.A(pi0299), .B(pi0200), .C(new_n7941_), .Y(new_n26836_));
  MX2X1    g24400(.A(new_n26836_), .B(new_n26673_), .S0(new_n2722_), .Y(new_n26837_));
  MX2X1    g24401(.A(pi1155), .B(new_n26673_), .S0(new_n2722_), .Y(new_n26838_));
  AND2X1   g24402(.A(new_n26838_), .B(new_n25053_), .Y(new_n26839_));
  OAI21X1  g24403(.A0(new_n26839_), .A1(new_n26837_), .B0(new_n12684_), .Y(new_n26840_));
  AOI21X1  g24404(.A0(new_n26840_), .A1(new_n26835_), .B0(new_n12706_), .Y(new_n26841_));
  OAI21X1  g24405(.A0(new_n25342_), .A1(new_n2722_), .B0(new_n26838_), .Y(new_n26842_));
  NAND2X1  g24406(.A(new_n26842_), .B(new_n12684_), .Y(new_n26843_));
  AND2X1   g24407(.A(pi1091), .B(pi0199), .Y(new_n26844_));
  AND2X1   g24408(.A(new_n26844_), .B(new_n2953_), .Y(new_n26845_));
  NOR3X1   g24409(.A(new_n26845_), .B(new_n26750_), .C(new_n12591_), .Y(new_n26846_));
  NOR2X1   g24410(.A(new_n26846_), .B(new_n12684_), .Y(new_n26847_));
  AOI21X1  g24411(.A0(new_n2722_), .A1(pi0243), .B0(pi1155), .Y(new_n26848_));
  OAI21X1  g24412(.A0(new_n8009_), .A1(pi0199), .B0(new_n26831_), .Y(new_n26849_));
  NAND2X1  g24413(.A(new_n26849_), .B(new_n26848_), .Y(new_n26850_));
  AOI21X1  g24414(.A0(new_n26850_), .A1(new_n26847_), .B0(pi1157), .Y(new_n26851_));
  AOI21X1  g24415(.A0(new_n26851_), .A1(new_n26843_), .B0(new_n26841_), .Y(new_n26852_));
  NAND2X1  g24416(.A(new_n26837_), .B(new_n12591_), .Y(new_n26853_));
  AOI21X1  g24417(.A0(new_n2722_), .A1(pi0243), .B0(new_n12591_), .Y(new_n26854_));
  AND2X1   g24418(.A(pi1091), .B(pi0200), .Y(new_n26855_));
  AND2X1   g24419(.A(new_n26855_), .B(new_n2953_), .Y(new_n26856_));
  INVX1    g24420(.A(new_n26856_), .Y(new_n26857_));
  AOI21X1  g24421(.A0(new_n26857_), .A1(new_n26854_), .B0(pi1156), .Y(new_n26858_));
  AOI22X1  g24422(.A0(new_n26858_), .A1(new_n26853_), .B0(new_n26847_), .B1(new_n26832_), .Y(new_n26859_));
  NOR2X1   g24423(.A(new_n26859_), .B(new_n12706_), .Y(new_n26860_));
  OR2X1    g24424(.A(new_n8547_), .B(new_n2722_), .Y(new_n26861_));
  AOI21X1  g24425(.A0(new_n26861_), .A1(new_n26848_), .B0(new_n26846_), .Y(new_n26862_));
  NOR4X1   g24426(.A(pi1156), .B(new_n2722_), .C(pi0299), .D(new_n8009_), .Y(new_n26863_));
  NOR2X1   g24427(.A(new_n26863_), .B(new_n26862_), .Y(new_n26864_));
  OAI21X1  g24428(.A0(new_n26864_), .A1(pi1157), .B0(new_n8548_), .Y(new_n26865_));
  OAI22X1  g24429(.A0(new_n26865_), .A1(new_n26860_), .B0(new_n26852_), .B1(new_n8548_), .Y(new_n26866_));
  NOR3X1   g24430(.A(new_n26833_), .B(new_n12706_), .C(new_n8548_), .Y(new_n26867_));
  AOI21X1  g24431(.A0(new_n26867_), .A1(new_n26840_), .B0(new_n23539_), .Y(new_n26868_));
  AND2X1   g24432(.A(pi1091), .B(pi0299), .Y(new_n26869_));
  INVX1    g24433(.A(new_n26869_), .Y(new_n26870_));
  AOI21X1  g24434(.A0(new_n26870_), .A1(new_n26864_), .B0(pi1157), .Y(new_n26871_));
  NAND2X1  g24435(.A(new_n25096_), .B(pi1091), .Y(new_n26872_));
  AOI22X1  g24436(.A0(new_n26872_), .A1(new_n26848_), .B0(new_n26857_), .B1(new_n26854_), .Y(new_n26873_));
  NOR2X1   g24437(.A(new_n26873_), .B(pi1156), .Y(new_n26874_));
  NOR3X1   g24438(.A(new_n26874_), .B(new_n12706_), .C(pi0211), .Y(new_n26875_));
  AOI21X1  g24439(.A0(new_n26875_), .A1(new_n26835_), .B0(new_n26871_), .Y(new_n26876_));
  AOI22X1  g24440(.A0(new_n26876_), .A1(new_n26868_), .B0(new_n26866_), .B1(new_n23539_), .Y(new_n26877_));
  OAI21X1  g24441(.A0(new_n26877_), .A1(new_n26781_), .B0(new_n6520_), .Y(new_n26878_));
  INVX1    g24442(.A(new_n26781_), .Y(new_n26879_));
  NOR3X1   g24443(.A(new_n26676_), .B(pi1091), .C(new_n3175_), .Y(new_n26880_));
  NOR4X1   g24444(.A(new_n26880_), .B(new_n26750_), .C(new_n12706_), .D(pi0211), .Y(new_n26881_));
  AOI21X1  g24445(.A0(new_n26744_), .A1(pi0243), .B0(new_n26881_), .Y(new_n26882_));
  OAI21X1  g24446(.A0(new_n26681_), .A1(pi0243), .B0(new_n26882_), .Y(new_n26883_));
  OR4X1    g24447(.A(new_n26689_), .B(new_n26679_), .C(pi1091), .D(new_n26673_), .Y(new_n26884_));
  MX2X1    g24448(.A(new_n12684_), .B(new_n12591_), .S0(new_n8548_), .Y(new_n26885_));
  INVX1    g24449(.A(new_n26885_), .Y(new_n26886_));
  OAI21X1  g24450(.A0(new_n26886_), .A1(new_n2722_), .B0(new_n23539_), .Y(new_n26887_));
  AOI21X1  g24451(.A0(new_n26689_), .A1(new_n26673_), .B0(new_n26887_), .Y(new_n26888_));
  AOI22X1  g24452(.A0(new_n26888_), .A1(new_n26884_), .B0(new_n26883_), .B1(pi0219), .Y(new_n26889_));
  AOI22X1  g24453(.A0(new_n26886_), .A1(new_n23539_), .B0(new_n25030_), .B1(pi1157), .Y(new_n26890_));
  MX2X1    g24454(.A(new_n26890_), .B(pi0243), .S0(new_n2722_), .Y(new_n26891_));
  OR2X1    g24455(.A(new_n26891_), .B(new_n26781_), .Y(new_n26892_));
  AND2X1   g24456(.A(new_n26892_), .B(po1038), .Y(new_n26893_));
  OAI21X1  g24457(.A0(new_n26889_), .A1(new_n26879_), .B0(new_n26893_), .Y(new_n26894_));
  INVX1    g24458(.A(pi0268), .Y(new_n26895_));
  INVX1    g24459(.A(pi0272), .Y(new_n26896_));
  INVX1    g24460(.A(pi0275), .Y(new_n26897_));
  INVX1    g24461(.A(pi0283), .Y(new_n26898_));
  NOR4X1   g24462(.A(new_n26898_), .B(new_n26897_), .C(new_n26896_), .D(new_n26895_), .Y(new_n26899_));
  AND2X1   g24463(.A(new_n26899_), .B(new_n26894_), .Y(new_n26900_));
  OAI21X1  g24464(.A0(new_n26878_), .A1(new_n26829_), .B0(new_n26900_), .Y(new_n26901_));
  NAND2X1  g24465(.A(new_n26877_), .B(new_n6520_), .Y(new_n26902_));
  AOI21X1  g24466(.A0(new_n26891_), .A1(po1038), .B0(new_n26899_), .Y(new_n26903_));
  AOI21X1  g24467(.A0(new_n26903_), .A1(new_n26902_), .B0(pi0230), .Y(new_n26904_));
  OR2X1    g24468(.A(new_n26890_), .B(new_n11776_), .Y(new_n26905_));
  OAI22X1  g24469(.A0(new_n8135_), .A1(pi1155), .B0(pi1156), .B1(new_n8009_), .Y(new_n26906_));
  AOI21X1  g24470(.A0(new_n25760_), .A1(pi0199), .B0(new_n26906_), .Y(new_n26907_));
  AOI21X1  g24471(.A0(new_n26907_), .A1(new_n11776_), .B0(new_n24954_), .Y(new_n26908_));
  AOI22X1  g24472(.A0(new_n26908_), .A1(new_n26905_), .B0(new_n26904_), .B1(new_n26901_), .Y(po0400));
  INVX1    g24473(.A(new_n25217_), .Y(new_n26910_));
  AOI22X1  g24474(.A0(new_n26340_), .A1(new_n26401_), .B0(new_n26321_), .B1(new_n26910_), .Y(new_n26911_));
  OAI21X1  g24475(.A0(new_n26911_), .A1(new_n26328_), .B0(pi0214), .Y(new_n26912_));
  NAND2X1  g24476(.A(new_n26912_), .B(new_n26394_), .Y(new_n26913_));
  INVX1    g24477(.A(new_n26328_), .Y(new_n26914_));
  OAI21X1  g24478(.A0(new_n26294_), .A1(new_n24960_), .B0(pi0212), .Y(new_n26915_));
  AOI21X1  g24479(.A0(new_n26911_), .A1(new_n24984_), .B0(new_n26915_), .Y(new_n26916_));
  AOI21X1  g24480(.A0(new_n26916_), .A1(new_n26914_), .B0(pi0219), .Y(new_n26917_));
  NOR3X1   g24481(.A(new_n26389_), .B(new_n25189_), .C(pi0211), .Y(new_n26918_));
  NOR2X1   g24482(.A(new_n26918_), .B(new_n26388_), .Y(new_n26919_));
  OAI21X1  g24483(.A0(new_n26919_), .A1(new_n26387_), .B0(new_n26363_), .Y(new_n26920_));
  AOI21X1  g24484(.A0(new_n26917_), .A1(new_n26913_), .B0(new_n26920_), .Y(new_n26921_));
  INVX1    g24485(.A(new_n26331_), .Y(new_n26922_));
  AND2X1   g24486(.A(new_n26916_), .B(new_n26922_), .Y(new_n26923_));
  AOI21X1  g24487(.A0(new_n26911_), .A1(pi0214), .B0(new_n26371_), .Y(new_n26924_));
  OR2X1    g24488(.A(new_n26924_), .B(pi0219), .Y(new_n26925_));
  OAI21X1  g24489(.A0(new_n25652_), .A1(new_n2953_), .B0(pi1147), .Y(new_n26926_));
  NOR2X1   g24490(.A(new_n26926_), .B(new_n26358_), .Y(new_n26927_));
  OAI21X1  g24491(.A0(new_n26925_), .A1(new_n26923_), .B0(new_n26927_), .Y(new_n26928_));
  NAND3X1  g24492(.A(new_n26928_), .B(new_n25653_), .C(new_n25003_), .Y(new_n26929_));
  OAI22X1  g24493(.A0(new_n26929_), .A1(new_n26921_), .B0(new_n26412_), .B1(new_n25003_), .Y(new_n26930_));
  NOR3X1   g24494(.A(new_n26244_), .B(new_n26224_), .C(pi1147), .Y(new_n26931_));
  NOR2X1   g24495(.A(new_n26931_), .B(new_n26227_), .Y(new_n26932_));
  OAI21X1  g24496(.A0(new_n26221_), .A1(new_n2953_), .B0(new_n26243_), .Y(new_n26933_));
  OAI21X1  g24497(.A0(new_n26233_), .A1(new_n25014_), .B0(new_n25253_), .Y(new_n26934_));
  AOI21X1  g24498(.A0(new_n26236_), .A1(new_n25014_), .B0(new_n26934_), .Y(new_n26935_));
  NAND2X1  g24499(.A(new_n26935_), .B(new_n26933_), .Y(new_n26936_));
  NOR2X1   g24500(.A(new_n26253_), .B(new_n25640_), .Y(new_n26937_));
  AOI21X1  g24501(.A0(new_n26937_), .A1(new_n26936_), .B0(po1038), .Y(new_n26938_));
  OAI21X1  g24502(.A0(new_n26938_), .A1(new_n26932_), .B0(pi0213), .Y(new_n26939_));
  AOI21X1  g24503(.A0(new_n25657_), .A1(new_n25003_), .B0(pi0209), .Y(new_n26940_));
  AOI22X1  g24504(.A0(new_n26940_), .A1(new_n26939_), .B0(new_n26930_), .B1(pi0209), .Y(new_n26941_));
  MX2X1    g24505(.A(new_n26941_), .B(pi0244), .S0(new_n24954_), .Y(po0401));
  NOR4X1   g24506(.A(new_n24957_), .B(new_n8034_), .C(new_n6520_), .D(new_n3165_), .Y(new_n26943_));
  NOR2X1   g24507(.A(new_n26943_), .B(pi1147), .Y(new_n26944_));
  OAI21X1  g24508(.A0(new_n26158_), .A1(new_n25969_), .B0(new_n26944_), .Y(new_n26945_));
  OR2X1    g24509(.A(new_n26639_), .B(pi0211), .Y(new_n26946_));
  OR2X1    g24510(.A(new_n26946_), .B(new_n24955_), .Y(new_n26947_));
  AOI21X1  g24511(.A0(new_n26947_), .A1(new_n26650_), .B0(po1038), .Y(new_n26948_));
  AND2X1   g24512(.A(new_n26282_), .B(pi0214), .Y(new_n26949_));
  OAI21X1  g24513(.A0(new_n26640_), .A1(pi0299), .B0(new_n26949_), .Y(new_n26950_));
  NAND2X1  g24514(.A(new_n26950_), .B(pi0212), .Y(new_n26951_));
  NOR4X1   g24515(.A(new_n26632_), .B(new_n26631_), .C(new_n25751_), .D(pi0299), .Y(new_n26952_));
  OAI21X1  g24516(.A0(new_n26952_), .A1(pi0211), .B0(new_n26644_), .Y(new_n26953_));
  NOR2X1   g24517(.A(new_n26953_), .B(pi0214), .Y(new_n26954_));
  AOI21X1  g24518(.A0(new_n26953_), .A1(new_n26645_), .B0(pi0219), .Y(new_n26955_));
  OAI21X1  g24519(.A0(new_n26954_), .A1(new_n26951_), .B0(new_n26955_), .Y(new_n26956_));
  AOI21X1  g24520(.A0(new_n26956_), .A1(new_n26948_), .B0(new_n26945_), .Y(new_n26957_));
  OR2X1    g24521(.A(new_n25955_), .B(new_n26091_), .Y(new_n26958_));
  NOR2X1   g24522(.A(new_n26958_), .B(new_n26943_), .Y(new_n26959_));
  MX2X1    g24523(.A(new_n26952_), .B(new_n26639_), .S0(pi0211), .Y(new_n26960_));
  MX2X1    g24524(.A(new_n26960_), .B(new_n26952_), .S0(new_n24984_), .Y(new_n26961_));
  NOR2X1   g24525(.A(new_n26961_), .B(new_n24961_), .Y(new_n26962_));
  OAI21X1  g24526(.A0(new_n26952_), .A1(new_n26646_), .B0(new_n23539_), .Y(new_n26963_));
  OAI21X1  g24527(.A0(new_n26963_), .A1(new_n26962_), .B0(new_n26948_), .Y(new_n26964_));
  AND2X1   g24528(.A(new_n26964_), .B(new_n26959_), .Y(new_n26965_));
  NOR3X1   g24529(.A(new_n26965_), .B(new_n26957_), .C(new_n26273_), .Y(new_n26966_));
  INVX1    g24530(.A(new_n26152_), .Y(new_n26967_));
  AOI21X1  g24531(.A0(new_n26967_), .A1(pi1147), .B0(new_n26959_), .Y(new_n26968_));
  INVX1    g24532(.A(new_n26968_), .Y(new_n26969_));
  AND2X1   g24533(.A(new_n26644_), .B(new_n26199_), .Y(new_n26970_));
  MX2X1    g24534(.A(new_n26970_), .B(new_n26960_), .S0(pi0214), .Y(new_n26971_));
  NOR2X1   g24535(.A(new_n26971_), .B(new_n24961_), .Y(new_n26972_));
  OAI21X1  g24536(.A0(new_n26970_), .A1(new_n26646_), .B0(new_n23539_), .Y(new_n26973_));
  OAI21X1  g24537(.A0(new_n26973_), .A1(new_n26972_), .B0(new_n26948_), .Y(new_n26974_));
  AND2X1   g24538(.A(new_n26974_), .B(new_n26969_), .Y(new_n26975_));
  INVX1    g24539(.A(new_n26944_), .Y(new_n26976_));
  AND2X1   g24540(.A(new_n26644_), .B(new_n24984_), .Y(new_n26977_));
  AOI21X1  g24541(.A0(new_n26649_), .A1(new_n24961_), .B0(pi0219), .Y(new_n26978_));
  OAI21X1  g24542(.A0(new_n26951_), .A1(new_n26977_), .B0(new_n26978_), .Y(new_n26979_));
  AOI21X1  g24543(.A0(new_n26979_), .A1(new_n26948_), .B0(new_n26976_), .Y(new_n26980_));
  NOR3X1   g24544(.A(new_n26980_), .B(new_n26975_), .C(pi1148), .Y(new_n26981_));
  OAI21X1  g24545(.A0(new_n26981_), .A1(new_n26966_), .B0(pi0213), .Y(new_n26982_));
  AOI21X1  g24546(.A0(new_n26653_), .A1(new_n26623_), .B0(pi0213), .Y(new_n26983_));
  NOR2X1   g24547(.A(new_n26983_), .B(pi0209), .Y(new_n26984_));
  INVX1    g24548(.A(new_n26945_), .Y(new_n26985_));
  AOI21X1  g24549(.A0(pi1146), .A1(pi0199), .B0(pi0200), .Y(new_n26986_));
  OR4X1    g24550(.A(new_n26986_), .B(new_n26310_), .C(pi0299), .D(new_n22803_), .Y(new_n26987_));
  OAI21X1  g24551(.A0(new_n25096_), .A1(new_n3165_), .B0(new_n26987_), .Y(new_n26988_));
  AND2X1   g24552(.A(new_n26988_), .B(pi0208), .Y(new_n26989_));
  NOR3X1   g24553(.A(pi1146), .B(pi0200), .C(new_n7941_), .Y(new_n26990_));
  NOR4X1   g24554(.A(new_n26990_), .B(new_n26310_), .C(pi0299), .D(new_n23109_), .Y(new_n26991_));
  NOR2X1   g24555(.A(new_n26991_), .B(pi0207), .Y(new_n26992_));
  NOR4X1   g24556(.A(new_n26992_), .B(new_n26990_), .C(new_n25054_), .D(new_n7896_), .Y(new_n26993_));
  AND2X1   g24557(.A(new_n26261_), .B(new_n23109_), .Y(new_n26994_));
  NOR3X1   g24558(.A(new_n26994_), .B(new_n26993_), .C(new_n26989_), .Y(new_n26995_));
  NOR2X1   g24559(.A(new_n26995_), .B(pi0299), .Y(new_n26996_));
  INVX1    g24560(.A(new_n26996_), .Y(new_n26997_));
  AOI21X1  g24561(.A0(new_n26997_), .A1(new_n24984_), .B0(pi0212), .Y(new_n26998_));
  INVX1    g24562(.A(new_n26998_), .Y(new_n26999_));
  NOR3X1   g24563(.A(new_n26986_), .B(new_n26310_), .C(pi0299), .Y(new_n27000_));
  OAI21X1  g24564(.A0(new_n25799_), .A1(new_n7896_), .B0(new_n27000_), .Y(new_n27001_));
  NOR2X1   g24565(.A(new_n27000_), .B(pi0299), .Y(new_n27002_));
  NOR2X1   g24566(.A(new_n27002_), .B(new_n26995_), .Y(new_n27003_));
  NOR2X1   g24567(.A(new_n27003_), .B(pi0299), .Y(new_n27004_));
  MX2X1    g24568(.A(new_n27004_), .B(new_n27001_), .S0(pi0211), .Y(new_n27005_));
  AND2X1   g24569(.A(new_n27005_), .B(new_n26997_), .Y(new_n27006_));
  OAI21X1  g24570(.A0(new_n27006_), .A1(new_n26999_), .B0(new_n23539_), .Y(new_n27007_));
  OAI21X1  g24571(.A0(new_n26995_), .A1(pi0299), .B0(new_n26949_), .Y(new_n27008_));
  AOI21X1  g24572(.A0(new_n27006_), .A1(new_n24984_), .B0(new_n24961_), .Y(new_n27009_));
  AOI21X1  g24573(.A0(new_n27009_), .A1(new_n27008_), .B0(new_n27007_), .Y(new_n27010_));
  AOI21X1  g24574(.A0(new_n26996_), .A1(new_n24994_), .B0(new_n23539_), .Y(new_n27011_));
  OAI21X1  g24575(.A0(new_n26995_), .A1(new_n24994_), .B0(new_n27011_), .Y(new_n27012_));
  NAND2X1  g24576(.A(new_n27012_), .B(new_n6520_), .Y(new_n27013_));
  OAI21X1  g24577(.A0(new_n27013_), .A1(new_n27010_), .B0(new_n26985_), .Y(new_n27014_));
  NOR2X1   g24578(.A(new_n26990_), .B(new_n25069_), .Y(new_n27015_));
  NOR2X1   g24579(.A(new_n27015_), .B(new_n7896_), .Y(new_n27016_));
  NOR4X1   g24580(.A(new_n26990_), .B(new_n26310_), .C(pi0299), .D(new_n22803_), .Y(new_n27017_));
  INVX1    g24581(.A(new_n27017_), .Y(new_n27018_));
  AOI21X1  g24582(.A0(new_n27018_), .A1(new_n26178_), .B0(new_n27016_), .Y(new_n27019_));
  OR2X1    g24583(.A(new_n27019_), .B(pi0214), .Y(new_n27020_));
  AND2X1   g24584(.A(new_n27020_), .B(new_n24961_), .Y(new_n27021_));
  NOR3X1   g24585(.A(new_n26986_), .B(new_n25268_), .C(pi0299), .Y(new_n27022_));
  AOI21X1  g24586(.A0(new_n27022_), .A1(new_n22803_), .B0(new_n26261_), .Y(new_n27023_));
  AOI21X1  g24587(.A0(new_n27023_), .A1(new_n27018_), .B0(new_n23109_), .Y(new_n27024_));
  INVX1    g24588(.A(new_n27024_), .Y(new_n27025_));
  AOI21X1  g24589(.A0(new_n27015_), .A1(new_n24980_), .B0(new_n26991_), .Y(new_n27026_));
  OAI21X1  g24590(.A0(new_n27025_), .A1(pi0299), .B0(new_n27026_), .Y(new_n27027_));
  OAI21X1  g24591(.A0(new_n27027_), .A1(pi0299), .B0(new_n27021_), .Y(new_n27028_));
  NAND2X1  g24592(.A(new_n27028_), .B(new_n23539_), .Y(new_n27029_));
  NOR2X1   g24593(.A(new_n27027_), .B(pi0299), .Y(new_n27030_));
  NOR3X1   g24594(.A(new_n27027_), .B(new_n26261_), .C(new_n25740_), .Y(new_n27031_));
  NOR3X1   g24595(.A(new_n27031_), .B(new_n27030_), .C(new_n24961_), .Y(new_n27032_));
  AOI21X1  g24596(.A0(new_n27019_), .A1(new_n24994_), .B0(new_n23539_), .Y(new_n27033_));
  OAI21X1  g24597(.A0(new_n27027_), .A1(new_n26261_), .B0(new_n24956_), .Y(new_n27034_));
  AOI21X1  g24598(.A0(new_n27034_), .A1(new_n27033_), .B0(po1038), .Y(new_n27035_));
  OAI21X1  g24599(.A0(new_n27032_), .A1(new_n27029_), .B0(new_n27035_), .Y(new_n27036_));
  AOI21X1  g24600(.A0(new_n27036_), .A1(new_n26959_), .B0(new_n26273_), .Y(new_n27037_));
  OAI22X1  g24601(.A0(new_n27022_), .A1(new_n7896_), .B0(new_n27017_), .B1(new_n25259_), .Y(new_n27038_));
  AND2X1   g24602(.A(new_n27038_), .B(new_n26199_), .Y(new_n27039_));
  INVX1    g24603(.A(new_n27039_), .Y(new_n27040_));
  NOR2X1   g24604(.A(new_n27038_), .B(pi0214), .Y(new_n27041_));
  NOR2X1   g24605(.A(new_n27041_), .B(pi0212), .Y(new_n27042_));
  INVX1    g24606(.A(new_n27042_), .Y(new_n27043_));
  AOI21X1  g24607(.A0(new_n27040_), .A1(pi0214), .B0(new_n27043_), .Y(new_n27044_));
  OR2X1    g24608(.A(new_n27039_), .B(pi0214), .Y(new_n27045_));
  AND2X1   g24609(.A(new_n27022_), .B(new_n24980_), .Y(new_n27046_));
  NOR4X1   g24610(.A(new_n27046_), .B(new_n27024_), .C(new_n26994_), .D(pi0299), .Y(new_n27047_));
  NOR2X1   g24611(.A(new_n27047_), .B(new_n24984_), .Y(new_n27048_));
  NOR2X1   g24612(.A(new_n27030_), .B(pi0211), .Y(new_n27049_));
  OAI21X1  g24613(.A0(new_n27049_), .A1(new_n27019_), .B0(new_n27048_), .Y(new_n27050_));
  AND2X1   g24614(.A(new_n27050_), .B(pi0212), .Y(new_n27051_));
  AND2X1   g24615(.A(new_n27051_), .B(new_n27045_), .Y(new_n27052_));
  OAI21X1  g24616(.A0(new_n27052_), .A1(new_n27044_), .B0(new_n23539_), .Y(new_n27053_));
  AOI21X1  g24617(.A0(new_n25741_), .A1(new_n3165_), .B0(new_n26300_), .Y(new_n27054_));
  NOR3X1   g24618(.A(new_n27046_), .B(new_n27024_), .C(new_n26994_), .Y(new_n27055_));
  INVX1    g24619(.A(new_n27038_), .Y(new_n27056_));
  AOI21X1  g24620(.A0(new_n27056_), .A1(new_n25323_), .B0(new_n24956_), .Y(new_n27057_));
  AOI21X1  g24621(.A0(new_n27041_), .A1(new_n24961_), .B0(new_n23539_), .Y(new_n27058_));
  OAI21X1  g24622(.A0(new_n27057_), .A1(new_n27055_), .B0(new_n27058_), .Y(new_n27059_));
  AND2X1   g24623(.A(new_n27059_), .B(new_n6520_), .Y(new_n27060_));
  OAI21X1  g24624(.A0(new_n27054_), .A1(new_n27053_), .B0(new_n27060_), .Y(new_n27061_));
  OAI21X1  g24625(.A0(new_n26996_), .A1(new_n26542_), .B0(new_n26988_), .Y(new_n27062_));
  AND2X1   g24626(.A(new_n27062_), .B(new_n23539_), .Y(new_n27063_));
  OAI21X1  g24627(.A0(new_n27001_), .A1(new_n25323_), .B0(pi0219), .Y(new_n27064_));
  AOI21X1  g24628(.A0(new_n27001_), .A1(pi0211), .B0(new_n24955_), .Y(new_n27065_));
  AOI21X1  g24629(.A0(new_n27065_), .A1(new_n27003_), .B0(new_n27064_), .Y(new_n27066_));
  NOR3X1   g24630(.A(new_n27066_), .B(new_n27063_), .C(po1038), .Y(new_n27067_));
  OAI21X1  g24631(.A0(new_n27067_), .A1(new_n26976_), .B0(new_n26273_), .Y(new_n27068_));
  AOI21X1  g24632(.A0(new_n27061_), .A1(new_n26969_), .B0(new_n27068_), .Y(new_n27069_));
  AOI21X1  g24633(.A0(new_n27037_), .A1(new_n27014_), .B0(new_n27069_), .Y(new_n27070_));
  OR2X1    g24634(.A(new_n27070_), .B(new_n25003_), .Y(new_n27071_));
  NOR2X1   g24635(.A(new_n27004_), .B(new_n24984_), .Y(new_n27072_));
  OAI21X1  g24636(.A0(new_n26996_), .A1(new_n26233_), .B0(new_n27072_), .Y(new_n27073_));
  OAI21X1  g24637(.A0(new_n27001_), .A1(pi0214), .B0(new_n27073_), .Y(new_n27074_));
  NOR2X1   g24638(.A(new_n26616_), .B(new_n2953_), .Y(new_n27075_));
  INVX1    g24639(.A(new_n27075_), .Y(new_n27076_));
  AOI21X1  g24640(.A0(new_n27076_), .A1(new_n26997_), .B0(new_n24961_), .Y(new_n27077_));
  OAI21X1  g24641(.A0(new_n27000_), .A1(pi0299), .B0(new_n27077_), .Y(new_n27078_));
  NAND2X1  g24642(.A(new_n27078_), .B(new_n23539_), .Y(new_n27079_));
  AOI21X1  g24643(.A0(new_n27074_), .A1(new_n24961_), .B0(new_n27079_), .Y(new_n27080_));
  INVX1    g24644(.A(new_n26363_), .Y(new_n27081_));
  OAI21X1  g24645(.A0(new_n27004_), .A1(new_n25217_), .B0(new_n8548_), .Y(new_n27082_));
  AOI21X1  g24646(.A0(new_n27082_), .A1(new_n27065_), .B0(new_n27064_), .Y(new_n27083_));
  OR2X1    g24647(.A(new_n27083_), .B(new_n27081_), .Y(new_n27084_));
  OR2X1    g24648(.A(new_n27027_), .B(new_n26233_), .Y(new_n27085_));
  AOI21X1  g24649(.A0(new_n27085_), .A1(new_n27048_), .B0(new_n27041_), .Y(new_n27086_));
  INVX1    g24650(.A(new_n27047_), .Y(new_n27087_));
  INVX1    g24651(.A(new_n27027_), .Y(new_n27088_));
  AOI21X1  g24652(.A0(new_n27076_), .A1(new_n27088_), .B0(new_n24961_), .Y(new_n27089_));
  AOI21X1  g24653(.A0(new_n27089_), .A1(new_n27087_), .B0(pi0219), .Y(new_n27090_));
  OAI21X1  g24654(.A0(new_n27086_), .A1(pi0212), .B0(new_n27090_), .Y(new_n27091_));
  INVX1    g24655(.A(new_n27057_), .Y(new_n27092_));
  AOI21X1  g24656(.A0(new_n27088_), .A1(new_n25216_), .B0(new_n27047_), .Y(new_n27093_));
  OAI21X1  g24657(.A0(new_n27093_), .A1(pi0211), .B0(new_n27092_), .Y(new_n27094_));
  AND2X1   g24658(.A(new_n6520_), .B(pi1147), .Y(new_n27095_));
  INVX1    g24659(.A(new_n27095_), .Y(new_n27096_));
  AOI21X1  g24660(.A0(new_n27094_), .A1(new_n27058_), .B0(new_n27096_), .Y(new_n27097_));
  OR2X1    g24661(.A(new_n26622_), .B(pi1148), .Y(new_n27098_));
  AOI21X1  g24662(.A0(new_n27097_), .A1(new_n27091_), .B0(new_n27098_), .Y(new_n27099_));
  OAI21X1  g24663(.A0(new_n27084_), .A1(new_n27080_), .B0(new_n27099_), .Y(new_n27100_));
  AOI21X1  g24664(.A0(new_n26997_), .A1(new_n26234_), .B0(new_n26999_), .Y(new_n27101_));
  NOR3X1   g24665(.A(new_n27101_), .B(new_n27077_), .C(pi0219), .Y(new_n27102_));
  INVX1    g24666(.A(new_n27011_), .Y(new_n27103_));
  OR4X1    g24667(.A(new_n26994_), .B(new_n26993_), .C(new_n26989_), .D(pi0299), .Y(new_n27104_));
  AND2X1   g24668(.A(new_n27104_), .B(new_n24956_), .Y(new_n27105_));
  AOI21X1  g24669(.A0(new_n27105_), .A1(new_n26910_), .B0(new_n27103_), .Y(new_n27106_));
  OR4X1    g24670(.A(new_n27106_), .B(new_n27102_), .C(po1038), .D(pi1147), .Y(new_n27107_));
  OAI21X1  g24671(.A0(new_n27085_), .A1(new_n24984_), .B0(new_n27021_), .Y(new_n27108_));
  NOR2X1   g24672(.A(new_n27089_), .B(pi0219), .Y(new_n27109_));
  NAND2X1  g24673(.A(new_n27109_), .B(new_n27108_), .Y(new_n27110_));
  OAI21X1  g24674(.A0(new_n27027_), .A1(new_n25215_), .B0(new_n24956_), .Y(new_n27111_));
  AOI21X1  g24675(.A0(new_n27111_), .A1(new_n27033_), .B0(new_n27096_), .Y(new_n27112_));
  OR2X1    g24676(.A(new_n26622_), .B(new_n26273_), .Y(new_n27113_));
  AOI21X1  g24677(.A0(new_n27112_), .A1(new_n27110_), .B0(new_n27113_), .Y(new_n27114_));
  AOI21X1  g24678(.A0(new_n27114_), .A1(new_n27107_), .B0(pi0213), .Y(new_n27115_));
  AOI21X1  g24679(.A0(new_n27115_), .A1(new_n27100_), .B0(new_n23244_), .Y(new_n27116_));
  AOI22X1  g24680(.A0(new_n27116_), .A1(new_n27071_), .B0(new_n26984_), .B1(new_n26982_), .Y(new_n27117_));
  MX2X1    g24681(.A(new_n27117_), .B(pi0245), .S0(new_n24954_), .Y(po0402));
  OR4X1    g24682(.A(new_n26152_), .B(new_n26151_), .C(new_n26150_), .D(pi1150), .Y(new_n27119_));
  OR4X1    g24683(.A(new_n26116_), .B(new_n26114_), .C(new_n26111_), .D(new_n26471_), .Y(new_n27120_));
  NAND3X1  g24684(.A(new_n27120_), .B(new_n27119_), .C(pi1149), .Y(new_n27121_));
  OAI22X1  g24685(.A0(new_n26175_), .A1(new_n26170_), .B0(new_n26158_), .B1(new_n25929_), .Y(new_n27122_));
  AOI21X1  g24686(.A0(new_n26212_), .A1(new_n26471_), .B0(pi1149), .Y(new_n27123_));
  OAI21X1  g24687(.A0(new_n27122_), .A1(new_n26471_), .B0(new_n27123_), .Y(new_n27124_));
  AND2X1   g24688(.A(new_n27124_), .B(new_n27121_), .Y(new_n27125_));
  NOR3X1   g24689(.A(new_n26145_), .B(new_n26121_), .C(pi1150), .Y(new_n27126_));
  INVX1    g24690(.A(new_n27126_), .Y(new_n27127_));
  AOI21X1  g24691(.A0(new_n26108_), .A1(pi1150), .B0(new_n26147_), .Y(new_n27128_));
  NOR3X1   g24692(.A(new_n26182_), .B(new_n26471_), .C(pi1149), .Y(new_n27129_));
  AOI21X1  g24693(.A0(new_n27128_), .A1(new_n27127_), .B0(new_n27129_), .Y(new_n27130_));
  MX2X1    g24694(.A(new_n27130_), .B(new_n27125_), .S0(pi1148), .Y(new_n27131_));
  NOR2X1   g24695(.A(new_n27131_), .B(new_n25003_), .Y(new_n27132_));
  INVX1    g24696(.A(new_n26151_), .Y(new_n27133_));
  AND2X1   g24697(.A(new_n26193_), .B(new_n7941_), .Y(new_n27134_));
  NOR2X1   g24698(.A(new_n26261_), .B(new_n23539_), .Y(new_n27135_));
  NOR3X1   g24699(.A(new_n27135_), .B(new_n24957_), .C(po1038), .Y(new_n27136_));
  INVX1    g24700(.A(new_n27136_), .Y(new_n27137_));
  OAI21X1  g24701(.A0(new_n27134_), .A1(new_n27133_), .B0(new_n27137_), .Y(new_n27138_));
  NOR2X1   g24702(.A(new_n26194_), .B(new_n26112_), .Y(new_n27139_));
  OAI22X1  g24703(.A0(new_n26194_), .A1(pi0299), .B0(new_n26199_), .B1(pi1146), .Y(new_n27140_));
  AOI21X1  g24704(.A0(new_n27140_), .A1(new_n24962_), .B0(new_n27139_), .Y(new_n27141_));
  OAI21X1  g24705(.A0(new_n27141_), .A1(pi0219), .B0(new_n27138_), .Y(new_n27142_));
  OAI21X1  g24706(.A0(new_n26959_), .A1(new_n26985_), .B0(new_n27142_), .Y(new_n27143_));
  OAI22X1  g24707(.A0(new_n26205_), .A1(new_n26203_), .B0(new_n26196_), .B1(pi0219), .Y(new_n27144_));
  AOI21X1  g24708(.A0(new_n27144_), .A1(new_n26985_), .B0(pi1150), .Y(new_n27145_));
  NOR2X1   g24709(.A(new_n27136_), .B(new_n26259_), .Y(new_n27146_));
  OR2X1    g24710(.A(new_n26265_), .B(new_n24984_), .Y(new_n27147_));
  INVX1    g24711(.A(new_n26445_), .Y(new_n27148_));
  AOI21X1  g24712(.A0(new_n26439_), .A1(new_n24961_), .B0(pi0219), .Y(new_n27149_));
  NAND2X1  g24713(.A(new_n27149_), .B(new_n27148_), .Y(new_n27150_));
  AOI21X1  g24714(.A0(new_n26436_), .A1(new_n27147_), .B0(new_n27150_), .Y(new_n27151_));
  OAI21X1  g24715(.A0(new_n27151_), .A1(new_n27146_), .B0(new_n26959_), .Y(new_n27152_));
  INVX1    g24716(.A(new_n26167_), .Y(new_n27153_));
  NAND2X1  g24717(.A(new_n26264_), .B(pi0211), .Y(new_n27154_));
  AOI21X1  g24718(.A0(new_n26439_), .A1(new_n8548_), .B0(new_n24984_), .Y(new_n27155_));
  OAI21X1  g24719(.A0(new_n26172_), .A1(pi0214), .B0(pi0212), .Y(new_n27156_));
  AOI21X1  g24720(.A0(new_n27155_), .A1(new_n27154_), .B0(new_n27156_), .Y(new_n27157_));
  OAI22X1  g24721(.A0(new_n27157_), .A1(new_n27153_), .B0(new_n27136_), .B1(new_n26259_), .Y(new_n27158_));
  AOI21X1  g24722(.A0(new_n27158_), .A1(new_n26985_), .B0(new_n26471_), .Y(new_n27159_));
  AOI22X1  g24723(.A0(new_n27159_), .A1(new_n27152_), .B0(new_n27145_), .B1(new_n27143_), .Y(new_n27160_));
  AOI21X1  g24724(.A0(pi1146), .A1(pi0211), .B0(pi0219), .Y(new_n27161_));
  OR4X1    g24725(.A(new_n27161_), .B(new_n27135_), .C(new_n26543_), .D(new_n26208_), .Y(new_n27162_));
  AOI22X1  g24726(.A0(new_n27162_), .A1(new_n26944_), .B0(new_n27137_), .B1(new_n26969_), .Y(new_n27163_));
  AND2X1   g24727(.A(new_n26179_), .B(pi1150), .Y(new_n27164_));
  AND2X1   g24728(.A(new_n25827_), .B(pi1150), .Y(new_n27165_));
  NOR4X1   g24729(.A(new_n2953_), .B(new_n24984_), .C(pi0212), .D(new_n8548_), .Y(new_n27166_));
  NOR4X1   g24730(.A(new_n27166_), .B(new_n27165_), .C(new_n27054_), .D(pi0219), .Y(new_n27167_));
  AOI21X1  g24731(.A0(new_n27167_), .A1(new_n26969_), .B0(pi1148), .Y(new_n27168_));
  OAI21X1  g24732(.A0(new_n27164_), .A1(new_n27163_), .B0(new_n27168_), .Y(new_n27169_));
  OAI21X1  g24733(.A0(new_n27160_), .A1(new_n26273_), .B0(new_n27169_), .Y(new_n27170_));
  AOI21X1  g24734(.A0(new_n26293_), .A1(new_n26216_), .B0(new_n26124_), .Y(new_n27171_));
  AOI21X1  g24735(.A0(new_n26132_), .A1(new_n26207_), .B0(new_n26143_), .Y(new_n27172_));
  INVX1    g24736(.A(new_n27172_), .Y(new_n27173_));
  OAI21X1  g24737(.A0(new_n26142_), .A1(pi1146), .B0(new_n27173_), .Y(new_n27174_));
  AOI21X1  g24738(.A0(new_n27171_), .A1(new_n26141_), .B0(new_n27174_), .Y(new_n27175_));
  OAI22X1  g24739(.A0(new_n26125_), .A1(new_n26124_), .B0(new_n25831_), .B1(pi0212), .Y(new_n27176_));
  AOI21X1  g24740(.A0(new_n27176_), .A1(new_n23539_), .B0(new_n27172_), .Y(new_n27177_));
  OAI21X1  g24741(.A0(new_n26124_), .A1(pi1146), .B0(new_n27177_), .Y(new_n27178_));
  AOI21X1  g24742(.A0(new_n27178_), .A1(new_n26944_), .B0(pi1150), .Y(new_n27179_));
  OAI21X1  g24743(.A0(new_n27175_), .A1(new_n26968_), .B0(new_n27179_), .Y(new_n27180_));
  NAND2X1  g24744(.A(new_n26588_), .B(new_n24984_), .Y(new_n27181_));
  AOI21X1  g24745(.A0(new_n27181_), .A1(new_n26105_), .B0(pi0219), .Y(new_n27182_));
  OR2X1    g24746(.A(new_n26588_), .B(new_n26095_), .Y(new_n27183_));
  OAI21X1  g24747(.A0(new_n27183_), .A1(pi0212), .B0(new_n27182_), .Y(new_n27184_));
  NAND3X1  g24748(.A(new_n25851_), .B(new_n2953_), .C(pi0208), .Y(new_n27185_));
  NAND3X1  g24749(.A(new_n27185_), .B(new_n26262_), .C(new_n26098_), .Y(new_n27186_));
  OR4X1    g24750(.A(new_n26278_), .B(new_n8503_), .C(new_n5118_), .D(pi0057), .Y(new_n27187_));
  AOI22X1  g24751(.A0(new_n27183_), .A1(new_n27182_), .B0(new_n27137_), .B1(new_n27187_), .Y(new_n27188_));
  OAI21X1  g24752(.A0(new_n27186_), .A1(new_n27184_), .B0(new_n27188_), .Y(new_n27189_));
  OAI21X1  g24753(.A0(new_n26104_), .A1(new_n26281_), .B0(new_n23539_), .Y(new_n27190_));
  OAI21X1  g24754(.A0(new_n27190_), .A1(new_n26591_), .B0(new_n26279_), .Y(new_n27191_));
  AOI21X1  g24755(.A0(new_n27189_), .A1(new_n26094_), .B0(new_n27191_), .Y(new_n27192_));
  AOI21X1  g24756(.A0(new_n27189_), .A1(new_n26969_), .B0(new_n26471_), .Y(new_n27193_));
  OAI21X1  g24757(.A0(new_n27192_), .A1(new_n26976_), .B0(new_n27193_), .Y(new_n27194_));
  NAND3X1  g24758(.A(new_n27194_), .B(new_n27180_), .C(new_n26273_), .Y(new_n27195_));
  INVX1    g24759(.A(new_n26959_), .Y(new_n27196_));
  AND2X1   g24760(.A(new_n27196_), .B(new_n26945_), .Y(new_n27197_));
  OAI21X1  g24761(.A0(new_n25984_), .A1(new_n25884_), .B0(new_n26203_), .Y(new_n27198_));
  INVX1    g24762(.A(new_n27198_), .Y(new_n27199_));
  OAI21X1  g24763(.A0(new_n27199_), .A1(new_n26190_), .B0(new_n26945_), .Y(new_n27200_));
  NAND2X1  g24764(.A(new_n26949_), .B(new_n25883_), .Y(new_n27201_));
  AOI21X1  g24765(.A0(new_n27201_), .A1(new_n26202_), .B0(new_n26205_), .Y(new_n27202_));
  AOI22X1  g24766(.A0(new_n27202_), .A1(new_n27200_), .B0(new_n27137_), .B1(new_n27133_), .Y(new_n27203_));
  OAI21X1  g24767(.A0(new_n27203_), .A1(new_n27197_), .B0(new_n26471_), .Y(new_n27204_));
  NAND3X1  g24768(.A(new_n27162_), .B(new_n26985_), .C(new_n26303_), .Y(new_n27205_));
  OAI21X1  g24769(.A0(new_n26292_), .A1(new_n24984_), .B0(new_n26298_), .Y(new_n27206_));
  NOR2X1   g24770(.A(new_n26295_), .B(pi0219), .Y(new_n27207_));
  AOI21X1  g24771(.A0(new_n27207_), .A1(new_n27206_), .B0(new_n26290_), .Y(new_n27208_));
  INVX1    g24772(.A(new_n27208_), .Y(new_n27209_));
  AOI21X1  g24773(.A0(new_n26114_), .A1(pi1146), .B0(new_n27196_), .Y(new_n27210_));
  AOI21X1  g24774(.A0(new_n27210_), .A1(new_n27209_), .B0(new_n26471_), .Y(new_n27211_));
  AOI21X1  g24775(.A0(new_n27211_), .A1(new_n27205_), .B0(new_n26273_), .Y(new_n27212_));
  AOI21X1  g24776(.A0(new_n27212_), .A1(new_n27204_), .B0(new_n26147_), .Y(new_n27213_));
  AOI22X1  g24777(.A0(new_n27213_), .A1(new_n27195_), .B0(new_n27170_), .B1(new_n26147_), .Y(new_n27214_));
  OAI21X1  g24778(.A0(new_n27214_), .A1(pi0213), .B0(pi0209), .Y(new_n27215_));
  OAI21X1  g24779(.A0(new_n27001_), .A1(pi0214), .B0(new_n24961_), .Y(new_n27216_));
  NAND2X1  g24780(.A(new_n27001_), .B(new_n26199_), .Y(new_n27217_));
  AOI21X1  g24781(.A0(new_n27217_), .A1(pi0214), .B0(new_n27216_), .Y(new_n27218_));
  OAI21X1  g24782(.A0(new_n27005_), .A1(new_n24984_), .B0(pi0212), .Y(new_n27219_));
  AOI21X1  g24783(.A0(new_n27217_), .A1(new_n24984_), .B0(new_n27219_), .Y(new_n27220_));
  OAI21X1  g24784(.A0(new_n27220_), .A1(new_n27218_), .B0(new_n23539_), .Y(new_n27221_));
  AOI21X1  g24785(.A0(new_n27001_), .A1(pi0219), .B0(new_n27081_), .Y(new_n27222_));
  INVX1    g24786(.A(new_n27053_), .Y(new_n27223_));
  OAI21X1  g24787(.A0(new_n27056_), .A1(new_n23539_), .B0(new_n27095_), .Y(new_n27224_));
  NOR2X1   g24788(.A(new_n26121_), .B(pi1150), .Y(new_n27225_));
  OAI21X1  g24789(.A0(new_n27224_), .A1(new_n27223_), .B0(new_n27225_), .Y(new_n27226_));
  AOI21X1  g24790(.A0(new_n27222_), .A1(new_n27221_), .B0(new_n27226_), .Y(new_n27227_));
  AND2X1   g24791(.A(new_n27001_), .B(pi0219), .Y(new_n27228_));
  NOR2X1   g24792(.A(new_n27004_), .B(pi0214), .Y(new_n27229_));
  OAI22X1  g24793(.A0(new_n27229_), .A1(new_n27219_), .B0(new_n27216_), .B1(new_n27072_), .Y(new_n27230_));
  AOI21X1  g24794(.A0(new_n27230_), .A1(new_n23539_), .B0(new_n27228_), .Y(new_n27231_));
  OAI21X1  g24795(.A0(new_n27047_), .A1(pi0214), .B0(new_n27051_), .Y(new_n27232_));
  OAI21X1  g24796(.A0(new_n27048_), .A1(new_n27043_), .B0(new_n27232_), .Y(new_n27233_));
  MX2X1    g24797(.A(new_n27233_), .B(new_n27038_), .S0(pi0219), .Y(new_n27234_));
  AOI21X1  g24798(.A0(new_n27234_), .A1(pi1147), .B0(po1038), .Y(new_n27235_));
  OAI21X1  g24799(.A0(new_n27231_), .A1(pi1147), .B0(new_n27235_), .Y(new_n27236_));
  NOR2X1   g24800(.A(new_n25955_), .B(new_n26471_), .Y(new_n27237_));
  AOI21X1  g24801(.A0(new_n27237_), .A1(new_n27236_), .B0(new_n27227_), .Y(new_n27238_));
  NAND2X1  g24802(.A(new_n26379_), .B(pi1150), .Y(new_n27239_));
  AOI21X1  g24803(.A0(new_n27003_), .A1(new_n26091_), .B0(new_n11777_), .Y(new_n27240_));
  NAND2X1  g24804(.A(new_n27038_), .B(pi1147), .Y(new_n27241_));
  INVX1    g24805(.A(new_n27001_), .Y(new_n27242_));
  AOI21X1  g24806(.A0(new_n27239_), .A1(new_n27242_), .B0(pi1147), .Y(new_n27243_));
  NOR2X1   g24807(.A(new_n27243_), .B(po1038), .Y(new_n27244_));
  AOI21X1  g24808(.A0(new_n27244_), .A1(new_n27241_), .B0(pi1149), .Y(new_n27245_));
  OAI21X1  g24809(.A0(new_n27240_), .A1(new_n27239_), .B0(new_n27245_), .Y(new_n27246_));
  OAI21X1  g24810(.A0(new_n27238_), .A1(new_n26147_), .B0(new_n27246_), .Y(new_n27247_));
  OAI21X1  g24811(.A0(new_n27105_), .A1(new_n27103_), .B0(new_n26363_), .Y(new_n27248_));
  OR4X1    g24812(.A(new_n27242_), .B(new_n26996_), .C(new_n9544_), .D(new_n24984_), .Y(new_n27249_));
  AOI21X1  g24813(.A0(new_n27249_), .A1(new_n27009_), .B0(new_n27007_), .Y(new_n27250_));
  OR2X1    g24814(.A(new_n27250_), .B(new_n27248_), .Y(new_n27251_));
  INVX1    g24815(.A(new_n27033_), .Y(new_n27252_));
  NOR3X1   g24816(.A(new_n27030_), .B(new_n24955_), .C(pi0211), .Y(new_n27253_));
  OAI21X1  g24817(.A0(new_n27253_), .A1(new_n27252_), .B0(new_n27095_), .Y(new_n27254_));
  NOR2X1   g24818(.A(new_n27049_), .B(new_n27019_), .Y(new_n27255_));
  INVX1    g24819(.A(new_n27255_), .Y(new_n27256_));
  NOR3X1   g24820(.A(new_n27027_), .B(new_n9544_), .C(new_n24984_), .Y(new_n27257_));
  NOR2X1   g24821(.A(new_n27257_), .B(new_n24961_), .Y(new_n27258_));
  OAI21X1  g24822(.A0(new_n27256_), .A1(pi0214), .B0(new_n27258_), .Y(new_n27259_));
  AOI21X1  g24823(.A0(new_n27256_), .A1(new_n27021_), .B0(pi0219), .Y(new_n27260_));
  AOI21X1  g24824(.A0(new_n27260_), .A1(new_n27259_), .B0(new_n27254_), .Y(new_n27261_));
  NOR3X1   g24825(.A(new_n27261_), .B(new_n26159_), .C(new_n26471_), .Y(new_n27262_));
  NAND2X1  g24826(.A(new_n27258_), .B(new_n27020_), .Y(new_n27263_));
  AOI21X1  g24827(.A0(new_n27019_), .A1(new_n24961_), .B0(pi0219), .Y(new_n27264_));
  AOI21X1  g24828(.A0(new_n27264_), .A1(new_n27263_), .B0(new_n27254_), .Y(new_n27265_));
  NOR3X1   g24829(.A(new_n26996_), .B(new_n26542_), .C(pi0219), .Y(new_n27266_));
  NOR2X1   g24830(.A(new_n25970_), .B(pi1150), .Y(new_n27267_));
  OAI21X1  g24831(.A0(new_n27266_), .A1(new_n27248_), .B0(new_n27267_), .Y(new_n27268_));
  OAI21X1  g24832(.A0(new_n27268_), .A1(new_n27265_), .B0(new_n26147_), .Y(new_n27269_));
  AOI21X1  g24833(.A0(new_n27262_), .A1(new_n27251_), .B0(new_n27269_), .Y(new_n27270_));
  NOR2X1   g24834(.A(new_n27030_), .B(new_n24961_), .Y(new_n27271_));
  OAI22X1  g24835(.A0(new_n27253_), .A1(new_n27252_), .B0(new_n27271_), .B1(new_n27029_), .Y(new_n27272_));
  NOR2X1   g24836(.A(new_n25235_), .B(new_n5117_), .Y(new_n27273_));
  NOR3X1   g24837(.A(new_n27273_), .B(new_n26091_), .C(pi0057), .Y(new_n27274_));
  OAI21X1  g24838(.A0(new_n27272_), .A1(new_n5118_), .B0(new_n27274_), .Y(new_n27275_));
  NAND4X1  g24839(.A(new_n26996_), .B(new_n25848_), .C(new_n24994_), .D(new_n5117_), .Y(new_n27276_));
  AOI21X1  g24840(.A0(new_n26995_), .A1(new_n2953_), .B0(new_n25235_), .Y(new_n27277_));
  NOR4X1   g24841(.A(new_n27277_), .B(new_n27273_), .C(pi1147), .D(pi0057), .Y(new_n27278_));
  AOI22X1  g24842(.A0(new_n27278_), .A1(new_n27276_), .B0(new_n25235_), .B1(pi0057), .Y(new_n27279_));
  AOI21X1  g24843(.A0(new_n27279_), .A1(new_n27275_), .B0(new_n26471_), .Y(new_n27280_));
  OR2X1    g24844(.A(new_n27217_), .B(new_n26996_), .Y(new_n27281_));
  OAI21X1  g24845(.A0(new_n27281_), .A1(new_n27072_), .B0(pi0212), .Y(new_n27282_));
  AOI21X1  g24846(.A0(new_n27249_), .A1(new_n26998_), .B0(pi0219), .Y(new_n27283_));
  AOI21X1  g24847(.A0(new_n27283_), .A1(new_n27282_), .B0(new_n27248_), .Y(new_n27284_));
  OR4X1    g24848(.A(new_n26554_), .B(new_n5118_), .C(new_n26091_), .D(pi0057), .Y(new_n27285_));
  NOR2X1   g24849(.A(new_n26152_), .B(pi1150), .Y(new_n27286_));
  OAI21X1  g24850(.A0(new_n27285_), .A1(new_n27272_), .B0(new_n27286_), .Y(new_n27287_));
  OAI21X1  g24851(.A0(new_n27287_), .A1(new_n27284_), .B0(pi1149), .Y(new_n27288_));
  OAI21X1  g24852(.A0(new_n27288_), .A1(new_n27280_), .B0(pi1148), .Y(new_n27289_));
  OAI21X1  g24853(.A0(new_n27289_), .A1(new_n27270_), .B0(pi0213), .Y(new_n27290_));
  AOI21X1  g24854(.A0(new_n27247_), .A1(new_n26273_), .B0(new_n27290_), .Y(new_n27291_));
  OAI21X1  g24855(.A0(new_n27070_), .A1(pi0213), .B0(new_n23244_), .Y(new_n27292_));
  OAI22X1  g24856(.A0(new_n27292_), .A1(new_n27291_), .B0(new_n27215_), .B1(new_n27132_), .Y(new_n27293_));
  NOR2X1   g24857(.A(pi0246), .B(pi0230), .Y(new_n27294_));
  AOI21X1  g24858(.A0(new_n27293_), .A1(pi0230), .B0(new_n27294_), .Y(po0403));
  NAND2X1  g24859(.A(new_n26502_), .B(new_n26091_), .Y(new_n27296_));
  OR2X1    g24860(.A(new_n26093_), .B(new_n25996_), .Y(new_n27297_));
  NOR2X1   g24861(.A(new_n26121_), .B(new_n25837_), .Y(new_n27298_));
  INVX1    g24862(.A(new_n27298_), .Y(new_n27299_));
  AOI21X1  g24863(.A0(new_n27184_), .A1(new_n27297_), .B0(new_n27299_), .Y(new_n27300_));
  NOR2X1   g24864(.A(new_n26152_), .B(new_n25837_), .Y(new_n27301_));
  INVX1    g24865(.A(new_n27301_), .Y(new_n27302_));
  AOI21X1  g24866(.A0(new_n27183_), .A1(new_n27182_), .B0(new_n26572_), .Y(new_n27303_));
  OR2X1    g24867(.A(new_n26140_), .B(new_n26127_), .Y(new_n27304_));
  AOI21X1  g24868(.A0(new_n27304_), .A1(new_n27173_), .B0(new_n26152_), .Y(new_n27305_));
  AOI21X1  g24869(.A0(new_n27305_), .A1(new_n25837_), .B0(new_n26091_), .Y(new_n27306_));
  OAI21X1  g24870(.A0(new_n27303_), .A1(new_n27302_), .B0(new_n27306_), .Y(new_n27307_));
  AND2X1   g24871(.A(new_n27307_), .B(new_n26147_), .Y(new_n27308_));
  OAI21X1  g24872(.A0(new_n27300_), .A1(new_n27296_), .B0(new_n27308_), .Y(new_n27309_));
  OAI21X1  g24873(.A0(new_n27199_), .A1(new_n26205_), .B0(new_n26558_), .Y(new_n27310_));
  INVX1    g24874(.A(new_n27310_), .Y(new_n27311_));
  AND2X1   g24875(.A(new_n26558_), .B(new_n26191_), .Y(new_n27312_));
  NOR4X1   g24876(.A(new_n27312_), .B(new_n27311_), .C(new_n25955_), .D(pi1151), .Y(new_n27313_));
  OAI21X1  g24877(.A0(new_n27208_), .A1(new_n26503_), .B0(new_n26091_), .Y(new_n27314_));
  NOR2X1   g24878(.A(new_n26513_), .B(new_n26091_), .Y(new_n27315_));
  OR4X1    g24879(.A(new_n26151_), .B(new_n26114_), .C(new_n26111_), .D(pi1151), .Y(new_n27316_));
  AOI21X1  g24880(.A0(new_n27316_), .A1(new_n27315_), .B0(new_n26147_), .Y(new_n27317_));
  OAI21X1  g24881(.A0(new_n27314_), .A1(new_n27313_), .B0(new_n27317_), .Y(new_n27318_));
  NAND3X1  g24882(.A(new_n27318_), .B(new_n27309_), .C(pi1150), .Y(new_n27319_));
  NOR2X1   g24883(.A(new_n25815_), .B(new_n24961_), .Y(new_n27320_));
  OAI21X1  g24884(.A0(new_n27320_), .A1(new_n27150_), .B0(new_n26174_), .Y(new_n27321_));
  AND2X1   g24885(.A(new_n27321_), .B(new_n26484_), .Y(new_n27322_));
  NOR2X1   g24886(.A(new_n26187_), .B(new_n24963_), .Y(new_n27323_));
  NOR4X1   g24887(.A(new_n27323_), .B(new_n26534_), .C(new_n26195_), .D(po1038), .Y(new_n27324_));
  NOR4X1   g24888(.A(new_n27324_), .B(new_n26211_), .C(new_n26111_), .D(pi1151), .Y(new_n27325_));
  NOR3X1   g24889(.A(new_n27325_), .B(new_n27322_), .C(new_n26091_), .Y(new_n27326_));
  INVX1    g24890(.A(new_n26259_), .Y(new_n27327_));
  AOI21X1  g24891(.A0(new_n26436_), .A1(new_n26435_), .B0(new_n27150_), .Y(new_n27328_));
  OAI21X1  g24892(.A0(new_n27328_), .A1(new_n27327_), .B0(new_n25969_), .Y(new_n27329_));
  NOR2X1   g24893(.A(new_n27329_), .B(new_n25837_), .Y(new_n27330_));
  NOR3X1   g24894(.A(new_n27324_), .B(new_n25955_), .C(pi1151), .Y(new_n27331_));
  OR2X1    g24895(.A(new_n27331_), .B(pi1147), .Y(new_n27332_));
  OAI21X1  g24896(.A0(new_n27332_), .A1(new_n27330_), .B0(pi1149), .Y(new_n27333_));
  INVX1    g24897(.A(new_n26180_), .Y(new_n27334_));
  OR2X1    g24898(.A(new_n27334_), .B(new_n26120_), .Y(new_n27335_));
  AOI21X1  g24899(.A0(new_n27335_), .A1(new_n25837_), .B0(pi1147), .Y(new_n27336_));
  AND2X1   g24900(.A(new_n26451_), .B(new_n25996_), .Y(new_n27337_));
  OAI21X1  g24901(.A0(new_n27337_), .A1(new_n27299_), .B0(new_n27336_), .Y(new_n27338_));
  NOR2X1   g24902(.A(new_n27302_), .B(new_n26601_), .Y(new_n27339_));
  NOR3X1   g24903(.A(new_n26152_), .B(new_n26150_), .C(pi1151), .Y(new_n27340_));
  NOR3X1   g24904(.A(new_n27340_), .B(new_n27339_), .C(new_n26091_), .Y(new_n27341_));
  NOR2X1   g24905(.A(new_n27341_), .B(pi1149), .Y(new_n27342_));
  AOI21X1  g24906(.A0(new_n27342_), .A1(new_n27338_), .B0(pi1150), .Y(new_n27343_));
  OAI21X1  g24907(.A0(new_n27333_), .A1(new_n27326_), .B0(new_n27343_), .Y(new_n27344_));
  AOI21X1  g24908(.A0(new_n27344_), .A1(new_n27319_), .B0(new_n26273_), .Y(new_n27345_));
  NOR2X1   g24909(.A(new_n26465_), .B(new_n26176_), .Y(new_n27346_));
  NOR2X1   g24910(.A(new_n26159_), .B(pi1151), .Y(new_n27347_));
  INVX1    g24911(.A(new_n27347_), .Y(new_n27348_));
  NOR2X1   g24912(.A(new_n27348_), .B(new_n26211_), .Y(new_n27349_));
  NOR3X1   g24913(.A(new_n27349_), .B(new_n27346_), .C(new_n26091_), .Y(new_n27350_));
  AOI21X1  g24914(.A0(new_n26259_), .A1(new_n26169_), .B0(new_n26225_), .Y(new_n27351_));
  NOR2X1   g24915(.A(new_n26225_), .B(pi1151), .Y(new_n27352_));
  AND2X1   g24916(.A(new_n27352_), .B(new_n26525_), .Y(new_n27353_));
  OR2X1    g24917(.A(new_n27353_), .B(pi1147), .Y(new_n27354_));
  AOI21X1  g24918(.A0(new_n27351_), .A1(pi1151), .B0(new_n27354_), .Y(new_n27355_));
  NOR3X1   g24919(.A(new_n27355_), .B(new_n27350_), .C(pi1150), .Y(new_n27356_));
  NOR3X1   g24920(.A(new_n26545_), .B(new_n26465_), .C(new_n26302_), .Y(new_n27357_));
  NOR2X1   g24921(.A(new_n26210_), .B(new_n26206_), .Y(new_n27358_));
  NOR3X1   g24922(.A(new_n27358_), .B(new_n26159_), .C(pi1151), .Y(new_n27359_));
  NOR3X1   g24923(.A(new_n27359_), .B(new_n27357_), .C(new_n26091_), .Y(new_n27360_));
  NOR3X1   g24924(.A(new_n26302_), .B(new_n26225_), .C(new_n25837_), .Y(new_n27361_));
  OR2X1    g24925(.A(new_n27361_), .B(pi1147), .Y(new_n27362_));
  AOI21X1  g24926(.A0(new_n27352_), .A1(new_n27310_), .B0(new_n27362_), .Y(new_n27363_));
  NOR3X1   g24927(.A(new_n27363_), .B(new_n27360_), .C(new_n26471_), .Y(new_n27364_));
  OAI21X1  g24928(.A0(new_n27364_), .A1(new_n27356_), .B0(pi1149), .Y(new_n27365_));
  OR2X1    g24929(.A(new_n25970_), .B(new_n25837_), .Y(new_n27366_));
  OR2X1    g24930(.A(new_n27190_), .B(new_n26591_), .Y(new_n27367_));
  AOI21X1  g24931(.A0(new_n27303_), .A1(new_n27367_), .B0(new_n27366_), .Y(new_n27368_));
  NOR3X1   g24932(.A(new_n27177_), .B(new_n25970_), .C(pi1151), .Y(new_n27369_));
  NOR3X1   g24933(.A(new_n27369_), .B(new_n27368_), .C(new_n26091_), .Y(new_n27370_));
  OAI21X1  g24934(.A0(new_n26241_), .A1(pi1151), .B0(new_n26091_), .Y(new_n27371_));
  NOR2X1   g24935(.A(new_n26093_), .B(new_n25837_), .Y(new_n27372_));
  OAI21X1  g24936(.A0(new_n27372_), .A1(new_n27371_), .B0(pi1150), .Y(new_n27373_));
  AOI21X1  g24937(.A0(new_n26543_), .A1(new_n25995_), .B0(new_n26600_), .Y(new_n27374_));
  NOR2X1   g24938(.A(new_n27374_), .B(new_n27366_), .Y(new_n27375_));
  AOI21X1  g24939(.A0(new_n26544_), .A1(new_n26209_), .B0(new_n26509_), .Y(new_n27376_));
  NOR3X1   g24940(.A(new_n27376_), .B(new_n27375_), .C(new_n26091_), .Y(new_n27377_));
  AND2X1   g24941(.A(pi1151), .B(new_n26091_), .Y(new_n27378_));
  NAND4X1  g24942(.A(new_n27378_), .B(new_n25259_), .C(new_n11776_), .D(new_n8130_), .Y(new_n27379_));
  NAND2X1  g24943(.A(new_n27379_), .B(new_n26471_), .Y(new_n27380_));
  OAI22X1  g24944(.A0(new_n27380_), .A1(new_n27377_), .B0(new_n27373_), .B1(new_n27370_), .Y(new_n27381_));
  AOI21X1  g24945(.A0(new_n27381_), .A1(new_n26147_), .B0(pi1148), .Y(new_n27382_));
  AND2X1   g24946(.A(new_n27382_), .B(new_n27365_), .Y(new_n27383_));
  OAI21X1  g24947(.A0(new_n27383_), .A1(new_n27345_), .B0(new_n25003_), .Y(new_n27384_));
  AOI21X1  g24948(.A0(new_n26517_), .A1(pi0213), .B0(new_n23244_), .Y(new_n27385_));
  NOR2X1   g24949(.A(new_n26225_), .B(new_n25837_), .Y(new_n27386_));
  NAND2X1  g24950(.A(new_n26550_), .B(pi1147), .Y(new_n27387_));
  AOI21X1  g24951(.A0(new_n27386_), .A1(new_n27310_), .B0(new_n27387_), .Y(new_n27388_));
  AOI21X1  g24952(.A0(new_n26124_), .A1(new_n26582_), .B0(po1038), .Y(new_n27389_));
  OAI21X1  g24953(.A0(new_n26133_), .A1(new_n26582_), .B0(new_n27389_), .Y(new_n27390_));
  AND2X1   g24954(.A(new_n27390_), .B(new_n26416_), .Y(new_n27391_));
  INVX1    g24955(.A(new_n27391_), .Y(new_n27392_));
  OAI21X1  g24956(.A0(new_n27392_), .A1(new_n27371_), .B0(new_n26471_), .Y(new_n27393_));
  OR2X1    g24957(.A(new_n27393_), .B(new_n27388_), .Y(new_n27394_));
  AOI21X1  g24958(.A0(new_n26143_), .A1(new_n26138_), .B0(new_n26503_), .Y(new_n27395_));
  NOR3X1   g24959(.A(new_n27312_), .B(new_n27311_), .C(new_n26503_), .Y(new_n27396_));
  AOI21X1  g24960(.A0(new_n26558_), .A1(new_n26191_), .B0(new_n26444_), .Y(new_n27397_));
  NOR3X1   g24961(.A(new_n27397_), .B(new_n27396_), .C(new_n26091_), .Y(new_n27398_));
  NOR2X1   g24962(.A(new_n27398_), .B(new_n26471_), .Y(new_n27399_));
  OAI21X1  g24963(.A0(new_n27395_), .A1(new_n27296_), .B0(new_n27399_), .Y(new_n27400_));
  AOI21X1  g24964(.A0(new_n27400_), .A1(new_n27394_), .B0(pi1149), .Y(new_n27401_));
  AOI21X1  g24965(.A0(new_n27303_), .A1(new_n27367_), .B0(new_n26509_), .Y(new_n27402_));
  OAI21X1  g24966(.A0(new_n26158_), .A1(new_n25929_), .B0(new_n27191_), .Y(new_n27403_));
  OAI21X1  g24967(.A0(new_n27403_), .A1(new_n25837_), .B0(new_n26091_), .Y(new_n27404_));
  OR4X1    g24968(.A(new_n26545_), .B(new_n26302_), .C(new_n26159_), .D(new_n25837_), .Y(new_n27405_));
  OAI21X1  g24969(.A0(new_n26288_), .A1(po1038), .B0(new_n27376_), .Y(new_n27406_));
  NAND3X1  g24970(.A(new_n27406_), .B(new_n27405_), .C(pi1147), .Y(new_n27407_));
  AND2X1   g24971(.A(new_n27407_), .B(new_n26471_), .Y(new_n27408_));
  OAI21X1  g24972(.A0(new_n27404_), .A1(new_n27402_), .B0(new_n27408_), .Y(new_n27409_));
  INVX1    g24973(.A(new_n26490_), .Y(new_n27410_));
  NAND2X1  g24974(.A(new_n26284_), .B(new_n26100_), .Y(new_n27411_));
  AOI21X1  g24975(.A0(new_n27411_), .A1(new_n26279_), .B0(new_n26485_), .Y(new_n27412_));
  NOR2X1   g24976(.A(new_n27412_), .B(pi1147), .Y(new_n27413_));
  OAI21X1  g24977(.A0(new_n27303_), .A1(new_n27410_), .B0(new_n27413_), .Y(new_n27414_));
  OAI21X1  g24978(.A0(new_n26554_), .A1(new_n26553_), .B0(new_n26967_), .Y(new_n27415_));
  OAI21X1  g24979(.A0(new_n27415_), .A1(pi1151), .B0(new_n27315_), .Y(new_n27416_));
  NAND3X1  g24980(.A(new_n27416_), .B(new_n27414_), .C(pi1150), .Y(new_n27417_));
  AOI21X1  g24981(.A0(new_n27417_), .A1(new_n27409_), .B0(new_n26147_), .Y(new_n27418_));
  NOR3X1   g24982(.A(new_n27418_), .B(new_n27401_), .C(new_n26273_), .Y(new_n27419_));
  NOR2X1   g24983(.A(new_n27346_), .B(new_n26091_), .Y(new_n27420_));
  NAND3X1  g24984(.A(new_n26529_), .B(new_n26450_), .C(new_n23539_), .Y(new_n27421_));
  NAND2X1  g24985(.A(new_n27421_), .B(new_n26174_), .Y(new_n27422_));
  OAI21X1  g24986(.A0(new_n27422_), .A1(new_n26170_), .B0(new_n26478_), .Y(new_n27423_));
  AND2X1   g24987(.A(new_n27423_), .B(new_n27420_), .Y(new_n27424_));
  NOR3X1   g24988(.A(new_n26092_), .B(new_n25842_), .C(new_n8074_), .Y(new_n27425_));
  NOR3X1   g24989(.A(new_n27425_), .B(new_n27374_), .C(new_n26465_), .Y(new_n27426_));
  OAI21X1  g24990(.A0(new_n27374_), .A1(new_n26509_), .B0(new_n26091_), .Y(new_n27427_));
  OAI21X1  g24991(.A0(new_n27427_), .A1(new_n27426_), .B0(new_n26471_), .Y(new_n27428_));
  OR2X1    g24992(.A(new_n27322_), .B(new_n26091_), .Y(new_n27429_));
  AOI21X1  g24993(.A0(new_n27421_), .A1(new_n26174_), .B0(new_n26152_), .Y(new_n27430_));
  AOI21X1  g24994(.A0(new_n27430_), .A1(new_n25837_), .B0(new_n27429_), .Y(new_n27431_));
  OAI21X1  g24995(.A0(new_n26092_), .A1(new_n25842_), .B0(new_n26484_), .Y(new_n27432_));
  NOR2X1   g24996(.A(new_n27432_), .B(new_n26601_), .Y(new_n27433_));
  OAI21X1  g24997(.A0(new_n26601_), .A1(new_n27410_), .B0(new_n26091_), .Y(new_n27434_));
  OAI21X1  g24998(.A0(new_n27434_), .A1(new_n27433_), .B0(pi1150), .Y(new_n27435_));
  OAI22X1  g24999(.A0(new_n27435_), .A1(new_n27431_), .B0(new_n27428_), .B1(new_n27424_), .Y(new_n27436_));
  INVX1    g25000(.A(new_n26121_), .Y(new_n27437_));
  OAI21X1  g25001(.A0(new_n26536_), .A1(new_n26197_), .B0(new_n27437_), .Y(new_n27438_));
  OR2X1    g25002(.A(new_n27324_), .B(new_n26503_), .Y(new_n27439_));
  AND2X1   g25003(.A(new_n27439_), .B(pi1147), .Y(new_n27440_));
  OAI21X1  g25004(.A0(new_n27438_), .A1(pi1151), .B0(new_n27440_), .Y(new_n27441_));
  AOI21X1  g25005(.A0(new_n26603_), .A1(new_n11777_), .B0(new_n25837_), .Y(new_n27442_));
  INVX1    g25006(.A(new_n27442_), .Y(new_n27443_));
  AOI21X1  g25007(.A0(new_n27443_), .A1(new_n27336_), .B0(new_n26471_), .Y(new_n27444_));
  OAI21X1  g25008(.A0(new_n26381_), .A1(new_n6520_), .B0(new_n26525_), .Y(new_n27445_));
  OAI21X1  g25009(.A0(new_n27134_), .A1(new_n27133_), .B0(new_n25837_), .Y(new_n27446_));
  NAND3X1  g25010(.A(new_n27446_), .B(new_n27445_), .C(pi1147), .Y(new_n27447_));
  AOI21X1  g25011(.A0(new_n27378_), .A1(new_n26181_), .B0(pi1150), .Y(new_n27448_));
  AOI22X1  g25012(.A0(new_n27448_), .A1(new_n27447_), .B0(new_n27444_), .B1(new_n27441_), .Y(new_n27449_));
  OAI21X1  g25013(.A0(new_n27449_), .A1(pi1149), .B0(new_n26273_), .Y(new_n27450_));
  AOI21X1  g25014(.A0(new_n27436_), .A1(pi1149), .B0(new_n27450_), .Y(new_n27451_));
  OAI21X1  g25015(.A0(new_n27451_), .A1(new_n27419_), .B0(pi0213), .Y(new_n27452_));
  AOI21X1  g25016(.A0(new_n26215_), .A1(new_n25003_), .B0(pi0209), .Y(new_n27453_));
  AOI22X1  g25017(.A0(new_n27453_), .A1(new_n27452_), .B0(new_n27385_), .B1(new_n27384_), .Y(new_n27454_));
  MX2X1    g25018(.A(new_n27454_), .B(pi0247), .S0(new_n24954_), .Y(po0404));
  NOR2X1   g25019(.A(new_n27303_), .B(new_n27302_), .Y(new_n27456_));
  OAI21X1  g25020(.A0(new_n26601_), .A1(new_n27410_), .B0(pi1152), .Y(new_n27457_));
  NOR2X1   g25021(.A(new_n27457_), .B(new_n27456_), .Y(new_n27458_));
  OR2X1    g25022(.A(new_n27340_), .B(pi1152), .Y(new_n27459_));
  AOI21X1  g25023(.A0(new_n27305_), .A1(pi1151), .B0(new_n27459_), .Y(new_n27460_));
  NOR3X1   g25024(.A(new_n27460_), .B(new_n27458_), .C(pi1150), .Y(new_n27461_));
  AOI21X1  g25025(.A0(new_n26110_), .A1(new_n25323_), .B0(pi1151), .Y(new_n27462_));
  NOR2X1   g25026(.A(new_n26513_), .B(new_n25289_), .Y(new_n27463_));
  INVX1    g25027(.A(new_n27463_), .Y(new_n27464_));
  AOI21X1  g25028(.A0(new_n27462_), .A1(new_n27321_), .B0(new_n27464_), .Y(new_n27465_));
  OR4X1    g25029(.A(new_n26151_), .B(new_n26114_), .C(new_n26111_), .D(new_n25837_), .Y(new_n27466_));
  NAND2X1  g25030(.A(new_n27466_), .B(new_n25289_), .Y(new_n27467_));
  OAI21X1  g25031(.A0(new_n27467_), .A1(new_n27325_), .B0(pi1150), .Y(new_n27468_));
  OAI21X1  g25032(.A0(new_n27468_), .A1(new_n27465_), .B0(pi1148), .Y(new_n27469_));
  OAI21X1  g25033(.A0(new_n27299_), .A1(new_n26145_), .B0(new_n25289_), .Y(new_n27470_));
  AOI21X1  g25034(.A0(new_n27335_), .A1(new_n25837_), .B0(new_n27470_), .Y(new_n27471_));
  OAI21X1  g25035(.A0(new_n27337_), .A1(new_n26444_), .B0(pi1152), .Y(new_n27472_));
  OAI21X1  g25036(.A0(new_n27472_), .A1(new_n27300_), .B0(new_n26471_), .Y(new_n27473_));
  NOR2X1   g25037(.A(new_n27473_), .B(new_n27471_), .Y(new_n27474_));
  NOR2X1   g25038(.A(new_n27329_), .B(pi1151), .Y(new_n27475_));
  OAI21X1  g25039(.A0(new_n27208_), .A1(new_n26503_), .B0(pi1152), .Y(new_n27476_));
  NOR2X1   g25040(.A(new_n27476_), .B(new_n27475_), .Y(new_n27477_));
  OR2X1    g25041(.A(new_n27331_), .B(pi1152), .Y(new_n27478_));
  OAI21X1  g25042(.A0(new_n27478_), .A1(new_n27396_), .B0(pi1150), .Y(new_n27479_));
  OAI21X1  g25043(.A0(new_n27479_), .A1(new_n27477_), .B0(new_n26273_), .Y(new_n27480_));
  OAI22X1  g25044(.A0(new_n27480_), .A1(new_n27474_), .B0(new_n27469_), .B1(new_n27461_), .Y(new_n27481_));
  NAND2X1  g25045(.A(new_n27481_), .B(pi1149), .Y(new_n27482_));
  INVX1    g25046(.A(new_n26176_), .Y(new_n27483_));
  AOI21X1  g25047(.A0(new_n27347_), .A1(new_n27483_), .B0(new_n25289_), .Y(new_n27484_));
  NOR3X1   g25048(.A(new_n27358_), .B(new_n26159_), .C(new_n25837_), .Y(new_n27485_));
  NOR3X1   g25049(.A(new_n27485_), .B(new_n27349_), .C(pi1152), .Y(new_n27486_));
  AOI21X1  g25050(.A0(new_n27484_), .A1(new_n27405_), .B0(new_n27486_), .Y(new_n27487_));
  NOR2X1   g25051(.A(new_n27374_), .B(new_n26509_), .Y(new_n27488_));
  OAI21X1  g25052(.A0(new_n27488_), .A1(new_n27368_), .B0(pi1152), .Y(new_n27489_));
  NOR3X1   g25053(.A(new_n27177_), .B(new_n25970_), .C(new_n25837_), .Y(new_n27490_));
  OAI21X1  g25054(.A0(new_n27490_), .A1(new_n27376_), .B0(new_n25289_), .Y(new_n27491_));
  AND2X1   g25055(.A(new_n27491_), .B(new_n26471_), .Y(new_n27492_));
  AOI21X1  g25056(.A0(new_n27492_), .A1(new_n27489_), .B0(new_n26273_), .Y(new_n27493_));
  OAI21X1  g25057(.A0(new_n27487_), .A1(new_n26471_), .B0(new_n27493_), .Y(new_n27494_));
  OR2X1    g25058(.A(new_n27361_), .B(new_n25289_), .Y(new_n27495_));
  AOI21X1  g25059(.A0(new_n27351_), .A1(new_n25837_), .B0(new_n27495_), .Y(new_n27496_));
  OR2X1    g25060(.A(new_n27353_), .B(pi1152), .Y(new_n27497_));
  AOI21X1  g25061(.A0(new_n27386_), .A1(new_n27310_), .B0(new_n27497_), .Y(new_n27498_));
  NOR3X1   g25062(.A(new_n27498_), .B(new_n27496_), .C(new_n26471_), .Y(new_n27499_));
  AND2X1   g25063(.A(new_n25289_), .B(pi1151), .Y(new_n27500_));
  NOR2X1   g25064(.A(new_n26179_), .B(pi1151), .Y(new_n27501_));
  OAI21X1  g25065(.A0(new_n26093_), .A1(new_n25837_), .B0(pi1152), .Y(new_n27502_));
  OAI21X1  g25066(.A0(new_n27502_), .A1(new_n27501_), .B0(new_n26471_), .Y(new_n27503_));
  AOI21X1  g25067(.A0(new_n27500_), .A1(new_n26241_), .B0(new_n27503_), .Y(new_n27504_));
  OAI21X1  g25068(.A0(new_n27504_), .A1(new_n27499_), .B0(new_n26273_), .Y(new_n27505_));
  NAND3X1  g25069(.A(new_n27505_), .B(new_n27494_), .C(new_n26147_), .Y(new_n27506_));
  AOI21X1  g25070(.A0(new_n27506_), .A1(new_n27482_), .B0(pi0213), .Y(new_n27507_));
  OAI21X1  g25071(.A0(new_n26145_), .A1(new_n26121_), .B0(new_n27500_), .Y(new_n27508_));
  AOI21X1  g25072(.A0(new_n26180_), .A1(new_n26157_), .B0(pi1151), .Y(new_n27509_));
  AOI21X1  g25073(.A0(new_n27509_), .A1(new_n26274_), .B0(new_n25289_), .Y(new_n27510_));
  OAI21X1  g25074(.A0(new_n26503_), .A1(new_n26107_), .B0(new_n27510_), .Y(new_n27511_));
  AND2X1   g25075(.A(new_n27511_), .B(new_n26471_), .Y(new_n27512_));
  AOI21X1  g25076(.A0(new_n27347_), .A1(new_n27483_), .B0(new_n27464_), .Y(new_n27513_));
  AOI21X1  g25077(.A0(new_n26153_), .A1(pi1151), .B0(pi1152), .Y(new_n27514_));
  INVX1    g25078(.A(new_n27514_), .Y(new_n27515_));
  NOR2X1   g25079(.A(new_n27515_), .B(new_n26510_), .Y(new_n27516_));
  NOR3X1   g25080(.A(new_n27516_), .B(new_n27513_), .C(new_n26471_), .Y(new_n27517_));
  AOI21X1  g25081(.A0(new_n27512_), .A1(new_n27508_), .B0(new_n27517_), .Y(new_n27518_));
  AND2X1   g25082(.A(new_n27518_), .B(pi0213), .Y(new_n27519_));
  OR2X1    g25083(.A(new_n27519_), .B(new_n23244_), .Y(new_n27520_));
  NOR2X1   g25084(.A(new_n26241_), .B(pi1151), .Y(new_n27521_));
  INVX1    g25085(.A(new_n27395_), .Y(new_n27522_));
  AOI21X1  g25086(.A0(new_n27392_), .A1(new_n25837_), .B0(new_n25289_), .Y(new_n27523_));
  AOI21X1  g25087(.A0(new_n27523_), .A1(new_n27522_), .B0(pi1150), .Y(new_n27524_));
  OAI21X1  g25088(.A0(new_n27470_), .A1(new_n27521_), .B0(new_n27524_), .Y(new_n27525_));
  OAI21X1  g25089(.A0(new_n27303_), .A1(new_n27302_), .B0(new_n25289_), .Y(new_n27526_));
  OR2X1    g25090(.A(new_n27526_), .B(new_n27402_), .Y(new_n27527_));
  NOR2X1   g25091(.A(new_n27412_), .B(new_n25289_), .Y(new_n27528_));
  OAI21X1  g25092(.A0(new_n27403_), .A1(pi1151), .B0(new_n27528_), .Y(new_n27529_));
  AND2X1   g25093(.A(new_n27529_), .B(pi1150), .Y(new_n27530_));
  AOI21X1  g25094(.A0(new_n27530_), .A1(new_n27527_), .B0(new_n26147_), .Y(new_n27531_));
  NOR3X1   g25095(.A(new_n27425_), .B(new_n27374_), .C(new_n27348_), .Y(new_n27532_));
  NOR3X1   g25096(.A(new_n27532_), .B(new_n27433_), .C(new_n25289_), .Y(new_n27533_));
  NOR3X1   g25097(.A(new_n27488_), .B(new_n27339_), .C(pi1152), .Y(new_n27534_));
  NOR3X1   g25098(.A(new_n27534_), .B(new_n27533_), .C(new_n26471_), .Y(new_n27535_));
  NOR3X1   g25099(.A(new_n27509_), .B(new_n27442_), .C(new_n25289_), .Y(new_n27536_));
  INVX1    g25100(.A(new_n27500_), .Y(new_n27537_));
  OAI21X1  g25101(.A0(new_n27537_), .A1(new_n27335_), .B0(new_n26471_), .Y(new_n27538_));
  OAI21X1  g25102(.A0(new_n27538_), .A1(new_n27536_), .B0(new_n26147_), .Y(new_n27539_));
  OAI21X1  g25103(.A0(new_n27539_), .A1(new_n27535_), .B0(new_n26273_), .Y(new_n27540_));
  AOI21X1  g25104(.A0(new_n27531_), .A1(new_n27525_), .B0(new_n27540_), .Y(new_n27541_));
  INVX1    g25105(.A(new_n27322_), .Y(new_n27542_));
  NAND2X1  g25106(.A(new_n27484_), .B(new_n27542_), .Y(new_n27543_));
  NAND2X1  g25107(.A(new_n27430_), .B(pi1151), .Y(new_n27544_));
  NAND3X1  g25108(.A(new_n27544_), .B(new_n27423_), .C(new_n25289_), .Y(new_n27545_));
  NAND3X1  g25109(.A(new_n27545_), .B(new_n27543_), .C(pi1150), .Y(new_n27546_));
  AND2X1   g25110(.A(new_n27446_), .B(new_n25289_), .Y(new_n27547_));
  OAI21X1  g25111(.A0(new_n27438_), .A1(new_n25837_), .B0(new_n27547_), .Y(new_n27548_));
  AOI21X1  g25112(.A0(new_n27352_), .A1(new_n26525_), .B0(new_n25289_), .Y(new_n27549_));
  AOI21X1  g25113(.A0(new_n27549_), .A1(new_n27439_), .B0(pi1150), .Y(new_n27550_));
  AOI21X1  g25114(.A0(new_n27550_), .A1(new_n27548_), .B0(pi1149), .Y(new_n27551_));
  INVX1    g25115(.A(new_n27396_), .Y(new_n27552_));
  AOI21X1  g25116(.A0(new_n27352_), .A1(new_n27310_), .B0(new_n25289_), .Y(new_n27553_));
  INVX1    g25117(.A(new_n26551_), .Y(new_n27554_));
  AOI21X1  g25118(.A0(new_n26558_), .A1(new_n26191_), .B0(new_n27299_), .Y(new_n27555_));
  OAI21X1  g25119(.A0(new_n27555_), .A1(new_n27554_), .B0(new_n26471_), .Y(new_n27556_));
  AOI21X1  g25120(.A0(new_n27553_), .A1(new_n27552_), .B0(new_n27556_), .Y(new_n27557_));
  AOI21X1  g25121(.A0(new_n27347_), .A1(new_n26546_), .B0(new_n27464_), .Y(new_n27558_));
  NOR2X1   g25122(.A(new_n27415_), .B(new_n25837_), .Y(new_n27559_));
  NAND2X1  g25123(.A(new_n27406_), .B(new_n25289_), .Y(new_n27560_));
  OAI21X1  g25124(.A0(new_n27560_), .A1(new_n27559_), .B0(pi1150), .Y(new_n27561_));
  OAI21X1  g25125(.A0(new_n27561_), .A1(new_n27558_), .B0(pi1149), .Y(new_n27562_));
  OAI21X1  g25126(.A0(new_n27562_), .A1(new_n27557_), .B0(pi1148), .Y(new_n27563_));
  AOI21X1  g25127(.A0(new_n27551_), .A1(new_n27546_), .B0(new_n27563_), .Y(new_n27564_));
  NOR3X1   g25128(.A(new_n27564_), .B(new_n27541_), .C(new_n25003_), .Y(new_n27565_));
  OAI21X1  g25129(.A0(new_n27131_), .A1(pi0213), .B0(new_n23244_), .Y(new_n27566_));
  OAI22X1  g25130(.A0(new_n27566_), .A1(new_n27565_), .B0(new_n27520_), .B1(new_n27507_), .Y(new_n27567_));
  NOR2X1   g25131(.A(pi0248), .B(pi0230), .Y(new_n27568_));
  AOI21X1  g25132(.A0(new_n27567_), .A1(pi0230), .B0(new_n27568_), .Y(po0405));
  NAND2X1  g25133(.A(new_n27518_), .B(new_n25003_), .Y(new_n27570_));
  AND2X1   g25134(.A(new_n25254_), .B(pi0299), .Y(new_n27571_));
  NOR3X1   g25135(.A(new_n27571_), .B(new_n26195_), .C(new_n25888_), .Y(new_n27572_));
  NOR3X1   g25136(.A(new_n27571_), .B(new_n26195_), .C(pi0214), .Y(new_n27573_));
  NOR2X1   g25137(.A(new_n26194_), .B(new_n25984_), .Y(new_n27574_));
  OR2X1    g25138(.A(new_n26524_), .B(new_n24984_), .Y(new_n27575_));
  OAI21X1  g25139(.A0(new_n27575_), .A1(new_n27574_), .B0(pi0212), .Y(new_n27576_));
  OAI22X1  g25140(.A0(new_n27576_), .A1(new_n27573_), .B0(new_n27572_), .B1(pi0212), .Y(new_n27577_));
  OAI21X1  g25141(.A0(new_n26194_), .A1(new_n23539_), .B0(new_n5117_), .Y(new_n27578_));
  AOI21X1  g25142(.A0(new_n27577_), .A1(new_n23539_), .B0(new_n27578_), .Y(new_n27579_));
  NOR3X1   g25143(.A(new_n25256_), .B(new_n25016_), .C(new_n5117_), .Y(new_n27580_));
  OR4X1    g25144(.A(new_n27580_), .B(new_n27579_), .C(pi1151), .D(pi0057), .Y(new_n27581_));
  NOR2X1   g25145(.A(new_n25257_), .B(new_n2436_), .Y(new_n27582_));
  MX2X1    g25146(.A(new_n25883_), .B(new_n25254_), .S0(pi0299), .Y(new_n27583_));
  NAND3X1  g25147(.A(new_n25883_), .B(new_n25872_), .C(pi0214), .Y(new_n27584_));
  NAND2X1  g25148(.A(new_n27584_), .B(pi0212), .Y(new_n27585_));
  AOI21X1  g25149(.A0(new_n27583_), .A1(new_n24984_), .B0(new_n27585_), .Y(new_n27586_));
  AND2X1   g25150(.A(new_n27583_), .B(pi0214), .Y(new_n27587_));
  OR2X1    g25151(.A(new_n25888_), .B(pi0212), .Y(new_n27588_));
  OAI21X1  g25152(.A0(new_n27588_), .A1(new_n27587_), .B0(new_n23539_), .Y(new_n27589_));
  AOI21X1  g25153(.A0(new_n25883_), .A1(pi0219), .B0(new_n5118_), .Y(new_n27590_));
  OAI21X1  g25154(.A0(new_n27589_), .A1(new_n27586_), .B0(new_n27590_), .Y(new_n27591_));
  NOR3X1   g25155(.A(new_n27580_), .B(new_n25837_), .C(pi0057), .Y(new_n27592_));
  AOI21X1  g25156(.A0(new_n27592_), .A1(new_n27591_), .B0(new_n27582_), .Y(new_n27593_));
  AOI21X1  g25157(.A0(new_n27593_), .A1(new_n27581_), .B0(pi1152), .Y(new_n27594_));
  NAND2X1  g25158(.A(new_n26520_), .B(new_n26519_), .Y(new_n27595_));
  NAND2X1  g25159(.A(new_n27595_), .B(new_n26161_), .Y(new_n27596_));
  OAI21X1  g25160(.A0(new_n27571_), .A1(new_n25815_), .B0(new_n24984_), .Y(new_n27597_));
  AND2X1   g25161(.A(new_n27597_), .B(pi0212), .Y(new_n27598_));
  OAI21X1  g25162(.A0(new_n27571_), .A1(new_n27148_), .B0(new_n27149_), .Y(new_n27599_));
  AOI21X1  g25163(.A0(new_n27598_), .A1(new_n27596_), .B0(new_n27599_), .Y(new_n27600_));
  NOR3X1   g25164(.A(new_n27600_), .B(new_n26175_), .C(pi1151), .Y(new_n27601_));
  OR2X1    g25165(.A(new_n26115_), .B(pi0219), .Y(new_n27602_));
  NOR2X1   g25166(.A(new_n25254_), .B(new_n2953_), .Y(new_n27603_));
  NAND2X1  g25167(.A(new_n27603_), .B(new_n25014_), .Y(new_n27604_));
  OAI21X1  g25168(.A0(new_n25291_), .A1(new_n24961_), .B0(new_n27604_), .Y(new_n27605_));
  AOI21X1  g25169(.A0(new_n27605_), .A1(new_n26112_), .B0(new_n27602_), .Y(new_n27606_));
  OAI21X1  g25170(.A0(new_n26289_), .A1(new_n26209_), .B0(pi1151), .Y(new_n27607_));
  OAI21X1  g25171(.A0(new_n27607_), .A1(new_n27606_), .B0(new_n25294_), .Y(new_n27608_));
  OAI21X1  g25172(.A0(new_n27608_), .A1(new_n27601_), .B0(pi1150), .Y(new_n27609_));
  NOR3X1   g25173(.A(new_n26131_), .B(new_n25361_), .C(pi0211), .Y(new_n27610_));
  NOR3X1   g25174(.A(new_n26131_), .B(new_n25139_), .C(new_n8548_), .Y(new_n27611_));
  NOR3X1   g25175(.A(new_n27611_), .B(new_n27610_), .C(new_n25516_), .Y(new_n27612_));
  OAI21X1  g25176(.A0(new_n26123_), .A1(new_n25854_), .B0(new_n25419_), .Y(new_n27613_));
  OAI21X1  g25177(.A0(new_n26583_), .A1(new_n25014_), .B0(new_n27613_), .Y(new_n27614_));
  OAI21X1  g25178(.A0(new_n27614_), .A1(new_n27612_), .B0(new_n23539_), .Y(new_n27615_));
  AND2X1   g25179(.A(new_n26143_), .B(pi1151), .Y(new_n27616_));
  AOI21X1  g25180(.A0(new_n27603_), .A1(new_n25014_), .B0(new_n25871_), .Y(new_n27617_));
  NOR3X1   g25181(.A(new_n27617_), .B(new_n25838_), .C(new_n25256_), .Y(new_n27618_));
  INVX1    g25182(.A(new_n27618_), .Y(new_n27619_));
  NAND2X1  g25183(.A(new_n27619_), .B(new_n25258_), .Y(new_n27620_));
  AOI21X1  g25184(.A0(new_n27616_), .A1(new_n27615_), .B0(new_n27620_), .Y(new_n27621_));
  NOR4X1   g25185(.A(new_n27571_), .B(new_n25840_), .C(new_n25831_), .D(pi0212), .Y(new_n27622_));
  OAI21X1  g25186(.A0(new_n27603_), .A1(new_n26589_), .B0(pi0212), .Y(new_n27623_));
  AOI21X1  g25187(.A0(new_n26575_), .A1(pi0214), .B0(new_n27623_), .Y(new_n27624_));
  OAI21X1  g25188(.A0(new_n25868_), .A1(pi0212), .B0(new_n23539_), .Y(new_n27625_));
  NOR3X1   g25189(.A(new_n27625_), .B(new_n27624_), .C(new_n27622_), .Y(new_n27626_));
  NOR4X1   g25190(.A(new_n27626_), .B(new_n26278_), .C(po1038), .D(new_n25837_), .Y(new_n27627_));
  NAND2X1  g25191(.A(new_n27374_), .B(new_n25837_), .Y(new_n27628_));
  NAND3X1  g25192(.A(new_n27628_), .B(new_n27619_), .C(new_n25294_), .Y(new_n27629_));
  OAI21X1  g25193(.A0(new_n27629_), .A1(new_n27627_), .B0(new_n26471_), .Y(new_n27630_));
  OAI22X1  g25194(.A0(new_n27630_), .A1(new_n27621_), .B0(new_n27609_), .B1(new_n27594_), .Y(new_n27631_));
  AOI21X1  g25195(.A0(new_n27631_), .A1(pi0213), .B0(pi0209), .Y(new_n27632_));
  NOR3X1   g25196(.A(new_n25532_), .B(new_n25402_), .C(pi0207), .Y(new_n27633_));
  NOR3X1   g25197(.A(new_n25415_), .B(new_n25139_), .C(new_n22803_), .Y(new_n27634_));
  NOR2X1   g25198(.A(new_n27634_), .B(new_n23109_), .Y(new_n27635_));
  INVX1    g25199(.A(new_n27635_), .Y(new_n27636_));
  OAI22X1  g25200(.A0(new_n27636_), .A1(new_n27633_), .B0(new_n25533_), .B1(new_n25122_), .Y(new_n27637_));
  AND2X1   g25201(.A(new_n27637_), .B(pi0211), .Y(new_n27638_));
  AOI22X1  g25202(.A0(new_n27638_), .A1(pi0214), .B0(new_n25417_), .B1(new_n25740_), .Y(new_n27639_));
  INVX1    g25203(.A(new_n27639_), .Y(new_n27640_));
  AOI21X1  g25204(.A0(new_n27640_), .A1(new_n24961_), .B0(pi0219), .Y(new_n27641_));
  MX2X1    g25205(.A(new_n27637_), .B(new_n25417_), .S0(pi0211), .Y(new_n27642_));
  INVX1    g25206(.A(new_n27638_), .Y(new_n27643_));
  AOI21X1  g25207(.A0(new_n25417_), .A1(new_n8548_), .B0(pi0214), .Y(new_n27644_));
  AOI21X1  g25208(.A0(new_n27644_), .A1(new_n27643_), .B0(new_n24961_), .Y(new_n27645_));
  OAI21X1  g25209(.A0(new_n27642_), .A1(new_n24984_), .B0(new_n27645_), .Y(new_n27646_));
  AOI21X1  g25210(.A0(new_n27646_), .A1(new_n27641_), .B0(new_n25418_), .Y(new_n27647_));
  NOR3X1   g25211(.A(new_n25416_), .B(po1038), .C(pi1152), .Y(new_n27648_));
  OAI22X1  g25212(.A0(new_n27648_), .A1(new_n27500_), .B0(new_n27647_), .B1(new_n27299_), .Y(new_n27649_));
  NAND2X1  g25213(.A(new_n25341_), .B(pi0214), .Y(new_n27650_));
  AOI21X1  g25214(.A0(new_n27650_), .A1(new_n25388_), .B0(pi0219), .Y(new_n27651_));
  AOI21X1  g25215(.A0(new_n25341_), .A1(new_n24984_), .B0(new_n24961_), .Y(new_n27652_));
  OAI21X1  g25216(.A0(new_n25356_), .A1(new_n24984_), .B0(new_n27652_), .Y(new_n27653_));
  OAI21X1  g25217(.A0(new_n25446_), .A1(new_n23539_), .B0(new_n6520_), .Y(new_n27654_));
  AOI21X1  g25218(.A0(new_n27653_), .A1(new_n27651_), .B0(new_n27654_), .Y(new_n27655_));
  AOI21X1  g25219(.A0(new_n26582_), .A1(new_n25354_), .B0(po1038), .Y(new_n27656_));
  OAI21X1  g25220(.A0(new_n26582_), .A1(new_n25356_), .B0(new_n27656_), .Y(new_n27657_));
  AOI21X1  g25221(.A0(new_n27657_), .A1(new_n27352_), .B0(new_n25289_), .Y(new_n27658_));
  OAI21X1  g25222(.A0(new_n27655_), .A1(new_n26503_), .B0(new_n27658_), .Y(new_n27659_));
  AOI21X1  g25223(.A0(new_n27659_), .A1(new_n27649_), .B0(pi1150), .Y(new_n27660_));
  OAI21X1  g25224(.A0(new_n25416_), .A1(new_n25323_), .B0(pi0219), .Y(new_n27661_));
  AOI21X1  g25225(.A0(new_n27642_), .A1(new_n25323_), .B0(new_n27661_), .Y(new_n27662_));
  OR2X1    g25226(.A(new_n27662_), .B(po1038), .Y(new_n27663_));
  OAI21X1  g25227(.A0(new_n27637_), .A1(new_n24984_), .B0(new_n27645_), .Y(new_n27664_));
  AOI21X1  g25228(.A0(new_n27664_), .A1(new_n27641_), .B0(new_n27663_), .Y(new_n27665_));
  OR2X1    g25229(.A(new_n27665_), .B(new_n27302_), .Y(new_n27666_));
  OAI21X1  g25230(.A0(new_n25416_), .A1(pi0212), .B0(new_n23539_), .Y(new_n27667_));
  AOI21X1  g25231(.A0(new_n27640_), .A1(pi0212), .B0(new_n27667_), .Y(new_n27668_));
  OAI21X1  g25232(.A0(new_n27668_), .A1(new_n27663_), .B0(new_n26478_), .Y(new_n27669_));
  NAND3X1  g25233(.A(new_n27669_), .B(new_n27666_), .C(new_n25289_), .Y(new_n27670_));
  INVX1    g25234(.A(new_n25359_), .Y(new_n27671_));
  MX2X1    g25235(.A(new_n25356_), .B(new_n25446_), .S0(new_n24984_), .Y(new_n27672_));
  MX2X1    g25236(.A(new_n25354_), .B(new_n25341_), .S0(pi0211), .Y(new_n27673_));
  NOR2X1   g25237(.A(new_n27673_), .B(new_n24984_), .Y(new_n27674_));
  AND2X1   g25238(.A(new_n25356_), .B(new_n24984_), .Y(new_n27675_));
  OR2X1    g25239(.A(new_n27675_), .B(new_n24961_), .Y(new_n27676_));
  OAI22X1  g25240(.A0(new_n27676_), .A1(new_n27674_), .B0(new_n27672_), .B1(pi0212), .Y(new_n27677_));
  AOI21X1  g25241(.A0(new_n27677_), .A1(new_n23539_), .B0(new_n27671_), .Y(new_n27678_));
  OAI21X1  g25242(.A0(new_n25341_), .A1(new_n24961_), .B0(new_n27651_), .Y(new_n27679_));
  AOI21X1  g25243(.A0(new_n27679_), .A1(new_n25359_), .B0(new_n26485_), .Y(new_n27680_));
  NOR2X1   g25244(.A(new_n27680_), .B(new_n25289_), .Y(new_n27681_));
  OAI21X1  g25245(.A0(new_n27678_), .A1(new_n27348_), .B0(new_n27681_), .Y(new_n27682_));
  AOI21X1  g25246(.A0(new_n27682_), .A1(new_n27670_), .B0(new_n26471_), .Y(new_n27683_));
  OAI21X1  g25247(.A0(new_n27683_), .A1(new_n27660_), .B0(new_n25003_), .Y(new_n27684_));
  AOI21X1  g25248(.A0(new_n25422_), .A1(pi0213), .B0(new_n23244_), .Y(new_n27685_));
  AOI22X1  g25249(.A0(new_n27685_), .A1(new_n27684_), .B0(new_n27632_), .B1(new_n27570_), .Y(new_n27686_));
  MX2X1    g25250(.A(new_n27686_), .B(pi0249), .S0(new_n24954_), .Y(po0406));
  NOR4X1   g25251(.A(new_n7832_), .B(new_n3138_), .C(new_n3256_), .D(new_n2487_), .Y(new_n27688_));
  OAI21X1  g25252(.A0(new_n27688_), .A1(new_n5087_), .B0(new_n3095_), .Y(new_n27689_));
  NAND3X1  g25253(.A(new_n5813_), .B(new_n3026_), .C(pi0075), .Y(new_n27690_));
  NAND3X1  g25254(.A(new_n6756_), .B(new_n7846_), .C(new_n3156_), .Y(new_n27691_));
  AOI21X1  g25255(.A0(new_n27690_), .A1(new_n27689_), .B0(new_n27691_), .Y(po0407));
  NOR3X1   g25256(.A(pi0476), .B(new_n8009_), .C(pi0199), .Y(new_n27693_));
  AOI21X1  g25257(.A0(new_n8130_), .A1(pi0897), .B0(new_n27693_), .Y(new_n27694_));
  INVX1    g25258(.A(pi1053), .Y(new_n27695_));
  AOI21X1  g25259(.A0(pi1039), .A1(pi0200), .B0(pi0199), .Y(new_n27696_));
  OAI21X1  g25260(.A0(new_n27695_), .A1(pi0200), .B0(new_n27696_), .Y(new_n27697_));
  MX2X1    g25261(.A(new_n27697_), .B(pi0251), .S0(new_n27694_), .Y(po0408));
  OAI21X1  g25262(.A0(new_n5033_), .A1(new_n5031_), .B0(new_n8624_), .Y(new_n27699_));
  INVX1    g25263(.A(pi1001), .Y(new_n27700_));
  OR2X1    g25264(.A(pi0984), .B(pi0979), .Y(new_n27701_));
  OR2X1    g25265(.A(new_n27701_), .B(new_n27700_), .Y(new_n27702_));
  NOR4X1   g25266(.A(new_n27702_), .B(new_n5243_), .C(new_n5041_), .D(new_n5038_), .Y(new_n27703_));
  AND2X1   g25267(.A(new_n2756_), .B(pi1092), .Y(new_n27704_));
  OAI21X1  g25268(.A0(new_n27703_), .A1(pi0252), .B0(new_n27704_), .Y(new_n27705_));
  MX2X1    g25269(.A(new_n5256_), .B(new_n5257_), .S0(new_n27705_), .Y(new_n27706_));
  OAI21X1  g25270(.A0(new_n27706_), .A1(new_n6270_), .B0(new_n27699_), .Y(new_n27707_));
  MX2X1    g25271(.A(new_n27706_), .B(new_n8625_), .S0(new_n5052_), .Y(new_n27708_));
  OAI21X1  g25272(.A0(new_n27708_), .A1(new_n5070_), .B0(pi0299), .Y(new_n27709_));
  AOI21X1  g25273(.A0(new_n27707_), .A1(new_n5070_), .B0(new_n27709_), .Y(new_n27710_));
  OAI21X1  g25274(.A0(new_n27708_), .A1(new_n5050_), .B0(new_n2953_), .Y(new_n27711_));
  AOI21X1  g25275(.A0(new_n27707_), .A1(new_n5050_), .B0(new_n27711_), .Y(new_n27712_));
  OR4X1    g25276(.A(new_n27712_), .B(new_n27710_), .C(new_n9590_), .D(new_n9580_), .Y(new_n27713_));
  AOI21X1  g25277(.A0(new_n8624_), .A1(new_n8245_), .B0(new_n6748_), .Y(new_n27714_));
  OR4X1    g25278(.A(new_n27702_), .B(new_n5038_), .C(new_n2959_), .D(pi0038), .Y(new_n27715_));
  OR4X1    g25279(.A(new_n27715_), .B(new_n24938_), .C(new_n14758_), .D(new_n7698_), .Y(new_n27716_));
  OAI21X1  g25280(.A0(new_n27716_), .A1(new_n5243_), .B0(new_n3053_), .Y(new_n27717_));
  AND2X1   g25281(.A(pi1092), .B(new_n2436_), .Y(new_n27718_));
  OAI21X1  g25282(.A0(new_n8623_), .A1(new_n2436_), .B0(new_n6748_), .Y(new_n27719_));
  AOI21X1  g25283(.A0(new_n27718_), .A1(new_n27717_), .B0(new_n27719_), .Y(new_n27720_));
  AOI21X1  g25284(.A0(new_n27714_), .A1(new_n27713_), .B0(new_n27720_), .Y(po0409));
  NOR4X1   g25285(.A(new_n25096_), .B(new_n25021_), .C(new_n9544_), .D(po1038), .Y(new_n27722_));
  AOI21X1  g25286(.A0(new_n5117_), .A1(new_n2436_), .B0(pi0211), .Y(new_n27723_));
  AND2X1   g25287(.A(new_n27723_), .B(pi0219), .Y(new_n27724_));
  NOR2X1   g25288(.A(new_n27724_), .B(new_n27722_), .Y(new_n27725_));
  INVX1    g25289(.A(new_n27725_), .Y(new_n27726_));
  AOI21X1  g25290(.A0(new_n27726_), .A1(pi1153), .B0(pi1151), .Y(new_n27727_));
  INVX1    g25291(.A(new_n8075_), .Y(new_n27728_));
  NOR2X1   g25292(.A(new_n25055_), .B(new_n25054_), .Y(new_n27729_));
  OAI22X1  g25293(.A0(new_n25084_), .A1(new_n27728_), .B0(new_n27729_), .B1(new_n8548_), .Y(new_n27730_));
  INVX1    g25294(.A(new_n27730_), .Y(new_n27731_));
  OAI22X1  g25295(.A0(new_n8502_), .A1(pi1153), .B0(pi0299), .B1(new_n8009_), .Y(new_n27732_));
  AOI21X1  g25296(.A0(new_n27732_), .A1(new_n25030_), .B0(po1038), .Y(new_n27733_));
  AND2X1   g25297(.A(new_n23539_), .B(pi0211), .Y(new_n27734_));
  OAI21X1  g25298(.A0(new_n25607_), .A1(new_n27734_), .B0(pi1151), .Y(new_n27735_));
  AOI21X1  g25299(.A0(new_n27733_), .A1(new_n27731_), .B0(new_n27735_), .Y(new_n27736_));
  OAI21X1  g25300(.A0(new_n27736_), .A1(new_n27727_), .B0(new_n25289_), .Y(new_n27737_));
  NOR4X1   g25301(.A(new_n25107_), .B(new_n12494_), .C(new_n23539_), .D(pi0211), .Y(new_n27738_));
  NOR4X1   g25302(.A(new_n27738_), .B(new_n25088_), .C(new_n8549_), .D(pi1151), .Y(new_n27739_));
  MX2X1    g25303(.A(pi0200), .B(pi0211), .S0(pi0299), .Y(new_n27740_));
  NOR2X1   g25304(.A(new_n27740_), .B(new_n12494_), .Y(new_n27741_));
  MX2X1    g25305(.A(new_n23539_), .B(new_n7941_), .S0(new_n2953_), .Y(new_n27742_));
  NOR3X1   g25306(.A(new_n27742_), .B(new_n27741_), .C(new_n25837_), .Y(new_n27743_));
  OR2X1    g25307(.A(new_n27743_), .B(po1038), .Y(new_n27744_));
  AOI21X1  g25308(.A0(new_n8075_), .A1(new_n25837_), .B0(new_n25606_), .Y(new_n27745_));
  AOI21X1  g25309(.A0(new_n27745_), .A1(po1038), .B0(new_n25289_), .Y(new_n27746_));
  OAI21X1  g25310(.A0(new_n27744_), .A1(new_n27739_), .B0(new_n27746_), .Y(new_n27747_));
  AOI21X1  g25311(.A0(new_n27747_), .A1(new_n27737_), .B0(new_n24954_), .Y(new_n27748_));
  NOR2X1   g25312(.A(new_n26698_), .B(new_n26697_), .Y(new_n27749_));
  INVX1    g25313(.A(new_n27749_), .Y(new_n27750_));
  INVX1    g25314(.A(new_n26736_), .Y(new_n27751_));
  OAI21X1  g25315(.A0(new_n27751_), .A1(new_n27750_), .B0(pi1153), .Y(new_n27752_));
  NOR2X1   g25316(.A(new_n26756_), .B(pi1153), .Y(new_n27753_));
  NOR2X1   g25317(.A(new_n27753_), .B(pi0219), .Y(new_n27754_));
  NAND2X1  g25318(.A(new_n27754_), .B(new_n27752_), .Y(new_n27755_));
  AOI21X1  g25319(.A0(new_n26701_), .A1(new_n26682_), .B0(new_n26716_), .Y(new_n27756_));
  INVX1    g25320(.A(new_n27756_), .Y(new_n27757_));
  AOI21X1  g25321(.A0(new_n26698_), .A1(new_n8548_), .B0(new_n27757_), .Y(new_n27758_));
  INVX1    g25322(.A(new_n26726_), .Y(new_n27759_));
  NOR2X1   g25323(.A(new_n27759_), .B(new_n26697_), .Y(new_n27760_));
  AND2X1   g25324(.A(new_n27760_), .B(new_n27758_), .Y(new_n27761_));
  OR2X1    g25325(.A(new_n27761_), .B(new_n12494_), .Y(new_n27762_));
  NOR2X1   g25326(.A(new_n26815_), .B(pi1153), .Y(new_n27763_));
  INVX1    g25327(.A(new_n27763_), .Y(new_n27764_));
  NAND3X1  g25328(.A(new_n27764_), .B(new_n27762_), .C(pi0219), .Y(new_n27765_));
  NAND3X1  g25329(.A(new_n27765_), .B(new_n27755_), .C(pi0253), .Y(new_n27766_));
  NOR2X1   g25330(.A(new_n26754_), .B(new_n26704_), .Y(new_n27767_));
  INVX1    g25331(.A(new_n27767_), .Y(new_n27768_));
  INVX1    g25332(.A(new_n26815_), .Y(new_n27769_));
  NOR3X1   g25333(.A(new_n27769_), .B(new_n26706_), .C(pi0211), .Y(new_n27770_));
  OAI21X1  g25334(.A0(new_n27770_), .A1(new_n26707_), .B0(pi1153), .Y(new_n27771_));
  NAND3X1  g25335(.A(new_n27771_), .B(new_n27768_), .C(pi0219), .Y(new_n27772_));
  INVX1    g25336(.A(new_n26715_), .Y(new_n27773_));
  INVX1    g25337(.A(new_n26716_), .Y(new_n27774_));
  NAND3X1  g25338(.A(new_n27774_), .B(new_n27773_), .C(pi1153), .Y(new_n27775_));
  NOR3X1   g25339(.A(new_n26754_), .B(new_n26716_), .C(pi1153), .Y(new_n27776_));
  INVX1    g25340(.A(new_n27776_), .Y(new_n27777_));
  NAND3X1  g25341(.A(new_n27777_), .B(new_n27775_), .C(new_n23539_), .Y(new_n27778_));
  NAND3X1  g25342(.A(new_n27778_), .B(new_n27772_), .C(new_n26778_), .Y(new_n27779_));
  AOI21X1  g25343(.A0(new_n27779_), .A1(new_n27766_), .B0(po1038), .Y(new_n27780_));
  INVX1    g25344(.A(new_n26689_), .Y(new_n27781_));
  AOI21X1  g25345(.A0(new_n26690_), .A1(new_n2722_), .B0(pi0219), .Y(new_n27782_));
  INVX1    g25346(.A(new_n27782_), .Y(new_n27783_));
  AOI21X1  g25347(.A0(new_n27781_), .A1(new_n8548_), .B0(new_n27783_), .Y(new_n27784_));
  NOR4X1   g25348(.A(new_n27784_), .B(new_n26680_), .C(new_n6520_), .D(pi0219), .Y(new_n27785_));
  AND2X1   g25349(.A(pi1091), .B(pi0219), .Y(new_n27786_));
  INVX1    g25350(.A(new_n27786_), .Y(new_n27787_));
  NOR2X1   g25351(.A(new_n27787_), .B(new_n25015_), .Y(new_n27788_));
  NOR3X1   g25352(.A(new_n27788_), .B(new_n27782_), .C(new_n26744_), .Y(new_n27789_));
  NOR2X1   g25353(.A(new_n27789_), .B(new_n26778_), .Y(new_n27790_));
  AOI21X1  g25354(.A0(new_n26744_), .A1(pi0211), .B0(new_n23539_), .Y(new_n27791_));
  OAI21X1  g25355(.A0(new_n26680_), .A1(pi0211), .B0(new_n27791_), .Y(new_n27792_));
  NOR2X1   g25356(.A(new_n26689_), .B(pi0219), .Y(new_n27793_));
  NOR2X1   g25357(.A(new_n27793_), .B(new_n27788_), .Y(new_n27794_));
  AOI21X1  g25358(.A0(new_n27794_), .A1(new_n27792_), .B0(pi0253), .Y(new_n27795_));
  OR2X1    g25359(.A(new_n27795_), .B(new_n6520_), .Y(new_n27796_));
  OAI21X1  g25360(.A0(new_n27796_), .A1(new_n27790_), .B0(pi1151), .Y(new_n27797_));
  NOR2X1   g25361(.A(new_n27797_), .B(new_n27785_), .Y(new_n27798_));
  INVX1    g25362(.A(new_n27798_), .Y(new_n27799_));
  INVX1    g25363(.A(new_n27758_), .Y(new_n27800_));
  OR2X1    g25364(.A(new_n26720_), .B(new_n26716_), .Y(new_n27801_));
  AND2X1   g25365(.A(new_n27801_), .B(new_n12494_), .Y(new_n27802_));
  NOR3X1   g25366(.A(new_n27802_), .B(new_n27800_), .C(new_n26715_), .Y(new_n27803_));
  MX2X1    g25367(.A(new_n27803_), .B(new_n26786_), .S0(pi0219), .Y(new_n27804_));
  AOI21X1  g25368(.A0(new_n27804_), .A1(new_n27772_), .B0(pi0253), .Y(new_n27805_));
  NOR2X1   g25369(.A(new_n26720_), .B(new_n26697_), .Y(new_n27806_));
  INVX1    g25370(.A(new_n27770_), .Y(new_n27807_));
  AOI21X1  g25371(.A0(new_n27807_), .A1(new_n27750_), .B0(new_n27783_), .Y(new_n27808_));
  OAI21X1  g25372(.A0(new_n27802_), .A1(new_n27806_), .B0(new_n27808_), .Y(new_n27809_));
  NOR3X1   g25373(.A(new_n26710_), .B(new_n26697_), .C(new_n23539_), .Y(new_n27810_));
  OAI21X1  g25374(.A0(new_n27762_), .A1(new_n26794_), .B0(new_n27810_), .Y(new_n27811_));
  AOI21X1  g25375(.A0(new_n27811_), .A1(new_n27809_), .B0(new_n26778_), .Y(new_n27812_));
  NOR3X1   g25376(.A(new_n27812_), .B(new_n27805_), .C(po1038), .Y(new_n27813_));
  OAI22X1  g25377(.A0(new_n27813_), .A1(pi1151), .B0(new_n27799_), .B1(new_n27780_), .Y(new_n27814_));
  NOR2X1   g25378(.A(new_n27796_), .B(new_n27790_), .Y(new_n27815_));
  INVX1    g25379(.A(new_n27793_), .Y(new_n27816_));
  AOI21X1  g25380(.A0(new_n26681_), .A1(new_n8548_), .B0(new_n27816_), .Y(new_n27817_));
  NOR2X1   g25381(.A(new_n27817_), .B(new_n27783_), .Y(new_n27818_));
  NOR2X1   g25382(.A(new_n26680_), .B(new_n23539_), .Y(new_n27819_));
  NOR2X1   g25383(.A(new_n27819_), .B(new_n6520_), .Y(new_n27820_));
  INVX1    g25384(.A(new_n27820_), .Y(new_n27821_));
  NOR2X1   g25385(.A(new_n27821_), .B(new_n27818_), .Y(new_n27822_));
  AOI21X1  g25386(.A0(new_n27822_), .A1(new_n26681_), .B0(new_n27815_), .Y(new_n27823_));
  AOI21X1  g25387(.A0(new_n27823_), .A1(new_n27814_), .B0(new_n25289_), .Y(new_n27824_));
  NAND2X1  g25388(.A(new_n27771_), .B(new_n27768_), .Y(new_n27825_));
  AOI22X1  g25389(.A0(new_n27808_), .A1(new_n27778_), .B0(new_n27825_), .B1(pi0219), .Y(new_n27826_));
  OAI21X1  g25390(.A0(new_n27826_), .A1(new_n26706_), .B0(new_n26778_), .Y(new_n27827_));
  OAI21X1  g25391(.A0(new_n26716_), .A1(new_n26701_), .B0(pi1153), .Y(new_n27828_));
  AND2X1   g25392(.A(new_n27782_), .B(new_n27758_), .Y(new_n27829_));
  AND2X1   g25393(.A(new_n27829_), .B(new_n27828_), .Y(new_n27830_));
  AOI21X1  g25394(.A0(new_n27760_), .A1(new_n27758_), .B0(new_n26782_), .Y(new_n27831_));
  OAI21X1  g25395(.A0(new_n26820_), .A1(pi1153), .B0(pi0219), .Y(new_n27832_));
  AOI21X1  g25396(.A0(new_n27831_), .A1(pi1153), .B0(new_n27832_), .Y(new_n27833_));
  OAI21X1  g25397(.A0(new_n27833_), .A1(new_n27830_), .B0(pi0253), .Y(new_n27834_));
  NAND3X1  g25398(.A(new_n27834_), .B(new_n27827_), .C(new_n6520_), .Y(new_n27835_));
  NAND3X1  g25399(.A(new_n27825_), .B(new_n26696_), .C(pi0219), .Y(new_n27836_));
  NOR2X1   g25400(.A(new_n26728_), .B(pi1153), .Y(new_n27837_));
  OR4X1    g25401(.A(new_n27837_), .B(new_n26757_), .C(new_n26706_), .D(pi0219), .Y(new_n27838_));
  AND2X1   g25402(.A(new_n27838_), .B(new_n26778_), .Y(new_n27839_));
  AOI21X1  g25403(.A0(new_n27768_), .A1(new_n2722_), .B0(pi1153), .Y(new_n27840_));
  NOR3X1   g25404(.A(new_n26720_), .B(new_n26716_), .C(pi0219), .Y(new_n27841_));
  NOR4X1   g25405(.A(new_n27841_), .B(new_n27840_), .C(new_n27761_), .D(new_n26794_), .Y(new_n27842_));
  OAI21X1  g25406(.A0(new_n27842_), .A1(new_n26778_), .B0(new_n6520_), .Y(new_n27843_));
  AOI21X1  g25407(.A0(new_n27839_), .A1(new_n27836_), .B0(new_n27843_), .Y(new_n27844_));
  OAI21X1  g25408(.A0(new_n27796_), .A1(new_n27790_), .B0(new_n25837_), .Y(new_n27845_));
  OAI21X1  g25409(.A0(new_n27845_), .A1(new_n27844_), .B0(new_n25289_), .Y(new_n27846_));
  AOI21X1  g25410(.A0(new_n27835_), .A1(new_n27798_), .B0(new_n27846_), .Y(new_n27847_));
  OAI21X1  g25411(.A0(new_n27847_), .A1(new_n27824_), .B0(new_n26899_), .Y(new_n27848_));
  NOR2X1   g25412(.A(new_n26834_), .B(pi1153), .Y(new_n27849_));
  OAI21X1  g25413(.A0(new_n26856_), .A1(new_n12494_), .B0(new_n25030_), .Y(new_n27850_));
  OAI22X1  g25414(.A0(new_n27850_), .A1(new_n27849_), .B0(new_n27731_), .B1(new_n2722_), .Y(new_n27851_));
  NAND2X1  g25415(.A(new_n27851_), .B(pi0253), .Y(new_n27852_));
  OAI21X1  g25416(.A0(new_n27741_), .A1(new_n9546_), .B0(pi1091), .Y(new_n27853_));
  AOI21X1  g25417(.A0(new_n27853_), .A1(new_n26778_), .B0(po1038), .Y(new_n27854_));
  OAI22X1  g25418(.A0(new_n5118_), .A1(pi0057), .B0(pi1091), .B1(pi0253), .Y(new_n27855_));
  AND2X1   g25419(.A(pi1091), .B(pi0211), .Y(new_n27856_));
  INVX1    g25420(.A(new_n27856_), .Y(new_n27857_));
  AND2X1   g25421(.A(new_n12494_), .B(pi1091), .Y(new_n27858_));
  INVX1    g25422(.A(new_n27858_), .Y(new_n27859_));
  OAI21X1  g25423(.A0(new_n27859_), .A1(new_n23539_), .B0(new_n27857_), .Y(new_n27860_));
  OAI21X1  g25424(.A0(new_n27860_), .A1(new_n27855_), .B0(pi1151), .Y(new_n27861_));
  AOI21X1  g25425(.A0(new_n27854_), .A1(new_n27852_), .B0(new_n27861_), .Y(new_n27862_));
  NOR3X1   g25426(.A(new_n27855_), .B(new_n27788_), .C(new_n23539_), .Y(new_n27863_));
  AND2X1   g25427(.A(pi1153), .B(pi1091), .Y(new_n27864_));
  AND2X1   g25428(.A(new_n27864_), .B(new_n27722_), .Y(new_n27865_));
  AND2X1   g25429(.A(new_n2722_), .B(pi0253), .Y(new_n27866_));
  NOR4X1   g25430(.A(new_n27866_), .B(new_n27865_), .C(new_n27863_), .D(pi1151), .Y(new_n27867_));
  OAI21X1  g25431(.A0(new_n27867_), .A1(new_n27862_), .B0(new_n25289_), .Y(new_n27868_));
  AND2X1   g25432(.A(new_n26861_), .B(new_n12494_), .Y(new_n27869_));
  NOR3X1   g25433(.A(new_n25039_), .B(new_n2722_), .C(pi0299), .Y(new_n27870_));
  OAI21X1  g25434(.A0(new_n27870_), .A1(new_n12494_), .B0(new_n25030_), .Y(new_n27871_));
  OR2X1    g25435(.A(new_n27871_), .B(new_n27869_), .Y(new_n27872_));
  INVX1    g25436(.A(new_n27734_), .Y(new_n27873_));
  NOR4X1   g25437(.A(new_n25088_), .B(new_n27873_), .C(new_n2722_), .D(pi0299), .Y(new_n27874_));
  NOR2X1   g25438(.A(new_n27874_), .B(new_n26778_), .Y(new_n27875_));
  NOR3X1   g25439(.A(new_n25107_), .B(new_n12494_), .C(new_n2722_), .Y(new_n27876_));
  OR2X1    g25440(.A(pi1153), .B(pi0199), .Y(new_n27877_));
  NOR4X1   g25441(.A(new_n27877_), .B(new_n2722_), .C(pi0299), .D(new_n8009_), .Y(new_n27878_));
  OR4X1    g25442(.A(new_n27878_), .B(new_n27876_), .C(new_n23539_), .D(pi0211), .Y(new_n27879_));
  NOR4X1   g25443(.A(new_n25055_), .B(new_n25048_), .C(new_n2722_), .D(pi0299), .Y(new_n27880_));
  NOR3X1   g25444(.A(new_n27880_), .B(new_n26869_), .C(new_n8548_), .Y(new_n27881_));
  NOR2X1   g25445(.A(new_n27881_), .B(pi0253), .Y(new_n27882_));
  AOI22X1  g25446(.A0(new_n27882_), .A1(new_n27879_), .B0(new_n27875_), .B1(new_n27872_), .Y(new_n27883_));
  XOR2X1   g25447(.A(pi0219), .B(new_n8548_), .Y(new_n27884_));
  INVX1    g25448(.A(new_n27884_), .Y(new_n27885_));
  NOR3X1   g25449(.A(new_n27885_), .B(new_n27880_), .C(new_n27866_), .Y(new_n27886_));
  OR4X1    g25450(.A(new_n27886_), .B(new_n27883_), .C(po1038), .D(pi1151), .Y(new_n27887_));
  OAI21X1  g25451(.A0(pi1091), .A1(new_n26778_), .B0(new_n27740_), .Y(new_n27888_));
  AOI21X1  g25452(.A0(new_n27888_), .A1(new_n27859_), .B0(new_n27742_), .Y(new_n27889_));
  OAI21X1  g25453(.A0(pi1091), .A1(pi0253), .B0(new_n6520_), .Y(new_n27890_));
  OAI22X1  g25454(.A0(new_n27890_), .A1(new_n27889_), .B0(new_n27855_), .B1(new_n27788_), .Y(new_n27891_));
  NOR3X1   g25455(.A(new_n2722_), .B(pi0219), .C(pi0211), .Y(new_n27892_));
  NOR3X1   g25456(.A(new_n27892_), .B(new_n27855_), .C(new_n27788_), .Y(new_n27893_));
  OR2X1    g25457(.A(new_n27893_), .B(new_n25289_), .Y(new_n27894_));
  AOI21X1  g25458(.A0(new_n27891_), .A1(pi1151), .B0(new_n27894_), .Y(new_n27895_));
  AOI21X1  g25459(.A0(new_n27895_), .A1(new_n27887_), .B0(new_n26899_), .Y(new_n27896_));
  AOI21X1  g25460(.A0(new_n27896_), .A1(new_n27868_), .B0(pi0230), .Y(new_n27897_));
  AOI21X1  g25461(.A0(new_n27897_), .A1(new_n27848_), .B0(new_n27748_), .Y(po0410));
  OAI22X1  g25462(.A0(new_n25053_), .A1(pi1153), .B0(new_n25039_), .B1(pi0299), .Y(new_n27899_));
  OAI22X1  g25463(.A0(new_n25393_), .A1(new_n25135_), .B0(new_n27899_), .B1(new_n12615_), .Y(new_n27900_));
  OAI22X1  g25464(.A0(new_n25346_), .A1(new_n27734_), .B0(new_n25031_), .B1(new_n2953_), .Y(new_n27901_));
  AOI22X1  g25465(.A0(new_n27901_), .A1(new_n25326_), .B0(new_n27900_), .B1(new_n27734_), .Y(new_n27902_));
  MX2X1    g25466(.A(new_n25830_), .B(new_n25628_), .S0(pi0219), .Y(new_n27903_));
  AOI21X1  g25467(.A0(new_n27903_), .A1(po1038), .B0(pi1152), .Y(new_n27904_));
  OAI21X1  g25468(.A0(new_n27902_), .A1(po1038), .B0(new_n27904_), .Y(new_n27905_));
  AND2X1   g25469(.A(pi1154), .B(pi0211), .Y(new_n27906_));
  OAI21X1  g25470(.A0(new_n25372_), .A1(new_n25045_), .B0(new_n27906_), .Y(new_n27907_));
  INVX1    g25471(.A(new_n27907_), .Y(new_n27908_));
  NOR2X1   g25472(.A(new_n25412_), .B(pi1154), .Y(new_n27909_));
  NOR3X1   g25473(.A(new_n27909_), .B(new_n27908_), .C(new_n25328_), .Y(new_n27910_));
  OR2X1    g25474(.A(new_n27910_), .B(new_n23539_), .Y(new_n27911_));
  OR2X1    g25475(.A(new_n12615_), .B(pi0200), .Y(new_n27912_));
  AOI22X1  g25476(.A0(new_n27912_), .A1(new_n25086_), .B0(new_n26186_), .B1(new_n25372_), .Y(new_n27913_));
  OR2X1    g25477(.A(new_n27913_), .B(pi0219), .Y(new_n27914_));
  AND2X1   g25478(.A(new_n27914_), .B(new_n6520_), .Y(new_n27915_));
  AND2X1   g25479(.A(new_n27915_), .B(new_n27911_), .Y(new_n27916_));
  NOR3X1   g25480(.A(pi1153), .B(pi0219), .C(new_n8548_), .Y(new_n27917_));
  OAI21X1  g25481(.A0(new_n27917_), .A1(new_n26085_), .B0(pi1152), .Y(new_n27918_));
  OAI21X1  g25482(.A0(new_n27918_), .A1(new_n27916_), .B0(new_n27905_), .Y(new_n27919_));
  AOI21X1  g25483(.A0(new_n27803_), .A1(new_n12494_), .B0(new_n26756_), .Y(new_n27920_));
  NOR3X1   g25484(.A(new_n27800_), .B(new_n26701_), .C(new_n12615_), .Y(new_n27921_));
  AOI21X1  g25485(.A0(new_n27921_), .A1(new_n27752_), .B0(new_n26779_), .Y(new_n27922_));
  OAI21X1  g25486(.A0(new_n27920_), .A1(pi1154), .B0(new_n27922_), .Y(new_n27923_));
  AOI21X1  g25487(.A0(new_n26706_), .A1(new_n26692_), .B0(new_n26821_), .Y(new_n27924_));
  AND2X1   g25488(.A(new_n27924_), .B(pi1154), .Y(new_n27925_));
  NOR3X1   g25489(.A(new_n26689_), .B(new_n2953_), .C(new_n8548_), .Y(new_n27926_));
  OAI21X1  g25490(.A0(new_n27926_), .A1(new_n26706_), .B0(new_n12494_), .Y(new_n27927_));
  AND2X1   g25491(.A(new_n27927_), .B(new_n26779_), .Y(new_n27928_));
  OAI21X1  g25492(.A0(new_n27925_), .A1(new_n26755_), .B0(new_n27928_), .Y(new_n27929_));
  AOI21X1  g25493(.A0(new_n27929_), .A1(new_n27923_), .B0(pi0219), .Y(new_n27930_));
  OAI21X1  g25494(.A0(new_n27761_), .A1(new_n12494_), .B0(pi1154), .Y(new_n27931_));
  AOI21X1  g25495(.A0(new_n26821_), .A1(new_n12494_), .B0(pi1154), .Y(new_n27932_));
  OAI21X1  g25496(.A0(new_n26815_), .A1(new_n12494_), .B0(new_n27932_), .Y(new_n27933_));
  AND2X1   g25497(.A(new_n27933_), .B(pi0254), .Y(new_n27934_));
  OAI21X1  g25498(.A0(new_n27931_), .A1(new_n27831_), .B0(new_n27934_), .Y(new_n27935_));
  INVX1    g25499(.A(new_n25628_), .Y(new_n27936_));
  AOI21X1  g25500(.A0(new_n27924_), .A1(new_n27764_), .B0(new_n27936_), .Y(new_n27937_));
  OAI21X1  g25501(.A0(new_n26680_), .A1(pi0200), .B0(new_n27937_), .Y(new_n27938_));
  NOR2X1   g25502(.A(new_n26745_), .B(pi1153), .Y(new_n27939_));
  NOR4X1   g25503(.A(new_n27939_), .B(new_n26754_), .C(new_n26704_), .D(new_n26701_), .Y(new_n27940_));
  NOR2X1   g25504(.A(new_n27940_), .B(pi1154), .Y(new_n27941_));
  OAI21X1  g25505(.A0(new_n27768_), .A1(new_n26706_), .B0(new_n27941_), .Y(new_n27942_));
  AND2X1   g25506(.A(new_n26707_), .B(pi1153), .Y(new_n27943_));
  OR4X1    g25507(.A(new_n27943_), .B(new_n26807_), .C(new_n12615_), .D(new_n8548_), .Y(new_n27944_));
  NAND4X1  g25508(.A(new_n27944_), .B(new_n27942_), .C(new_n27938_), .D(new_n26779_), .Y(new_n27945_));
  AOI21X1  g25509(.A0(new_n27945_), .A1(new_n27935_), .B0(new_n23539_), .Y(new_n27946_));
  NOR3X1   g25510(.A(new_n27946_), .B(new_n27930_), .C(new_n26778_), .Y(new_n27947_));
  OR2X1    g25511(.A(new_n26845_), .B(new_n12494_), .Y(new_n27948_));
  AND2X1   g25512(.A(new_n27948_), .B(new_n12615_), .Y(new_n27949_));
  AOI21X1  g25513(.A0(new_n25376_), .A1(new_n8548_), .B0(new_n27849_), .Y(new_n27950_));
  INVX1    g25514(.A(new_n27906_), .Y(new_n27951_));
  NOR4X1   g25515(.A(new_n25400_), .B(new_n25053_), .C(new_n27951_), .D(new_n2722_), .Y(new_n27952_));
  AOI21X1  g25516(.A0(new_n27950_), .A1(new_n27949_), .B0(new_n27952_), .Y(new_n27953_));
  AND2X1   g25517(.A(pi1091), .B(new_n8548_), .Y(new_n27954_));
  AOI21X1  g25518(.A0(new_n27954_), .A1(pi1154), .B0(new_n27786_), .Y(new_n27955_));
  OAI22X1  g25519(.A0(new_n27955_), .A1(new_n27910_), .B0(new_n27953_), .B1(pi0219), .Y(new_n27956_));
  AND2X1   g25520(.A(new_n27956_), .B(pi0254), .Y(new_n27957_));
  NOR2X1   g25521(.A(new_n25412_), .B(new_n23539_), .Y(new_n27958_));
  OAI21X1  g25522(.A0(new_n27740_), .A1(new_n12615_), .B0(new_n27958_), .Y(new_n27959_));
  AND2X1   g25523(.A(new_n27959_), .B(new_n27914_), .Y(new_n27960_));
  AOI21X1  g25524(.A0(new_n27960_), .A1(pi1091), .B0(pi0254), .Y(new_n27961_));
  OAI21X1  g25525(.A0(new_n27961_), .A1(new_n27957_), .B0(new_n26778_), .Y(new_n27962_));
  NAND2X1  g25526(.A(new_n27962_), .B(new_n6520_), .Y(new_n27963_));
  OAI21X1  g25527(.A0(new_n26880_), .A1(pi0211), .B0(new_n27819_), .Y(new_n27964_));
  AND2X1   g25528(.A(new_n26689_), .B(new_n23539_), .Y(new_n27965_));
  INVX1    g25529(.A(new_n27965_), .Y(new_n27966_));
  NAND2X1  g25530(.A(new_n25474_), .B(pi1091), .Y(new_n27967_));
  AOI21X1  g25531(.A0(new_n27858_), .A1(new_n27734_), .B0(new_n26779_), .Y(new_n27968_));
  NAND4X1  g25532(.A(new_n27968_), .B(new_n27967_), .C(new_n27966_), .D(new_n27964_), .Y(new_n27969_));
  OAI21X1  g25533(.A0(new_n12494_), .A1(new_n2722_), .B0(new_n27817_), .Y(new_n27970_));
  NAND4X1  g25534(.A(new_n27970_), .B(new_n27967_), .C(new_n27792_), .D(new_n26779_), .Y(new_n27971_));
  NAND3X1  g25535(.A(new_n27971_), .B(new_n27969_), .C(pi0253), .Y(new_n27972_));
  AOI22X1  g25536(.A0(new_n5117_), .A1(new_n2436_), .B0(new_n2722_), .B1(new_n26779_), .Y(new_n27973_));
  OAI21X1  g25537(.A0(new_n27903_), .A1(new_n2722_), .B0(new_n27973_), .Y(new_n27974_));
  OAI21X1  g25538(.A0(new_n5118_), .A1(pi0057), .B0(new_n27892_), .Y(new_n27975_));
  AND2X1   g25539(.A(new_n27975_), .B(new_n27974_), .Y(new_n27976_));
  OAI21X1  g25540(.A0(new_n6520_), .A1(new_n26778_), .B0(new_n27976_), .Y(new_n27977_));
  AOI21X1  g25541(.A0(new_n27977_), .A1(new_n27972_), .B0(new_n25289_), .Y(new_n27978_));
  OAI21X1  g25542(.A0(new_n27963_), .A1(new_n27947_), .B0(new_n27978_), .Y(new_n27979_));
  NOR4X1   g25543(.A(new_n26706_), .B(new_n26704_), .C(new_n26695_), .D(pi1154), .Y(new_n27980_));
  NOR3X1   g25544(.A(new_n26720_), .B(new_n26710_), .C(pi1153), .Y(new_n27981_));
  NOR3X1   g25545(.A(new_n27981_), .B(new_n27980_), .C(new_n27760_), .Y(new_n27982_));
  OAI21X1  g25546(.A0(new_n26794_), .A1(new_n27936_), .B0(pi0219), .Y(new_n27983_));
  NOR3X1   g25547(.A(new_n27981_), .B(new_n27770_), .C(new_n27749_), .Y(new_n27984_));
  NOR4X1   g25548(.A(new_n26700_), .B(new_n26691_), .C(new_n12615_), .D(pi0299), .Y(new_n27985_));
  OR2X1    g25549(.A(new_n27985_), .B(pi0219), .Y(new_n27986_));
  OAI22X1  g25550(.A0(new_n27986_), .A1(new_n27984_), .B0(new_n27983_), .B1(new_n27982_), .Y(new_n27987_));
  AOI21X1  g25551(.A0(new_n27764_), .A1(new_n26787_), .B0(new_n27951_), .Y(new_n27988_));
  OR4X1    g25552(.A(new_n27988_), .B(new_n27941_), .C(new_n27937_), .D(new_n23539_), .Y(new_n27989_));
  NOR3X1   g25553(.A(new_n26754_), .B(new_n26716_), .C(new_n26701_), .Y(new_n27990_));
  OAI21X1  g25554(.A0(new_n26728_), .A1(pi1153), .B0(new_n27990_), .Y(new_n27991_));
  NAND2X1  g25555(.A(new_n27991_), .B(new_n12615_), .Y(new_n27992_));
  NOR2X1   g25556(.A(new_n26757_), .B(new_n26706_), .Y(new_n27993_));
  NOR2X1   g25557(.A(new_n27993_), .B(new_n12615_), .Y(new_n27994_));
  AOI21X1  g25558(.A0(new_n26702_), .A1(pi1154), .B0(new_n26698_), .Y(new_n27995_));
  OAI21X1  g25559(.A0(new_n27995_), .A1(pi0211), .B0(new_n23539_), .Y(new_n27996_));
  AOI21X1  g25560(.A0(new_n27994_), .A1(new_n27991_), .B0(new_n27996_), .Y(new_n27997_));
  AOI21X1  g25561(.A0(new_n27997_), .A1(new_n27992_), .B0(pi0254), .Y(new_n27998_));
  AOI22X1  g25562(.A0(new_n27998_), .A1(new_n27989_), .B0(new_n27987_), .B1(pi0254), .Y(new_n27999_));
  AND2X1   g25563(.A(new_n27858_), .B(new_n26836_), .Y(new_n28000_));
  AOI21X1  g25564(.A0(new_n27948_), .A1(new_n12615_), .B0(new_n8548_), .Y(new_n28001_));
  OAI21X1  g25565(.A0(new_n28000_), .A1(new_n27876_), .B0(new_n28001_), .Y(new_n28002_));
  OAI21X1  g25566(.A0(new_n25346_), .A1(new_n2722_), .B0(pi1154), .Y(new_n28003_));
  AOI21X1  g25567(.A0(new_n27864_), .A1(new_n8547_), .B0(pi1154), .Y(new_n28004_));
  NOR2X1   g25568(.A(new_n28004_), .B(pi0211), .Y(new_n28005_));
  NAND2X1  g25569(.A(new_n28005_), .B(new_n28003_), .Y(new_n28006_));
  AOI21X1  g25570(.A0(new_n28006_), .A1(new_n28002_), .B0(pi0219), .Y(new_n28007_));
  NOR2X1   g25571(.A(new_n28003_), .B(new_n8548_), .Y(new_n28008_));
  NOR3X1   g25572(.A(new_n25096_), .B(pi1153), .C(new_n2722_), .Y(new_n28009_));
  NOR3X1   g25573(.A(new_n28009_), .B(new_n27876_), .C(new_n27936_), .Y(new_n28010_));
  NOR4X1   g25574(.A(new_n28010_), .B(new_n28008_), .C(new_n28004_), .D(new_n23539_), .Y(new_n28011_));
  OR2X1    g25575(.A(new_n28011_), .B(new_n28007_), .Y(new_n28012_));
  OAI21X1  g25576(.A0(pi0219), .A1(new_n8548_), .B0(pi1091), .Y(new_n28013_));
  OAI21X1  g25577(.A0(new_n28013_), .A1(new_n25324_), .B0(new_n12615_), .Y(new_n28014_));
  OAI21X1  g25578(.A0(new_n26836_), .A1(new_n2722_), .B0(new_n12494_), .Y(new_n28015_));
  OAI21X1  g25579(.A0(new_n27870_), .A1(new_n12494_), .B0(new_n28015_), .Y(new_n28016_));
  AOI21X1  g25580(.A0(new_n25039_), .A1(new_n2953_), .B0(new_n2722_), .Y(new_n28017_));
  INVX1    g25581(.A(new_n28017_), .Y(new_n28018_));
  AOI21X1  g25582(.A0(new_n28018_), .A1(new_n28016_), .B0(new_n27885_), .Y(new_n28019_));
  OAI21X1  g25583(.A0(new_n27871_), .A1(new_n26872_), .B0(pi1154), .Y(new_n28020_));
  OAI21X1  g25584(.A0(new_n28020_), .A1(new_n28019_), .B0(new_n28014_), .Y(new_n28021_));
  AND2X1   g25585(.A(new_n12615_), .B(pi1091), .Y(new_n28022_));
  NAND2X1  g25586(.A(new_n28022_), .B(new_n25135_), .Y(new_n28023_));
  AOI21X1  g25587(.A0(new_n28023_), .A1(new_n28016_), .B0(new_n27873_), .Y(new_n28024_));
  NOR2X1   g25588(.A(new_n28024_), .B(new_n26779_), .Y(new_n28025_));
  AOI22X1  g25589(.A0(new_n28025_), .A1(new_n28021_), .B0(new_n28012_), .B1(new_n26779_), .Y(new_n28026_));
  AOI21X1  g25590(.A0(new_n28026_), .A1(new_n26778_), .B0(po1038), .Y(new_n28027_));
  OAI21X1  g25591(.A0(new_n27999_), .A1(new_n26778_), .B0(new_n28027_), .Y(new_n28028_));
  OAI21X1  g25592(.A0(new_n6520_), .A1(new_n26778_), .B0(new_n27974_), .Y(new_n28029_));
  NOR2X1   g25593(.A(new_n27969_), .B(new_n27818_), .Y(new_n28030_));
  NOR2X1   g25594(.A(new_n27784_), .B(pi0219), .Y(new_n28031_));
  OAI21X1  g25595(.A0(new_n27971_), .A1(new_n28031_), .B0(pi0253), .Y(new_n28032_));
  OAI21X1  g25596(.A0(new_n28032_), .A1(new_n28030_), .B0(new_n28029_), .Y(new_n28033_));
  NAND3X1  g25597(.A(new_n28033_), .B(new_n28028_), .C(new_n25289_), .Y(new_n28034_));
  NAND3X1  g25598(.A(new_n28034_), .B(new_n27979_), .C(new_n26899_), .Y(new_n28035_));
  AND2X1   g25599(.A(new_n27974_), .B(new_n25289_), .Y(new_n28036_));
  OAI21X1  g25600(.A0(new_n28026_), .A1(po1038), .B0(new_n28036_), .Y(new_n28037_));
  OR4X1    g25601(.A(new_n27961_), .B(new_n27957_), .C(new_n5118_), .D(pi0057), .Y(new_n28038_));
  AND2X1   g25602(.A(new_n27976_), .B(pi1152), .Y(new_n28039_));
  AOI21X1  g25603(.A0(new_n28039_), .A1(new_n28038_), .B0(new_n26899_), .Y(new_n28040_));
  AOI21X1  g25604(.A0(new_n28040_), .A1(new_n28037_), .B0(pi0230), .Y(new_n28041_));
  AOI22X1  g25605(.A0(new_n28041_), .A1(new_n28035_), .B0(new_n27919_), .B1(pi0230), .Y(po0411));
  MX2X1    g25606(.A(pi1049), .B(pi1036), .S0(pi0200), .Y(new_n28043_));
  MX2X1    g25607(.A(new_n28043_), .B(pi0255), .S0(new_n27694_), .Y(po0412));
  MX2X1    g25608(.A(pi1048), .B(pi1070), .S0(pi0200), .Y(new_n28045_));
  MX2X1    g25609(.A(new_n28045_), .B(pi0256), .S0(new_n27694_), .Y(po0413));
  MX2X1    g25610(.A(pi1084), .B(pi1065), .S0(pi0200), .Y(new_n28047_));
  MX2X1    g25611(.A(new_n28047_), .B(pi0257), .S0(new_n27694_), .Y(po0414));
  MX2X1    g25612(.A(pi1072), .B(pi1062), .S0(pi0200), .Y(new_n28049_));
  MX2X1    g25613(.A(new_n28049_), .B(pi0258), .S0(new_n27694_), .Y(po0415));
  MX2X1    g25614(.A(pi1059), .B(pi1069), .S0(pi0200), .Y(new_n28051_));
  MX2X1    g25615(.A(new_n28051_), .B(pi0259), .S0(new_n27694_), .Y(po0416));
  INVX1    g25616(.A(pi1044), .Y(new_n28053_));
  AOI21X1  g25617(.A0(pi1067), .A1(pi0200), .B0(pi0199), .Y(new_n28054_));
  OAI21X1  g25618(.A0(new_n28053_), .A1(pi0200), .B0(new_n28054_), .Y(new_n28055_));
  MX2X1    g25619(.A(new_n28055_), .B(pi0260), .S0(new_n27694_), .Y(po0417));
  INVX1    g25620(.A(pi1037), .Y(new_n28057_));
  AOI21X1  g25621(.A0(pi1040), .A1(pi0200), .B0(pi0199), .Y(new_n28058_));
  OAI21X1  g25622(.A0(new_n28057_), .A1(pi0200), .B0(new_n28058_), .Y(new_n28059_));
  MX2X1    g25623(.A(new_n28059_), .B(pi0261), .S0(new_n27694_), .Y(po0418));
  MX2X1    g25624(.A(new_n3706_), .B(pi0262), .S0(new_n2756_), .Y(new_n28061_));
  OR2X1    g25625(.A(new_n28061_), .B(pi0228), .Y(new_n28062_));
  AOI21X1  g25626(.A0(pi0262), .A1(pi0123), .B0(new_n3013_), .Y(new_n28063_));
  OAI21X1  g25627(.A0(pi1142), .A1(pi0123), .B0(new_n28063_), .Y(new_n28064_));
  AND2X1   g25628(.A(new_n28064_), .B(new_n28062_), .Y(new_n28065_));
  INVX1    g25629(.A(new_n28065_), .Y(new_n28066_));
  INVX1    g25630(.A(new_n26603_), .Y(new_n28067_));
  INVX1    g25631(.A(pi0123), .Y(new_n28068_));
  MX2X1    g25632(.A(pi1093), .B(new_n28068_), .S0(pi0228), .Y(new_n28069_));
  OAI22X1  g25633(.A0(new_n28069_), .A1(pi0262), .B0(new_n28067_), .B1(new_n2953_), .Y(new_n28070_));
  AOI21X1  g25634(.A0(new_n28069_), .A1(pi0199), .B0(new_n25666_), .Y(new_n28071_));
  OAI21X1  g25635(.A0(new_n28071_), .A1(new_n28070_), .B0(new_n28066_), .Y(new_n28072_));
  NOR3X1   g25636(.A(new_n28069_), .B(pi0262), .C(pi0207), .Y(new_n28073_));
  OAI22X1  g25637(.A0(new_n28073_), .A1(pi0208), .B0(new_n28067_), .B1(new_n2953_), .Y(new_n28074_));
  AND2X1   g25638(.A(new_n28074_), .B(new_n28072_), .Y(new_n28075_));
  INVX1    g25639(.A(new_n28069_), .Y(new_n28076_));
  OAI21X1  g25640(.A0(new_n28076_), .A1(new_n25851_), .B0(new_n2953_), .Y(new_n28077_));
  OAI21X1  g25641(.A0(new_n28077_), .A1(new_n28065_), .B0(pi0208), .Y(new_n28078_));
  AOI21X1  g25642(.A0(new_n28070_), .A1(pi0299), .B0(new_n28078_), .Y(new_n28079_));
  OR2X1    g25643(.A(new_n28079_), .B(po1038), .Y(new_n28080_));
  AOI21X1  g25644(.A0(new_n28064_), .A1(new_n28062_), .B0(new_n6520_), .Y(new_n28081_));
  OAI21X1  g25645(.A0(new_n28076_), .A1(new_n26603_), .B0(new_n28081_), .Y(new_n28082_));
  OAI21X1  g25646(.A0(new_n28080_), .A1(new_n28075_), .B0(new_n28082_), .Y(po0419));
  AND2X1   g25647(.A(pi0254), .B(pi0253), .Y(new_n28084_));
  AND2X1   g25648(.A(new_n28084_), .B(pi0267), .Y(new_n28085_));
  INVX1    g25649(.A(new_n28085_), .Y(new_n28086_));
  NOR3X1   g25650(.A(new_n26706_), .B(new_n26698_), .C(pi1155), .Y(new_n28087_));
  NOR3X1   g25651(.A(new_n28087_), .B(new_n26717_), .C(new_n12615_), .Y(new_n28088_));
  AOI21X1  g25652(.A0(new_n26728_), .A1(new_n12591_), .B0(pi1154), .Y(new_n28089_));
  OR4X1    g25653(.A(new_n26754_), .B(new_n26716_), .C(new_n26701_), .D(new_n12591_), .Y(new_n28090_));
  NAND2X1  g25654(.A(new_n28090_), .B(new_n28089_), .Y(new_n28091_));
  NOR3X1   g25655(.A(new_n26716_), .B(new_n26706_), .C(pi1155), .Y(new_n28092_));
  NOR3X1   g25656(.A(new_n28092_), .B(new_n26717_), .C(new_n12615_), .Y(new_n28093_));
  OAI21X1  g25657(.A0(new_n28093_), .A1(new_n27985_), .B0(new_n12684_), .Y(new_n28094_));
  AOI22X1  g25658(.A0(new_n28094_), .A1(new_n28091_), .B0(new_n27993_), .B1(pi1156), .Y(new_n28095_));
  OAI21X1  g25659(.A0(new_n28095_), .A1(new_n28088_), .B0(pi0211), .Y(new_n28096_));
  NOR4X1   g25660(.A(new_n26754_), .B(new_n26701_), .C(new_n26698_), .D(new_n12591_), .Y(new_n28097_));
  NOR3X1   g25661(.A(new_n28097_), .B(new_n26742_), .C(pi1154), .Y(new_n28098_));
  OR4X1    g25662(.A(new_n28098_), .B(new_n28093_), .C(new_n27985_), .D(pi1156), .Y(new_n28099_));
  INVX1    g25663(.A(new_n28093_), .Y(new_n28100_));
  OAI21X1  g25664(.A0(new_n26757_), .A1(new_n26706_), .B0(new_n28098_), .Y(new_n28101_));
  AND2X1   g25665(.A(new_n28101_), .B(pi1156), .Y(new_n28102_));
  AOI21X1  g25666(.A0(new_n28102_), .A1(new_n28100_), .B0(pi0211), .Y(new_n28103_));
  AOI21X1  g25667(.A0(new_n28103_), .A1(new_n28099_), .B0(pi0219), .Y(new_n28104_));
  INVX1    g25668(.A(pi0263), .Y(new_n28105_));
  INVX1    g25669(.A(new_n26754_), .Y(new_n28106_));
  AOI21X1  g25670(.A0(new_n26711_), .A1(new_n26709_), .B0(new_n26812_), .Y(new_n28107_));
  MX2X1    g25671(.A(new_n26708_), .B(new_n12615_), .S0(new_n26702_), .Y(new_n28108_));
  NOR2X1   g25672(.A(new_n28108_), .B(new_n28107_), .Y(new_n28109_));
  AOI21X1  g25673(.A0(new_n28109_), .A1(new_n28106_), .B0(pi1156), .Y(new_n28110_));
  NOR2X1   g25674(.A(new_n27924_), .B(new_n12591_), .Y(new_n28111_));
  NOR2X1   g25675(.A(new_n27769_), .B(new_n26706_), .Y(new_n28112_));
  OAI21X1  g25676(.A0(new_n28112_), .A1(pi1155), .B0(new_n12615_), .Y(new_n28113_));
  NOR2X1   g25677(.A(new_n28113_), .B(new_n28111_), .Y(new_n28114_));
  AND2X1   g25678(.A(pi1156), .B(new_n8548_), .Y(new_n28115_));
  OAI21X1  g25679(.A0(new_n28107_), .A1(new_n12615_), .B0(new_n28115_), .Y(new_n28116_));
  NOR2X1   g25680(.A(new_n28116_), .B(new_n28114_), .Y(new_n28117_));
  AND2X1   g25681(.A(pi1156), .B(pi0211), .Y(new_n28118_));
  INVX1    g25682(.A(new_n28118_), .Y(new_n28119_));
  OAI21X1  g25683(.A0(new_n28109_), .A1(new_n28119_), .B0(pi0219), .Y(new_n28120_));
  NOR3X1   g25684(.A(new_n28120_), .B(new_n28117_), .C(new_n28110_), .Y(new_n28121_));
  OR2X1    g25685(.A(new_n28121_), .B(new_n28105_), .Y(new_n28122_));
  AOI21X1  g25686(.A0(new_n28104_), .A1(new_n28096_), .B0(new_n28122_), .Y(new_n28123_));
  NOR4X1   g25687(.A(new_n27767_), .B(new_n26755_), .C(pi1155), .D(pi1091), .Y(new_n28124_));
  INVX1    g25688(.A(new_n28124_), .Y(new_n28125_));
  AOI21X1  g25689(.A0(new_n27750_), .A1(pi1155), .B0(pi1154), .Y(new_n28126_));
  AOI21X1  g25690(.A0(new_n28126_), .A1(new_n28125_), .B0(pi1156), .Y(new_n28127_));
  INVX1    g25691(.A(new_n28127_), .Y(new_n28128_));
  OR2X1    g25692(.A(new_n26702_), .B(new_n26698_), .Y(new_n28129_));
  AOI21X1  g25693(.A0(new_n26757_), .A1(pi1155), .B0(new_n12615_), .Y(new_n28130_));
  INVX1    g25694(.A(new_n28130_), .Y(new_n28131_));
  NOR2X1   g25695(.A(new_n28131_), .B(new_n28129_), .Y(new_n28132_));
  NOR3X1   g25696(.A(new_n27767_), .B(pi1155), .C(pi1091), .Y(new_n28133_));
  INVX1    g25697(.A(new_n28133_), .Y(new_n28134_));
  AOI21X1  g25698(.A0(new_n26789_), .A1(pi1155), .B0(pi1154), .Y(new_n28135_));
  AND2X1   g25699(.A(new_n28135_), .B(new_n28134_), .Y(new_n28136_));
  OR2X1    g25700(.A(new_n28136_), .B(new_n28132_), .Y(new_n28137_));
  OAI21X1  g25701(.A0(new_n26689_), .A1(new_n2953_), .B0(new_n27806_), .Y(new_n28138_));
  OAI21X1  g25702(.A0(new_n27759_), .A1(pi1155), .B0(new_n28138_), .Y(new_n28139_));
  AOI21X1  g25703(.A0(new_n28139_), .A1(new_n12615_), .B0(new_n12684_), .Y(new_n28140_));
  OAI21X1  g25704(.A0(new_n26685_), .A1(pi1091), .B0(new_n8009_), .Y(new_n28141_));
  AOI22X1  g25705(.A0(new_n28135_), .A1(new_n26726_), .B0(new_n28132_), .B1(new_n28141_), .Y(new_n28142_));
  AOI21X1  g25706(.A0(new_n28142_), .A1(new_n28140_), .B0(pi0211), .Y(new_n28143_));
  OAI21X1  g25707(.A0(new_n28137_), .A1(new_n28128_), .B0(new_n28143_), .Y(new_n28144_));
  OAI21X1  g25708(.A0(new_n28131_), .A1(new_n27751_), .B0(new_n28140_), .Y(new_n28145_));
  NAND2X1  g25709(.A(new_n28130_), .B(new_n27756_), .Y(new_n28146_));
  AOI21X1  g25710(.A0(new_n28146_), .A1(new_n28127_), .B0(new_n8548_), .Y(new_n28147_));
  AOI21X1  g25711(.A0(new_n28147_), .A1(new_n28145_), .B0(pi0219), .Y(new_n28148_));
  INVX1    g25712(.A(new_n26701_), .Y(new_n28149_));
  NAND2X1  g25713(.A(new_n26820_), .B(pi1154), .Y(new_n28150_));
  AOI21X1  g25714(.A0(new_n26697_), .A1(pi1155), .B0(new_n28150_), .Y(new_n28151_));
  AOI22X1  g25715(.A0(new_n28151_), .A1(new_n28149_), .B0(new_n28135_), .B1(new_n26726_), .Y(new_n28152_));
  NOR2X1   g25716(.A(new_n28152_), .B(new_n28119_), .Y(new_n28153_));
  AOI21X1  g25717(.A0(new_n28135_), .A1(new_n28134_), .B0(new_n28151_), .Y(new_n28154_));
  OAI21X1  g25718(.A0(new_n27768_), .A1(pi1154), .B0(new_n26783_), .Y(new_n28155_));
  INVX1    g25719(.A(new_n28115_), .Y(new_n28156_));
  AOI21X1  g25720(.A0(new_n26697_), .A1(pi1155), .B0(new_n28156_), .Y(new_n28157_));
  AOI21X1  g25721(.A0(new_n28157_), .A1(new_n28155_), .B0(new_n23539_), .Y(new_n28158_));
  OAI21X1  g25722(.A0(new_n28154_), .A1(pi1156), .B0(new_n28158_), .Y(new_n28159_));
  OAI21X1  g25723(.A0(new_n28159_), .A1(new_n28153_), .B0(new_n28105_), .Y(new_n28160_));
  AOI21X1  g25724(.A0(new_n28148_), .A1(new_n28144_), .B0(new_n28160_), .Y(new_n28161_));
  NOR3X1   g25725(.A(new_n28161_), .B(new_n28123_), .C(new_n28086_), .Y(new_n28162_));
  OAI21X1  g25726(.A0(new_n25377_), .A1(new_n12591_), .B0(new_n26856_), .Y(new_n28163_));
  OAI21X1  g25727(.A0(new_n28018_), .A1(pi1154), .B0(new_n28163_), .Y(new_n28164_));
  INVX1    g25728(.A(new_n28164_), .Y(new_n28165_));
  AOI21X1  g25729(.A0(new_n28165_), .A1(new_n26870_), .B0(new_n28119_), .Y(new_n28166_));
  OR2X1    g25730(.A(new_n12591_), .B(pi0199), .Y(new_n28167_));
  AOI21X1  g25731(.A0(new_n28167_), .A1(new_n25082_), .B0(new_n12615_), .Y(new_n28168_));
  NOR3X1   g25732(.A(new_n28168_), .B(new_n28156_), .C(new_n2722_), .Y(new_n28169_));
  OAI21X1  g25733(.A0(new_n25111_), .A1(pi1154), .B0(new_n28169_), .Y(new_n28170_));
  AOI21X1  g25734(.A0(new_n25342_), .A1(pi1154), .B0(new_n2722_), .Y(new_n28171_));
  NOR2X1   g25735(.A(new_n25059_), .B(pi1156), .Y(new_n28172_));
  AOI21X1  g25736(.A0(new_n28172_), .A1(new_n28171_), .B0(new_n23539_), .Y(new_n28173_));
  AND2X1   g25737(.A(new_n28173_), .B(new_n28170_), .Y(new_n28174_));
  INVX1    g25738(.A(new_n28174_), .Y(new_n28175_));
  OAI21X1  g25739(.A0(pi1154), .A1(pi0199), .B0(new_n25053_), .Y(new_n28176_));
  NAND2X1  g25740(.A(new_n28176_), .B(new_n27856_), .Y(new_n28177_));
  OAI22X1  g25741(.A0(new_n28177_), .A1(new_n25157_), .B0(new_n28165_), .B1(pi0211), .Y(new_n28178_));
  AND2X1   g25742(.A(new_n28178_), .B(pi1156), .Y(new_n28179_));
  OAI21X1  g25743(.A0(new_n25135_), .A1(new_n12591_), .B0(new_n28171_), .Y(new_n28180_));
  INVX1    g25744(.A(new_n28180_), .Y(new_n28181_));
  AOI21X1  g25745(.A0(new_n8132_), .A1(pi1154), .B0(new_n25059_), .Y(new_n28182_));
  AOI22X1  g25746(.A0(new_n28182_), .A1(new_n27954_), .B0(new_n28181_), .B1(pi0211), .Y(new_n28183_));
  OAI21X1  g25747(.A0(new_n28183_), .A1(pi1156), .B0(new_n23539_), .Y(new_n28184_));
  OAI22X1  g25748(.A0(new_n28184_), .A1(new_n28179_), .B0(new_n28175_), .B1(new_n28166_), .Y(new_n28185_));
  NOR2X1   g25749(.A(new_n8131_), .B(pi1155), .Y(new_n28186_));
  NOR3X1   g25750(.A(new_n28186_), .B(new_n25111_), .C(pi1154), .Y(new_n28187_));
  AOI21X1  g25751(.A0(new_n25087_), .A1(pi1155), .B0(new_n25053_), .Y(new_n28188_));
  OAI21X1  g25752(.A0(new_n28188_), .A1(new_n12615_), .B0(pi1156), .Y(new_n28189_));
  AOI21X1  g25753(.A0(new_n28181_), .A1(new_n12684_), .B0(new_n8548_), .Y(new_n28190_));
  OAI21X1  g25754(.A0(new_n28189_), .A1(new_n28187_), .B0(new_n28190_), .Y(new_n28191_));
  OAI22X1  g25755(.A0(new_n25731_), .A1(new_n25064_), .B0(new_n8131_), .B1(new_n12615_), .Y(new_n28192_));
  AOI21X1  g25756(.A0(new_n28192_), .A1(new_n8548_), .B0(pi0219), .Y(new_n28193_));
  AND2X1   g25757(.A(new_n28193_), .B(new_n28191_), .Y(new_n28194_));
  INVX1    g25758(.A(new_n28194_), .Y(new_n28195_));
  OAI21X1  g25759(.A0(new_n25062_), .A1(new_n12615_), .B0(pi1156), .Y(new_n28196_));
  AND2X1   g25760(.A(new_n28196_), .B(new_n2953_), .Y(new_n28197_));
  NOR4X1   g25761(.A(new_n25062_), .B(new_n8130_), .C(pi1154), .D(pi0299), .Y(new_n28198_));
  NOR3X1   g25762(.A(new_n28198_), .B(new_n28197_), .C(new_n25984_), .Y(new_n28199_));
  INVX1    g25763(.A(new_n28182_), .Y(new_n28200_));
  AOI21X1  g25764(.A0(new_n28197_), .A1(new_n28200_), .B0(new_n23539_), .Y(new_n28201_));
  OAI21X1  g25765(.A0(new_n28199_), .A1(new_n12684_), .B0(new_n28201_), .Y(new_n28202_));
  AND2X1   g25766(.A(pi1091), .B(pi0263), .Y(new_n28203_));
  AND2X1   g25767(.A(new_n28203_), .B(new_n28202_), .Y(new_n28204_));
  AOI22X1  g25768(.A0(new_n28204_), .A1(new_n28195_), .B0(new_n28185_), .B1(new_n28105_), .Y(new_n28205_));
  OAI21X1  g25769(.A0(new_n28205_), .A1(new_n28085_), .B0(new_n6520_), .Y(new_n28206_));
  INVX1    g25770(.A(new_n26899_), .Y(new_n28207_));
  INVX1    g25771(.A(new_n27964_), .Y(new_n28208_));
  NAND2X1  g25772(.A(new_n26680_), .B(pi0211), .Y(new_n28209_));
  MX2X1    g25773(.A(new_n28022_), .B(new_n12591_), .S0(pi0211), .Y(new_n28210_));
  AOI21X1  g25774(.A0(new_n28210_), .A1(new_n28209_), .B0(new_n26689_), .Y(new_n28211_));
  NOR2X1   g25775(.A(new_n28211_), .B(pi0219), .Y(new_n28212_));
  NOR3X1   g25776(.A(new_n28212_), .B(new_n28208_), .C(pi0263), .Y(new_n28213_));
  INVX1    g25777(.A(new_n27792_), .Y(new_n28214_));
  INVX1    g25778(.A(new_n27954_), .Y(new_n28215_));
  OAI22X1  g25779(.A0(new_n28215_), .A1(new_n12615_), .B0(new_n12591_), .B1(new_n8548_), .Y(new_n28216_));
  AOI21X1  g25780(.A0(new_n28216_), .A1(new_n28209_), .B0(new_n27816_), .Y(new_n28217_));
  NOR3X1   g25781(.A(new_n28217_), .B(new_n28214_), .C(new_n28105_), .Y(new_n28218_));
  AOI21X1  g25782(.A0(pi1156), .A1(new_n8548_), .B0(new_n23539_), .Y(new_n28219_));
  AOI21X1  g25783(.A0(new_n28219_), .A1(pi1091), .B0(new_n28086_), .Y(new_n28220_));
  OAI21X1  g25784(.A0(new_n28218_), .A1(new_n28213_), .B0(new_n28220_), .Y(new_n28221_));
  AOI21X1  g25785(.A0(pi1155), .A1(pi0211), .B0(pi0219), .Y(new_n28222_));
  AOI21X1  g25786(.A0(new_n28222_), .A1(new_n27936_), .B0(new_n28219_), .Y(new_n28223_));
  MX2X1    g25787(.A(new_n28223_), .B(new_n28105_), .S0(new_n2722_), .Y(new_n28224_));
  AOI21X1  g25788(.A0(new_n28224_), .A1(new_n28086_), .B0(new_n6520_), .Y(new_n28225_));
  AOI21X1  g25789(.A0(new_n28225_), .A1(new_n28221_), .B0(new_n28207_), .Y(new_n28226_));
  OAI21X1  g25790(.A0(new_n28206_), .A1(new_n28162_), .B0(new_n28226_), .Y(new_n28227_));
  OAI21X1  g25791(.A0(new_n28224_), .A1(new_n6520_), .B0(new_n28207_), .Y(new_n28228_));
  AOI21X1  g25792(.A0(new_n28205_), .A1(new_n6520_), .B0(new_n28228_), .Y(new_n28229_));
  NOR2X1   g25793(.A(new_n28229_), .B(pi0230), .Y(new_n28230_));
  INVX1    g25794(.A(new_n28193_), .Y(new_n28231_));
  NOR3X1   g25795(.A(new_n25064_), .B(new_n25060_), .C(new_n8503_), .Y(new_n28232_));
  NOR3X1   g25796(.A(new_n25450_), .B(new_n25062_), .C(pi0299), .Y(new_n28233_));
  OAI21X1  g25797(.A0(new_n28232_), .A1(pi1156), .B0(new_n28233_), .Y(new_n28234_));
  AOI21X1  g25798(.A0(new_n28234_), .A1(new_n25100_), .B0(new_n8548_), .Y(new_n28235_));
  AOI21X1  g25799(.A0(new_n25984_), .A1(pi1156), .B0(new_n23539_), .Y(new_n28236_));
  AOI21X1  g25800(.A0(new_n28236_), .A1(new_n28234_), .B0(po1038), .Y(new_n28237_));
  OAI21X1  g25801(.A0(new_n28235_), .A1(new_n28231_), .B0(new_n28237_), .Y(new_n28238_));
  AOI21X1  g25802(.A0(new_n28223_), .A1(po1038), .B0(new_n24954_), .Y(new_n28239_));
  AOI22X1  g25803(.A0(new_n28239_), .A1(new_n28238_), .B0(new_n28230_), .B1(new_n28227_), .Y(po0420));
  NOR2X1   g25804(.A(new_n26684_), .B(new_n7734_), .Y(new_n28241_));
  INVX1    g25805(.A(new_n28241_), .Y(new_n28242_));
  AOI21X1  g25806(.A0(new_n28242_), .A1(pi0264), .B0(pi1091), .Y(new_n28243_));
  OAI21X1  g25807(.A0(new_n28242_), .A1(pi0796), .B0(new_n28243_), .Y(new_n28244_));
  NAND2X1  g25808(.A(pi1141), .B(pi1091), .Y(new_n28245_));
  AND2X1   g25809(.A(new_n28245_), .B(new_n28244_), .Y(new_n28246_));
  AND2X1   g25810(.A(pi1142), .B(pi1091), .Y(new_n28247_));
  INVX1    g25811(.A(new_n28247_), .Y(new_n28248_));
  NAND2X1  g25812(.A(new_n28248_), .B(new_n28244_), .Y(new_n28249_));
  AOI21X1  g25813(.A0(new_n28249_), .A1(pi0200), .B0(pi0199), .Y(new_n28250_));
  OAI21X1  g25814(.A0(new_n28246_), .A1(pi0200), .B0(new_n28250_), .Y(new_n28251_));
  INVX1    g25815(.A(new_n26675_), .Y(new_n28252_));
  AOI21X1  g25816(.A0(new_n28252_), .A1(pi0264), .B0(pi1091), .Y(new_n28253_));
  OAI21X1  g25817(.A0(new_n28252_), .A1(pi0796), .B0(new_n28253_), .Y(new_n28254_));
  AND2X1   g25818(.A(pi1143), .B(pi1091), .Y(new_n28255_));
  AOI21X1  g25819(.A0(new_n28255_), .A1(new_n8009_), .B0(new_n7941_), .Y(new_n28256_));
  AOI21X1  g25820(.A0(new_n28256_), .A1(new_n28254_), .B0(new_n11777_), .Y(new_n28257_));
  AOI21X1  g25821(.A0(new_n28249_), .A1(pi0211), .B0(pi0219), .Y(new_n28258_));
  OAI21X1  g25822(.A0(new_n28246_), .A1(pi0211), .B0(new_n28258_), .Y(new_n28259_));
  AOI21X1  g25823(.A0(new_n27954_), .A1(new_n24964_), .B0(new_n23539_), .Y(new_n28260_));
  AOI21X1  g25824(.A0(new_n28260_), .A1(new_n28254_), .B0(new_n11776_), .Y(new_n28261_));
  AOI22X1  g25825(.A0(new_n28261_), .A1(new_n28259_), .B0(new_n28257_), .B1(new_n28251_), .Y(new_n28262_));
  AOI21X1  g25826(.A0(pi1142), .A1(pi0211), .B0(pi0219), .Y(new_n28263_));
  OAI21X1  g25827(.A0(new_n3847_), .A1(pi0211), .B0(new_n28263_), .Y(new_n28264_));
  AOI22X1  g25828(.A0(new_n28264_), .A1(new_n25652_), .B0(new_n6520_), .B1(new_n2953_), .Y(new_n28265_));
  OR2X1    g25829(.A(new_n3847_), .B(pi0199), .Y(new_n28266_));
  AOI21X1  g25830(.A0(new_n28266_), .A1(new_n25634_), .B0(new_n24976_), .Y(new_n28267_));
  OAI21X1  g25831(.A0(new_n28267_), .A1(new_n11777_), .B0(pi0230), .Y(new_n28268_));
  OAI22X1  g25832(.A0(new_n28268_), .A1(new_n28265_), .B0(new_n28262_), .B1(pi0230), .Y(po0421));
  AOI21X1  g25833(.A0(new_n28242_), .A1(pi0265), .B0(pi1091), .Y(new_n28270_));
  OAI21X1  g25834(.A0(new_n28242_), .A1(pi0819), .B0(new_n28270_), .Y(new_n28271_));
  AND2X1   g25835(.A(new_n28271_), .B(new_n28248_), .Y(new_n28272_));
  OAI21X1  g25836(.A0(new_n3495_), .A1(new_n2722_), .B0(new_n28271_), .Y(new_n28273_));
  AOI21X1  g25837(.A0(new_n28273_), .A1(pi0200), .B0(pi0199), .Y(new_n28274_));
  OAI21X1  g25838(.A0(new_n28272_), .A1(pi0200), .B0(new_n28274_), .Y(new_n28275_));
  AOI21X1  g25839(.A0(new_n28252_), .A1(pi0265), .B0(pi1091), .Y(new_n28276_));
  OAI21X1  g25840(.A0(new_n28252_), .A1(pi0819), .B0(new_n28276_), .Y(new_n28277_));
  AND2X1   g25841(.A(pi1144), .B(pi1091), .Y(new_n28278_));
  AOI21X1  g25842(.A0(new_n28278_), .A1(new_n8009_), .B0(new_n7941_), .Y(new_n28279_));
  AOI21X1  g25843(.A0(new_n28279_), .A1(new_n28277_), .B0(new_n11777_), .Y(new_n28280_));
  AOI21X1  g25844(.A0(new_n28273_), .A1(pi0211), .B0(pi0219), .Y(new_n28281_));
  OAI21X1  g25845(.A0(new_n28272_), .A1(pi0211), .B0(new_n28281_), .Y(new_n28282_));
  AOI21X1  g25846(.A0(pi1091), .A1(new_n8548_), .B0(new_n23539_), .Y(new_n28283_));
  OR2X1    g25847(.A(new_n28283_), .B(new_n26621_), .Y(new_n28284_));
  AOI21X1  g25848(.A0(new_n28284_), .A1(new_n28277_), .B0(new_n11776_), .Y(new_n28285_));
  AOI22X1  g25849(.A0(new_n28285_), .A1(new_n28282_), .B0(new_n28280_), .B1(new_n28275_), .Y(new_n28286_));
  INVX1    g25850(.A(new_n26621_), .Y(new_n28287_));
  AOI21X1  g25851(.A0(pi1143), .A1(pi0211), .B0(pi0219), .Y(new_n28288_));
  OAI21X1  g25852(.A0(new_n3706_), .A1(pi0211), .B0(new_n28288_), .Y(new_n28289_));
  AOI21X1  g25853(.A0(new_n28289_), .A1(new_n28287_), .B0(new_n11776_), .Y(new_n28290_));
  OR2X1    g25854(.A(new_n3706_), .B(pi0199), .Y(new_n28291_));
  AOI21X1  g25855(.A0(new_n26624_), .A1(new_n28291_), .B0(new_n24971_), .Y(new_n28292_));
  OAI21X1  g25856(.A0(new_n28292_), .A1(new_n11777_), .B0(pi0230), .Y(new_n28293_));
  OAI22X1  g25857(.A0(new_n28293_), .A1(new_n28290_), .B0(new_n28286_), .B1(pi0230), .Y(po0422));
  AND2X1   g25858(.A(pi1136), .B(new_n8548_), .Y(new_n28295_));
  OAI22X1  g25859(.A0(new_n28295_), .A1(new_n23539_), .B0(pi1135), .B1(new_n8548_), .Y(new_n28296_));
  NOR2X1   g25860(.A(new_n28296_), .B(new_n8075_), .Y(new_n28297_));
  AOI21X1  g25861(.A0(pi1135), .A1(new_n7941_), .B0(new_n8009_), .Y(new_n28298_));
  AOI21X1  g25862(.A0(pi1136), .A1(pi0199), .B0(pi0200), .Y(new_n28299_));
  NOR3X1   g25863(.A(new_n28299_), .B(new_n28298_), .C(pi0299), .Y(new_n28300_));
  AOI21X1  g25864(.A0(new_n28297_), .A1(pi0299), .B0(new_n28300_), .Y(new_n28301_));
  AOI21X1  g25865(.A0(new_n28297_), .A1(po1038), .B0(new_n24954_), .Y(new_n28302_));
  OAI21X1  g25866(.A0(new_n28301_), .A1(po1038), .B0(new_n28302_), .Y(new_n28303_));
  INVX1    g25867(.A(pi0948), .Y(new_n28304_));
  AOI21X1  g25868(.A0(new_n28241_), .A1(new_n28304_), .B0(pi1091), .Y(new_n28305_));
  OAI21X1  g25869(.A0(new_n28241_), .A1(pi0266), .B0(new_n28305_), .Y(new_n28306_));
  AND2X1   g25870(.A(new_n28306_), .B(new_n7941_), .Y(new_n28307_));
  NAND2X1  g25871(.A(pi1136), .B(pi1091), .Y(new_n28308_));
  AOI21X1  g25872(.A0(new_n26675_), .A1(new_n28304_), .B0(pi1091), .Y(new_n28309_));
  OAI21X1  g25873(.A0(new_n26675_), .A1(pi0266), .B0(new_n28309_), .Y(new_n28310_));
  AND2X1   g25874(.A(new_n28310_), .B(pi0199), .Y(new_n28311_));
  AOI21X1  g25875(.A0(new_n28311_), .A1(new_n28308_), .B0(new_n28307_), .Y(new_n28312_));
  INVX1    g25876(.A(pi1135), .Y(new_n28313_));
  OAI21X1  g25877(.A0(new_n28313_), .A1(new_n2722_), .B0(new_n28307_), .Y(new_n28314_));
  AOI21X1  g25878(.A0(new_n28310_), .A1(pi0199), .B0(new_n8009_), .Y(new_n28315_));
  AOI22X1  g25879(.A0(new_n28315_), .A1(new_n28314_), .B0(new_n28312_), .B1(new_n8009_), .Y(new_n28316_));
  AOI21X1  g25880(.A0(new_n28295_), .A1(new_n27954_), .B0(new_n23539_), .Y(new_n28317_));
  AOI21X1  g25881(.A0(new_n28317_), .A1(new_n28310_), .B0(new_n11776_), .Y(new_n28318_));
  AND2X1   g25882(.A(new_n28306_), .B(new_n23539_), .Y(new_n28319_));
  OAI21X1  g25883(.A0(new_n27857_), .A1(new_n28313_), .B0(new_n28319_), .Y(new_n28320_));
  AOI21X1  g25884(.A0(new_n28320_), .A1(new_n28318_), .B0(pi0230), .Y(new_n28321_));
  OAI21X1  g25885(.A0(new_n28316_), .A1(new_n11777_), .B0(new_n28321_), .Y(new_n28322_));
  AOI21X1  g25886(.A0(new_n28322_), .A1(new_n28303_), .B0(pi1134), .Y(new_n28323_));
  NOR3X1   g25887(.A(pi1136), .B(pi0200), .C(new_n7941_), .Y(new_n28324_));
  NOR4X1   g25888(.A(new_n28324_), .B(new_n28298_), .C(po1038), .D(pi0299), .Y(new_n28325_));
  OAI21X1  g25889(.A0(new_n28296_), .A1(new_n11776_), .B0(pi0230), .Y(new_n28326_));
  AND2X1   g25890(.A(new_n28315_), .B(new_n28314_), .Y(new_n28327_));
  INVX1    g25891(.A(new_n28327_), .Y(new_n28328_));
  AND2X1   g25892(.A(pi1091), .B(new_n7941_), .Y(new_n28329_));
  OAI21X1  g25893(.A0(new_n28329_), .A1(new_n28312_), .B0(new_n8009_), .Y(new_n28330_));
  AOI21X1  g25894(.A0(new_n28330_), .A1(new_n28328_), .B0(new_n11777_), .Y(new_n28331_));
  INVX1    g25895(.A(new_n28318_), .Y(new_n28332_));
  OAI21X1  g25896(.A0(pi1135), .A1(new_n8548_), .B0(pi1091), .Y(new_n28333_));
  AND2X1   g25897(.A(new_n28333_), .B(new_n28319_), .Y(new_n28334_));
  OAI21X1  g25898(.A0(new_n28334_), .A1(new_n28332_), .B0(new_n24954_), .Y(new_n28335_));
  OAI22X1  g25899(.A0(new_n28335_), .A1(new_n28331_), .B0(new_n28326_), .B1(new_n28325_), .Y(new_n28336_));
  AOI21X1  g25900(.A0(new_n28336_), .A1(pi1134), .B0(new_n28323_), .Y(po0423));
  INVX1    g25901(.A(new_n28084_), .Y(new_n28338_));
  NOR3X1   g25902(.A(new_n27939_), .B(new_n27768_), .C(new_n26706_), .Y(new_n28339_));
  INVX1    g25903(.A(new_n28339_), .Y(new_n28340_));
  NAND3X1  g25904(.A(new_n28340_), .B(new_n26808_), .C(new_n12615_), .Y(new_n28341_));
  OR4X1    g25905(.A(new_n27943_), .B(new_n26787_), .C(new_n12591_), .D(new_n12615_), .Y(new_n28342_));
  AOI21X1  g25906(.A0(new_n28342_), .A1(new_n28341_), .B0(new_n8548_), .Y(new_n28343_));
  NOR3X1   g25907(.A(new_n26710_), .B(new_n26706_), .C(new_n12494_), .Y(new_n28344_));
  OR4X1    g25908(.A(new_n28344_), .B(new_n28112_), .C(new_n12591_), .D(pi0211), .Y(new_n28345_));
  OR2X1    g25909(.A(new_n28345_), .B(new_n27925_), .Y(new_n28346_));
  OR4X1    g25910(.A(new_n26754_), .B(new_n26704_), .C(new_n26701_), .D(new_n12615_), .Y(new_n28347_));
  NAND3X1  g25911(.A(new_n28347_), .B(new_n28340_), .C(new_n12591_), .Y(new_n28348_));
  NAND3X1  g25912(.A(new_n28348_), .B(new_n28346_), .C(new_n26780_), .Y(new_n28349_));
  AOI21X1  g25913(.A0(new_n27777_), .A1(new_n27757_), .B0(new_n26789_), .Y(new_n28350_));
  NOR2X1   g25914(.A(new_n28350_), .B(new_n12615_), .Y(new_n28351_));
  OR2X1    g25915(.A(new_n26820_), .B(pi1154), .Y(new_n28352_));
  OAI21X1  g25916(.A0(new_n28352_), .A1(new_n27840_), .B0(new_n12591_), .Y(new_n28353_));
  NOR2X1   g25917(.A(new_n28353_), .B(new_n28351_), .Y(new_n28354_));
  AOI21X1  g25918(.A0(new_n27760_), .A1(new_n27758_), .B0(new_n26794_), .Y(new_n28355_));
  AND2X1   g25919(.A(new_n27828_), .B(pi1155), .Y(new_n28356_));
  OAI21X1  g25920(.A0(new_n27768_), .A1(pi1154), .B0(new_n26697_), .Y(new_n28357_));
  NAND2X1  g25921(.A(new_n28357_), .B(new_n28356_), .Y(new_n28358_));
  OAI21X1  g25922(.A0(new_n28358_), .A1(new_n28355_), .B0(pi0267), .Y(new_n28359_));
  OAI22X1  g25923(.A0(new_n28359_), .A1(new_n28354_), .B0(new_n28349_), .B1(new_n28343_), .Y(new_n28360_));
  NAND2X1  g25924(.A(new_n28360_), .B(pi0219), .Y(new_n28361_));
  OAI21X1  g25925(.A0(new_n28350_), .A1(new_n27750_), .B0(new_n28111_), .Y(new_n28362_));
  OAI21X1  g25926(.A0(new_n27753_), .A1(pi1154), .B0(pi1155), .Y(new_n28363_));
  AOI22X1  g25927(.A0(new_n28363_), .A1(new_n26735_), .B0(new_n28362_), .B1(pi1154), .Y(new_n28364_));
  NOR3X1   g25928(.A(new_n28339_), .B(new_n27990_), .C(pi1155), .Y(new_n28365_));
  NOR3X1   g25929(.A(new_n28365_), .B(new_n28364_), .C(new_n8548_), .Y(new_n28366_));
  OAI21X1  g25930(.A0(new_n26755_), .A1(new_n12494_), .B0(new_n12591_), .Y(new_n28367_));
  NOR3X1   g25931(.A(new_n28367_), .B(new_n27837_), .C(new_n26706_), .Y(new_n28368_));
  OR2X1    g25932(.A(new_n28344_), .B(new_n27993_), .Y(new_n28369_));
  AND2X1   g25933(.A(new_n28369_), .B(pi1155), .Y(new_n28370_));
  NOR3X1   g25934(.A(new_n28370_), .B(new_n28368_), .C(pi1154), .Y(new_n28371_));
  AOI21X1  g25935(.A0(new_n28106_), .A1(new_n26764_), .B0(pi1153), .Y(new_n28372_));
  NOR2X1   g25936(.A(new_n28097_), .B(new_n12615_), .Y(new_n28373_));
  OAI21X1  g25937(.A0(new_n28372_), .A1(new_n28367_), .B0(new_n28373_), .Y(new_n28374_));
  OAI21X1  g25938(.A0(new_n28374_), .A1(new_n28370_), .B0(new_n8548_), .Y(new_n28375_));
  OAI21X1  g25939(.A0(new_n28375_), .A1(new_n28371_), .B0(new_n26780_), .Y(new_n28376_));
  OAI21X1  g25940(.A0(new_n26766_), .A1(pi1153), .B0(new_n26757_), .Y(new_n28377_));
  NOR3X1   g25941(.A(new_n26698_), .B(new_n26697_), .C(pi1155), .Y(new_n28378_));
  INVX1    g25942(.A(new_n28356_), .Y(new_n28379_));
  OAI21X1  g25943(.A0(new_n28379_), .A1(new_n28138_), .B0(pi1154), .Y(new_n28380_));
  AOI21X1  g25944(.A0(new_n28378_), .A1(new_n28377_), .B0(new_n28380_), .Y(new_n28381_));
  NOR2X1   g25945(.A(new_n27776_), .B(pi1154), .Y(new_n28382_));
  AOI21X1  g25946(.A0(new_n28382_), .A1(new_n28129_), .B0(pi1155), .Y(new_n28383_));
  NOR4X1   g25947(.A(new_n28383_), .B(new_n27776_), .C(new_n26736_), .D(pi1154), .Y(new_n28384_));
  OAI21X1  g25948(.A0(new_n28384_), .A1(new_n28381_), .B0(pi0211), .Y(new_n28385_));
  OAI21X1  g25949(.A0(new_n28377_), .A1(new_n12615_), .B0(new_n28383_), .Y(new_n28386_));
  OR2X1    g25950(.A(new_n27981_), .B(new_n26764_), .Y(new_n28387_));
  AOI21X1  g25951(.A0(new_n26697_), .A1(pi1154), .B0(new_n12591_), .Y(new_n28388_));
  AOI21X1  g25952(.A0(new_n28388_), .A1(new_n28387_), .B0(pi0211), .Y(new_n28389_));
  AOI21X1  g25953(.A0(new_n28389_), .A1(new_n28386_), .B0(new_n26780_), .Y(new_n28390_));
  AOI21X1  g25954(.A0(new_n28390_), .A1(new_n28385_), .B0(pi0219), .Y(new_n28391_));
  OAI21X1  g25955(.A0(new_n28376_), .A1(new_n28366_), .B0(new_n28391_), .Y(new_n28392_));
  AOI21X1  g25956(.A0(new_n28392_), .A1(new_n28361_), .B0(new_n28338_), .Y(new_n28393_));
  AOI21X1  g25957(.A0(new_n26857_), .A1(pi1153), .B0(new_n12591_), .Y(new_n28394_));
  NOR3X1   g25958(.A(new_n25415_), .B(pi1155), .C(new_n2722_), .Y(new_n28395_));
  AOI21X1  g25959(.A0(new_n28394_), .A1(new_n28015_), .B0(new_n28395_), .Y(new_n28396_));
  NOR2X1   g25960(.A(new_n28396_), .B(pi1154), .Y(new_n28397_));
  INVX1    g25961(.A(new_n27869_), .Y(new_n28398_));
  AND2X1   g25962(.A(new_n27948_), .B(new_n12591_), .Y(new_n28399_));
  AOI22X1  g25963(.A0(new_n28399_), .A1(new_n28398_), .B0(new_n28394_), .B1(new_n28017_), .Y(new_n28400_));
  OAI21X1  g25964(.A0(new_n28400_), .A1(new_n12615_), .B0(new_n23539_), .Y(new_n28401_));
  NOR4X1   g25965(.A(new_n27849_), .B(new_n25377_), .C(new_n12591_), .D(new_n2722_), .Y(new_n28402_));
  NOR3X1   g25966(.A(new_n25334_), .B(pi0299), .C(pi0199), .Y(new_n28403_));
  NOR4X1   g25967(.A(new_n28403_), .B(new_n28402_), .C(new_n12615_), .D(new_n2722_), .Y(new_n28404_));
  NAND2X1  g25968(.A(new_n25342_), .B(pi1153), .Y(new_n28405_));
  AND2X1   g25969(.A(new_n28405_), .B(new_n28022_), .Y(new_n28406_));
  OAI21X1  g25970(.A0(new_n25803_), .A1(new_n12591_), .B0(new_n28406_), .Y(new_n28407_));
  NAND2X1  g25971(.A(new_n28407_), .B(pi0219), .Y(new_n28408_));
  OAI22X1  g25972(.A0(new_n28408_), .A1(new_n28404_), .B0(new_n28401_), .B1(new_n28397_), .Y(new_n28409_));
  MX2X1    g25973(.A(new_n25336_), .B(new_n25107_), .S0(pi1155), .Y(new_n28410_));
  NOR4X1   g25974(.A(new_n25350_), .B(new_n25268_), .C(new_n12591_), .D(pi0299), .Y(new_n28411_));
  NOR3X1   g25975(.A(new_n28411_), .B(new_n12615_), .C(new_n2722_), .Y(new_n28412_));
  OAI21X1  g25976(.A0(new_n28410_), .A1(new_n9545_), .B0(new_n28412_), .Y(new_n28413_));
  OAI22X1  g25977(.A0(new_n26836_), .A1(new_n2722_), .B0(new_n25096_), .B1(pi1155), .Y(new_n28414_));
  AOI21X1  g25978(.A0(new_n28414_), .A1(new_n28406_), .B0(new_n8548_), .Y(new_n28415_));
  AOI22X1  g25979(.A0(new_n28415_), .A1(new_n28413_), .B0(new_n28409_), .B1(new_n8548_), .Y(new_n28416_));
  NOR3X1   g25980(.A(new_n25336_), .B(pi1155), .C(new_n2722_), .Y(new_n28417_));
  OR4X1    g25981(.A(new_n28417_), .B(new_n28402_), .C(new_n12615_), .D(new_n8548_), .Y(new_n28418_));
  AOI21X1  g25982(.A0(new_n25082_), .A1(new_n12615_), .B0(new_n25118_), .Y(new_n28419_));
  NAND3X1  g25983(.A(new_n28419_), .B(new_n25399_), .C(pi1091), .Y(new_n28420_));
  AOI21X1  g25984(.A0(new_n28420_), .A1(new_n8548_), .B0(pi0219), .Y(new_n28421_));
  OR2X1    g25985(.A(new_n28402_), .B(new_n12615_), .Y(new_n28422_));
  NOR4X1   g25986(.A(new_n25335_), .B(pi1155), .C(new_n2722_), .D(pi0299), .Y(new_n28423_));
  OR2X1    g25987(.A(new_n28423_), .B(new_n28422_), .Y(new_n28424_));
  OR4X1    g25988(.A(new_n25377_), .B(new_n25351_), .C(new_n12591_), .D(new_n12615_), .Y(new_n28425_));
  AOI21X1  g25989(.A0(new_n28425_), .A1(new_n28424_), .B0(new_n8548_), .Y(new_n28426_));
  OAI21X1  g25990(.A0(new_n25096_), .A1(pi1155), .B0(new_n28022_), .Y(new_n28427_));
  OAI21X1  g25991(.A0(new_n28427_), .A1(new_n25803_), .B0(new_n8548_), .Y(new_n28428_));
  AOI21X1  g25992(.A0(new_n28424_), .A1(pi1154), .B0(new_n28428_), .Y(new_n28429_));
  NOR3X1   g25993(.A(new_n28429_), .B(new_n28426_), .C(new_n23539_), .Y(new_n28430_));
  AOI21X1  g25994(.A0(new_n28421_), .A1(new_n28418_), .B0(new_n28430_), .Y(new_n28431_));
  NOR2X1   g25995(.A(new_n25415_), .B(pi1155), .Y(new_n28432_));
  AOI22X1  g25996(.A0(new_n27864_), .A1(new_n25053_), .B0(new_n27858_), .B1(new_n26836_), .Y(new_n28433_));
  NOR2X1   g25997(.A(new_n28433_), .B(new_n28432_), .Y(new_n28434_));
  OR2X1    g25998(.A(pi1154), .B(new_n8548_), .Y(new_n28435_));
  OAI21X1  g25999(.A0(new_n28435_), .A1(new_n28434_), .B0(new_n26780_), .Y(new_n28436_));
  OAI22X1  g26000(.A0(new_n28436_), .A1(new_n28431_), .B0(new_n28416_), .B1(new_n26780_), .Y(new_n28437_));
  AND2X1   g26001(.A(new_n28437_), .B(new_n28338_), .Y(new_n28438_));
  OR2X1    g26002(.A(new_n28438_), .B(po1038), .Y(new_n28439_));
  NOR3X1   g26003(.A(new_n27965_), .B(new_n28208_), .C(new_n26780_), .Y(new_n28440_));
  NOR3X1   g26004(.A(new_n26689_), .B(new_n26679_), .C(pi1091), .Y(new_n28441_));
  OR2X1    g26005(.A(new_n28441_), .B(pi0267), .Y(new_n28442_));
  OAI21X1  g26006(.A0(new_n28442_), .A1(new_n28214_), .B0(new_n28084_), .Y(new_n28443_));
  AND2X1   g26007(.A(pi1155), .B(new_n8548_), .Y(new_n28444_));
  OR2X1    g26008(.A(new_n27906_), .B(pi0219), .Y(new_n28445_));
  OAI22X1  g26009(.A0(new_n28445_), .A1(new_n25015_), .B0(new_n28444_), .B1(new_n23539_), .Y(new_n28446_));
  NOR3X1   g26010(.A(new_n28084_), .B(pi1091), .C(pi0267), .Y(new_n28447_));
  AOI21X1  g26011(.A0(new_n28446_), .A1(pi1091), .B0(new_n28447_), .Y(new_n28448_));
  OAI21X1  g26012(.A0(new_n28443_), .A1(new_n28440_), .B0(new_n28448_), .Y(new_n28449_));
  AOI21X1  g26013(.A0(new_n28449_), .A1(po1038), .B0(new_n28207_), .Y(new_n28450_));
  OAI21X1  g26014(.A0(new_n28439_), .A1(new_n28393_), .B0(new_n28450_), .Y(new_n28451_));
  MX2X1    g26015(.A(new_n28446_), .B(new_n26780_), .S0(new_n2722_), .Y(new_n28452_));
  AOI21X1  g26016(.A0(new_n28452_), .A1(po1038), .B0(new_n26899_), .Y(new_n28453_));
  OAI21X1  g26017(.A0(new_n28437_), .A1(po1038), .B0(new_n28453_), .Y(new_n28454_));
  AND2X1   g26018(.A(new_n28454_), .B(new_n24954_), .Y(new_n28455_));
  NOR2X1   g26019(.A(new_n25351_), .B(new_n23539_), .Y(new_n28456_));
  INVX1    g26020(.A(new_n25336_), .Y(new_n28457_));
  OAI21X1  g26021(.A0(new_n28405_), .A1(pi1155), .B0(new_n12615_), .Y(new_n28458_));
  NOR4X1   g26022(.A(new_n25344_), .B(new_n12591_), .C(pi0299), .D(pi0200), .Y(new_n28459_));
  AOI21X1  g26023(.A0(new_n28458_), .A1(new_n28457_), .B0(new_n28459_), .Y(new_n28460_));
  OAI21X1  g26024(.A0(new_n28460_), .A1(new_n28456_), .B0(pi0211), .Y(new_n28461_));
  AOI21X1  g26025(.A0(pi1154), .A1(new_n7941_), .B0(new_n8009_), .Y(new_n28462_));
  NOR3X1   g26026(.A(new_n28462_), .B(new_n25350_), .C(new_n25108_), .Y(new_n28463_));
  OAI21X1  g26027(.A0(new_n28463_), .A1(new_n25024_), .B0(pi0219), .Y(new_n28464_));
  NAND3X1  g26028(.A(new_n28419_), .B(new_n25399_), .C(new_n23539_), .Y(new_n28465_));
  NAND3X1  g26029(.A(new_n28465_), .B(new_n28464_), .C(new_n8548_), .Y(new_n28466_));
  AND2X1   g26030(.A(new_n28466_), .B(new_n6520_), .Y(new_n28467_));
  OAI21X1  g26031(.A0(new_n28446_), .A1(new_n6520_), .B0(pi0230), .Y(new_n28468_));
  AOI21X1  g26032(.A0(new_n28467_), .A1(new_n28461_), .B0(new_n28468_), .Y(new_n28469_));
  AOI21X1  g26033(.A0(new_n28455_), .A1(new_n28451_), .B0(new_n28469_), .Y(po0424));
  AND2X1   g26034(.A(pi0283), .B(pi0272), .Y(new_n28471_));
  AND2X1   g26035(.A(new_n28471_), .B(pi0275), .Y(new_n28472_));
  INVX1    g26036(.A(new_n27784_), .Y(new_n28473_));
  AOI21X1  g26037(.A0(new_n27807_), .A1(new_n26708_), .B0(new_n23539_), .Y(new_n28474_));
  AOI22X1  g26038(.A0(new_n28474_), .A1(new_n26786_), .B0(new_n27829_), .B1(new_n27773_), .Y(new_n28475_));
  AOI21X1  g26039(.A0(new_n27760_), .A1(new_n27758_), .B0(po1038), .Y(new_n28476_));
  AOI22X1  g26040(.A0(new_n28476_), .A1(new_n28475_), .B0(new_n27820_), .B1(new_n28473_), .Y(new_n28477_));
  INVX1    g26041(.A(new_n28477_), .Y(new_n28478_));
  AOI21X1  g26042(.A0(new_n26756_), .A1(new_n23539_), .B0(po1038), .Y(new_n28479_));
  OAI21X1  g26043(.A0(new_n27769_), .A1(new_n23539_), .B0(new_n28479_), .Y(new_n28480_));
  INVX1    g26044(.A(new_n28480_), .Y(new_n28481_));
  AOI21X1  g26045(.A0(new_n27966_), .A1(new_n27820_), .B0(new_n28481_), .Y(new_n28482_));
  INVX1    g26046(.A(new_n28482_), .Y(new_n28483_));
  MX2X1    g26047(.A(new_n28483_), .B(new_n28478_), .S0(new_n25837_), .Y(new_n28484_));
  NOR3X1   g26048(.A(new_n27817_), .B(new_n28214_), .C(new_n6520_), .Y(new_n28485_));
  NAND3X1  g26049(.A(new_n27964_), .B(new_n27783_), .C(po1038), .Y(new_n28486_));
  NAND2X1  g26050(.A(new_n28486_), .B(new_n28485_), .Y(new_n28487_));
  NOR2X1   g26051(.A(new_n26704_), .B(new_n23539_), .Y(new_n28488_));
  OAI21X1  g26052(.A0(new_n28488_), .A1(new_n27808_), .B0(new_n26709_), .Y(new_n28489_));
  OR4X1    g26053(.A(new_n28489_), .B(new_n26754_), .C(new_n5118_), .D(pi0057), .Y(new_n28490_));
  NAND3X1  g26054(.A(new_n28490_), .B(new_n28487_), .C(new_n25837_), .Y(new_n28491_));
  NOR3X1   g26055(.A(new_n26744_), .B(new_n6520_), .C(new_n23539_), .Y(new_n28492_));
  OR2X1    g26056(.A(new_n28492_), .B(new_n27793_), .Y(new_n28493_));
  AOI21X1  g26057(.A0(new_n28479_), .A1(new_n26746_), .B0(new_n28493_), .Y(new_n28494_));
  AOI21X1  g26058(.A0(new_n28483_), .A1(new_n26681_), .B0(new_n28494_), .Y(new_n28495_));
  AOI21X1  g26059(.A0(new_n28495_), .A1(pi1151), .B0(pi0268), .Y(new_n28496_));
  AOI22X1  g26060(.A0(new_n28496_), .A1(new_n28491_), .B0(new_n28484_), .B1(pi0268), .Y(new_n28497_));
  OR2X1    g26061(.A(new_n28497_), .B(pi1152), .Y(new_n28498_));
  AND2X1   g26062(.A(new_n27964_), .B(po1038), .Y(new_n28499_));
  INVX1    g26063(.A(new_n28499_), .Y(new_n28500_));
  NOR2X1   g26064(.A(new_n27841_), .B(new_n26782_), .Y(new_n28501_));
  OAI21X1  g26065(.A0(new_n28501_), .A1(new_n28475_), .B0(new_n6520_), .Y(new_n28502_));
  NOR2X1   g26066(.A(new_n27831_), .B(new_n26744_), .Y(new_n28503_));
  OAI22X1  g26067(.A0(new_n28503_), .A1(new_n28502_), .B0(new_n28500_), .B1(new_n27784_), .Y(new_n28504_));
  INVX1    g26068(.A(new_n28504_), .Y(new_n28505_));
  NOR2X1   g26069(.A(new_n26677_), .B(pi1091), .Y(new_n28506_));
  INVX1    g26070(.A(new_n28506_), .Y(new_n28507_));
  AND2X1   g26071(.A(new_n28476_), .B(new_n28507_), .Y(new_n28508_));
  AOI21X1  g26072(.A0(new_n28499_), .A1(new_n27966_), .B0(new_n28481_), .Y(new_n28509_));
  INVX1    g26073(.A(new_n28509_), .Y(new_n28510_));
  NOR2X1   g26074(.A(new_n28510_), .B(new_n28508_), .Y(new_n28511_));
  INVX1    g26075(.A(new_n28511_), .Y(new_n28512_));
  AOI21X1  g26076(.A0(new_n28512_), .A1(pi1151), .B0(new_n26895_), .Y(new_n28513_));
  OAI21X1  g26077(.A0(new_n28505_), .A1(pi1151), .B0(new_n28513_), .Y(new_n28514_));
  AOI21X1  g26078(.A0(new_n28489_), .A1(new_n27807_), .B0(po1038), .Y(new_n28515_));
  NOR2X1   g26079(.A(new_n28515_), .B(new_n28485_), .Y(new_n28516_));
  NOR3X1   g26080(.A(new_n26716_), .B(new_n26715_), .C(pi0219), .Y(new_n28517_));
  OAI21X1  g26081(.A0(new_n28517_), .A1(new_n28474_), .B0(new_n6520_), .Y(new_n28518_));
  NOR3X1   g26082(.A(new_n28214_), .B(new_n28031_), .C(new_n6520_), .Y(new_n28519_));
  INVX1    g26083(.A(new_n28519_), .Y(new_n28520_));
  NAND3X1  g26084(.A(new_n28520_), .B(new_n28518_), .C(new_n28487_), .Y(new_n28521_));
  AOI21X1  g26085(.A0(new_n28521_), .A1(pi1151), .B0(pi0268), .Y(new_n28522_));
  OAI21X1  g26086(.A0(new_n28516_), .A1(pi1151), .B0(new_n28522_), .Y(new_n28523_));
  NAND3X1  g26087(.A(new_n28523_), .B(new_n28514_), .C(pi1152), .Y(new_n28524_));
  AOI21X1  g26088(.A0(new_n28524_), .A1(new_n28498_), .B0(new_n26471_), .Y(new_n28525_));
  AND2X1   g26089(.A(new_n27792_), .B(po1038), .Y(new_n28526_));
  INVX1    g26090(.A(new_n28518_), .Y(new_n28527_));
  OAI21X1  g26091(.A0(new_n26706_), .A1(new_n26698_), .B0(new_n23539_), .Y(new_n28528_));
  AND2X1   g26092(.A(new_n28528_), .B(new_n26696_), .Y(new_n28529_));
  AOI22X1  g26093(.A0(new_n28529_), .A1(new_n28527_), .B0(new_n28526_), .B1(new_n27816_), .Y(new_n28530_));
  OAI21X1  g26094(.A0(new_n28475_), .A1(po1038), .B0(new_n28520_), .Y(new_n28531_));
  AOI21X1  g26095(.A0(new_n28531_), .A1(pi1151), .B0(new_n25289_), .Y(new_n28532_));
  OAI21X1  g26096(.A0(new_n28530_), .A1(pi1151), .B0(new_n28532_), .Y(new_n28533_));
  AOI21X1  g26097(.A0(new_n28031_), .A1(po1038), .B0(new_n28492_), .Y(new_n28534_));
  AND2X1   g26098(.A(new_n28534_), .B(new_n28502_), .Y(new_n28535_));
  INVX1    g26099(.A(new_n28535_), .Y(new_n28536_));
  AOI21X1  g26100(.A0(new_n28494_), .A1(new_n25837_), .B0(pi1152), .Y(new_n28537_));
  OAI21X1  g26101(.A0(new_n28536_), .A1(new_n25837_), .B0(new_n28537_), .Y(new_n28538_));
  AOI21X1  g26102(.A0(new_n28538_), .A1(new_n28533_), .B0(pi0268), .Y(new_n28539_));
  NOR3X1   g26103(.A(new_n28208_), .B(new_n27818_), .C(new_n6520_), .Y(new_n28540_));
  NOR2X1   g26104(.A(new_n28355_), .B(new_n23539_), .Y(new_n28541_));
  OAI21X1  g26105(.A0(new_n28541_), .A1(new_n27808_), .B0(new_n27806_), .Y(new_n28542_));
  AOI21X1  g26106(.A0(new_n28542_), .A1(new_n6520_), .B0(new_n28540_), .Y(new_n28543_));
  OR4X1    g26107(.A(new_n28541_), .B(new_n27841_), .C(new_n5118_), .D(pi0057), .Y(new_n28544_));
  AND2X1   g26108(.A(new_n28544_), .B(new_n28486_), .Y(new_n28545_));
  INVX1    g26109(.A(new_n28545_), .Y(new_n28546_));
  OAI21X1  g26110(.A0(new_n28546_), .A1(pi1151), .B0(pi1152), .Y(new_n28547_));
  AOI21X1  g26111(.A0(new_n28543_), .A1(pi1151), .B0(new_n28547_), .Y(new_n28548_));
  INVX1    g26112(.A(new_n27822_), .Y(new_n28549_));
  OR2X1    g26113(.A(new_n27810_), .B(po1038), .Y(new_n28550_));
  OAI21X1  g26114(.A0(new_n28550_), .A1(new_n27808_), .B0(new_n28549_), .Y(new_n28551_));
  NOR2X1   g26115(.A(new_n28551_), .B(new_n25837_), .Y(new_n28552_));
  NOR2X1   g26116(.A(new_n28482_), .B(new_n26681_), .Y(new_n28553_));
  OAI21X1  g26117(.A0(new_n28553_), .A1(pi1151), .B0(new_n25289_), .Y(new_n28554_));
  OAI21X1  g26118(.A0(new_n28554_), .A1(new_n28552_), .B0(pi0268), .Y(new_n28555_));
  OAI21X1  g26119(.A0(new_n28555_), .A1(new_n28548_), .B0(new_n26471_), .Y(new_n28556_));
  NOR2X1   g26120(.A(new_n28556_), .B(new_n28539_), .Y(new_n28557_));
  OAI21X1  g26121(.A0(new_n28557_), .A1(new_n28525_), .B0(new_n28472_), .Y(new_n28558_));
  INVX1    g26122(.A(new_n28472_), .Y(new_n28559_));
  NAND2X1  g26123(.A(pi1152), .B(pi0268), .Y(new_n28560_));
  NOR4X1   g26124(.A(new_n5118_), .B(pi0299), .C(pi0199), .D(pi0057), .Y(new_n28561_));
  NOR2X1   g26125(.A(new_n28561_), .B(new_n26180_), .Y(new_n28562_));
  AOI22X1  g26126(.A0(new_n25053_), .A1(new_n6520_), .B0(new_n11777_), .B1(new_n8548_), .Y(new_n28563_));
  OAI21X1  g26127(.A0(new_n28563_), .A1(new_n25289_), .B0(new_n28562_), .Y(new_n28564_));
  AOI21X1  g26128(.A0(new_n28563_), .A1(new_n25837_), .B0(new_n26471_), .Y(new_n28565_));
  AND2X1   g26129(.A(new_n28565_), .B(new_n28564_), .Y(new_n28566_));
  AOI22X1  g26130(.A0(new_n27884_), .A1(new_n11777_), .B0(new_n25107_), .B1(new_n6520_), .Y(new_n28567_));
  NOR2X1   g26131(.A(new_n28567_), .B(new_n25837_), .Y(new_n28568_));
  MX2X1    g26132(.A(new_n8550_), .B(new_n27873_), .S0(po1038), .Y(new_n28569_));
  OR2X1    g26133(.A(new_n28569_), .B(new_n25837_), .Y(new_n28570_));
  AOI21X1  g26134(.A0(new_n28570_), .A1(new_n25289_), .B0(pi1150), .Y(new_n28571_));
  OAI21X1  g26135(.A0(new_n27726_), .A1(pi1151), .B0(new_n28571_), .Y(new_n28572_));
  AOI21X1  g26136(.A0(new_n28568_), .A1(pi1152), .B0(new_n28572_), .Y(new_n28573_));
  AOI21X1  g26137(.A0(new_n28566_), .A1(new_n28560_), .B0(new_n28573_), .Y(new_n28574_));
  AOI21X1  g26138(.A0(new_n28566_), .A1(pi1152), .B0(new_n2722_), .Y(new_n28575_));
  OAI22X1  g26139(.A0(new_n28575_), .A1(new_n26895_), .B0(new_n28574_), .B1(new_n2722_), .Y(new_n28576_));
  AOI21X1  g26140(.A0(new_n28576_), .A1(new_n28559_), .B0(pi0230), .Y(new_n28577_));
  NOR3X1   g26141(.A(new_n28573_), .B(new_n28566_), .C(new_n24954_), .Y(new_n28578_));
  AOI21X1  g26142(.A0(new_n28577_), .A1(new_n28558_), .B0(new_n28578_), .Y(po0425));
  AOI21X1  g26143(.A0(pi1137), .A1(new_n7941_), .B0(new_n8009_), .Y(new_n28580_));
  NAND2X1  g26144(.A(pi1138), .B(pi0199), .Y(new_n28581_));
  AOI21X1  g26145(.A0(pi1136), .A1(new_n7941_), .B0(pi0200), .Y(new_n28582_));
  AOI21X1  g26146(.A0(new_n28582_), .A1(new_n28581_), .B0(new_n28580_), .Y(new_n28583_));
  AND2X1   g26147(.A(pi1138), .B(new_n8548_), .Y(new_n28584_));
  MX2X1    g26148(.A(pi1136), .B(pi1137), .S0(pi0211), .Y(new_n28585_));
  MX2X1    g26149(.A(new_n28585_), .B(new_n28584_), .S0(pi0219), .Y(new_n28586_));
  MX2X1    g26150(.A(new_n28586_), .B(new_n28583_), .S0(new_n11776_), .Y(new_n28587_));
  INVX1    g26151(.A(new_n28561_), .Y(new_n28588_));
  INVX1    g26152(.A(new_n26855_), .Y(new_n28589_));
  OAI22X1  g26153(.A0(new_n28308_), .A1(pi0200), .B0(new_n28589_), .B1(new_n4422_), .Y(new_n28590_));
  AND2X1   g26154(.A(new_n28585_), .B(pi1091), .Y(new_n28591_));
  OAI22X1  g26155(.A0(new_n28591_), .A1(new_n27334_), .B0(new_n28590_), .B1(new_n28588_), .Y(new_n28592_));
  AOI21X1  g26156(.A0(new_n28242_), .A1(pi0269), .B0(pi1091), .Y(new_n28593_));
  OAI21X1  g26157(.A0(new_n28242_), .A1(pi0817), .B0(new_n28593_), .Y(new_n28594_));
  AOI21X1  g26158(.A0(new_n28252_), .A1(pi0269), .B0(pi1091), .Y(new_n28595_));
  OAI21X1  g26159(.A0(new_n28252_), .A1(pi0817), .B0(new_n28595_), .Y(new_n28596_));
  AOI21X1  g26160(.A0(new_n6520_), .A1(new_n2953_), .B0(new_n23539_), .Y(new_n28597_));
  OAI21X1  g26161(.A0(new_n28215_), .A1(new_n4281_), .B0(new_n28597_), .Y(new_n28598_));
  AND2X1   g26162(.A(pi1091), .B(new_n8009_), .Y(new_n28599_));
  INVX1    g26163(.A(new_n28599_), .Y(new_n28600_));
  OAI21X1  g26164(.A0(new_n28600_), .A1(new_n4281_), .B0(pi0199), .Y(new_n28601_));
  OAI21X1  g26165(.A0(new_n28601_), .A1(new_n11777_), .B0(new_n28598_), .Y(new_n28602_));
  AOI22X1  g26166(.A0(new_n28602_), .A1(new_n28596_), .B0(new_n28594_), .B1(new_n28592_), .Y(new_n28603_));
  MX2X1    g26167(.A(new_n28603_), .B(new_n28587_), .S0(pi0230), .Y(po0426));
  INVX1    g26168(.A(pi0805), .Y(new_n28605_));
  NAND2X1  g26169(.A(new_n26675_), .B(new_n28605_), .Y(new_n28606_));
  AOI21X1  g26170(.A0(new_n28252_), .A1(pi0270), .B0(pi1091), .Y(new_n28607_));
  NAND3X1  g26171(.A(pi1141), .B(pi1091), .C(new_n8548_), .Y(new_n28608_));
  NAND2X1  g26172(.A(new_n28608_), .B(new_n28597_), .Y(new_n28609_));
  OAI21X1  g26173(.A0(new_n28245_), .A1(pi0200), .B0(pi0199), .Y(new_n28610_));
  OR4X1    g26174(.A(new_n28610_), .B(new_n5118_), .C(pi0299), .D(pi0057), .Y(new_n28611_));
  AOI22X1  g26175(.A0(new_n28611_), .A1(new_n28609_), .B0(new_n28607_), .B1(new_n28606_), .Y(new_n28612_));
  INVX1    g26176(.A(pi0270), .Y(new_n28613_));
  OAI21X1  g26177(.A0(new_n28241_), .A1(new_n28613_), .B0(new_n2722_), .Y(new_n28614_));
  AOI21X1  g26178(.A0(new_n28241_), .A1(new_n28605_), .B0(new_n28614_), .Y(new_n28615_));
  MX2X1    g26179(.A(pi1139), .B(pi1140), .S0(pi0211), .Y(new_n28616_));
  NAND2X1  g26180(.A(new_n28616_), .B(pi1091), .Y(new_n28617_));
  AND2X1   g26181(.A(pi1140), .B(pi1091), .Y(new_n28618_));
  AOI22X1  g26182(.A0(new_n28618_), .A1(pi0200), .B0(new_n28599_), .B1(pi1139), .Y(new_n28619_));
  AOI22X1  g26183(.A0(new_n28619_), .A1(new_n28561_), .B0(new_n28617_), .B1(new_n26180_), .Y(new_n28620_));
  OAI21X1  g26184(.A0(new_n28620_), .A1(new_n28615_), .B0(new_n24954_), .Y(new_n28621_));
  AND2X1   g26185(.A(pi1141), .B(new_n8548_), .Y(new_n28622_));
  MX2X1    g26186(.A(new_n28616_), .B(new_n28622_), .S0(pi0219), .Y(new_n28623_));
  AND2X1   g26187(.A(pi1140), .B(new_n7941_), .Y(new_n28624_));
  AND2X1   g26188(.A(pi1141), .B(pi0199), .Y(new_n28625_));
  OAI21X1  g26189(.A0(new_n4035_), .A1(pi0199), .B0(new_n8009_), .Y(new_n28626_));
  OAI22X1  g26190(.A0(new_n28626_), .A1(new_n28625_), .B0(new_n28624_), .B1(new_n8009_), .Y(new_n28627_));
  AOI21X1  g26191(.A0(new_n28627_), .A1(new_n11776_), .B0(new_n24954_), .Y(new_n28628_));
  OAI21X1  g26192(.A0(new_n28623_), .A1(new_n11776_), .B0(new_n28628_), .Y(new_n28629_));
  OAI21X1  g26193(.A0(new_n28621_), .A1(new_n28612_), .B0(new_n28629_), .Y(po0427));
  MX2X1    g26194(.A(new_n26880_), .B(new_n28506_), .S0(pi0271), .Y(new_n28631_));
  INVX1    g26195(.A(new_n28631_), .Y(new_n28632_));
  AND2X1   g26196(.A(new_n26685_), .B(new_n2722_), .Y(new_n28633_));
  MX2X1    g26197(.A(new_n28633_), .B(new_n26686_), .S0(new_n26688_), .Y(new_n28634_));
  AND2X1   g26198(.A(pi1146), .B(pi1091), .Y(new_n28635_));
  NAND2X1  g26199(.A(new_n28635_), .B(new_n8548_), .Y(new_n28636_));
  OAI21X1  g26200(.A0(new_n28635_), .A1(new_n28634_), .B0(new_n28636_), .Y(new_n28637_));
  AOI21X1  g26201(.A0(new_n26222_), .A1(pi1091), .B0(pi0219), .Y(new_n28638_));
  AOI22X1  g26202(.A0(new_n28638_), .A1(new_n28637_), .B0(new_n28632_), .B1(pi0219), .Y(new_n28639_));
  OR2X1    g26203(.A(new_n26091_), .B(pi0211), .Y(new_n28640_));
  OAI22X1  g26204(.A0(new_n28640_), .A1(new_n27787_), .B0(po1038), .B1(pi0299), .Y(new_n28641_));
  NOR2X1   g26205(.A(new_n28635_), .B(new_n28634_), .Y(new_n28642_));
  MX2X1    g26206(.A(new_n28642_), .B(new_n28632_), .S0(pi0199), .Y(new_n28643_));
  AND2X1   g26207(.A(pi1145), .B(pi1091), .Y(new_n28644_));
  OR2X1    g26208(.A(new_n28644_), .B(pi0199), .Y(new_n28645_));
  OAI22X1  g26209(.A0(new_n28645_), .A1(new_n28634_), .B0(new_n28631_), .B1(new_n7941_), .Y(new_n28646_));
  AOI21X1  g26210(.A0(new_n26844_), .A1(pi1147), .B0(pi0200), .Y(new_n28647_));
  AOI22X1  g26211(.A0(new_n28647_), .A1(new_n28646_), .B0(new_n28643_), .B1(pi0200), .Y(new_n28648_));
  OAI22X1  g26212(.A0(new_n28648_), .A1(new_n11777_), .B0(new_n28641_), .B1(new_n28639_), .Y(new_n28649_));
  AOI21X1  g26213(.A0(new_n26282_), .A1(new_n26230_), .B0(pi0219), .Y(new_n28650_));
  AOI21X1  g26214(.A0(pi1145), .A1(new_n7941_), .B0(pi0200), .Y(new_n28651_));
  NOR3X1   g26215(.A(new_n28651_), .B(new_n26310_), .C(pi0299), .Y(new_n28652_));
  NOR4X1   g26216(.A(new_n25096_), .B(new_n25021_), .C(new_n9544_), .D(new_n26091_), .Y(new_n28653_));
  OR2X1    g26217(.A(new_n28653_), .B(new_n28652_), .Y(new_n28654_));
  OAI21X1  g26218(.A0(new_n28654_), .A1(new_n28650_), .B0(new_n6520_), .Y(new_n28655_));
  AOI22X1  g26219(.A0(new_n28640_), .A1(pi0219), .B0(new_n27161_), .B1(new_n26252_), .Y(new_n28656_));
  AOI21X1  g26220(.A0(new_n28656_), .A1(po1038), .B0(new_n24954_), .Y(new_n28657_));
  AOI22X1  g26221(.A0(new_n28657_), .A1(new_n28655_), .B0(new_n28649_), .B1(new_n24954_), .Y(po0428));
  OAI21X1  g26222(.A0(new_n28483_), .A1(pi1150), .B0(pi1149), .Y(new_n28659_));
  AOI21X1  g26223(.A0(new_n28511_), .A1(pi1150), .B0(new_n28659_), .Y(new_n28660_));
  OAI21X1  g26224(.A0(new_n28478_), .A1(pi1150), .B0(new_n26147_), .Y(new_n28661_));
  AOI21X1  g26225(.A0(new_n28505_), .A1(pi1150), .B0(new_n28661_), .Y(new_n28662_));
  OAI21X1  g26226(.A0(new_n28662_), .A1(new_n28660_), .B0(pi1148), .Y(new_n28663_));
  OAI21X1  g26227(.A0(new_n28553_), .A1(pi1150), .B0(new_n26147_), .Y(new_n28664_));
  AOI21X1  g26228(.A0(new_n28545_), .A1(pi1150), .B0(new_n28664_), .Y(new_n28665_));
  OAI21X1  g26229(.A0(new_n28551_), .A1(pi1150), .B0(pi1149), .Y(new_n28666_));
  AOI21X1  g26230(.A0(new_n28543_), .A1(pi1150), .B0(new_n28666_), .Y(new_n28667_));
  OAI21X1  g26231(.A0(new_n28667_), .A1(new_n28665_), .B0(new_n26273_), .Y(new_n28668_));
  AND2X1   g26232(.A(new_n28668_), .B(pi0283), .Y(new_n28669_));
  INVX1    g26233(.A(new_n28562_), .Y(new_n28670_));
  MX2X1    g26234(.A(new_n9547_), .B(new_n27728_), .S0(po1038), .Y(new_n28671_));
  AOI21X1  g26235(.A0(new_n28671_), .A1(new_n26471_), .B0(new_n28563_), .Y(new_n28672_));
  AOI21X1  g26236(.A0(new_n26471_), .A1(pi1149), .B0(new_n28563_), .Y(new_n28673_));
  OAI22X1  g26237(.A0(new_n28673_), .A1(new_n28670_), .B0(new_n28672_), .B1(pi1149), .Y(new_n28674_));
  AOI21X1  g26238(.A0(new_n28674_), .A1(pi1091), .B0(new_n26273_), .Y(new_n28675_));
  AOI21X1  g26239(.A0(new_n27726_), .A1(pi1150), .B0(pi1149), .Y(new_n28676_));
  AND2X1   g26240(.A(new_n28676_), .B(pi1091), .Y(new_n28677_));
  INVX1    g26241(.A(new_n28567_), .Y(new_n28678_));
  AOI21X1  g26242(.A0(new_n28678_), .A1(pi1091), .B0(new_n26471_), .Y(new_n28679_));
  OAI22X1  g26243(.A0(new_n28013_), .A1(new_n11776_), .B0(new_n26849_), .B1(po1038), .Y(new_n28680_));
  OAI21X1  g26244(.A0(new_n28680_), .A1(pi1150), .B0(pi1149), .Y(new_n28681_));
  OAI21X1  g26245(.A0(new_n28681_), .A1(new_n28679_), .B0(new_n26273_), .Y(new_n28682_));
  OAI21X1  g26246(.A0(new_n28682_), .A1(new_n28677_), .B0(new_n26898_), .Y(new_n28683_));
  OAI21X1  g26247(.A0(new_n28683_), .A1(new_n28675_), .B0(pi0272), .Y(new_n28684_));
  AOI21X1  g26248(.A0(new_n28669_), .A1(new_n28663_), .B0(new_n28684_), .Y(new_n28685_));
  NAND2X1  g26249(.A(new_n28521_), .B(pi1150), .Y(new_n28686_));
  OR2X1    g26250(.A(new_n28495_), .B(pi1150), .Y(new_n28687_));
  AND2X1   g26251(.A(new_n28687_), .B(pi1149), .Y(new_n28688_));
  OAI21X1  g26252(.A0(new_n28515_), .A1(new_n28485_), .B0(pi1150), .Y(new_n28689_));
  AOI21X1  g26253(.A0(new_n28490_), .A1(new_n28487_), .B0(pi1150), .Y(new_n28690_));
  NOR2X1   g26254(.A(new_n28690_), .B(pi1149), .Y(new_n28691_));
  AOI22X1  g26255(.A0(new_n28691_), .A1(new_n28689_), .B0(new_n28688_), .B1(new_n28686_), .Y(new_n28692_));
  OAI21X1  g26256(.A0(new_n28531_), .A1(new_n26471_), .B0(pi1149), .Y(new_n28693_));
  AOI21X1  g26257(.A0(new_n28536_), .A1(new_n26471_), .B0(new_n28693_), .Y(new_n28694_));
  OAI21X1  g26258(.A0(new_n28494_), .A1(pi1150), .B0(new_n26147_), .Y(new_n28695_));
  AOI21X1  g26259(.A0(new_n28530_), .A1(pi1150), .B0(new_n28695_), .Y(new_n28696_));
  OR2X1    g26260(.A(new_n28696_), .B(pi1148), .Y(new_n28697_));
  OAI22X1  g26261(.A0(new_n28697_), .A1(new_n28694_), .B0(new_n28692_), .B1(new_n26273_), .Y(new_n28698_));
  OR2X1    g26262(.A(new_n11776_), .B(pi0211), .Y(new_n28699_));
  AOI21X1  g26263(.A0(new_n25044_), .A1(new_n6520_), .B0(new_n26180_), .Y(new_n28700_));
  AOI21X1  g26264(.A0(new_n28700_), .A1(new_n28699_), .B0(new_n26471_), .Y(new_n28701_));
  NOR3X1   g26265(.A(new_n28701_), .B(new_n28670_), .C(new_n26147_), .Y(new_n28702_));
  OAI21X1  g26266(.A0(new_n28672_), .A1(pi1149), .B0(pi1148), .Y(new_n28703_));
  NOR3X1   g26267(.A(new_n28703_), .B(new_n28702_), .C(new_n2722_), .Y(new_n28704_));
  OAI21X1  g26268(.A0(new_n28569_), .A1(pi1150), .B0(pi1149), .Y(new_n28705_));
  AOI21X1  g26269(.A0(new_n28567_), .A1(pi1150), .B0(new_n28705_), .Y(new_n28706_));
  OR4X1    g26270(.A(new_n28706_), .B(new_n28676_), .C(pi1148), .D(new_n2722_), .Y(new_n28707_));
  NAND2X1  g26271(.A(new_n28707_), .B(new_n26898_), .Y(new_n28708_));
  OAI21X1  g26272(.A0(new_n28708_), .A1(new_n28704_), .B0(new_n26896_), .Y(new_n28709_));
  AOI21X1  g26273(.A0(new_n28698_), .A1(pi0283), .B0(new_n28709_), .Y(new_n28710_));
  NOR3X1   g26274(.A(new_n28710_), .B(new_n28685_), .C(pi0230), .Y(new_n28711_));
  OR2X1    g26275(.A(new_n28569_), .B(pi1150), .Y(new_n28712_));
  AOI21X1  g26276(.A0(new_n28701_), .A1(new_n28567_), .B0(new_n26147_), .Y(new_n28713_));
  AND2X1   g26277(.A(new_n28713_), .B(new_n28712_), .Y(new_n28714_));
  NOR3X1   g26278(.A(new_n28714_), .B(new_n28676_), .C(pi1148), .Y(new_n28715_));
  OAI21X1  g26279(.A0(new_n28703_), .A1(new_n28702_), .B0(pi0230), .Y(new_n28716_));
  NOR2X1   g26280(.A(new_n28716_), .B(new_n28715_), .Y(new_n28717_));
  NOR2X1   g26281(.A(new_n28717_), .B(new_n28711_), .Y(po0429));
  MX2X1    g26282(.A(new_n26703_), .B(new_n26678_), .S0(pi0273), .Y(new_n28719_));
  INVX1    g26283(.A(new_n28719_), .Y(new_n28720_));
  NOR3X1   g26284(.A(new_n26685_), .B(pi1091), .C(new_n26688_), .Y(new_n28721_));
  OAI21X1  g26285(.A0(new_n28721_), .A1(pi0273), .B0(new_n26690_), .Y(new_n28722_));
  AOI21X1  g26286(.A0(new_n28635_), .A1(new_n8548_), .B0(pi0219), .Y(new_n28723_));
  AOI22X1  g26287(.A0(new_n28723_), .A1(new_n28722_), .B0(new_n28720_), .B1(pi0219), .Y(new_n28724_));
  AND2X1   g26288(.A(new_n28724_), .B(pi0299), .Y(new_n28725_));
  AOI21X1  g26289(.A0(new_n28635_), .A1(new_n8009_), .B0(pi0199), .Y(new_n28726_));
  NAND2X1  g26290(.A(new_n28726_), .B(new_n28722_), .Y(new_n28727_));
  AOI21X1  g26291(.A0(new_n28720_), .A1(pi0199), .B0(pi0299), .Y(new_n28728_));
  AND2X1   g26292(.A(new_n28728_), .B(new_n28727_), .Y(new_n28729_));
  OR2X1    g26293(.A(new_n28729_), .B(new_n28725_), .Y(new_n28730_));
  OR2X1    g26294(.A(new_n26813_), .B(new_n8549_), .Y(new_n28731_));
  AOI21X1  g26295(.A0(new_n28731_), .A1(pi1091), .B0(new_n28730_), .Y(new_n28732_));
  OAI22X1  g26296(.A0(new_n28732_), .A1(po1038), .B0(new_n28549_), .B1(new_n2722_), .Y(new_n28733_));
  NAND2X1  g26297(.A(new_n28724_), .B(po1038), .Y(new_n28734_));
  AOI21X1  g26298(.A0(new_n28730_), .A1(new_n26363_), .B0(pi1148), .Y(new_n28735_));
  NOR3X1   g26299(.A(new_n2722_), .B(new_n23539_), .C(pi0211), .Y(new_n28736_));
  OAI21X1  g26300(.A0(new_n28736_), .A1(new_n28724_), .B0(pi0299), .Y(new_n28737_));
  INVX1    g26301(.A(new_n26845_), .Y(new_n28738_));
  AOI21X1  g26302(.A0(new_n28643_), .A1(pi0200), .B0(new_n28738_), .Y(new_n28739_));
  AOI21X1  g26303(.A0(new_n28728_), .A1(new_n28727_), .B0(new_n28739_), .Y(new_n28740_));
  AOI21X1  g26304(.A0(new_n28740_), .A1(new_n28737_), .B0(po1038), .Y(new_n28741_));
  AND2X1   g26305(.A(new_n27786_), .B(new_n27723_), .Y(new_n28742_));
  NOR3X1   g26306(.A(new_n28742_), .B(new_n28741_), .C(new_n26273_), .Y(new_n28743_));
  OAI21X1  g26307(.A0(new_n28743_), .A1(new_n28735_), .B0(new_n28734_), .Y(new_n28744_));
  AOI21X1  g26308(.A0(new_n28733_), .A1(pi1147), .B0(new_n28744_), .Y(new_n28745_));
  OAI21X1  g26309(.A0(new_n26261_), .A1(pi0211), .B0(new_n26180_), .Y(new_n28746_));
  OAI21X1  g26310(.A0(new_n8135_), .A1(pi1146), .B0(new_n28561_), .Y(new_n28747_));
  AOI21X1  g26311(.A0(new_n28747_), .A1(new_n28746_), .B0(new_n26091_), .Y(new_n28748_));
  OR2X1    g26312(.A(new_n27095_), .B(new_n3165_), .Y(new_n28749_));
  OAI21X1  g26313(.A0(new_n28749_), .A1(new_n28671_), .B0(new_n26273_), .Y(new_n28750_));
  NOR2X1   g26314(.A(new_n28750_), .B(new_n28748_), .Y(new_n28751_));
  NAND2X1  g26315(.A(new_n26180_), .B(pi1147), .Y(new_n28752_));
  AOI22X1  g26316(.A0(new_n28752_), .A1(new_n28699_), .B0(new_n8075_), .B1(new_n3165_), .Y(new_n28753_));
  OAI21X1  g26317(.A0(new_n26091_), .A1(pi0199), .B0(pi0200), .Y(new_n28754_));
  OAI21X1  g26318(.A0(new_n8135_), .A1(pi1146), .B0(new_n28754_), .Y(new_n28755_));
  OAI21X1  g26319(.A0(new_n28755_), .A1(new_n11777_), .B0(pi1148), .Y(new_n28756_));
  OAI21X1  g26320(.A0(new_n28756_), .A1(new_n28753_), .B0(pi0230), .Y(new_n28757_));
  OAI22X1  g26321(.A0(new_n28757_), .A1(new_n28751_), .B0(new_n28745_), .B1(pi0230), .Y(po0430));
  NAND2X1  g26322(.A(pi1144), .B(pi1091), .Y(new_n28759_));
  AOI21X1  g26323(.A0(new_n28242_), .A1(pi0274), .B0(pi1091), .Y(new_n28760_));
  OAI21X1  g26324(.A0(new_n28242_), .A1(pi0659), .B0(new_n28760_), .Y(new_n28761_));
  AOI21X1  g26325(.A0(new_n28761_), .A1(new_n28759_), .B0(new_n8009_), .Y(new_n28762_));
  INVX1    g26326(.A(new_n28761_), .Y(new_n28763_));
  OAI21X1  g26327(.A0(new_n28763_), .A1(new_n28255_), .B0(new_n8009_), .Y(new_n28764_));
  NAND2X1  g26328(.A(new_n28764_), .B(new_n7941_), .Y(new_n28765_));
  AOI21X1  g26329(.A0(new_n28252_), .A1(pi0274), .B0(pi1091), .Y(new_n28766_));
  OAI21X1  g26330(.A0(new_n28252_), .A1(pi0659), .B0(new_n28766_), .Y(new_n28767_));
  AOI21X1  g26331(.A0(new_n28644_), .A1(new_n8009_), .B0(new_n7941_), .Y(new_n28768_));
  AOI21X1  g26332(.A0(new_n28768_), .A1(new_n28767_), .B0(new_n11777_), .Y(new_n28769_));
  OAI21X1  g26333(.A0(new_n28765_), .A1(new_n28762_), .B0(new_n28769_), .Y(new_n28770_));
  OAI21X1  g26334(.A0(new_n28763_), .A1(new_n28278_), .B0(pi0211), .Y(new_n28771_));
  OAI21X1  g26335(.A0(new_n28763_), .A1(new_n28255_), .B0(new_n8548_), .Y(new_n28772_));
  NAND3X1  g26336(.A(new_n28772_), .B(new_n28771_), .C(new_n23539_), .Y(new_n28773_));
  AOI21X1  g26337(.A0(new_n26222_), .A1(pi1091), .B0(new_n23539_), .Y(new_n28774_));
  AOI21X1  g26338(.A0(new_n28774_), .A1(new_n28767_), .B0(new_n11776_), .Y(new_n28775_));
  AOI21X1  g26339(.A0(new_n28775_), .A1(new_n28773_), .B0(pi0230), .Y(new_n28776_));
  AND2X1   g26340(.A(pi1144), .B(pi0211), .Y(new_n28777_));
  NOR3X1   g26341(.A(new_n28777_), .B(new_n24964_), .C(pi0219), .Y(new_n28778_));
  OR2X1    g26342(.A(new_n28778_), .B(new_n26223_), .Y(new_n28779_));
  AND2X1   g26343(.A(new_n25638_), .B(new_n2953_), .Y(new_n28780_));
  INVX1    g26344(.A(new_n28780_), .Y(new_n28781_));
  AOI22X1  g26345(.A0(new_n25751_), .A1(new_n8548_), .B0(pi0299), .B1(new_n23539_), .Y(new_n28782_));
  AOI21X1  g26346(.A0(pi1143), .A1(new_n7941_), .B0(new_n26322_), .Y(new_n28783_));
  OAI22X1  g26347(.A0(new_n28783_), .A1(new_n28781_), .B0(new_n28782_), .B1(new_n28778_), .Y(new_n28784_));
  AOI21X1  g26348(.A0(new_n28784_), .A1(new_n6520_), .B0(new_n24954_), .Y(new_n28785_));
  AOI22X1  g26349(.A0(new_n28785_), .A1(new_n28779_), .B0(new_n28776_), .B1(new_n28770_), .Y(po0431));
  AOI21X1  g26350(.A0(new_n28569_), .A1(new_n25837_), .B0(new_n26471_), .Y(new_n28787_));
  OAI21X1  g26351(.A0(new_n28567_), .A1(new_n25837_), .B0(new_n28787_), .Y(new_n28788_));
  AOI21X1  g26352(.A0(new_n27726_), .A1(new_n26507_), .B0(pi1149), .Y(new_n28789_));
  NOR3X1   g26353(.A(new_n28561_), .B(new_n26180_), .C(new_n26147_), .Y(new_n28790_));
  OAI21X1  g26354(.A0(new_n28563_), .A1(new_n25837_), .B0(new_n28790_), .Y(new_n28791_));
  NAND3X1  g26355(.A(new_n28563_), .B(new_n26471_), .C(pi1149), .Y(new_n28792_));
  NAND2X1  g26356(.A(new_n28792_), .B(new_n28791_), .Y(new_n28793_));
  AOI21X1  g26357(.A0(new_n28789_), .A1(new_n28788_), .B0(new_n28793_), .Y(new_n28794_));
  OR2X1    g26358(.A(new_n28563_), .B(new_n25837_), .Y(new_n28795_));
  AOI22X1  g26359(.A0(new_n28790_), .A1(new_n28795_), .B0(new_n28568_), .B1(new_n26147_), .Y(new_n28796_));
  OR2X1    g26360(.A(new_n28563_), .B(new_n26147_), .Y(new_n28797_));
  AOI21X1  g26361(.A0(new_n28671_), .A1(new_n25837_), .B0(new_n28797_), .Y(new_n28798_));
  OR2X1    g26362(.A(new_n25837_), .B(pi1149), .Y(new_n28799_));
  OAI21X1  g26363(.A0(new_n28799_), .A1(new_n27725_), .B0(new_n26471_), .Y(new_n28800_));
  OAI22X1  g26364(.A0(new_n28800_), .A1(new_n28798_), .B0(new_n28796_), .B1(new_n26471_), .Y(new_n28801_));
  NOR3X1   g26365(.A(pi1151), .B(new_n26471_), .C(pi1149), .Y(new_n28802_));
  AOI22X1  g26366(.A0(new_n28802_), .A1(new_n28680_), .B0(new_n28801_), .B1(pi1091), .Y(new_n28803_));
  AOI21X1  g26367(.A0(new_n28794_), .A1(pi1091), .B0(pi0275), .Y(new_n28804_));
  NOR2X1   g26368(.A(new_n28804_), .B(new_n28471_), .Y(new_n28805_));
  OAI21X1  g26369(.A0(new_n28803_), .A1(new_n26897_), .B0(new_n28805_), .Y(new_n28806_));
  AND2X1   g26370(.A(new_n28530_), .B(new_n26471_), .Y(new_n28807_));
  OAI21X1  g26371(.A0(new_n28531_), .A1(new_n26471_), .B0(pi1151), .Y(new_n28808_));
  INVX1    g26372(.A(new_n28494_), .Y(new_n28809_));
  AOI21X1  g26373(.A0(new_n28809_), .A1(new_n26471_), .B0(pi1151), .Y(new_n28810_));
  OAI21X1  g26374(.A0(new_n28535_), .A1(new_n26471_), .B0(new_n28810_), .Y(new_n28811_));
  OAI21X1  g26375(.A0(new_n28808_), .A1(new_n28807_), .B0(new_n28811_), .Y(new_n28812_));
  AND2X1   g26376(.A(new_n28812_), .B(new_n26897_), .Y(new_n28813_));
  MX2X1    g26377(.A(new_n28545_), .B(new_n28543_), .S0(pi1150), .Y(new_n28814_));
  MX2X1    g26378(.A(new_n28553_), .B(new_n28551_), .S0(pi1150), .Y(new_n28815_));
  OAI21X1  g26379(.A0(new_n28815_), .A1(pi1151), .B0(pi0275), .Y(new_n28816_));
  AOI21X1  g26380(.A0(new_n28814_), .A1(pi1151), .B0(new_n28816_), .Y(new_n28817_));
  NOR3X1   g26381(.A(new_n28817_), .B(new_n28813_), .C(pi1149), .Y(new_n28818_));
  OAI21X1  g26382(.A0(new_n28477_), .A1(pi1151), .B0(new_n26471_), .Y(new_n28819_));
  AOI21X1  g26383(.A0(new_n28504_), .A1(pi1151), .B0(new_n28819_), .Y(new_n28820_));
  OAI21X1  g26384(.A0(new_n28482_), .A1(pi1151), .B0(pi1150), .Y(new_n28821_));
  AOI21X1  g26385(.A0(new_n28512_), .A1(pi1151), .B0(new_n28821_), .Y(new_n28822_));
  NOR3X1   g26386(.A(new_n28822_), .B(new_n28820_), .C(new_n26897_), .Y(new_n28823_));
  INVX1    g26387(.A(new_n28516_), .Y(new_n28824_));
  NAND2X1  g26388(.A(new_n28686_), .B(pi1151), .Y(new_n28825_));
  AOI21X1  g26389(.A0(new_n28824_), .A1(new_n26471_), .B0(new_n28825_), .Y(new_n28826_));
  OAI21X1  g26390(.A0(new_n28495_), .A1(new_n26471_), .B0(new_n25837_), .Y(new_n28827_));
  OAI21X1  g26391(.A0(new_n28827_), .A1(new_n28690_), .B0(new_n26897_), .Y(new_n28828_));
  OAI21X1  g26392(.A0(new_n28828_), .A1(new_n28826_), .B0(pi1149), .Y(new_n28829_));
  OAI21X1  g26393(.A0(new_n28829_), .A1(new_n28823_), .B0(new_n28471_), .Y(new_n28830_));
  OAI21X1  g26394(.A0(new_n28830_), .A1(new_n28818_), .B0(new_n28806_), .Y(new_n28831_));
  MX2X1    g26395(.A(new_n28831_), .B(new_n28794_), .S0(pi0230), .Y(po0432));
  OAI21X1  g26396(.A0(new_n28242_), .A1(new_n26683_), .B0(new_n3175_), .Y(new_n28833_));
  MX2X1    g26397(.A(new_n3346_), .B(new_n2439_), .S0(new_n8548_), .Y(new_n28834_));
  OAI21X1  g26398(.A0(new_n28834_), .A1(new_n2722_), .B0(new_n26180_), .Y(new_n28835_));
  AOI22X1  g26399(.A0(new_n28278_), .A1(new_n8009_), .B0(new_n26855_), .B1(pi1145), .Y(new_n28836_));
  NAND4X1  g26400(.A(new_n28836_), .B(new_n6520_), .C(new_n2953_), .D(new_n7941_), .Y(new_n28837_));
  AOI22X1  g26401(.A0(new_n28837_), .A1(new_n28835_), .B0(new_n28833_), .B1(new_n28633_), .Y(new_n28838_));
  AOI21X1  g26402(.A0(new_n26676_), .A1(new_n3175_), .B0(new_n28507_), .Y(new_n28839_));
  AOI21X1  g26403(.A0(new_n28635_), .A1(new_n8009_), .B0(new_n7941_), .Y(new_n28840_));
  AOI22X1  g26404(.A0(new_n28840_), .A1(new_n11776_), .B0(new_n28636_), .B1(new_n28597_), .Y(new_n28841_));
  OAI21X1  g26405(.A0(new_n28841_), .A1(new_n28839_), .B0(new_n24954_), .Y(new_n28842_));
  OAI21X1  g26406(.A0(new_n2439_), .A1(pi0199), .B0(new_n26986_), .Y(new_n28843_));
  AOI21X1  g26407(.A0(new_n28843_), .A1(new_n26315_), .B0(new_n11777_), .Y(new_n28844_));
  OAI22X1  g26408(.A0(new_n28834_), .A1(pi0219), .B0(new_n25031_), .B1(new_n3165_), .Y(new_n28845_));
  OAI21X1  g26409(.A0(new_n28845_), .A1(new_n11776_), .B0(pi0230), .Y(new_n28846_));
  OAI22X1  g26410(.A0(new_n28846_), .A1(new_n28844_), .B0(new_n28842_), .B1(new_n28838_), .Y(po0433));
  INVX1    g26411(.A(new_n28618_), .Y(new_n28848_));
  AOI21X1  g26412(.A0(new_n28242_), .A1(pi0277), .B0(pi1091), .Y(new_n28849_));
  OAI21X1  g26413(.A0(new_n28242_), .A1(pi0820), .B0(new_n28849_), .Y(new_n28850_));
  AND2X1   g26414(.A(new_n28850_), .B(new_n28848_), .Y(new_n28851_));
  NAND2X1  g26415(.A(new_n28850_), .B(new_n28245_), .Y(new_n28852_));
  AOI21X1  g26416(.A0(new_n28852_), .A1(pi0200), .B0(pi0199), .Y(new_n28853_));
  OAI21X1  g26417(.A0(new_n28851_), .A1(pi0200), .B0(new_n28853_), .Y(new_n28854_));
  AOI21X1  g26418(.A0(new_n28252_), .A1(pi0277), .B0(pi1091), .Y(new_n28855_));
  OAI21X1  g26419(.A0(new_n28252_), .A1(pi0820), .B0(new_n28855_), .Y(new_n28856_));
  AOI21X1  g26420(.A0(new_n28247_), .A1(new_n8009_), .B0(new_n7941_), .Y(new_n28857_));
  AOI21X1  g26421(.A0(new_n28857_), .A1(new_n28856_), .B0(new_n11777_), .Y(new_n28858_));
  AOI21X1  g26422(.A0(new_n28852_), .A1(pi0211), .B0(pi0219), .Y(new_n28859_));
  OAI21X1  g26423(.A0(new_n28851_), .A1(pi0211), .B0(new_n28859_), .Y(new_n28860_));
  OAI21X1  g26424(.A0(new_n3706_), .A1(pi0211), .B0(pi0219), .Y(new_n28861_));
  OAI21X1  g26425(.A0(new_n27954_), .A1(new_n23539_), .B0(new_n28861_), .Y(new_n28862_));
  AOI21X1  g26426(.A0(new_n28862_), .A1(new_n28856_), .B0(new_n11776_), .Y(new_n28863_));
  AOI22X1  g26427(.A0(new_n28863_), .A1(new_n28860_), .B0(new_n28858_), .B1(new_n28854_), .Y(new_n28864_));
  AOI21X1  g26428(.A0(pi1140), .A1(new_n8548_), .B0(pi0219), .Y(new_n28865_));
  OAI21X1  g26429(.A0(new_n3847_), .A1(new_n8548_), .B0(new_n28865_), .Y(new_n28866_));
  AOI21X1  g26430(.A0(new_n28866_), .A1(new_n28861_), .B0(new_n11776_), .Y(new_n28867_));
  INVX1    g26431(.A(new_n28624_), .Y(new_n28868_));
  AOI22X1  g26432(.A0(new_n28868_), .A1(new_n24969_), .B0(new_n28266_), .B1(pi0200), .Y(new_n28869_));
  OAI21X1  g26433(.A0(new_n28869_), .A1(new_n11777_), .B0(pi0230), .Y(new_n28870_));
  OAI22X1  g26434(.A0(new_n28870_), .A1(new_n28867_), .B0(new_n28864_), .B1(pi0230), .Y(po0434));
  INVX1    g26435(.A(pi0278), .Y(po1130));
  OAI21X1  g26436(.A0(new_n28252_), .A1(pi0976), .B0(new_n2722_), .Y(new_n28873_));
  AOI21X1  g26437(.A0(new_n28252_), .A1(po1130), .B0(new_n28873_), .Y(new_n28874_));
  NOR2X1   g26438(.A(pi1132), .B(new_n2722_), .Y(new_n28875_));
  NAND2X1  g26439(.A(new_n28241_), .B(pi0976), .Y(new_n28876_));
  AOI21X1  g26440(.A0(new_n28242_), .A1(pi0278), .B0(pi1091), .Y(new_n28877_));
  AOI21X1  g26441(.A0(new_n28877_), .A1(new_n28876_), .B0(new_n28875_), .Y(new_n28878_));
  OR2X1    g26442(.A(new_n28878_), .B(pi0199), .Y(new_n28879_));
  OAI21X1  g26443(.A0(new_n28874_), .A1(new_n7941_), .B0(new_n28879_), .Y(new_n28880_));
  INVX1    g26444(.A(pi1133), .Y(new_n28881_));
  AOI22X1  g26445(.A0(new_n28877_), .A1(new_n28876_), .B0(new_n28881_), .B1(pi1091), .Y(new_n28882_));
  MX2X1    g26446(.A(new_n28882_), .B(new_n28874_), .S0(pi0199), .Y(new_n28883_));
  OAI21X1  g26447(.A0(new_n28883_), .A1(new_n8009_), .B0(new_n2953_), .Y(new_n28884_));
  AOI21X1  g26448(.A0(new_n28880_), .A1(new_n8009_), .B0(new_n28884_), .Y(new_n28885_));
  MX2X1    g26449(.A(pi1132), .B(pi1133), .S0(pi0211), .Y(new_n28886_));
  INVX1    g26450(.A(new_n28886_), .Y(new_n28887_));
  AOI22X1  g26451(.A0(new_n28887_), .A1(pi1091), .B0(new_n28877_), .B1(new_n28876_), .Y(new_n28888_));
  MX2X1    g26452(.A(new_n28888_), .B(new_n28874_), .S0(pi0219), .Y(new_n28889_));
  AND2X1   g26453(.A(new_n28889_), .B(pi0299), .Y(new_n28890_));
  OAI21X1  g26454(.A0(new_n28890_), .A1(new_n28885_), .B0(new_n6520_), .Y(new_n28891_));
  AOI21X1  g26455(.A0(new_n28889_), .A1(po1038), .B0(pi0230), .Y(new_n28892_));
  NAND2X1  g26456(.A(new_n28886_), .B(new_n25947_), .Y(new_n28893_));
  AOI21X1  g26457(.A0(pi1132), .A1(new_n7941_), .B0(pi0200), .Y(new_n28894_));
  AOI21X1  g26458(.A0(pi1133), .A1(new_n7941_), .B0(new_n8009_), .Y(new_n28895_));
  OR2X1    g26459(.A(new_n28895_), .B(pi0299), .Y(new_n28896_));
  OAI22X1  g26460(.A0(new_n28896_), .A1(new_n28894_), .B0(new_n28887_), .B1(new_n25633_), .Y(new_n28897_));
  AOI21X1  g26461(.A0(new_n28897_), .A1(new_n6520_), .B0(new_n24954_), .Y(new_n28898_));
  AOI22X1  g26462(.A0(new_n28898_), .A1(new_n28893_), .B0(new_n28892_), .B1(new_n28891_), .Y(new_n28899_));
  OAI21X1  g26463(.A0(new_n28886_), .A1(pi0219), .B0(new_n26110_), .Y(new_n28900_));
  NOR3X1   g26464(.A(pi1132), .B(pi0200), .C(pi0199), .Y(new_n28901_));
  AOI22X1  g26465(.A0(new_n28886_), .A1(new_n25021_), .B0(new_n25030_), .B1(pi0299), .Y(new_n28902_));
  OAI21X1  g26466(.A0(new_n28901_), .A1(new_n28896_), .B0(new_n28902_), .Y(new_n28903_));
  AOI21X1  g26467(.A0(new_n28903_), .A1(new_n6520_), .B0(new_n24954_), .Y(new_n28904_));
  INVX1    g26468(.A(new_n26844_), .Y(new_n28905_));
  AND2X1   g26469(.A(new_n28880_), .B(new_n8009_), .Y(new_n28906_));
  AOI21X1  g26470(.A0(new_n28906_), .A1(new_n28905_), .B0(new_n28884_), .Y(new_n28907_));
  NOR4X1   g26471(.A(new_n2722_), .B(new_n2953_), .C(new_n23539_), .D(pi0211), .Y(new_n28908_));
  OR2X1    g26472(.A(new_n28908_), .B(new_n28890_), .Y(new_n28909_));
  OAI21X1  g26473(.A0(new_n28909_), .A1(new_n28907_), .B0(new_n6520_), .Y(new_n28910_));
  INVX1    g26474(.A(new_n28742_), .Y(new_n28911_));
  AND2X1   g26475(.A(new_n28892_), .B(new_n28911_), .Y(new_n28912_));
  AOI22X1  g26476(.A0(new_n28912_), .A1(new_n28910_), .B0(new_n28904_), .B1(new_n28900_), .Y(new_n28913_));
  MX2X1    g26477(.A(new_n28913_), .B(new_n28899_), .S0(new_n4755_), .Y(po0435));
  NOR2X1   g26478(.A(new_n26675_), .B(pi0279), .Y(new_n28915_));
  OAI21X1  g26479(.A0(new_n28252_), .A1(pi0958), .B0(new_n2722_), .Y(new_n28916_));
  OAI22X1  g26480(.A0(new_n28916_), .A1(new_n28915_), .B0(new_n28600_), .B1(new_n28313_), .Y(new_n28917_));
  NAND2X1  g26481(.A(new_n28917_), .B(pi0199), .Y(new_n28918_));
  OAI21X1  g26482(.A0(new_n28241_), .A1(new_n4652_), .B0(new_n2722_), .Y(new_n28919_));
  AOI21X1  g26483(.A0(new_n28241_), .A1(pi0958), .B0(new_n28919_), .Y(new_n28920_));
  OAI21X1  g26484(.A0(new_n28600_), .A1(pi1133), .B0(new_n7941_), .Y(new_n28921_));
  OR2X1    g26485(.A(new_n28921_), .B(new_n28920_), .Y(new_n28922_));
  AOI21X1  g26486(.A0(new_n28922_), .A1(new_n28918_), .B0(new_n11777_), .Y(new_n28923_));
  NAND2X1  g26487(.A(new_n28923_), .B(new_n28589_), .Y(new_n28924_));
  AOI21X1  g26488(.A0(pi1133), .A1(new_n8548_), .B0(new_n2722_), .Y(new_n28925_));
  OAI21X1  g26489(.A0(new_n28925_), .A1(new_n28920_), .B0(new_n23539_), .Y(new_n28926_));
  AOI21X1  g26490(.A0(new_n27954_), .A1(pi1135), .B0(new_n23539_), .Y(new_n28927_));
  OAI21X1  g26491(.A0(new_n28916_), .A1(new_n28915_), .B0(new_n28927_), .Y(new_n28928_));
  NAND3X1  g26492(.A(new_n28928_), .B(new_n28926_), .C(new_n11777_), .Y(new_n28929_));
  AND2X1   g26493(.A(new_n28929_), .B(new_n24954_), .Y(new_n28930_));
  MX2X1    g26494(.A(new_n28313_), .B(new_n28881_), .S0(new_n7941_), .Y(new_n28931_));
  AOI21X1  g26495(.A0(new_n28881_), .A1(new_n8548_), .B0(pi0219), .Y(new_n28932_));
  AOI22X1  g26496(.A0(new_n28932_), .A1(new_n8548_), .B0(new_n25030_), .B1(pi1135), .Y(new_n28933_));
  OAI22X1  g26497(.A0(new_n28933_), .A1(new_n2953_), .B0(new_n28931_), .B1(new_n25054_), .Y(new_n28934_));
  OAI21X1  g26498(.A0(new_n28933_), .A1(new_n6520_), .B0(pi0230), .Y(new_n28935_));
  AOI21X1  g26499(.A0(new_n28934_), .A1(new_n6520_), .B0(new_n28935_), .Y(new_n28936_));
  AOI21X1  g26500(.A0(new_n28930_), .A1(new_n28924_), .B0(new_n28936_), .Y(new_n28937_));
  OAI21X1  g26501(.A0(new_n28313_), .A1(pi0200), .B0(pi0199), .Y(new_n28938_));
  OAI21X1  g26502(.A0(new_n8135_), .A1(pi1133), .B0(new_n28938_), .Y(new_n28939_));
  AOI21X1  g26503(.A0(new_n25030_), .A1(pi1135), .B0(new_n28932_), .Y(new_n28940_));
  MX2X1    g26504(.A(new_n28940_), .B(new_n28939_), .S0(new_n11776_), .Y(new_n28941_));
  AOI21X1  g26505(.A0(new_n28881_), .A1(new_n8548_), .B0(new_n2722_), .Y(new_n28942_));
  AOI21X1  g26506(.A0(new_n28942_), .A1(new_n26180_), .B0(new_n28923_), .Y(new_n28943_));
  AOI22X1  g26507(.A0(new_n28943_), .A1(new_n28930_), .B0(new_n28941_), .B1(pi0230), .Y(new_n28944_));
  MX2X1    g26508(.A(new_n28944_), .B(new_n28937_), .S0(new_n4755_), .Y(po0436));
  INVX1    g26509(.A(pi1136), .Y(new_n28946_));
  MX2X1    g26510(.A(new_n28946_), .B(new_n28313_), .S0(new_n8548_), .Y(new_n28947_));
  NAND2X1  g26511(.A(new_n28947_), .B(pi1091), .Y(new_n28948_));
  AOI21X1  g26512(.A0(new_n28241_), .A1(pi0914), .B0(pi1091), .Y(new_n28949_));
  OAI21X1  g26513(.A0(new_n28241_), .A1(pi0280), .B0(new_n28949_), .Y(new_n28950_));
  AOI21X1  g26514(.A0(new_n28950_), .A1(new_n28948_), .B0(pi0219), .Y(new_n28951_));
  AOI21X1  g26515(.A0(pi1137), .A1(new_n8548_), .B0(new_n23539_), .Y(new_n28952_));
  OR2X1    g26516(.A(new_n28952_), .B(new_n28283_), .Y(new_n28953_));
  AOI21X1  g26517(.A0(new_n28252_), .A1(pi0280), .B0(pi1091), .Y(new_n28954_));
  OAI21X1  g26518(.A0(new_n28252_), .A1(pi0914), .B0(new_n28954_), .Y(new_n28955_));
  AOI21X1  g26519(.A0(new_n28955_), .A1(new_n28953_), .B0(new_n28951_), .Y(new_n28956_));
  NAND3X1  g26520(.A(pi1137), .B(pi1091), .C(new_n8009_), .Y(new_n28957_));
  AOI21X1  g26521(.A0(new_n28957_), .A1(new_n28955_), .B0(new_n7941_), .Y(new_n28958_));
  INVX1    g26522(.A(new_n28950_), .Y(new_n28959_));
  AND2X1   g26523(.A(pi1136), .B(pi0200), .Y(new_n28960_));
  OAI21X1  g26524(.A0(new_n28313_), .A1(pi0200), .B0(pi1091), .Y(new_n28961_));
  OAI21X1  g26525(.A0(new_n28961_), .A1(new_n28960_), .B0(new_n7941_), .Y(new_n28962_));
  OAI21X1  g26526(.A0(new_n28962_), .A1(new_n28959_), .B0(new_n11776_), .Y(new_n28963_));
  OAI22X1  g26527(.A0(new_n28963_), .A1(new_n28958_), .B0(new_n28956_), .B1(new_n11776_), .Y(new_n28964_));
  AOI21X1  g26528(.A0(pi1136), .A1(new_n7941_), .B0(new_n8009_), .Y(new_n28965_));
  OAI21X1  g26529(.A0(new_n28313_), .A1(pi0199), .B0(new_n8009_), .Y(new_n28966_));
  AOI21X1  g26530(.A0(pi1137), .A1(pi0199), .B0(new_n28966_), .Y(new_n28967_));
  OR4X1    g26531(.A(new_n28967_), .B(new_n28965_), .C(po1038), .D(pi0299), .Y(new_n28968_));
  AOI21X1  g26532(.A0(new_n28947_), .A1(new_n23539_), .B0(new_n28952_), .Y(new_n28969_));
  AOI21X1  g26533(.A0(new_n28969_), .A1(new_n11777_), .B0(new_n24954_), .Y(new_n28970_));
  AOI22X1  g26534(.A0(new_n28970_), .A1(new_n28968_), .B0(new_n28964_), .B1(new_n24954_), .Y(po0437));
  AOI21X1  g26535(.A0(pi1138), .A1(new_n7941_), .B0(new_n8009_), .Y(new_n28972_));
  NAND2X1  g26536(.A(pi1139), .B(pi0199), .Y(new_n28973_));
  AOI21X1  g26537(.A0(pi1137), .A1(new_n7941_), .B0(pi0200), .Y(new_n28974_));
  AOI21X1  g26538(.A0(new_n28974_), .A1(new_n28973_), .B0(new_n28972_), .Y(new_n28975_));
  AND2X1   g26539(.A(pi1139), .B(new_n8548_), .Y(new_n28976_));
  MX2X1    g26540(.A(pi1137), .B(pi1138), .S0(pi0211), .Y(new_n28977_));
  MX2X1    g26541(.A(new_n28977_), .B(new_n28976_), .S0(pi0219), .Y(new_n28978_));
  MX2X1    g26542(.A(new_n28978_), .B(new_n28975_), .S0(new_n11776_), .Y(new_n28979_));
  AOI21X1  g26543(.A0(new_n28242_), .A1(pi0281), .B0(pi1091), .Y(new_n28980_));
  OAI21X1  g26544(.A0(new_n28242_), .A1(pi0830), .B0(new_n28980_), .Y(new_n28981_));
  AND2X1   g26545(.A(new_n28977_), .B(pi1091), .Y(new_n28982_));
  OAI21X1  g26546(.A0(new_n28589_), .A1(new_n4281_), .B0(new_n28957_), .Y(new_n28983_));
  OAI22X1  g26547(.A0(new_n28983_), .A1(new_n28588_), .B0(new_n28982_), .B1(new_n27334_), .Y(new_n28984_));
  AOI21X1  g26548(.A0(new_n28252_), .A1(pi0281), .B0(pi1091), .Y(new_n28985_));
  OAI21X1  g26549(.A0(new_n28252_), .A1(pi0830), .B0(new_n28985_), .Y(new_n28986_));
  OAI21X1  g26550(.A0(new_n28215_), .A1(new_n4035_), .B0(new_n28597_), .Y(new_n28987_));
  OAI21X1  g26551(.A0(new_n28600_), .A1(new_n4035_), .B0(pi0199), .Y(new_n28988_));
  OAI21X1  g26552(.A0(new_n28988_), .A1(new_n11777_), .B0(new_n28987_), .Y(new_n28989_));
  AOI22X1  g26553(.A0(new_n28989_), .A1(new_n28986_), .B0(new_n28984_), .B1(new_n28981_), .Y(new_n28990_));
  MX2X1    g26554(.A(new_n28990_), .B(new_n28979_), .S0(pi0230), .Y(po0438));
  AOI21X1  g26555(.A0(pi1139), .A1(new_n7941_), .B0(new_n8009_), .Y(new_n28992_));
  NAND2X1  g26556(.A(pi1140), .B(pi0199), .Y(new_n28993_));
  AOI21X1  g26557(.A0(pi1138), .A1(new_n7941_), .B0(pi0200), .Y(new_n28994_));
  AOI21X1  g26558(.A0(new_n28994_), .A1(new_n28993_), .B0(new_n28992_), .Y(new_n28995_));
  AND2X1   g26559(.A(pi1140), .B(new_n8548_), .Y(new_n28996_));
  MX2X1    g26560(.A(pi1138), .B(pi1139), .S0(pi0211), .Y(new_n28997_));
  MX2X1    g26561(.A(new_n28997_), .B(new_n28996_), .S0(pi0219), .Y(new_n28998_));
  MX2X1    g26562(.A(new_n28998_), .B(new_n28995_), .S0(new_n11776_), .Y(new_n28999_));
  AOI21X1  g26563(.A0(new_n28242_), .A1(pi0282), .B0(pi1091), .Y(new_n29000_));
  OAI21X1  g26564(.A0(new_n28242_), .A1(pi0836), .B0(new_n29000_), .Y(new_n29001_));
  AND2X1   g26565(.A(new_n28997_), .B(pi1091), .Y(new_n29002_));
  OAI22X1  g26566(.A0(new_n28600_), .A1(new_n4281_), .B0(new_n28589_), .B1(new_n4035_), .Y(new_n29003_));
  OAI22X1  g26567(.A0(new_n29003_), .A1(new_n28588_), .B0(new_n29002_), .B1(new_n27334_), .Y(new_n29004_));
  AOI21X1  g26568(.A0(new_n28252_), .A1(pi0282), .B0(pi1091), .Y(new_n29005_));
  OAI21X1  g26569(.A0(new_n28252_), .A1(pi0836), .B0(new_n29005_), .Y(new_n29006_));
  OAI21X1  g26570(.A0(new_n28215_), .A1(new_n3988_), .B0(new_n28597_), .Y(new_n29007_));
  OAI21X1  g26571(.A0(new_n28848_), .A1(pi0200), .B0(pi0199), .Y(new_n29008_));
  OAI21X1  g26572(.A0(new_n29008_), .A1(new_n11777_), .B0(new_n29007_), .Y(new_n29009_));
  AOI22X1  g26573(.A0(new_n29009_), .A1(new_n29006_), .B0(new_n29004_), .B1(new_n29001_), .Y(new_n29010_));
  MX2X1    g26574(.A(new_n29010_), .B(new_n28999_), .S0(pi0230), .Y(po0439));
  OR2X1    g26575(.A(new_n28671_), .B(new_n26091_), .Y(new_n29012_));
  NAND3X1  g26576(.A(new_n29012_), .B(new_n28678_), .C(pi1149), .Y(new_n29013_));
  OAI21X1  g26577(.A0(new_n28561_), .A1(new_n26180_), .B0(pi1147), .Y(new_n29014_));
  NAND3X1  g26578(.A(new_n29014_), .B(new_n28569_), .C(new_n26147_), .Y(new_n29015_));
  NAND3X1  g26579(.A(new_n29015_), .B(new_n29013_), .C(pi1148), .Y(new_n29016_));
  OAI22X1  g26580(.A0(new_n28671_), .A1(new_n26091_), .B0(new_n27725_), .B1(new_n26147_), .Y(new_n29017_));
  AOI21X1  g26581(.A0(new_n29017_), .A1(new_n26273_), .B0(new_n24954_), .Y(new_n29018_));
  OAI21X1  g26582(.A0(new_n28546_), .A1(pi1147), .B0(new_n26273_), .Y(new_n29019_));
  AOI21X1  g26583(.A0(new_n28505_), .A1(pi1147), .B0(new_n29019_), .Y(new_n29020_));
  AND2X1   g26584(.A(new_n28543_), .B(new_n26091_), .Y(new_n29021_));
  OAI21X1  g26585(.A0(new_n28512_), .A1(new_n26091_), .B0(pi1148), .Y(new_n29022_));
  OAI21X1  g26586(.A0(new_n29022_), .A1(new_n29021_), .B0(pi1149), .Y(new_n29023_));
  AND2X1   g26587(.A(new_n28477_), .B(pi1147), .Y(new_n29024_));
  OAI21X1  g26588(.A0(new_n28553_), .A1(pi1147), .B0(new_n26273_), .Y(new_n29025_));
  OR2X1    g26589(.A(new_n29025_), .B(new_n29024_), .Y(new_n29026_));
  AOI21X1  g26590(.A0(new_n28482_), .A1(pi1147), .B0(new_n26273_), .Y(new_n29027_));
  OAI21X1  g26591(.A0(new_n28551_), .A1(pi1147), .B0(new_n29027_), .Y(new_n29028_));
  AND2X1   g26592(.A(new_n29028_), .B(new_n26147_), .Y(new_n29029_));
  AOI21X1  g26593(.A0(new_n29029_), .A1(new_n29026_), .B0(new_n26898_), .Y(new_n29030_));
  OAI21X1  g26594(.A0(new_n29023_), .A1(new_n29020_), .B0(new_n29030_), .Y(new_n29031_));
  AOI21X1  g26595(.A0(new_n28530_), .A1(new_n26091_), .B0(new_n26147_), .Y(new_n29032_));
  OAI21X1  g26596(.A0(new_n28824_), .A1(new_n26091_), .B0(new_n29032_), .Y(new_n29033_));
  NAND3X1  g26597(.A(new_n28490_), .B(new_n28487_), .C(pi1147), .Y(new_n29034_));
  AOI21X1  g26598(.A0(new_n28809_), .A1(new_n26091_), .B0(pi1149), .Y(new_n29035_));
  AOI21X1  g26599(.A0(new_n29035_), .A1(new_n29034_), .B0(pi1148), .Y(new_n29036_));
  NAND2X1  g26600(.A(new_n29036_), .B(new_n29033_), .Y(new_n29037_));
  AOI21X1  g26601(.A0(new_n28495_), .A1(pi1147), .B0(pi1149), .Y(new_n29038_));
  OAI21X1  g26602(.A0(new_n28535_), .A1(pi1147), .B0(new_n29038_), .Y(new_n29039_));
  OR2X1    g26603(.A(new_n28531_), .B(pi1147), .Y(new_n29040_));
  NAND4X1  g26604(.A(new_n28520_), .B(new_n28518_), .C(new_n28487_), .D(pi1147), .Y(new_n29041_));
  AND2X1   g26605(.A(new_n29041_), .B(pi1149), .Y(new_n29042_));
  AOI21X1  g26606(.A0(new_n29042_), .A1(new_n29040_), .B0(new_n26273_), .Y(new_n29043_));
  AOI21X1  g26607(.A0(new_n29043_), .A1(new_n29039_), .B0(pi0283), .Y(new_n29044_));
  AOI21X1  g26608(.A0(new_n29044_), .A1(new_n29037_), .B0(pi0230), .Y(new_n29045_));
  AOI22X1  g26609(.A0(new_n29045_), .A1(new_n29031_), .B0(new_n29018_), .B1(new_n29016_), .Y(po0440));
  NAND2X1  g26610(.A(new_n28069_), .B(pi1143), .Y(new_n29047_));
  OAI22X1  g26611(.A0(new_n29047_), .A1(new_n26182_), .B0(new_n28069_), .B1(pi0284), .Y(po0441));
  INVX1    g26612(.A(pi0285), .Y(new_n29049_));
  INVX1    g26613(.A(pi0288), .Y(new_n29050_));
  INVX1    g26614(.A(pi0289), .Y(new_n29051_));
  INVX1    g26615(.A(pi0286), .Y(new_n29052_));
  NOR4X1   g26616(.A(new_n7853_), .B(new_n9249_), .C(new_n3131_), .D(new_n29052_), .Y(new_n29053_));
  INVX1    g26617(.A(new_n29053_), .Y(new_n29054_));
  NOR4X1   g26618(.A(new_n29054_), .B(new_n29051_), .C(new_n29050_), .D(new_n29049_), .Y(new_n29055_));
  NOR2X1   g26619(.A(new_n7853_), .B(new_n3131_), .Y(new_n29056_));
  NOR3X1   g26620(.A(new_n29054_), .B(new_n29051_), .C(new_n29050_), .Y(new_n29057_));
  AOI21X1  g26621(.A0(new_n29056_), .A1(pi0285), .B0(new_n29057_), .Y(new_n29058_));
  OR4X1    g26622(.A(new_n29058_), .B(new_n29055_), .C(new_n5118_), .D(pi0057), .Y(new_n29059_));
  INVX1    g26623(.A(new_n29057_), .Y(new_n29060_));
  NOR3X1   g26624(.A(new_n10212_), .B(pi0288), .C(pi0286), .Y(new_n29061_));
  AOI21X1  g26625(.A0(new_n29061_), .A1(new_n29051_), .B0(new_n29049_), .Y(new_n29062_));
  OAI21X1  g26626(.A0(new_n29060_), .A1(po1038), .B0(new_n29062_), .Y(new_n29063_));
  AOI21X1  g26627(.A0(new_n29063_), .A1(new_n29059_), .B0(pi0793), .Y(po0442));
  NOR3X1   g26628(.A(pi0289), .B(pi0286), .C(pi0285), .Y(new_n29065_));
  NOR2X1   g26629(.A(new_n29065_), .B(pi0288), .Y(new_n29066_));
  INVX1    g26630(.A(new_n29056_), .Y(new_n29067_));
  AOI21X1  g26631(.A0(new_n29067_), .A1(new_n9249_), .B0(new_n29052_), .Y(new_n29068_));
  NOR3X1   g26632(.A(new_n29056_), .B(new_n10212_), .C(pi0286), .Y(new_n29069_));
  OAI21X1  g26633(.A0(new_n29069_), .A1(new_n29068_), .B0(new_n29066_), .Y(new_n29070_));
  OAI21X1  g26634(.A0(new_n29067_), .A1(new_n9249_), .B0(new_n29052_), .Y(new_n29071_));
  NOR2X1   g26635(.A(new_n29053_), .B(new_n29050_), .Y(new_n29072_));
  AOI21X1  g26636(.A0(new_n29072_), .A1(new_n29071_), .B0(po1038), .Y(new_n29073_));
  INVX1    g26637(.A(pi0793), .Y(new_n29074_));
  NAND4X1  g26638(.A(new_n29066_), .B(new_n6256_), .C(new_n5938_), .D(new_n2722_), .Y(new_n29075_));
  AND2X1   g26639(.A(new_n29075_), .B(pi0286), .Y(new_n29076_));
  OAI21X1  g26640(.A0(new_n29075_), .A1(pi0286), .B0(po1038), .Y(new_n29077_));
  OAI21X1  g26641(.A0(new_n29077_), .A1(new_n29076_), .B0(new_n29074_), .Y(new_n29078_));
  AOI21X1  g26642(.A0(new_n29073_), .A1(new_n29070_), .B0(new_n29078_), .Y(po0443));
  AOI21X1  g26643(.A0(pi0457), .A1(new_n7862_), .B0(pi0332), .Y(po0444));
  OAI21X1  g26644(.A0(new_n9249_), .A1(new_n29050_), .B0(new_n29075_), .Y(new_n29081_));
  NOR3X1   g26645(.A(new_n7853_), .B(po1038), .C(new_n3131_), .Y(po0637));
  OAI21X1  g26646(.A0(po0637), .A1(new_n29081_), .B0(new_n29074_), .Y(new_n29083_));
  AOI21X1  g26647(.A0(po0637), .A1(new_n29081_), .B0(new_n29083_), .Y(po0445));
  NAND2X1  g26648(.A(new_n29072_), .B(new_n29051_), .Y(new_n29085_));
  OR2X1    g26649(.A(pi0289), .B(new_n29049_), .Y(new_n29086_));
  OR4X1    g26650(.A(new_n29086_), .B(new_n29056_), .C(new_n10212_), .D(pi0286), .Y(new_n29087_));
  OR2X1    g26651(.A(new_n29069_), .B(new_n29051_), .Y(new_n29088_));
  NAND3X1  g26652(.A(new_n29088_), .B(new_n29087_), .C(new_n29050_), .Y(new_n29089_));
  NAND3X1  g26653(.A(new_n29089_), .B(new_n29085_), .C(new_n29060_), .Y(new_n29090_));
  NOR2X1   g26654(.A(new_n29061_), .B(new_n29051_), .Y(new_n29091_));
  NOR4X1   g26655(.A(new_n29086_), .B(new_n10212_), .C(pi0288), .D(pi0286), .Y(new_n29092_));
  OR2X1    g26656(.A(new_n29092_), .B(new_n6520_), .Y(new_n29093_));
  OAI21X1  g26657(.A0(new_n29093_), .A1(new_n29091_), .B0(new_n29074_), .Y(new_n29094_));
  AOI21X1  g26658(.A0(new_n29090_), .A1(new_n6520_), .B0(new_n29094_), .Y(po0446));
  MX2X1    g26659(.A(pi1048), .B(pi0290), .S0(pi0476), .Y(po0447));
  MX2X1    g26660(.A(pi1049), .B(pi0291), .S0(pi0476), .Y(po0448));
  MX2X1    g26661(.A(pi1084), .B(pi0292), .S0(pi0476), .Y(po0449));
  MX2X1    g26662(.A(pi1059), .B(pi0293), .S0(pi0476), .Y(po0450));
  MX2X1    g26663(.A(pi1072), .B(pi0294), .S0(pi0476), .Y(po0451));
  MX2X1    g26664(.A(pi1053), .B(pi0295), .S0(pi0476), .Y(po0452));
  MX2X1    g26665(.A(pi1037), .B(pi0296), .S0(pi0476), .Y(po0453));
  MX2X1    g26666(.A(pi1044), .B(pi0297), .S0(pi0476), .Y(po0454));
  MX2X1    g26667(.A(pi1044), .B(pi0298), .S0(pi0478), .Y(po0455));
  NOR3X1   g26668(.A(new_n3003_), .B(new_n2555_), .C(new_n3112_), .Y(new_n29105_));
  NOR4X1   g26669(.A(new_n9776_), .B(new_n8284_), .C(new_n2506_), .D(pi0054), .Y(new_n29106_));
  AND2X1   g26670(.A(new_n8435_), .B(new_n3109_), .Y(new_n29107_));
  OAI21X1  g26671(.A0(new_n29106_), .A1(new_n29105_), .B0(new_n29107_), .Y(new_n29108_));
  AOI21X1  g26672(.A0(new_n29108_), .A1(new_n2959_), .B0(new_n8433_), .Y(po0456));
  INVX1    g26673(.A(pi0300), .Y(new_n29110_));
  AND2X1   g26674(.A(new_n3153_), .B(pi0057), .Y(new_n29111_));
  NAND4X1  g26675(.A(new_n29111_), .B(new_n7604_), .C(new_n3148_), .D(new_n3130_), .Y(new_n29112_));
  NOR2X1   g26676(.A(new_n29112_), .B(pi0312), .Y(new_n29113_));
  AOI21X1  g26677(.A0(new_n29113_), .A1(new_n29110_), .B0(pi0055), .Y(new_n29114_));
  OAI21X1  g26678(.A0(new_n29113_), .A1(new_n29110_), .B0(new_n29114_), .Y(po0457));
  INVX1    g26679(.A(pi0301), .Y(new_n29116_));
  AND2X1   g26680(.A(new_n29114_), .B(new_n29116_), .Y(new_n29117_));
  OR2X1    g26681(.A(new_n29116_), .B(pi0055), .Y(new_n29118_));
  NOR4X1   g26682(.A(new_n29118_), .B(new_n29112_), .C(pi0312), .D(pi0300), .Y(new_n29119_));
  OR2X1    g26683(.A(new_n29119_), .B(new_n29117_), .Y(po0458));
  NOR4X1   g26684(.A(new_n5118_), .B(new_n4781_), .C(new_n2962_), .D(pi0057), .Y(new_n29121_));
  INVX1    g26685(.A(new_n29121_), .Y(new_n29122_));
  INVX1    g26686(.A(pi0937), .Y(new_n29123_));
  NOR2X1   g26687(.A(pi0223), .B(pi0222), .Y(new_n29124_));
  OAI22X1  g26688(.A0(new_n29124_), .A1(new_n29123_), .B0(new_n23896_), .B1(new_n26674_), .Y(new_n29125_));
  OR2X1    g26689(.A(new_n29125_), .B(new_n29122_), .Y(new_n29126_));
  NOR3X1   g26690(.A(new_n11776_), .B(new_n10137_), .C(pi0215), .Y(new_n29127_));
  INVX1    g26691(.A(new_n29127_), .Y(new_n29128_));
  AOI21X1  g26692(.A0(new_n29128_), .A1(new_n29126_), .B0(new_n22797_), .Y(new_n29129_));
  AOI21X1  g26693(.A0(new_n11777_), .A1(new_n4827_), .B0(new_n29121_), .Y(new_n29130_));
  AND2X1   g26694(.A(new_n29130_), .B(new_n26273_), .Y(new_n29131_));
  NOR3X1   g26695(.A(pi0221), .B(new_n2438_), .C(pi0215), .Y(new_n29132_));
  NOR4X1   g26696(.A(new_n2721_), .B(new_n2437_), .C(pi0216), .D(pi0215), .Y(new_n29133_));
  AOI22X1  g26697(.A0(new_n29133_), .A1(new_n29123_), .B0(new_n29132_), .B1(new_n26674_), .Y(new_n29134_));
  OAI22X1  g26698(.A0(new_n29134_), .A1(new_n11776_), .B0(new_n29126_), .B1(new_n2970_), .Y(new_n29135_));
  NOR3X1   g26699(.A(new_n29135_), .B(new_n29131_), .C(new_n29129_), .Y(po0459));
  MX2X1    g26700(.A(pi1049), .B(pi0303), .S0(pi0478), .Y(po0460));
  MX2X1    g26701(.A(pi1048), .B(pi0304), .S0(pi0478), .Y(po0461));
  MX2X1    g26702(.A(pi1084), .B(pi0305), .S0(pi0478), .Y(po0462));
  MX2X1    g26703(.A(pi1059), .B(pi0306), .S0(pi0478), .Y(po0463));
  MX2X1    g26704(.A(pi1053), .B(pi0307), .S0(pi0478), .Y(po0464));
  MX2X1    g26705(.A(pi1037), .B(pi0308), .S0(pi0478), .Y(po0465));
  MX2X1    g26706(.A(pi1072), .B(pi0309), .S0(pi0478), .Y(po0466));
  AND2X1   g26707(.A(new_n29130_), .B(pi1147), .Y(new_n29144_));
  OR4X1    g26708(.A(new_n11776_), .B(new_n4770_), .C(new_n10136_), .D(pi0215), .Y(new_n29145_));
  NOR3X1   g26709(.A(new_n26688_), .B(pi0221), .C(new_n2438_), .Y(new_n29146_));
  AOI21X1  g26710(.A0(new_n3037_), .A1(pi0934), .B0(new_n29146_), .Y(new_n29147_));
  INVX1    g26711(.A(pi0934), .Y(new_n29148_));
  AOI22X1  g26712(.A0(new_n3163_), .A1(new_n26688_), .B0(new_n29148_), .B1(pi0222), .Y(new_n29149_));
  AOI21X1  g26713(.A0(new_n29149_), .A1(new_n29121_), .B0(new_n29127_), .Y(new_n29150_));
  OAI21X1  g26714(.A0(new_n29147_), .A1(new_n29145_), .B0(new_n29150_), .Y(new_n29151_));
  OAI21X1  g26715(.A0(new_n29151_), .A1(new_n29144_), .B0(new_n22718_), .Y(new_n29152_));
  NAND3X1  g26716(.A(new_n29147_), .B(new_n11777_), .C(new_n4827_), .Y(new_n29153_));
  OAI21X1  g26717(.A0(new_n29149_), .A1(new_n29122_), .B0(pi1147), .Y(new_n29154_));
  AOI21X1  g26718(.A0(new_n11776_), .A1(new_n3008_), .B0(new_n29154_), .Y(new_n29155_));
  NAND2X1  g26719(.A(new_n29121_), .B(new_n2971_), .Y(new_n29156_));
  AOI21X1  g26720(.A0(new_n29156_), .A1(new_n29145_), .B0(pi1147), .Y(new_n29157_));
  AOI22X1  g26721(.A0(new_n29157_), .A1(new_n29151_), .B0(new_n29155_), .B1(new_n29153_), .Y(new_n29158_));
  OAI21X1  g26722(.A0(new_n29158_), .A1(new_n22718_), .B0(new_n29152_), .Y(po0467));
  NOR2X1   g26723(.A(pi0311), .B(pi0055), .Y(new_n29160_));
  MX2X1    g26724(.A(new_n29160_), .B(pi0311), .S0(new_n29119_), .Y(po0468));
  XOR2X1   g26725(.A(new_n29112_), .B(pi0312), .Y(new_n29162_));
  NOR2X1   g26726(.A(new_n29162_), .B(pi0055), .Y(po0469));
  INVX1    g26727(.A(pi0313), .Y(new_n29164_));
  NOR2X1   g26728(.A(new_n9799_), .B(new_n7843_), .Y(new_n29165_));
  OAI21X1  g26729(.A0(new_n9803_), .A1(new_n5922_), .B0(new_n7669_), .Y(new_n29166_));
  NOR2X1   g26730(.A(new_n29166_), .B(new_n29165_), .Y(new_n29167_));
  MX2X1    g26731(.A(new_n29167_), .B(new_n29164_), .S0(pi0954), .Y(po0470));
  INVX1    g26732(.A(new_n5319_), .Y(new_n29169_));
  OAI21X1  g26733(.A0(new_n8436_), .A1(new_n29169_), .B0(new_n11215_), .Y(new_n29170_));
  OAI21X1  g26734(.A0(new_n11018_), .A1(new_n2959_), .B0(new_n3277_), .Y(new_n29171_));
  AOI21X1  g26735(.A0(new_n11119_), .A1(new_n2959_), .B0(new_n29171_), .Y(new_n29172_));
  NOR4X1   g26736(.A(new_n5118_), .B(new_n3139_), .C(new_n3136_), .D(pi0057), .Y(new_n29173_));
  OAI21X1  g26737(.A0(new_n29172_), .A1(new_n11207_), .B0(new_n29173_), .Y(new_n29174_));
  NAND2X1  g26738(.A(new_n10434_), .B(new_n10432_), .Y(new_n29175_));
  AOI21X1  g26739(.A0(new_n29174_), .A1(new_n29170_), .B0(new_n29175_), .Y(po0471));
  OR4X1    g26740(.A(new_n7853_), .B(po1038), .C(new_n3131_), .D(pi0340), .Y(new_n29177_));
  MX2X1    g26741(.A(pi1080), .B(pi0315), .S0(new_n29177_), .Y(po0472));
  MX2X1    g26742(.A(pi1047), .B(pi0316), .S0(new_n29177_), .Y(po0473));
  OR4X1    g26743(.A(new_n7853_), .B(po1038), .C(new_n3131_), .D(pi0330), .Y(new_n29180_));
  MX2X1    g26744(.A(pi1078), .B(pi0317), .S0(new_n29180_), .Y(po0474));
  OR4X1    g26745(.A(new_n7853_), .B(po1038), .C(new_n3131_), .D(pi0341), .Y(new_n29182_));
  MX2X1    g26746(.A(pi1074), .B(pi0318), .S0(new_n29182_), .Y(po0475));
  MX2X1    g26747(.A(pi1072), .B(pi0319), .S0(new_n29182_), .Y(po0476));
  MX2X1    g26748(.A(pi1048), .B(pi0320), .S0(new_n29177_), .Y(po0477));
  MX2X1    g26749(.A(pi1058), .B(pi0321), .S0(new_n29177_), .Y(po0478));
  MX2X1    g26750(.A(pi1051), .B(pi0322), .S0(new_n29177_), .Y(po0479));
  MX2X1    g26751(.A(pi1065), .B(pi0323), .S0(new_n29177_), .Y(po0480));
  MX2X1    g26752(.A(pi1086), .B(pi0324), .S0(new_n29182_), .Y(po0481));
  MX2X1    g26753(.A(pi1063), .B(pi0325), .S0(new_n29182_), .Y(po0482));
  MX2X1    g26754(.A(pi1057), .B(pi0326), .S0(new_n29182_), .Y(po0483));
  MX2X1    g26755(.A(pi1040), .B(pi0327), .S0(new_n29177_), .Y(po0484));
  MX2X1    g26756(.A(pi1058), .B(pi0328), .S0(new_n29182_), .Y(po0485));
  MX2X1    g26757(.A(pi1043), .B(pi0329), .S0(new_n29182_), .Y(po0486));
  NOR3X1   g26758(.A(new_n6520_), .B(new_n2781_), .C(new_n2755_), .Y(new_n29195_));
  INVX1    g26759(.A(new_n29195_), .Y(new_n29196_));
  NOR2X1   g26760(.A(new_n2781_), .B(new_n2755_), .Y(new_n29197_));
  NAND2X1  g26761(.A(new_n29197_), .B(new_n6520_), .Y(new_n29198_));
  MX2X1    g26762(.A(pi0330), .B(pi0340), .S0(new_n29056_), .Y(new_n29199_));
  OAI22X1  g26763(.A0(new_n29199_), .A1(new_n29198_), .B0(new_n29196_), .B1(pi0330), .Y(po0487));
  MX2X1    g26764(.A(pi0331), .B(pi0341), .S0(new_n29056_), .Y(new_n29201_));
  OAI22X1  g26765(.A0(new_n29201_), .A1(new_n29198_), .B0(new_n29196_), .B1(pi0331), .Y(po0488));
  NOR3X1   g26766(.A(new_n8256_), .B(new_n8284_), .C(pi0332), .Y(new_n29203_));
  AOI21X1  g26767(.A0(new_n9570_), .A1(new_n8256_), .B0(new_n5908_), .Y(new_n29204_));
  NOR2X1   g26768(.A(new_n29204_), .B(pi0070), .Y(new_n29205_));
  NOR3X1   g26769(.A(new_n29205_), .B(new_n7260_), .C(new_n2445_), .Y(new_n29206_));
  OAI21X1  g26770(.A0(new_n29206_), .A1(new_n29203_), .B0(new_n2959_), .Y(new_n29207_));
  AOI21X1  g26771(.A0(new_n7863_), .A1(pi0039), .B0(pi0038), .Y(new_n29208_));
  AOI21X1  g26772(.A0(new_n29208_), .A1(new_n29207_), .B0(new_n24863_), .Y(po0489));
  MX2X1    g26773(.A(pi1040), .B(pi0333), .S0(new_n29182_), .Y(po0490));
  MX2X1    g26774(.A(pi1065), .B(pi0334), .S0(new_n29182_), .Y(po0491));
  MX2X1    g26775(.A(pi1069), .B(pi0335), .S0(new_n29182_), .Y(po0492));
  MX2X1    g26776(.A(pi1070), .B(pi0336), .S0(new_n29180_), .Y(po0493));
  MX2X1    g26777(.A(pi1044), .B(pi0337), .S0(new_n29180_), .Y(po0494));
  MX2X1    g26778(.A(pi1072), .B(pi0338), .S0(new_n29180_), .Y(po0495));
  MX2X1    g26779(.A(pi1086), .B(pi0339), .S0(new_n29180_), .Y(po0496));
  OR2X1    g26780(.A(new_n29056_), .B(pi0340), .Y(new_n29217_));
  NOR3X1   g26781(.A(new_n7853_), .B(new_n3131_), .C(pi0331), .Y(new_n29218_));
  NOR2X1   g26782(.A(new_n29218_), .B(new_n29198_), .Y(new_n29219_));
  AOI22X1  g26783(.A0(new_n29219_), .A1(new_n29217_), .B0(new_n29195_), .B1(pi0340), .Y(po0497));
  OAI21X1  g26784(.A0(po0637), .A1(pi0341), .B0(new_n29180_), .Y(new_n29221_));
  AND2X1   g26785(.A(new_n29221_), .B(new_n29197_), .Y(po0498));
  MX2X1    g26786(.A(pi1049), .B(pi0342), .S0(new_n29177_), .Y(po0499));
  MX2X1    g26787(.A(pi1062), .B(pi0343), .S0(new_n29177_), .Y(po0500));
  MX2X1    g26788(.A(pi1069), .B(pi0344), .S0(new_n29177_), .Y(po0501));
  MX2X1    g26789(.A(pi1039), .B(pi0345), .S0(new_n29177_), .Y(po0502));
  MX2X1    g26790(.A(pi1067), .B(pi0346), .S0(new_n29177_), .Y(po0503));
  MX2X1    g26791(.A(pi1055), .B(pi0347), .S0(new_n29177_), .Y(po0504));
  MX2X1    g26792(.A(pi1087), .B(pi0348), .S0(new_n29177_), .Y(po0505));
  MX2X1    g26793(.A(pi1043), .B(pi0349), .S0(new_n29177_), .Y(po0506));
  MX2X1    g26794(.A(pi1035), .B(pi0350), .S0(new_n29177_), .Y(po0507));
  MX2X1    g26795(.A(pi1079), .B(pi0351), .S0(new_n29177_), .Y(po0508));
  MX2X1    g26796(.A(pi1078), .B(pi0352), .S0(new_n29177_), .Y(po0509));
  MX2X1    g26797(.A(pi1063), .B(pi0353), .S0(new_n29177_), .Y(po0510));
  MX2X1    g26798(.A(pi1045), .B(pi0354), .S0(new_n29177_), .Y(po0511));
  MX2X1    g26799(.A(pi1084), .B(pi0355), .S0(new_n29177_), .Y(po0512));
  MX2X1    g26800(.A(pi1081), .B(pi0356), .S0(new_n29177_), .Y(po0513));
  MX2X1    g26801(.A(pi1076), .B(pi0357), .S0(new_n29177_), .Y(po0514));
  MX2X1    g26802(.A(pi1071), .B(pi0358), .S0(new_n29177_), .Y(po0515));
  MX2X1    g26803(.A(pi1068), .B(pi0359), .S0(new_n29177_), .Y(po0516));
  MX2X1    g26804(.A(pi1042), .B(pi0360), .S0(new_n29177_), .Y(po0517));
  MX2X1    g26805(.A(pi1059), .B(pi0361), .S0(new_n29177_), .Y(po0518));
  MX2X1    g26806(.A(pi1070), .B(pi0362), .S0(new_n29177_), .Y(po0519));
  MX2X1    g26807(.A(pi1049), .B(pi0363), .S0(new_n29180_), .Y(po0520));
  MX2X1    g26808(.A(pi1062), .B(pi0364), .S0(new_n29180_), .Y(po0521));
  MX2X1    g26809(.A(pi1065), .B(pi0365), .S0(new_n29180_), .Y(po0522));
  MX2X1    g26810(.A(pi1069), .B(pi0366), .S0(new_n29180_), .Y(po0523));
  MX2X1    g26811(.A(pi1039), .B(pi0367), .S0(new_n29180_), .Y(po0524));
  MX2X1    g26812(.A(pi1067), .B(pi0368), .S0(new_n29180_), .Y(po0525));
  MX2X1    g26813(.A(pi1080), .B(pi0369), .S0(new_n29180_), .Y(po0526));
  MX2X1    g26814(.A(pi1055), .B(pi0370), .S0(new_n29180_), .Y(po0527));
  MX2X1    g26815(.A(pi1051), .B(pi0371), .S0(new_n29180_), .Y(po0528));
  MX2X1    g26816(.A(pi1048), .B(pi0372), .S0(new_n29180_), .Y(po0529));
  MX2X1    g26817(.A(pi1087), .B(pi0373), .S0(new_n29180_), .Y(po0530));
  MX2X1    g26818(.A(pi1035), .B(pi0374), .S0(new_n29180_), .Y(po0531));
  MX2X1    g26819(.A(pi1047), .B(pi0375), .S0(new_n29180_), .Y(po0532));
  MX2X1    g26820(.A(pi1079), .B(pi0376), .S0(new_n29180_), .Y(po0533));
  MX2X1    g26821(.A(pi1074), .B(pi0377), .S0(new_n29180_), .Y(po0534));
  MX2X1    g26822(.A(pi1063), .B(pi0378), .S0(new_n29180_), .Y(po0535));
  MX2X1    g26823(.A(pi1045), .B(pi0379), .S0(new_n29180_), .Y(po0536));
  MX2X1    g26824(.A(pi1084), .B(pi0380), .S0(new_n29180_), .Y(po0537));
  MX2X1    g26825(.A(pi1081), .B(pi0381), .S0(new_n29180_), .Y(po0538));
  MX2X1    g26826(.A(pi1076), .B(pi0382), .S0(new_n29180_), .Y(po0539));
  MX2X1    g26827(.A(pi1071), .B(pi0383), .S0(new_n29180_), .Y(po0540));
  MX2X1    g26828(.A(pi1068), .B(pi0384), .S0(new_n29180_), .Y(po0541));
  MX2X1    g26829(.A(pi1042), .B(pi0385), .S0(new_n29180_), .Y(po0542));
  MX2X1    g26830(.A(pi1059), .B(pi0386), .S0(new_n29180_), .Y(po0543));
  MX2X1    g26831(.A(pi1053), .B(pi0387), .S0(new_n29180_), .Y(po0544));
  MX2X1    g26832(.A(pi1037), .B(pi0388), .S0(new_n29180_), .Y(po0545));
  MX2X1    g26833(.A(pi1036), .B(pi0389), .S0(new_n29180_), .Y(po0546));
  MX2X1    g26834(.A(pi1049), .B(pi0390), .S0(new_n29182_), .Y(po0547));
  MX2X1    g26835(.A(pi1062), .B(pi0391), .S0(new_n29182_), .Y(po0548));
  MX2X1    g26836(.A(pi1039), .B(pi0392), .S0(new_n29182_), .Y(po0549));
  MX2X1    g26837(.A(pi1067), .B(pi0393), .S0(new_n29182_), .Y(po0550));
  MX2X1    g26838(.A(pi1080), .B(pi0394), .S0(new_n29182_), .Y(po0551));
  MX2X1    g26839(.A(pi1055), .B(pi0395), .S0(new_n29182_), .Y(po0552));
  MX2X1    g26840(.A(pi1051), .B(pi0396), .S0(new_n29182_), .Y(po0553));
  MX2X1    g26841(.A(pi1048), .B(pi0397), .S0(new_n29182_), .Y(po0554));
  MX2X1    g26842(.A(pi1087), .B(pi0398), .S0(new_n29182_), .Y(po0555));
  MX2X1    g26843(.A(pi1047), .B(pi0399), .S0(new_n29182_), .Y(po0556));
  MX2X1    g26844(.A(pi1035), .B(pi0400), .S0(new_n29182_), .Y(po0557));
  MX2X1    g26845(.A(pi1079), .B(pi0401), .S0(new_n29182_), .Y(po0558));
  MX2X1    g26846(.A(pi1078), .B(pi0402), .S0(new_n29182_), .Y(po0559));
  MX2X1    g26847(.A(pi1045), .B(pi0403), .S0(new_n29182_), .Y(po0560));
  MX2X1    g26848(.A(pi1084), .B(pi0404), .S0(new_n29182_), .Y(po0561));
  MX2X1    g26849(.A(pi1081), .B(pi0405), .S0(new_n29182_), .Y(po0562));
  MX2X1    g26850(.A(pi1076), .B(pi0406), .S0(new_n29182_), .Y(po0563));
  MX2X1    g26851(.A(pi1071), .B(pi0407), .S0(new_n29182_), .Y(po0564));
  MX2X1    g26852(.A(pi1068), .B(pi0408), .S0(new_n29182_), .Y(po0565));
  MX2X1    g26853(.A(pi1042), .B(pi0409), .S0(new_n29182_), .Y(po0566));
  MX2X1    g26854(.A(pi1059), .B(pi0410), .S0(new_n29182_), .Y(po0567));
  MX2X1    g26855(.A(pi1053), .B(pi0411), .S0(new_n29182_), .Y(po0568));
  MX2X1    g26856(.A(pi1037), .B(pi0412), .S0(new_n29182_), .Y(po0569));
  MX2X1    g26857(.A(pi1036), .B(pi0413), .S0(new_n29182_), .Y(po0570));
  OR4X1    g26858(.A(new_n7853_), .B(po1038), .C(new_n3131_), .D(pi0331), .Y(new_n29295_));
  MX2X1    g26859(.A(pi1049), .B(pi0414), .S0(new_n29295_), .Y(po0571));
  MX2X1    g26860(.A(pi1062), .B(pi0415), .S0(new_n29295_), .Y(po0572));
  MX2X1    g26861(.A(pi1069), .B(pi0416), .S0(new_n29295_), .Y(po0573));
  MX2X1    g26862(.A(pi1039), .B(pi0417), .S0(new_n29295_), .Y(po0574));
  MX2X1    g26863(.A(pi1067), .B(pi0418), .S0(new_n29295_), .Y(po0575));
  MX2X1    g26864(.A(pi1080), .B(pi0419), .S0(new_n29295_), .Y(po0576));
  MX2X1    g26865(.A(pi1055), .B(pi0420), .S0(new_n29295_), .Y(po0577));
  MX2X1    g26866(.A(pi1051), .B(pi0421), .S0(new_n29295_), .Y(po0578));
  MX2X1    g26867(.A(pi1048), .B(pi0422), .S0(new_n29295_), .Y(po0579));
  MX2X1    g26868(.A(pi1087), .B(pi0423), .S0(new_n29295_), .Y(po0580));
  MX2X1    g26869(.A(pi1047), .B(pi0424), .S0(new_n29295_), .Y(po0581));
  MX2X1    g26870(.A(pi1035), .B(pi0425), .S0(new_n29295_), .Y(po0582));
  MX2X1    g26871(.A(pi1079), .B(pi0426), .S0(new_n29295_), .Y(po0583));
  MX2X1    g26872(.A(pi1078), .B(pi0427), .S0(new_n29295_), .Y(po0584));
  MX2X1    g26873(.A(pi1045), .B(pi0428), .S0(new_n29295_), .Y(po0585));
  MX2X1    g26874(.A(pi1084), .B(pi0429), .S0(new_n29295_), .Y(po0586));
  MX2X1    g26875(.A(pi1076), .B(pi0430), .S0(new_n29295_), .Y(po0587));
  MX2X1    g26876(.A(pi1071), .B(pi0431), .S0(new_n29295_), .Y(po0588));
  MX2X1    g26877(.A(pi1068), .B(pi0432), .S0(new_n29295_), .Y(po0589));
  MX2X1    g26878(.A(pi1042), .B(pi0433), .S0(new_n29295_), .Y(po0590));
  MX2X1    g26879(.A(pi1059), .B(pi0434), .S0(new_n29295_), .Y(po0591));
  MX2X1    g26880(.A(pi1053), .B(pi0435), .S0(new_n29295_), .Y(po0592));
  MX2X1    g26881(.A(pi1037), .B(pi0436), .S0(new_n29295_), .Y(po0593));
  MX2X1    g26882(.A(pi1070), .B(pi0437), .S0(new_n29295_), .Y(po0594));
  MX2X1    g26883(.A(pi1036), .B(pi0438), .S0(new_n29295_), .Y(po0595));
  MX2X1    g26884(.A(pi1057), .B(pi0439), .S0(new_n29180_), .Y(po0596));
  MX2X1    g26885(.A(pi1043), .B(pi0440), .S0(new_n29180_), .Y(po0597));
  MX2X1    g26886(.A(pi1044), .B(pi0441), .S0(new_n29177_), .Y(po0598));
  MX2X1    g26887(.A(pi1058), .B(pi0442), .S0(new_n29180_), .Y(po0599));
  MX2X1    g26888(.A(pi1044), .B(pi0443), .S0(new_n29295_), .Y(po0600));
  MX2X1    g26889(.A(pi1072), .B(pi0444), .S0(new_n29295_), .Y(po0601));
  MX2X1    g26890(.A(pi1081), .B(pi0445), .S0(new_n29295_), .Y(po0602));
  MX2X1    g26891(.A(pi1086), .B(pi0446), .S0(new_n29295_), .Y(po0603));
  MX2X1    g26892(.A(pi1040), .B(pi0447), .S0(new_n29180_), .Y(po0604));
  MX2X1    g26893(.A(pi1074), .B(pi0448), .S0(new_n29295_), .Y(po0605));
  MX2X1    g26894(.A(pi1057), .B(pi0449), .S0(new_n29295_), .Y(po0606));
  MX2X1    g26895(.A(pi1036), .B(pi0450), .S0(new_n29177_), .Y(po0607));
  MX2X1    g26896(.A(pi1063), .B(pi0451), .S0(new_n29295_), .Y(po0608));
  MX2X1    g26897(.A(pi1053), .B(pi0452), .S0(new_n29177_), .Y(po0609));
  MX2X1    g26898(.A(pi1040), .B(pi0453), .S0(new_n29295_), .Y(po0610));
  MX2X1    g26899(.A(pi1043), .B(pi0454), .S0(new_n29295_), .Y(po0611));
  MX2X1    g26900(.A(pi1037), .B(pi0455), .S0(new_n29177_), .Y(po0612));
  MX2X1    g26901(.A(pi1044), .B(pi0456), .S0(new_n29182_), .Y(po0613));
  INVX1    g26902(.A(pi0821), .Y(new_n29339_));
  NAND4X1  g26903(.A(pi0601), .B(pi0600), .C(pi0597), .D(pi0594), .Y(new_n29340_));
  INVX1    g26904(.A(pi0595), .Y(new_n29341_));
  INVX1    g26905(.A(pi0804), .Y(new_n29342_));
  INVX1    g26906(.A(pi0810), .Y(new_n29343_));
  NAND3X1  g26907(.A(new_n29343_), .B(new_n29342_), .C(new_n29341_), .Y(new_n29344_));
  INVX1    g26908(.A(pi0596), .Y(new_n29345_));
  INVX1    g26909(.A(pi0599), .Y(new_n29346_));
  AOI21X1  g26910(.A0(pi0810), .A1(new_n29346_), .B0(new_n29345_), .Y(new_n29347_));
  AND2X1   g26911(.A(pi0815), .B(pi0595), .Y(new_n29348_));
  OAI21X1  g26912(.A0(new_n29347_), .A1(new_n29342_), .B0(new_n29348_), .Y(new_n29349_));
  AOI21X1  g26913(.A0(new_n29349_), .A1(new_n29344_), .B0(new_n29340_), .Y(new_n29350_));
  AOI21X1  g26914(.A0(new_n29343_), .A1(pi0600), .B0(new_n29342_), .Y(new_n29351_));
  AOI21X1  g26915(.A0(new_n29343_), .A1(new_n29342_), .B0(pi0601), .Y(new_n29352_));
  NOR3X1   g26916(.A(new_n29352_), .B(new_n29351_), .C(pi0815), .Y(new_n29353_));
  OAI21X1  g26917(.A0(new_n29353_), .A1(new_n29350_), .B0(pi0605), .Y(new_n29354_));
  INVX1    g26918(.A(pi0815), .Y(new_n29355_));
  INVX1    g26919(.A(pi0594), .Y(new_n29356_));
  INVX1    g26920(.A(pi0600), .Y(new_n29357_));
  INVX1    g26921(.A(pi0990), .Y(new_n29358_));
  NOR3X1   g26922(.A(new_n29358_), .B(new_n29357_), .C(new_n29356_), .Y(new_n29359_));
  NAND3X1  g26923(.A(new_n29359_), .B(new_n29351_), .C(new_n29355_), .Y(new_n29360_));
  AOI21X1  g26924(.A0(new_n29360_), .A1(new_n29354_), .B0(new_n29339_), .Y(po0614));
  MX2X1    g26925(.A(pi1072), .B(pi0458), .S0(new_n29177_), .Y(po0615));
  MX2X1    g26926(.A(pi1058), .B(pi0459), .S0(new_n29295_), .Y(po0616));
  MX2X1    g26927(.A(pi1086), .B(pi0460), .S0(new_n29177_), .Y(po0617));
  MX2X1    g26928(.A(pi1057), .B(pi0461), .S0(new_n29177_), .Y(po0618));
  MX2X1    g26929(.A(pi1074), .B(pi0462), .S0(new_n29177_), .Y(po0619));
  MX2X1    g26930(.A(pi1070), .B(pi0463), .S0(new_n29182_), .Y(po0620));
  MX2X1    g26931(.A(pi1065), .B(pi0464), .S0(new_n29295_), .Y(po0621));
  OR2X1    g26932(.A(new_n4782_), .B(new_n4771_), .Y(new_n29369_));
  AND2X1   g26933(.A(new_n29369_), .B(pi0926), .Y(new_n29370_));
  OAI21X1  g26934(.A0(new_n8519_), .A1(new_n8516_), .B0(new_n26673_), .Y(new_n29371_));
  OAI21X1  g26935(.A0(new_n29369_), .A1(new_n12706_), .B0(new_n29371_), .Y(new_n29372_));
  AOI22X1  g26936(.A0(new_n29124_), .A1(new_n2953_), .B0(new_n4898_), .B1(new_n2437_), .Y(new_n29373_));
  AOI21X1  g26937(.A0(pi1157), .A1(new_n26673_), .B0(new_n29373_), .Y(new_n29374_));
  OAI21X1  g26938(.A0(new_n8534_), .A1(pi0216), .B0(new_n3285_), .Y(new_n29375_));
  INVX1    g26939(.A(pi0926), .Y(new_n29376_));
  NOR3X1   g26940(.A(new_n12706_), .B(new_n29376_), .C(pi0243), .Y(new_n29377_));
  AOI22X1  g26941(.A0(new_n29377_), .A1(new_n29375_), .B0(new_n29374_), .B1(new_n29371_), .Y(new_n29378_));
  OAI21X1  g26942(.A0(new_n29372_), .A1(new_n29370_), .B0(new_n29378_), .Y(new_n29379_));
  AOI21X1  g26943(.A0(new_n29132_), .A1(new_n26673_), .B0(new_n6520_), .Y(new_n29380_));
  AOI22X1  g26944(.A0(new_n29133_), .A1(pi0926), .B0(new_n4828_), .B1(pi1157), .Y(new_n29381_));
  AOI22X1  g26945(.A0(new_n29381_), .A1(new_n29380_), .B0(new_n29379_), .B1(new_n6520_), .Y(po0622));
  NOR2X1   g26946(.A(new_n29132_), .B(new_n6520_), .Y(new_n29383_));
  NOR4X1   g26947(.A(new_n8519_), .B(new_n8516_), .C(new_n5118_), .D(pi0057), .Y(new_n29384_));
  NOR2X1   g26948(.A(new_n29384_), .B(new_n29383_), .Y(new_n29385_));
  OR2X1    g26949(.A(new_n29385_), .B(pi0943), .Y(new_n29386_));
  NAND3X1  g26950(.A(new_n29156_), .B(new_n29145_), .C(pi0943), .Y(new_n29387_));
  AOI21X1  g26951(.A0(new_n29387_), .A1(new_n29386_), .B0(pi1151), .Y(new_n29388_));
  NOR2X1   g26952(.A(new_n29386_), .B(new_n29130_), .Y(new_n29389_));
  MX2X1    g26953(.A(new_n3269_), .B(new_n3008_), .S0(new_n11776_), .Y(new_n29390_));
  NAND3X1  g26954(.A(new_n29390_), .B(pi1151), .C(pi0943), .Y(new_n29391_));
  MX2X1    g26955(.A(new_n29373_), .B(new_n3037_), .S0(po1038), .Y(new_n29392_));
  OAI21X1  g26956(.A0(new_n29392_), .A1(pi0275), .B0(new_n29391_), .Y(new_n29393_));
  NOR3X1   g26957(.A(new_n29393_), .B(new_n29389_), .C(new_n29388_), .Y(po0623));
  NOR4X1   g26958(.A(new_n27701_), .B(new_n27700_), .C(pi0287), .D(new_n2549_), .Y(new_n29395_));
  AOI21X1  g26959(.A0(new_n29395_), .A1(po0950), .B0(new_n7668_), .Y(new_n29396_));
  NOR3X1   g26960(.A(new_n9754_), .B(new_n9753_), .C(new_n2472_), .Y(new_n29397_));
  NOR3X1   g26961(.A(new_n11899_), .B(new_n8284_), .C(new_n6789_), .Y(new_n29398_));
  OAI21X1  g26962(.A0(new_n29397_), .A1(pi0102), .B0(new_n29398_), .Y(new_n29399_));
  NOR3X1   g26963(.A(new_n29399_), .B(new_n2603_), .C(pi0098), .Y(new_n29400_));
  INVX1    g26964(.A(new_n29400_), .Y(new_n29401_));
  XOR2X1   g26965(.A(new_n29401_), .B(new_n29395_), .Y(new_n29402_));
  MX2X1    g26966(.A(new_n29401_), .B(new_n29402_), .S0(new_n5895_), .Y(new_n29403_));
  NOR2X1   g26967(.A(new_n29403_), .B(new_n5985_), .Y(new_n29404_));
  OAI21X1  g26968(.A0(new_n29402_), .A1(new_n8259_), .B0(pi1091), .Y(new_n29405_));
  NOR2X1   g26969(.A(new_n29403_), .B(pi1093), .Y(new_n29406_));
  MX2X1    g26970(.A(new_n29401_), .B(new_n29402_), .S0(new_n5939_), .Y(new_n29407_));
  OAI21X1  g26971(.A0(new_n29407_), .A1(new_n2756_), .B0(new_n2722_), .Y(new_n29408_));
  OAI22X1  g26972(.A0(new_n29408_), .A1(new_n29406_), .B0(new_n29405_), .B1(new_n29404_), .Y(new_n29409_));
  NOR3X1   g26973(.A(new_n8436_), .B(new_n29169_), .C(new_n3092_), .Y(new_n29410_));
  AOI21X1  g26974(.A0(new_n29410_), .A1(new_n29409_), .B0(new_n29396_), .Y(po0624));
  NOR4X1   g26975(.A(new_n9580_), .B(new_n7605_), .C(pi0039), .D(new_n2996_), .Y(new_n29412_));
  OAI22X1  g26976(.A0(new_n29412_), .A1(new_n5860_), .B0(new_n8477_), .B1(new_n7690_), .Y(po0625));
  AND2X1   g26977(.A(new_n29369_), .B(pi0942), .Y(new_n29414_));
  OAI21X1  g26978(.A0(new_n8519_), .A1(new_n8516_), .B0(new_n28105_), .Y(new_n29415_));
  OAI21X1  g26979(.A0(new_n29369_), .A1(new_n12684_), .B0(new_n29415_), .Y(new_n29416_));
  AOI21X1  g26980(.A0(pi1156), .A1(new_n28105_), .B0(new_n29373_), .Y(new_n29417_));
  INVX1    g26981(.A(pi0942), .Y(new_n29418_));
  NOR3X1   g26982(.A(new_n12684_), .B(new_n29418_), .C(pi0263), .Y(new_n29419_));
  AOI22X1  g26983(.A0(new_n29419_), .A1(new_n29375_), .B0(new_n29417_), .B1(new_n29415_), .Y(new_n29420_));
  OAI21X1  g26984(.A0(new_n29416_), .A1(new_n29414_), .B0(new_n29420_), .Y(new_n29421_));
  AOI21X1  g26985(.A0(new_n29132_), .A1(new_n28105_), .B0(new_n6520_), .Y(new_n29422_));
  AOI22X1  g26986(.A0(new_n29133_), .A1(pi0942), .B0(new_n4828_), .B1(pi1156), .Y(new_n29423_));
  AOI22X1  g26987(.A0(new_n29423_), .A1(new_n29422_), .B0(new_n29421_), .B1(new_n6520_), .Y(po0626));
  AND2X1   g26988(.A(new_n29369_), .B(pi0925), .Y(new_n29425_));
  OAI21X1  g26989(.A0(new_n8519_), .A1(new_n8516_), .B0(pi0267), .Y(new_n29426_));
  OAI21X1  g26990(.A0(new_n29369_), .A1(new_n12591_), .B0(new_n29426_), .Y(new_n29427_));
  AND2X1   g26991(.A(pi1155), .B(pi0267), .Y(new_n29428_));
  NOR2X1   g26992(.A(new_n29428_), .B(new_n29373_), .Y(new_n29429_));
  AND2X1   g26993(.A(new_n29428_), .B(pi0925), .Y(new_n29430_));
  AOI22X1  g26994(.A0(new_n29430_), .A1(new_n29375_), .B0(new_n29429_), .B1(new_n29426_), .Y(new_n29431_));
  OAI21X1  g26995(.A0(new_n29427_), .A1(new_n29425_), .B0(new_n29431_), .Y(new_n29432_));
  AOI21X1  g26996(.A0(new_n29132_), .A1(pi0267), .B0(new_n6520_), .Y(new_n29433_));
  AOI22X1  g26997(.A0(new_n29133_), .A1(pi0925), .B0(new_n4828_), .B1(pi1155), .Y(new_n29434_));
  AOI22X1  g26998(.A0(new_n29434_), .A1(new_n29433_), .B0(new_n29432_), .B1(new_n6520_), .Y(po0627));
  AND2X1   g26999(.A(new_n29369_), .B(pi0941), .Y(new_n29436_));
  OAI21X1  g27000(.A0(new_n8519_), .A1(new_n8516_), .B0(pi0253), .Y(new_n29437_));
  OAI21X1  g27001(.A0(new_n29369_), .A1(new_n12494_), .B0(new_n29437_), .Y(new_n29438_));
  AND2X1   g27002(.A(pi1153), .B(pi0253), .Y(new_n29439_));
  NOR2X1   g27003(.A(new_n29439_), .B(new_n29373_), .Y(new_n29440_));
  AND2X1   g27004(.A(new_n29439_), .B(pi0941), .Y(new_n29441_));
  AOI22X1  g27005(.A0(new_n29441_), .A1(new_n29375_), .B0(new_n29440_), .B1(new_n29437_), .Y(new_n29442_));
  OAI21X1  g27006(.A0(new_n29438_), .A1(new_n29436_), .B0(new_n29442_), .Y(new_n29443_));
  AOI21X1  g27007(.A0(new_n29132_), .A1(pi0253), .B0(new_n6520_), .Y(new_n29444_));
  AOI22X1  g27008(.A0(new_n29133_), .A1(pi0941), .B0(new_n4828_), .B1(pi1153), .Y(new_n29445_));
  AOI22X1  g27009(.A0(new_n29445_), .A1(new_n29444_), .B0(new_n29443_), .B1(new_n6520_), .Y(po0628));
  AND2X1   g27010(.A(new_n29369_), .B(pi0923), .Y(new_n29447_));
  OAI21X1  g27011(.A0(new_n8519_), .A1(new_n8516_), .B0(pi0254), .Y(new_n29448_));
  OAI21X1  g27012(.A0(new_n29369_), .A1(new_n12615_), .B0(new_n29448_), .Y(new_n29449_));
  AND2X1   g27013(.A(pi1154), .B(pi0254), .Y(new_n29450_));
  NOR2X1   g27014(.A(new_n29450_), .B(new_n29373_), .Y(new_n29451_));
  AND2X1   g27015(.A(new_n29450_), .B(pi0923), .Y(new_n29452_));
  AOI22X1  g27016(.A0(new_n29452_), .A1(new_n29375_), .B0(new_n29451_), .B1(new_n29448_), .Y(new_n29453_));
  OAI21X1  g27017(.A0(new_n29449_), .A1(new_n29447_), .B0(new_n29453_), .Y(new_n29454_));
  AOI21X1  g27018(.A0(new_n29132_), .A1(pi0254), .B0(new_n6520_), .Y(new_n29455_));
  AOI22X1  g27019(.A0(new_n29133_), .A1(pi0923), .B0(new_n4828_), .B1(pi1154), .Y(new_n29456_));
  AOI22X1  g27020(.A0(new_n29456_), .A1(new_n29455_), .B0(new_n29454_), .B1(new_n6520_), .Y(po0629));
  OR2X1    g27021(.A(new_n29385_), .B(pi0922), .Y(new_n29458_));
  NAND3X1  g27022(.A(new_n29156_), .B(new_n29145_), .C(pi0922), .Y(new_n29459_));
  AOI21X1  g27023(.A0(new_n29459_), .A1(new_n29458_), .B0(pi1152), .Y(new_n29460_));
  NOR2X1   g27024(.A(new_n29458_), .B(new_n29130_), .Y(new_n29461_));
  NAND3X1  g27025(.A(new_n29390_), .B(pi1152), .C(pi0922), .Y(new_n29462_));
  OAI21X1  g27026(.A0(new_n29392_), .A1(pi0268), .B0(new_n29462_), .Y(new_n29463_));
  NOR3X1   g27027(.A(new_n29463_), .B(new_n29461_), .C(new_n29460_), .Y(po0630));
  OR2X1    g27028(.A(new_n29385_), .B(pi0931), .Y(new_n29465_));
  NAND3X1  g27029(.A(new_n29156_), .B(new_n29145_), .C(pi0931), .Y(new_n29466_));
  AOI21X1  g27030(.A0(new_n29466_), .A1(new_n29465_), .B0(pi1150), .Y(new_n29467_));
  NOR2X1   g27031(.A(new_n29465_), .B(new_n29130_), .Y(new_n29468_));
  NAND3X1  g27032(.A(new_n29390_), .B(pi1150), .C(pi0931), .Y(new_n29469_));
  OAI21X1  g27033(.A0(new_n29392_), .A1(pi0272), .B0(new_n29469_), .Y(new_n29470_));
  NOR3X1   g27034(.A(new_n29470_), .B(new_n29468_), .C(new_n29467_), .Y(po0631));
  OR2X1    g27035(.A(new_n29385_), .B(pi0936), .Y(new_n29472_));
  NAND3X1  g27036(.A(new_n29156_), .B(new_n29145_), .C(pi0936), .Y(new_n29473_));
  AOI21X1  g27037(.A0(new_n29473_), .A1(new_n29472_), .B0(pi1149), .Y(new_n29474_));
  NOR2X1   g27038(.A(new_n29472_), .B(new_n29130_), .Y(new_n29475_));
  NAND3X1  g27039(.A(new_n29390_), .B(pi1149), .C(pi0936), .Y(new_n29476_));
  OAI21X1  g27040(.A0(new_n29392_), .A1(pi0283), .B0(new_n29476_), .Y(new_n29477_));
  NOR3X1   g27041(.A(new_n29477_), .B(new_n29475_), .C(new_n29474_), .Y(po0632));
  OR4X1    g27042(.A(new_n6520_), .B(pi0219), .C(new_n8548_), .D(new_n2663_), .Y(new_n29479_));
  OAI21X1  g27043(.A0(new_n8549_), .A1(new_n8547_), .B0(new_n7660_), .Y(new_n29480_));
  NOR3X1   g27044(.A(new_n29480_), .B(new_n2582_), .C(new_n2506_), .Y(new_n29481_));
  AOI21X1  g27045(.A0(new_n9534_), .A1(new_n8550_), .B0(new_n29481_), .Y(new_n29482_));
  NOR3X1   g27046(.A(new_n29482_), .B(new_n8284_), .C(new_n3131_), .Y(new_n29483_));
  AOI22X1  g27047(.A0(new_n29483_), .A1(new_n9540_), .B0(new_n8553_), .B1(pi0071), .Y(new_n29484_));
  OAI21X1  g27048(.A0(new_n29484_), .A1(po1038), .B0(new_n29479_), .Y(po0633));
  INVX1    g27049(.A(new_n29167_), .Y(po0634));
  NOR2X1   g27050(.A(new_n28671_), .B(new_n2663_), .Y(po0635));
  MX2X1    g27051(.A(pi0481), .B(pi0248), .S0(new_n22715_), .Y(po0638));
  MX2X1    g27052(.A(pi0482), .B(pi0249), .S0(new_n22728_), .Y(po0639));
  MX2X1    g27053(.A(pi0483), .B(pi0242), .S0(new_n22801_), .Y(po0640));
  MX2X1    g27054(.A(pi0484), .B(pi0249), .S0(new_n22801_), .Y(po0641));
  MX2X1    g27055(.A(pi0485), .B(pi0234), .S0(new_n23537_), .Y(po0642));
  MX2X1    g27056(.A(pi0486), .B(pi0244), .S0(new_n23537_), .Y(po0643));
  MX2X1    g27057(.A(pi0487), .B(pi0246), .S0(new_n22715_), .Y(po0644));
  INVX1    g27058(.A(pi0488), .Y(new_n29495_));
  MX2X1    g27059(.A(new_n29495_), .B(pi0239), .S0(new_n22715_), .Y(po0645));
  MX2X1    g27060(.A(pi0489), .B(pi0242), .S0(new_n23537_), .Y(po0646));
  MX2X1    g27061(.A(pi0490), .B(pi0241), .S0(new_n22801_), .Y(po0647));
  MX2X1    g27062(.A(pi0491), .B(pi0238), .S0(new_n22801_), .Y(po0648));
  MX2X1    g27063(.A(pi0492), .B(pi0240), .S0(new_n22801_), .Y(po0649));
  MX2X1    g27064(.A(pi0493), .B(pi0244), .S0(new_n22801_), .Y(po0650));
  INVX1    g27065(.A(pi0494), .Y(new_n29502_));
  MX2X1    g27066(.A(new_n29502_), .B(pi0239), .S0(new_n22801_), .Y(po0651));
  MX2X1    g27067(.A(pi0495), .B(pi0235), .S0(new_n22801_), .Y(po0652));
  MX2X1    g27068(.A(pi0496), .B(pi0249), .S0(new_n22795_), .Y(po0653));
  INVX1    g27069(.A(pi0497), .Y(new_n29506_));
  MX2X1    g27070(.A(new_n29506_), .B(pi0239), .S0(new_n22795_), .Y(po0654));
  MX2X1    g27071(.A(pi0498), .B(pi0238), .S0(new_n22728_), .Y(po0655));
  MX2X1    g27072(.A(pi0499), .B(pi0246), .S0(new_n22795_), .Y(po0656));
  MX2X1    g27073(.A(pi0500), .B(pi0241), .S0(new_n22795_), .Y(po0657));
  MX2X1    g27074(.A(pi0501), .B(pi0248), .S0(new_n22795_), .Y(po0658));
  MX2X1    g27075(.A(pi0502), .B(pi0247), .S0(new_n22795_), .Y(po0659));
  MX2X1    g27076(.A(pi0503), .B(pi0245), .S0(new_n22795_), .Y(po0660));
  MX2X1    g27077(.A(pi0504), .B(pi0242), .S0(new_n22792_), .Y(po0661));
  INVX1    g27078(.A(pi0505), .Y(new_n29515_));
  MX2X1    g27079(.A(new_n5120_), .B(new_n5219_), .S0(new_n11776_), .Y(new_n29516_));
  AND2X1   g27080(.A(new_n29516_), .B(new_n2990_), .Y(new_n29517_));
  AND2X1   g27081(.A(new_n29517_), .B(new_n22795_), .Y(new_n29518_));
  OR4X1    g27082(.A(new_n22791_), .B(new_n22790_), .C(new_n22713_), .D(new_n2990_), .Y(new_n29519_));
  NAND3X1  g27083(.A(new_n29515_), .B(pi0237), .C(new_n22718_), .Y(new_n29520_));
  OAI22X1  g27084(.A0(new_n29520_), .A1(new_n29519_), .B0(new_n29518_), .B1(new_n29515_), .Y(po0662));
  MX2X1    g27085(.A(pi0506), .B(pi0241), .S0(new_n22792_), .Y(po0663));
  MX2X1    g27086(.A(pi0507), .B(pi0238), .S0(new_n22792_), .Y(po0664));
  MX2X1    g27087(.A(pi0508), .B(pi0247), .S0(new_n22792_), .Y(po0665));
  MX2X1    g27088(.A(pi0509), .B(pi0245), .S0(new_n22792_), .Y(po0666));
  MX2X1    g27089(.A(pi0510), .B(pi0242), .S0(new_n22715_), .Y(po0667));
  NOR3X1   g27090(.A(po1038), .B(new_n5340_), .C(pi0299), .Y(new_n29527_));
  NOR3X1   g27091(.A(new_n29527_), .B(new_n22714_), .C(pi0234), .Y(new_n29528_));
  INVX1    g27092(.A(new_n29528_), .Y(new_n29529_));
  MX2X1    g27093(.A(pi0511), .B(new_n29529_), .S0(new_n22715_), .Y(po0668));
  MX2X1    g27094(.A(pi0512), .B(pi0235), .S0(new_n22715_), .Y(po0669));
  MX2X1    g27095(.A(pi0513), .B(pi0244), .S0(new_n22715_), .Y(po0670));
  MX2X1    g27096(.A(pi0514), .B(pi0245), .S0(new_n22715_), .Y(po0671));
  MX2X1    g27097(.A(pi0515), .B(pi0240), .S0(new_n22715_), .Y(po0672));
  MX2X1    g27098(.A(pi0516), .B(pi0247), .S0(new_n22715_), .Y(po0673));
  MX2X1    g27099(.A(pi0517), .B(pi0238), .S0(new_n22715_), .Y(po0674));
  INVX1    g27100(.A(pi0518), .Y(new_n29537_));
  AND2X1   g27101(.A(new_n29528_), .B(new_n22722_), .Y(new_n29538_));
  OR4X1    g27102(.A(new_n22714_), .B(new_n22713_), .C(new_n22712_), .D(new_n2990_), .Y(new_n29539_));
  NAND3X1  g27103(.A(new_n29537_), .B(pi0237), .C(new_n22718_), .Y(new_n29540_));
  OAI22X1  g27104(.A0(new_n29540_), .A1(new_n29539_), .B0(new_n29538_), .B1(new_n29537_), .Y(po0675));
  INVX1    g27105(.A(pi0519), .Y(new_n29542_));
  MX2X1    g27106(.A(new_n29542_), .B(pi0239), .S0(new_n22722_), .Y(po0676));
  MX2X1    g27107(.A(pi0520), .B(pi0246), .S0(new_n22722_), .Y(po0677));
  MX2X1    g27108(.A(pi0521), .B(pi0248), .S0(new_n22722_), .Y(po0678));
  MX2X1    g27109(.A(pi0522), .B(pi0238), .S0(new_n22722_), .Y(po0679));
  INVX1    g27110(.A(pi0523), .Y(new_n29547_));
  AND2X1   g27111(.A(new_n29528_), .B(new_n23553_), .Y(new_n29548_));
  NAND3X1  g27112(.A(new_n29547_), .B(new_n22797_), .C(pi0233), .Y(new_n29549_));
  OAI22X1  g27113(.A0(new_n29549_), .A1(new_n29539_), .B0(new_n29548_), .B1(new_n29547_), .Y(po0680));
  INVX1    g27114(.A(pi0524), .Y(new_n29551_));
  MX2X1    g27115(.A(new_n29551_), .B(pi0239), .S0(new_n23553_), .Y(po0681));
  MX2X1    g27116(.A(pi0525), .B(pi0245), .S0(new_n23553_), .Y(po0682));
  MX2X1    g27117(.A(pi0526), .B(pi0246), .S0(new_n23553_), .Y(po0683));
  MX2X1    g27118(.A(pi0527), .B(pi0247), .S0(new_n23553_), .Y(po0684));
  MX2X1    g27119(.A(pi0528), .B(pi0249), .S0(new_n23553_), .Y(po0685));
  MX2X1    g27120(.A(pi0529), .B(pi0238), .S0(new_n23553_), .Y(po0686));
  MX2X1    g27121(.A(pi0530), .B(pi0240), .S0(new_n23553_), .Y(po0687));
  MX2X1    g27122(.A(pi0531), .B(pi0235), .S0(new_n22728_), .Y(po0688));
  MX2X1    g27123(.A(pi0532), .B(pi0247), .S0(new_n22728_), .Y(po0689));
  MX2X1    g27124(.A(pi0533), .B(pi0235), .S0(new_n22792_), .Y(po0690));
  INVX1    g27125(.A(pi0534), .Y(new_n29562_));
  MX2X1    g27126(.A(new_n29562_), .B(pi0239), .S0(new_n22792_), .Y(po0691));
  MX2X1    g27127(.A(pi0535), .B(pi0240), .S0(new_n22792_), .Y(po0692));
  MX2X1    g27128(.A(pi0536), .B(pi0246), .S0(new_n22792_), .Y(po0693));
  MX2X1    g27129(.A(pi0537), .B(pi0248), .S0(new_n22792_), .Y(po0694));
  MX2X1    g27130(.A(pi0538), .B(pi0249), .S0(new_n22792_), .Y(po0695));
  MX2X1    g27131(.A(pi0539), .B(pi0242), .S0(new_n22795_), .Y(po0696));
  MX2X1    g27132(.A(pi0540), .B(pi0235), .S0(new_n22795_), .Y(po0697));
  MX2X1    g27133(.A(pi0541), .B(pi0244), .S0(new_n22795_), .Y(po0698));
  MX2X1    g27134(.A(pi0542), .B(pi0240), .S0(new_n22795_), .Y(po0699));
  MX2X1    g27135(.A(pi0543), .B(pi0238), .S0(new_n22795_), .Y(po0700));
  INVX1    g27136(.A(pi0544), .Y(new_n29573_));
  AND2X1   g27137(.A(new_n29517_), .B(new_n22801_), .Y(new_n29574_));
  NAND3X1  g27138(.A(new_n29573_), .B(new_n22797_), .C(pi0233), .Y(new_n29575_));
  OAI22X1  g27139(.A0(new_n29575_), .A1(new_n29519_), .B0(new_n29574_), .B1(new_n29573_), .Y(po0701));
  MX2X1    g27140(.A(pi0545), .B(pi0245), .S0(new_n22801_), .Y(po0702));
  MX2X1    g27141(.A(pi0546), .B(pi0246), .S0(new_n22801_), .Y(po0703));
  MX2X1    g27142(.A(pi0547), .B(pi0247), .S0(new_n22801_), .Y(po0704));
  MX2X1    g27143(.A(pi0548), .B(pi0248), .S0(new_n22801_), .Y(po0705));
  MX2X1    g27144(.A(pi0549), .B(pi0235), .S0(new_n23537_), .Y(po0706));
  INVX1    g27145(.A(pi0550), .Y(new_n29582_));
  MX2X1    g27146(.A(new_n29582_), .B(pi0239), .S0(new_n23537_), .Y(po0707));
  MX2X1    g27147(.A(pi0551), .B(pi0240), .S0(new_n23537_), .Y(po0708));
  MX2X1    g27148(.A(pi0552), .B(pi0247), .S0(new_n23537_), .Y(po0709));
  MX2X1    g27149(.A(pi0553), .B(pi0241), .S0(new_n23537_), .Y(po0710));
  MX2X1    g27150(.A(pi0554), .B(pi0248), .S0(new_n23537_), .Y(po0711));
  MX2X1    g27151(.A(pi0555), .B(pi0249), .S0(new_n23537_), .Y(po0712));
  MX2X1    g27152(.A(pi0556), .B(pi0242), .S0(new_n22728_), .Y(po0713));
  INVX1    g27153(.A(pi0557), .Y(new_n29590_));
  AND2X1   g27154(.A(new_n29517_), .B(new_n22792_), .Y(new_n29591_));
  NAND2X1  g27155(.A(new_n22589_), .B(new_n29590_), .Y(new_n29592_));
  OAI22X1  g27156(.A0(new_n29592_), .A1(new_n29519_), .B0(new_n29591_), .B1(new_n29590_), .Y(po0714));
  MX2X1    g27157(.A(pi0558), .B(pi0244), .S0(new_n22792_), .Y(po0715));
  MX2X1    g27158(.A(pi0559), .B(pi0241), .S0(new_n22715_), .Y(po0716));
  MX2X1    g27159(.A(pi0560), .B(pi0240), .S0(new_n22728_), .Y(po0717));
  MX2X1    g27160(.A(pi0561), .B(pi0247), .S0(new_n22722_), .Y(po0718));
  MX2X1    g27161(.A(pi0562), .B(pi0241), .S0(new_n22728_), .Y(po0719));
  MX2X1    g27162(.A(pi0563), .B(pi0246), .S0(new_n23537_), .Y(po0720));
  MX2X1    g27163(.A(pi0564), .B(pi0246), .S0(new_n22728_), .Y(po0721));
  MX2X1    g27164(.A(pi0565), .B(pi0248), .S0(new_n22728_), .Y(po0722));
  MX2X1    g27165(.A(pi0566), .B(pi0244), .S0(new_n22728_), .Y(po0723));
  AND2X1   g27166(.A(pi1092), .B(new_n5928_), .Y(new_n29603_));
  NOR4X1   g27167(.A(new_n14184_), .B(new_n14178_), .C(new_n23670_), .D(new_n5027_), .Y(new_n29604_));
  NOR3X1   g27168(.A(pi1093), .B(new_n2755_), .C(pi0567), .Y(new_n29605_));
  NOR3X1   g27169(.A(new_n29605_), .B(new_n29604_), .C(pi0789), .Y(new_n29606_));
  AND2X1   g27170(.A(new_n29604_), .B(new_n12637_), .Y(new_n29607_));
  OR2X1    g27171(.A(new_n29607_), .B(new_n29605_), .Y(new_n29608_));
  AOI21X1  g27172(.A0(new_n29604_), .A1(pi0619), .B0(new_n29605_), .Y(new_n29609_));
  OAI21X1  g27173(.A0(new_n29609_), .A1(new_n12638_), .B0(pi0789), .Y(new_n29610_));
  AOI21X1  g27174(.A0(new_n29608_), .A1(new_n12638_), .B0(new_n29610_), .Y(new_n29611_));
  NOR2X1   g27175(.A(new_n29611_), .B(new_n29606_), .Y(new_n29612_));
  NOR4X1   g27176(.A(new_n13569_), .B(new_n12219_), .C(new_n2740_), .D(new_n5029_), .Y(new_n29613_));
  NOR2X1   g27177(.A(new_n29613_), .B(new_n29605_), .Y(new_n29614_));
  AND2X1   g27178(.A(new_n29611_), .B(new_n16243_), .Y(new_n29615_));
  NOR4X1   g27179(.A(new_n29615_), .B(new_n29614_), .C(new_n12641_), .D(new_n12618_), .Y(new_n29616_));
  OAI21X1  g27180(.A0(new_n29616_), .A1(new_n29612_), .B0(new_n12842_), .Y(new_n29617_));
  NOR4X1   g27181(.A(new_n29611_), .B(new_n29606_), .C(new_n12767_), .D(new_n12690_), .Y(new_n29618_));
  NOR4X1   g27182(.A(new_n29614_), .B(new_n12659_), .C(new_n12641_), .D(new_n12618_), .Y(new_n29619_));
  AOI21X1  g27183(.A0(new_n29619_), .A1(pi0641), .B0(new_n29605_), .Y(new_n29620_));
  AOI21X1  g27184(.A0(new_n29619_), .A1(new_n12672_), .B0(new_n29605_), .Y(new_n29621_));
  OAI22X1  g27185(.A0(new_n29621_), .A1(new_n23014_), .B0(new_n29620_), .B1(new_n23011_), .Y(new_n29622_));
  OAI21X1  g27186(.A0(new_n29622_), .A1(new_n29618_), .B0(pi0788), .Y(new_n29623_));
  AOI21X1  g27187(.A0(new_n29623_), .A1(new_n29617_), .B0(new_n14273_), .Y(new_n29624_));
  MX2X1    g27188(.A(new_n29612_), .B(new_n29605_), .S0(new_n12841_), .Y(new_n29625_));
  NAND2X1  g27189(.A(new_n29625_), .B(new_n12867_), .Y(new_n29626_));
  INVX1    g27190(.A(new_n29605_), .Y(new_n29627_));
  OR2X1    g27191(.A(new_n29614_), .B(new_n13624_), .Y(new_n29628_));
  OAI21X1  g27192(.A0(new_n29628_), .A1(new_n12683_), .B0(new_n29627_), .Y(new_n29629_));
  AOI21X1  g27193(.A0(new_n29629_), .A1(pi1156), .B0(pi0629), .Y(new_n29630_));
  NAND2X1  g27194(.A(new_n29630_), .B(new_n29626_), .Y(new_n29631_));
  NAND2X1  g27195(.A(new_n29625_), .B(new_n12865_), .Y(new_n29632_));
  OAI21X1  g27196(.A0(new_n29628_), .A1(pi0628), .B0(new_n29627_), .Y(new_n29633_));
  AOI21X1  g27197(.A0(new_n29633_), .A1(new_n12684_), .B0(new_n12689_), .Y(new_n29634_));
  AOI21X1  g27198(.A0(new_n29634_), .A1(new_n29632_), .B0(new_n11884_), .Y(new_n29635_));
  AOI21X1  g27199(.A0(new_n29635_), .A1(new_n29631_), .B0(new_n29624_), .Y(new_n29636_));
  MX2X1    g27200(.A(new_n29625_), .B(new_n29605_), .S0(new_n12711_), .Y(new_n29637_));
  AOI21X1  g27201(.A0(new_n29637_), .A1(pi0647), .B0(pi1157), .Y(new_n29638_));
  OAI21X1  g27202(.A0(new_n29636_), .A1(pi0647), .B0(new_n29638_), .Y(new_n29639_));
  OR4X1    g27203(.A(new_n29614_), .B(new_n13639_), .C(new_n13624_), .D(new_n12705_), .Y(new_n29640_));
  NOR2X1   g27204(.A(new_n29605_), .B(new_n12706_), .Y(new_n29641_));
  AOI21X1  g27205(.A0(new_n29641_), .A1(new_n29640_), .B0(pi0630), .Y(new_n29642_));
  AOI21X1  g27206(.A0(new_n29637_), .A1(new_n12705_), .B0(new_n12706_), .Y(new_n29643_));
  OAI21X1  g27207(.A0(new_n29636_), .A1(new_n12705_), .B0(new_n29643_), .Y(new_n29644_));
  OR4X1    g27208(.A(new_n29614_), .B(new_n13639_), .C(new_n13624_), .D(pi0647), .Y(new_n29645_));
  NOR2X1   g27209(.A(new_n29605_), .B(pi1157), .Y(new_n29646_));
  AOI21X1  g27210(.A0(new_n29646_), .A1(new_n29645_), .B0(new_n12723_), .Y(new_n29647_));
  AOI22X1  g27211(.A0(new_n29647_), .A1(new_n29644_), .B0(new_n29642_), .B1(new_n29639_), .Y(new_n29648_));
  MX2X1    g27212(.A(new_n29648_), .B(new_n29636_), .S0(new_n11883_), .Y(new_n29649_));
  NOR4X1   g27213(.A(new_n29614_), .B(new_n13651_), .C(new_n13639_), .D(new_n13624_), .Y(new_n29650_));
  OR2X1    g27214(.A(new_n29650_), .B(new_n29605_), .Y(new_n29651_));
  AOI21X1  g27215(.A0(new_n29651_), .A1(pi0644), .B0(pi0715), .Y(new_n29652_));
  OAI21X1  g27216(.A0(new_n29649_), .A1(pi0644), .B0(new_n29652_), .Y(new_n29653_));
  NAND4X1  g27217(.A(new_n29625_), .B(new_n12736_), .C(new_n14123_), .D(new_n12743_), .Y(new_n29654_));
  NAND3X1  g27218(.A(new_n29654_), .B(new_n29627_), .C(pi0715), .Y(new_n29655_));
  AOI21X1  g27219(.A0(new_n29655_), .A1(new_n29653_), .B0(pi1160), .Y(new_n29656_));
  OAI21X1  g27220(.A0(new_n29651_), .A1(pi0644), .B0(pi0715), .Y(new_n29657_));
  AOI21X1  g27221(.A0(new_n29649_), .A1(pi0644), .B0(new_n29657_), .Y(new_n29658_));
  NAND4X1  g27222(.A(new_n29625_), .B(new_n12736_), .C(new_n14123_), .D(pi0644), .Y(new_n29659_));
  AOI21X1  g27223(.A0(new_n29659_), .A1(new_n29627_), .B0(pi0715), .Y(new_n29660_));
  OR2X1    g27224(.A(new_n29660_), .B(new_n11882_), .Y(new_n29661_));
  OAI21X1  g27225(.A0(new_n29661_), .A1(new_n29658_), .B0(pi0790), .Y(new_n29662_));
  OAI22X1  g27226(.A0(new_n29662_), .A1(new_n29656_), .B0(new_n29649_), .B1(pi0790), .Y(new_n29663_));
  MX2X1    g27227(.A(new_n29663_), .B(new_n29603_), .S0(new_n24954_), .Y(po0724));
  MX2X1    g27228(.A(pi0568), .B(pi0245), .S0(new_n22728_), .Y(po0725));
  INVX1    g27229(.A(pi0569), .Y(new_n29666_));
  MX2X1    g27230(.A(new_n29666_), .B(pi0239), .S0(new_n22728_), .Y(po0726));
  INVX1    g27231(.A(pi0570), .Y(new_n29668_));
  AND2X1   g27232(.A(new_n29528_), .B(new_n22728_), .Y(new_n29669_));
  NAND2X1  g27233(.A(new_n22725_), .B(new_n29668_), .Y(new_n29670_));
  OAI22X1  g27234(.A0(new_n29670_), .A1(new_n29539_), .B0(new_n29669_), .B1(new_n29668_), .Y(po0727));
  MX2X1    g27235(.A(pi0571), .B(pi0241), .S0(new_n23553_), .Y(po0728));
  MX2X1    g27236(.A(pi0572), .B(pi0244), .S0(new_n23553_), .Y(po0729));
  MX2X1    g27237(.A(pi0573), .B(pi0242), .S0(new_n23553_), .Y(po0730));
  MX2X1    g27238(.A(pi0574), .B(pi0241), .S0(new_n22722_), .Y(po0731));
  MX2X1    g27239(.A(pi0575), .B(pi0235), .S0(new_n23553_), .Y(po0732));
  MX2X1    g27240(.A(pi0576), .B(pi0248), .S0(new_n23553_), .Y(po0733));
  MX2X1    g27241(.A(pi0577), .B(pi0238), .S0(new_n23537_), .Y(po0734));
  MX2X1    g27242(.A(pi0578), .B(pi0249), .S0(new_n22722_), .Y(po0735));
  MX2X1    g27243(.A(pi0579), .B(pi0249), .S0(new_n22715_), .Y(po0736));
  MX2X1    g27244(.A(pi0580), .B(pi0245), .S0(new_n23537_), .Y(po0737));
  MX2X1    g27245(.A(pi0581), .B(pi0235), .S0(new_n22722_), .Y(po0738));
  MX2X1    g27246(.A(pi0582), .B(pi0240), .S0(new_n22722_), .Y(po0739));
  MX2X1    g27247(.A(pi0584), .B(pi0245), .S0(new_n22722_), .Y(po0741));
  MX2X1    g27248(.A(pi0585), .B(pi0244), .S0(new_n22722_), .Y(po0742));
  MX2X1    g27249(.A(pi0586), .B(pi0242), .S0(new_n22722_), .Y(po0743));
  OR4X1    g27250(.A(new_n23246_), .B(new_n14178_), .C(new_n12171_), .D(new_n24954_), .Y(new_n29687_));
  OR4X1    g27251(.A(new_n29687_), .B(new_n16294_), .C(new_n14185_), .D(new_n12841_), .Y(new_n29688_));
  OAI21X1  g27252(.A0(new_n22667_), .A1(pi0230), .B0(new_n29688_), .Y(po0744));
  NAND2X1  g27253(.A(new_n9046_), .B(new_n28068_), .Y(new_n29690_));
  OAI21X1  g27254(.A0(new_n29690_), .A1(pi0591), .B0(new_n29197_), .Y(new_n29691_));
  AOI21X1  g27255(.A0(new_n29690_), .A1(new_n9028_), .B0(new_n29691_), .Y(po0745));
  INVX1    g27256(.A(new_n29516_), .Y(new_n29693_));
  OR2X1    g27257(.A(new_n29693_), .B(pi0204), .Y(new_n29694_));
  NOR2X1   g27258(.A(new_n29527_), .B(new_n22714_), .Y(new_n29695_));
  AOI21X1  g27259(.A0(new_n29695_), .A1(new_n22588_), .B0(new_n22718_), .Y(new_n29696_));
  OR2X1    g27260(.A(new_n29693_), .B(pi0205), .Y(new_n29697_));
  AOI21X1  g27261(.A0(new_n29695_), .A1(new_n22717_), .B0(pi0233), .Y(new_n29698_));
  AOI22X1  g27262(.A0(new_n29698_), .A1(new_n29697_), .B0(new_n29696_), .B1(new_n29694_), .Y(new_n29699_));
  OR2X1    g27263(.A(new_n29693_), .B(pi0206), .Y(new_n29700_));
  AOI21X1  g27264(.A0(new_n29695_), .A1(new_n23551_), .B0(new_n22718_), .Y(new_n29701_));
  OR2X1    g27265(.A(new_n29693_), .B(pi0218), .Y(new_n29702_));
  AOI21X1  g27266(.A0(new_n29695_), .A1(new_n22724_), .B0(pi0233), .Y(new_n29703_));
  AOI22X1  g27267(.A0(new_n29703_), .A1(new_n29702_), .B0(new_n29701_), .B1(new_n29700_), .Y(new_n29704_));
  MX2X1    g27268(.A(new_n29704_), .B(new_n29699_), .S0(pi0237), .Y(po0746));
  NOR4X1   g27269(.A(new_n5096_), .B(new_n5251_), .C(new_n9028_), .D(pi0123), .Y(new_n29706_));
  AOI21X1  g27270(.A0(new_n9046_), .A1(new_n28068_), .B0(new_n6168_), .Y(new_n29707_));
  OR4X1    g27271(.A(new_n29707_), .B(new_n29706_), .C(new_n2781_), .D(new_n2755_), .Y(po0747));
  OAI21X1  g27272(.A0(new_n29690_), .A1(pi0592), .B0(new_n29197_), .Y(new_n29709_));
  AOI21X1  g27273(.A0(new_n29690_), .A1(new_n6074_), .B0(new_n29709_), .Y(po0748));
  OAI21X1  g27274(.A0(new_n29690_), .A1(pi0590), .B0(new_n29197_), .Y(new_n29711_));
  AOI21X1  g27275(.A0(new_n29690_), .A1(new_n6120_), .B0(new_n29711_), .Y(po0749));
  INVX1    g27276(.A(pi0517), .Y(new_n29713_));
  INVX1    g27277(.A(pi0509), .Y(new_n29714_));
  INVX1    g27278(.A(pi0533), .Y(new_n29715_));
  INVX1    g27279(.A(pi0537), .Y(new_n29716_));
  INVX1    g27280(.A(pi0249), .Y(new_n29717_));
  AOI21X1  g27281(.A0(new_n29516_), .A1(new_n2990_), .B0(pi0557), .Y(new_n29718_));
  AOI21X1  g27282(.A0(new_n29516_), .A1(pi0234), .B0(new_n29590_), .Y(new_n29719_));
  XOR2X1   g27283(.A(pi0536), .B(pi0246), .Y(new_n29720_));
  NOR4X1   g27284(.A(new_n29720_), .B(new_n29719_), .C(new_n29718_), .D(pi0538), .Y(new_n29721_));
  INVX1    g27285(.A(pi0538), .Y(new_n29722_));
  NOR4X1   g27286(.A(new_n29720_), .B(new_n29719_), .C(new_n29718_), .D(new_n29722_), .Y(new_n29723_));
  MX2X1    g27287(.A(new_n29723_), .B(new_n29721_), .S0(new_n29717_), .Y(new_n29724_));
  AOI21X1  g27288(.A0(new_n29724_), .A1(new_n29716_), .B0(pi0248), .Y(new_n29725_));
  INVX1    g27289(.A(pi0248), .Y(new_n29726_));
  AOI21X1  g27290(.A0(new_n29724_), .A1(pi0537), .B0(new_n29726_), .Y(new_n29727_));
  NOR2X1   g27291(.A(new_n29727_), .B(new_n29725_), .Y(new_n29728_));
  INVX1    g27292(.A(pi0241), .Y(new_n29729_));
  XOR2X1   g27293(.A(pi0506), .B(new_n29729_), .Y(new_n29730_));
  NAND2X1  g27294(.A(new_n29730_), .B(new_n29728_), .Y(new_n29731_));
  XOR2X1   g27295(.A(pi0535), .B(pi0240), .Y(new_n29732_));
  NOR3X1   g27296(.A(new_n29732_), .B(new_n29731_), .C(new_n29562_), .Y(new_n29733_));
  NOR3X1   g27297(.A(new_n29732_), .B(new_n29731_), .C(pi0534), .Y(new_n29734_));
  MX2X1    g27298(.A(new_n29734_), .B(new_n29733_), .S0(new_n3253_), .Y(new_n29735_));
  AOI21X1  g27299(.A0(new_n29735_), .A1(pi0504), .B0(new_n4894_), .Y(new_n29736_));
  INVX1    g27300(.A(pi0504), .Y(new_n29737_));
  AOI21X1  g27301(.A0(new_n29735_), .A1(new_n29737_), .B0(pi0242), .Y(new_n29738_));
  NOR3X1   g27302(.A(new_n29738_), .B(new_n29736_), .C(new_n29715_), .Y(new_n29739_));
  NOR3X1   g27303(.A(new_n29738_), .B(new_n29736_), .C(pi0533), .Y(new_n29740_));
  MX2X1    g27304(.A(new_n29740_), .B(new_n29739_), .S0(pi0235), .Y(new_n29741_));
  AOI21X1  g27305(.A0(new_n29741_), .A1(pi0558), .B0(new_n4697_), .Y(new_n29742_));
  INVX1    g27306(.A(pi0558), .Y(new_n29743_));
  AOI21X1  g27307(.A0(new_n29741_), .A1(new_n29743_), .B0(pi0244), .Y(new_n29744_));
  NOR3X1   g27308(.A(new_n29744_), .B(new_n29742_), .C(new_n29714_), .Y(new_n29745_));
  NOR3X1   g27309(.A(new_n29744_), .B(new_n29742_), .C(pi0509), .Y(new_n29746_));
  MX2X1    g27310(.A(new_n29746_), .B(new_n29745_), .S0(pi0245), .Y(new_n29747_));
  AOI21X1  g27311(.A0(new_n29747_), .A1(pi0508), .B0(new_n4117_), .Y(new_n29748_));
  INVX1    g27312(.A(pi0508), .Y(new_n29749_));
  NOR2X1   g27313(.A(new_n29745_), .B(new_n4550_), .Y(new_n29750_));
  NOR2X1   g27314(.A(new_n29739_), .B(new_n3392_), .Y(new_n29751_));
  NOR2X1   g27315(.A(new_n29733_), .B(pi0239), .Y(new_n29752_));
  INVX1    g27316(.A(pi0240), .Y(new_n29753_));
  XOR2X1   g27317(.A(pi0481), .B(pi0248), .Y(new_n29754_));
  INVX1    g27318(.A(pi0511), .Y(new_n29755_));
  NOR3X1   g27319(.A(new_n29527_), .B(new_n22714_), .C(new_n2990_), .Y(new_n29756_));
  INVX1    g27320(.A(pi0246), .Y(new_n29757_));
  XOR2X1   g27321(.A(pi0487), .B(new_n29757_), .Y(new_n29758_));
  OAI21X1  g27322(.A0(new_n29756_), .A1(new_n29755_), .B0(new_n29758_), .Y(new_n29759_));
  AOI21X1  g27323(.A0(new_n29529_), .A1(new_n29755_), .B0(new_n29759_), .Y(new_n29760_));
  XOR2X1   g27324(.A(pi0579), .B(new_n29717_), .Y(new_n29761_));
  NAND2X1  g27325(.A(new_n29761_), .B(new_n29760_), .Y(new_n29762_));
  NOR2X1   g27326(.A(new_n29762_), .B(new_n29754_), .Y(new_n29763_));
  AOI21X1  g27327(.A0(new_n29763_), .A1(pi0559), .B0(new_n29729_), .Y(new_n29764_));
  INVX1    g27328(.A(pi0559), .Y(new_n29765_));
  AOI21X1  g27329(.A0(new_n29763_), .A1(new_n29765_), .B0(pi0241), .Y(new_n29766_));
  NOR2X1   g27330(.A(new_n29766_), .B(new_n29764_), .Y(new_n29767_));
  AOI21X1  g27331(.A0(new_n29767_), .A1(pi0515), .B0(new_n29753_), .Y(new_n29768_));
  INVX1    g27332(.A(pi0515), .Y(new_n29769_));
  AOI21X1  g27333(.A0(new_n29760_), .A1(new_n29717_), .B0(pi0579), .Y(new_n29770_));
  OAI21X1  g27334(.A0(new_n29721_), .A1(pi0249), .B0(new_n29760_), .Y(new_n29771_));
  AOI21X1  g27335(.A0(new_n29771_), .A1(pi0579), .B0(new_n29770_), .Y(new_n29772_));
  OR2X1    g27336(.A(new_n29772_), .B(new_n29724_), .Y(new_n29773_));
  OAI21X1  g27337(.A0(new_n29762_), .A1(new_n29716_), .B0(new_n29726_), .Y(new_n29774_));
  AOI21X1  g27338(.A0(new_n29773_), .A1(new_n29716_), .B0(new_n29774_), .Y(new_n29775_));
  OR2X1    g27339(.A(new_n29775_), .B(new_n29727_), .Y(new_n29776_));
  OAI21X1  g27340(.A0(new_n29762_), .A1(pi0537), .B0(pi0248), .Y(new_n29777_));
  AOI21X1  g27341(.A0(new_n29773_), .A1(pi0537), .B0(new_n29777_), .Y(new_n29778_));
  OR2X1    g27342(.A(new_n29778_), .B(new_n29725_), .Y(new_n29779_));
  MX2X1    g27343(.A(new_n29776_), .B(new_n29779_), .S0(pi0481), .Y(new_n29780_));
  OR2X1    g27344(.A(new_n29780_), .B(pi0559), .Y(new_n29781_));
  AOI21X1  g27345(.A0(new_n29728_), .A1(pi0559), .B0(pi0241), .Y(new_n29782_));
  AOI21X1  g27346(.A0(new_n29782_), .A1(new_n29781_), .B0(new_n29764_), .Y(new_n29783_));
  OR2X1    g27347(.A(new_n29780_), .B(new_n29765_), .Y(new_n29784_));
  AOI21X1  g27348(.A0(new_n29728_), .A1(new_n29765_), .B0(new_n29729_), .Y(new_n29785_));
  AOI21X1  g27349(.A0(new_n29785_), .A1(new_n29784_), .B0(new_n29766_), .Y(new_n29786_));
  MX2X1    g27350(.A(new_n29783_), .B(new_n29786_), .S0(pi0506), .Y(new_n29787_));
  OAI21X1  g27351(.A0(new_n29731_), .A1(new_n29769_), .B0(new_n29753_), .Y(new_n29788_));
  AOI21X1  g27352(.A0(new_n29787_), .A1(new_n29769_), .B0(new_n29788_), .Y(new_n29789_));
  OR2X1    g27353(.A(new_n29789_), .B(new_n29768_), .Y(new_n29790_));
  AOI21X1  g27354(.A0(new_n29767_), .A1(new_n29769_), .B0(pi0240), .Y(new_n29791_));
  OAI21X1  g27355(.A0(new_n29731_), .A1(pi0515), .B0(pi0240), .Y(new_n29792_));
  AOI21X1  g27356(.A0(new_n29787_), .A1(pi0515), .B0(new_n29792_), .Y(new_n29793_));
  OR2X1    g27357(.A(new_n29793_), .B(new_n29791_), .Y(new_n29794_));
  MX2X1    g27358(.A(new_n29790_), .B(new_n29794_), .S0(pi0535), .Y(new_n29795_));
  OR2X1    g27359(.A(new_n29795_), .B(pi0534), .Y(new_n29796_));
  NOR2X1   g27360(.A(new_n29791_), .B(new_n29768_), .Y(new_n29797_));
  AOI21X1  g27361(.A0(new_n29797_), .A1(pi0534), .B0(new_n3253_), .Y(new_n29798_));
  AOI21X1  g27362(.A0(new_n29798_), .A1(new_n29796_), .B0(new_n29752_), .Y(new_n29799_));
  NOR2X1   g27363(.A(new_n29734_), .B(new_n3253_), .Y(new_n29800_));
  OR2X1    g27364(.A(new_n29795_), .B(new_n29562_), .Y(new_n29801_));
  AOI21X1  g27365(.A0(new_n29797_), .A1(new_n29562_), .B0(pi0239), .Y(new_n29802_));
  AOI21X1  g27366(.A0(new_n29802_), .A1(new_n29801_), .B0(new_n29800_), .Y(new_n29803_));
  MX2X1    g27367(.A(new_n29803_), .B(new_n29799_), .S0(new_n29495_), .Y(new_n29804_));
  XOR2X1   g27368(.A(pi0488), .B(pi0239), .Y(new_n29805_));
  NAND2X1  g27369(.A(new_n29805_), .B(new_n29797_), .Y(new_n29806_));
  OAI21X1  g27370(.A0(new_n29806_), .A1(new_n29737_), .B0(new_n4894_), .Y(new_n29807_));
  AOI21X1  g27371(.A0(new_n29804_), .A1(new_n29737_), .B0(new_n29807_), .Y(new_n29808_));
  OR2X1    g27372(.A(new_n29808_), .B(new_n29736_), .Y(new_n29809_));
  OAI21X1  g27373(.A0(new_n29806_), .A1(pi0504), .B0(pi0242), .Y(new_n29810_));
  AOI21X1  g27374(.A0(new_n29804_), .A1(pi0504), .B0(new_n29810_), .Y(new_n29811_));
  OR2X1    g27375(.A(new_n29811_), .B(new_n29738_), .Y(new_n29812_));
  MX2X1    g27376(.A(new_n29809_), .B(new_n29812_), .S0(pi0510), .Y(new_n29813_));
  OR2X1    g27377(.A(new_n29813_), .B(pi0533), .Y(new_n29814_));
  XOR2X1   g27378(.A(pi0510), .B(pi0242), .Y(new_n29815_));
  NOR2X1   g27379(.A(new_n29815_), .B(new_n29806_), .Y(new_n29816_));
  AOI21X1  g27380(.A0(new_n29816_), .A1(pi0533), .B0(pi0235), .Y(new_n29817_));
  AOI21X1  g27381(.A0(new_n29817_), .A1(new_n29814_), .B0(new_n29751_), .Y(new_n29818_));
  NOR2X1   g27382(.A(new_n29740_), .B(pi0235), .Y(new_n29819_));
  OR2X1    g27383(.A(new_n29813_), .B(new_n29715_), .Y(new_n29820_));
  AOI21X1  g27384(.A0(new_n29816_), .A1(new_n29715_), .B0(new_n3392_), .Y(new_n29821_));
  AOI21X1  g27385(.A0(new_n29821_), .A1(new_n29820_), .B0(new_n29819_), .Y(new_n29822_));
  MX2X1    g27386(.A(new_n29818_), .B(new_n29822_), .S0(pi0512), .Y(new_n29823_));
  XOR2X1   g27387(.A(pi0512), .B(pi0235), .Y(new_n29824_));
  NOR3X1   g27388(.A(new_n29824_), .B(new_n29815_), .C(new_n29806_), .Y(new_n29825_));
  INVX1    g27389(.A(new_n29825_), .Y(new_n29826_));
  OAI21X1  g27390(.A0(new_n29826_), .A1(new_n29743_), .B0(new_n4697_), .Y(new_n29827_));
  AOI21X1  g27391(.A0(new_n29823_), .A1(new_n29743_), .B0(new_n29827_), .Y(new_n29828_));
  OR2X1    g27392(.A(new_n29828_), .B(new_n29742_), .Y(new_n29829_));
  OAI21X1  g27393(.A0(new_n29826_), .A1(pi0558), .B0(pi0244), .Y(new_n29830_));
  AOI21X1  g27394(.A0(new_n29823_), .A1(pi0558), .B0(new_n29830_), .Y(new_n29831_));
  OR2X1    g27395(.A(new_n29831_), .B(new_n29744_), .Y(new_n29832_));
  MX2X1    g27396(.A(new_n29829_), .B(new_n29832_), .S0(pi0513), .Y(new_n29833_));
  OR2X1    g27397(.A(new_n29833_), .B(pi0509), .Y(new_n29834_));
  XOR2X1   g27398(.A(pi0513), .B(pi0244), .Y(new_n29835_));
  NOR4X1   g27399(.A(new_n29835_), .B(new_n29824_), .C(new_n29815_), .D(new_n29806_), .Y(new_n29836_));
  AOI21X1  g27400(.A0(new_n29836_), .A1(pi0509), .B0(pi0245), .Y(new_n29837_));
  AOI21X1  g27401(.A0(new_n29837_), .A1(new_n29834_), .B0(new_n29750_), .Y(new_n29838_));
  NOR2X1   g27402(.A(new_n29746_), .B(pi0245), .Y(new_n29839_));
  OR2X1    g27403(.A(new_n29833_), .B(new_n29714_), .Y(new_n29840_));
  AOI21X1  g27404(.A0(new_n29836_), .A1(new_n29714_), .B0(new_n4550_), .Y(new_n29841_));
  AOI21X1  g27405(.A0(new_n29841_), .A1(new_n29840_), .B0(new_n29839_), .Y(new_n29842_));
  MX2X1    g27406(.A(new_n29838_), .B(new_n29842_), .S0(pi0514), .Y(new_n29843_));
  XOR2X1   g27407(.A(pi0514), .B(new_n4550_), .Y(new_n29844_));
  NAND2X1  g27408(.A(new_n29844_), .B(new_n29836_), .Y(new_n29845_));
  OAI21X1  g27409(.A0(new_n29845_), .A1(new_n29749_), .B0(new_n4117_), .Y(new_n29846_));
  AOI21X1  g27410(.A0(new_n29843_), .A1(new_n29749_), .B0(new_n29846_), .Y(new_n29847_));
  OR2X1    g27411(.A(new_n29847_), .B(new_n29748_), .Y(new_n29848_));
  AOI21X1  g27412(.A0(new_n29747_), .A1(new_n29749_), .B0(pi0247), .Y(new_n29849_));
  OAI21X1  g27413(.A0(new_n29845_), .A1(pi0508), .B0(pi0247), .Y(new_n29850_));
  AOI21X1  g27414(.A0(new_n29843_), .A1(pi0508), .B0(new_n29850_), .Y(new_n29851_));
  OR2X1    g27415(.A(new_n29851_), .B(new_n29849_), .Y(new_n29852_));
  MX2X1    g27416(.A(new_n29848_), .B(new_n29852_), .S0(pi0516), .Y(new_n29853_));
  OAI21X1  g27417(.A0(new_n29853_), .A1(pi0238), .B0(new_n29713_), .Y(new_n29854_));
  NOR3X1   g27418(.A(new_n29849_), .B(new_n29748_), .C(pi0238), .Y(new_n29855_));
  XOR2X1   g27419(.A(pi0516), .B(new_n4117_), .Y(new_n29856_));
  NAND3X1  g27420(.A(new_n29856_), .B(new_n29844_), .C(new_n29836_), .Y(new_n29857_));
  OAI21X1  g27421(.A0(new_n29857_), .A1(new_n3578_), .B0(pi0517), .Y(new_n29858_));
  NOR2X1   g27422(.A(new_n29858_), .B(new_n29855_), .Y(new_n29859_));
  NOR2X1   g27423(.A(new_n29859_), .B(pi0507), .Y(new_n29860_));
  AND2X1   g27424(.A(new_n29860_), .B(new_n29854_), .Y(new_n29861_));
  OR2X1    g27425(.A(new_n29853_), .B(new_n3578_), .Y(new_n29862_));
  NOR3X1   g27426(.A(new_n29849_), .B(new_n29748_), .C(new_n3578_), .Y(new_n29863_));
  OAI21X1  g27427(.A0(new_n29857_), .A1(pi0238), .B0(new_n29713_), .Y(new_n29864_));
  OAI21X1  g27428(.A0(new_n29864_), .A1(new_n29863_), .B0(pi0507), .Y(new_n29865_));
  AOI21X1  g27429(.A0(new_n29862_), .A1(pi0517), .B0(new_n29865_), .Y(new_n29866_));
  OAI21X1  g27430(.A0(new_n29866_), .A1(new_n29861_), .B0(pi0233), .Y(new_n29867_));
  XOR2X1   g27431(.A(pi0542), .B(new_n29753_), .Y(new_n29868_));
  AOI21X1  g27432(.A0(new_n29516_), .A1(pi0234), .B0(new_n29515_), .Y(new_n29869_));
  AOI21X1  g27433(.A0(new_n29516_), .A1(new_n2990_), .B0(pi0505), .Y(new_n29870_));
  XOR2X1   g27434(.A(pi0501), .B(new_n29726_), .Y(new_n29871_));
  XOR2X1   g27435(.A(pi0499), .B(new_n29757_), .Y(new_n29872_));
  XOR2X1   g27436(.A(pi0496), .B(new_n29717_), .Y(new_n29873_));
  NAND3X1  g27437(.A(new_n29873_), .B(new_n29872_), .C(new_n29871_), .Y(new_n29874_));
  XOR2X1   g27438(.A(pi0500), .B(pi0241), .Y(new_n29875_));
  NOR4X1   g27439(.A(new_n29875_), .B(new_n29874_), .C(new_n29870_), .D(new_n29869_), .Y(new_n29876_));
  AND2X1   g27440(.A(new_n29876_), .B(new_n29868_), .Y(new_n29877_));
  AOI21X1  g27441(.A0(new_n29877_), .A1(pi0497), .B0(pi0239), .Y(new_n29878_));
  AOI21X1  g27442(.A0(new_n29877_), .A1(new_n29506_), .B0(new_n3253_), .Y(new_n29879_));
  NOR2X1   g27443(.A(new_n29879_), .B(new_n29878_), .Y(new_n29880_));
  AOI21X1  g27444(.A0(new_n29880_), .A1(pi0539), .B0(new_n4894_), .Y(new_n29881_));
  INVX1    g27445(.A(pi0539), .Y(new_n29882_));
  AOI21X1  g27446(.A0(new_n29880_), .A1(new_n29882_), .B0(pi0242), .Y(new_n29883_));
  NOR2X1   g27447(.A(new_n29883_), .B(new_n29881_), .Y(new_n29884_));
  AOI21X1  g27448(.A0(new_n29884_), .A1(pi0540), .B0(new_n3392_), .Y(new_n29885_));
  INVX1    g27449(.A(pi0540), .Y(new_n29886_));
  AOI21X1  g27450(.A0(new_n29884_), .A1(new_n29886_), .B0(pi0235), .Y(new_n29887_));
  NOR2X1   g27451(.A(new_n29887_), .B(new_n29885_), .Y(new_n29888_));
  XOR2X1   g27452(.A(pi0541), .B(new_n4697_), .Y(new_n29889_));
  NAND2X1  g27453(.A(new_n29889_), .B(new_n29888_), .Y(new_n29890_));
  XOR2X1   g27454(.A(pi0503), .B(pi0245), .Y(new_n29891_));
  NOR3X1   g27455(.A(new_n29891_), .B(new_n29890_), .C(pi0502), .Y(new_n29892_));
  AOI21X1  g27456(.A0(new_n29892_), .A1(pi0561), .B0(pi0247), .Y(new_n29893_));
  INVX1    g27457(.A(pi0585), .Y(new_n29894_));
  NOR2X1   g27458(.A(new_n29756_), .B(new_n29537_), .Y(new_n29895_));
  XOR2X1   g27459(.A(pi0521), .B(pi0248), .Y(new_n29896_));
  XOR2X1   g27460(.A(pi0520), .B(pi0246), .Y(new_n29897_));
  XOR2X1   g27461(.A(pi0574), .B(pi0241), .Y(new_n29898_));
  XOR2X1   g27462(.A(pi0578), .B(pi0249), .Y(new_n29899_));
  NOR4X1   g27463(.A(new_n29899_), .B(new_n29898_), .C(new_n29897_), .D(new_n29896_), .Y(new_n29900_));
  OAI21X1  g27464(.A0(new_n29528_), .A1(pi0518), .B0(new_n29900_), .Y(new_n29901_));
  NOR2X1   g27465(.A(new_n29901_), .B(new_n29895_), .Y(new_n29902_));
  AOI21X1  g27466(.A0(new_n29902_), .A1(pi0582), .B0(new_n29753_), .Y(new_n29903_));
  INVX1    g27467(.A(pi0582), .Y(new_n29904_));
  AOI21X1  g27468(.A0(new_n29902_), .A1(new_n29904_), .B0(pi0240), .Y(new_n29905_));
  XOR2X1   g27469(.A(pi0519), .B(new_n3253_), .Y(new_n29906_));
  XOR2X1   g27470(.A(pi0586), .B(pi0242), .Y(new_n29907_));
  OR4X1    g27471(.A(new_n29907_), .B(new_n29906_), .C(new_n29905_), .D(new_n29903_), .Y(new_n29908_));
  XOR2X1   g27472(.A(pi0581), .B(pi0235), .Y(new_n29909_));
  NOR3X1   g27473(.A(new_n29909_), .B(new_n29908_), .C(new_n29894_), .Y(new_n29910_));
  NOR3X1   g27474(.A(new_n29909_), .B(new_n29908_), .C(pi0585), .Y(new_n29911_));
  MX2X1    g27475(.A(new_n29911_), .B(new_n29910_), .S0(pi0244), .Y(new_n29912_));
  AOI21X1  g27476(.A0(new_n29912_), .A1(pi0584), .B0(new_n4550_), .Y(new_n29913_));
  INVX1    g27477(.A(pi0584), .Y(new_n29914_));
  NOR2X1   g27478(.A(new_n29910_), .B(new_n4697_), .Y(new_n29915_));
  INVX1    g27479(.A(pi0500), .Y(new_n29916_));
  NAND2X1  g27480(.A(pi0500), .B(pi0241), .Y(new_n29917_));
  OR4X1    g27481(.A(new_n29917_), .B(new_n29874_), .C(new_n29870_), .D(new_n29869_), .Y(new_n29918_));
  OAI21X1  g27482(.A0(new_n29901_), .A1(new_n29895_), .B0(new_n29918_), .Y(new_n29919_));
  AOI21X1  g27483(.A0(new_n29876_), .A1(new_n29916_), .B0(new_n29919_), .Y(new_n29920_));
  OR2X1    g27484(.A(new_n29920_), .B(pi0582), .Y(new_n29921_));
  AOI21X1  g27485(.A0(new_n29876_), .A1(pi0582), .B0(pi0240), .Y(new_n29922_));
  AOI21X1  g27486(.A0(new_n29922_), .A1(new_n29921_), .B0(new_n29903_), .Y(new_n29923_));
  OR2X1    g27487(.A(new_n29920_), .B(new_n29904_), .Y(new_n29924_));
  AOI21X1  g27488(.A0(new_n29876_), .A1(new_n29904_), .B0(new_n29753_), .Y(new_n29925_));
  AOI21X1  g27489(.A0(new_n29925_), .A1(new_n29924_), .B0(new_n29905_), .Y(new_n29926_));
  MX2X1    g27490(.A(new_n29923_), .B(new_n29926_), .S0(pi0542), .Y(new_n29927_));
  OR2X1    g27491(.A(new_n29905_), .B(new_n29903_), .Y(new_n29928_));
  OAI21X1  g27492(.A0(new_n29928_), .A1(new_n29506_), .B0(pi0239), .Y(new_n29929_));
  AOI21X1  g27493(.A0(new_n29927_), .A1(new_n29506_), .B0(new_n29929_), .Y(new_n29930_));
  OAI21X1  g27494(.A0(new_n29930_), .A1(new_n29878_), .B0(new_n29542_), .Y(new_n29931_));
  OAI21X1  g27495(.A0(new_n29928_), .A1(pi0497), .B0(new_n3253_), .Y(new_n29932_));
  AOI21X1  g27496(.A0(new_n29927_), .A1(pi0497), .B0(new_n29932_), .Y(new_n29933_));
  OAI21X1  g27497(.A0(new_n29933_), .A1(new_n29879_), .B0(pi0519), .Y(new_n29934_));
  NAND3X1  g27498(.A(new_n29934_), .B(new_n29931_), .C(new_n29882_), .Y(new_n29935_));
  NOR3X1   g27499(.A(new_n29906_), .B(new_n29905_), .C(new_n29903_), .Y(new_n29936_));
  AOI21X1  g27500(.A0(new_n29936_), .A1(pi0539), .B0(pi0242), .Y(new_n29937_));
  AOI21X1  g27501(.A0(new_n29937_), .A1(new_n29935_), .B0(new_n29881_), .Y(new_n29938_));
  NAND3X1  g27502(.A(new_n29934_), .B(new_n29931_), .C(pi0539), .Y(new_n29939_));
  AOI21X1  g27503(.A0(new_n29936_), .A1(new_n29882_), .B0(new_n4894_), .Y(new_n29940_));
  AOI21X1  g27504(.A0(new_n29940_), .A1(new_n29939_), .B0(new_n29883_), .Y(new_n29941_));
  MX2X1    g27505(.A(new_n29938_), .B(new_n29941_), .S0(pi0586), .Y(new_n29942_));
  OAI21X1  g27506(.A0(new_n29908_), .A1(new_n29886_), .B0(new_n3392_), .Y(new_n29943_));
  AOI21X1  g27507(.A0(new_n29942_), .A1(new_n29886_), .B0(new_n29943_), .Y(new_n29944_));
  OR2X1    g27508(.A(new_n29944_), .B(new_n29885_), .Y(new_n29945_));
  OAI21X1  g27509(.A0(new_n29908_), .A1(pi0540), .B0(pi0235), .Y(new_n29946_));
  AOI21X1  g27510(.A0(new_n29942_), .A1(pi0540), .B0(new_n29946_), .Y(new_n29947_));
  OR2X1    g27511(.A(new_n29947_), .B(new_n29887_), .Y(new_n29948_));
  MX2X1    g27512(.A(new_n29945_), .B(new_n29948_), .S0(pi0581), .Y(new_n29949_));
  OR2X1    g27513(.A(new_n29949_), .B(pi0585), .Y(new_n29950_));
  AOI21X1  g27514(.A0(new_n29888_), .A1(pi0585), .B0(pi0244), .Y(new_n29951_));
  AOI21X1  g27515(.A0(new_n29951_), .A1(new_n29950_), .B0(new_n29915_), .Y(new_n29952_));
  NOR2X1   g27516(.A(new_n29911_), .B(pi0244), .Y(new_n29953_));
  OR2X1    g27517(.A(new_n29949_), .B(new_n29894_), .Y(new_n29954_));
  AOI21X1  g27518(.A0(new_n29888_), .A1(new_n29894_), .B0(new_n4697_), .Y(new_n29955_));
  AOI21X1  g27519(.A0(new_n29955_), .A1(new_n29954_), .B0(new_n29953_), .Y(new_n29956_));
  MX2X1    g27520(.A(new_n29952_), .B(new_n29956_), .S0(pi0541), .Y(new_n29957_));
  OAI21X1  g27521(.A0(new_n29890_), .A1(new_n29914_), .B0(new_n4550_), .Y(new_n29958_));
  AOI21X1  g27522(.A0(new_n29957_), .A1(new_n29914_), .B0(new_n29958_), .Y(new_n29959_));
  NOR2X1   g27523(.A(new_n29959_), .B(new_n29913_), .Y(new_n29960_));
  AOI21X1  g27524(.A0(new_n29912_), .A1(new_n29914_), .B0(pi0245), .Y(new_n29961_));
  OAI21X1  g27525(.A0(new_n29890_), .A1(pi0584), .B0(pi0245), .Y(new_n29962_));
  AOI21X1  g27526(.A0(new_n29957_), .A1(pi0584), .B0(new_n29962_), .Y(new_n29963_));
  NOR2X1   g27527(.A(new_n29963_), .B(new_n29961_), .Y(new_n29964_));
  MX2X1    g27528(.A(new_n29960_), .B(new_n29964_), .S0(pi0503), .Y(new_n29965_));
  NOR2X1   g27529(.A(new_n29961_), .B(new_n29913_), .Y(new_n29966_));
  INVX1    g27530(.A(new_n29966_), .Y(new_n29967_));
  AOI21X1  g27531(.A0(new_n29967_), .A1(pi0502), .B0(pi0561), .Y(new_n29968_));
  OAI21X1  g27532(.A0(new_n29965_), .A1(pi0502), .B0(new_n29968_), .Y(new_n29969_));
  INVX1    g27533(.A(pi0561), .Y(new_n29970_));
  INVX1    g27534(.A(pi0502), .Y(new_n29971_));
  NOR3X1   g27535(.A(new_n29891_), .B(new_n29890_), .C(new_n29971_), .Y(new_n29972_));
  AOI21X1  g27536(.A0(new_n29972_), .A1(new_n29970_), .B0(new_n4117_), .Y(new_n29973_));
  AOI21X1  g27537(.A0(new_n29967_), .A1(new_n29971_), .B0(new_n29970_), .Y(new_n29974_));
  OAI21X1  g27538(.A0(new_n29965_), .A1(new_n29971_), .B0(new_n29974_), .Y(new_n29975_));
  AOI22X1  g27539(.A0(new_n29975_), .A1(new_n29973_), .B0(new_n29969_), .B1(new_n29893_), .Y(new_n29976_));
  AOI21X1  g27540(.A0(new_n29976_), .A1(new_n3578_), .B0(pi0522), .Y(new_n29977_));
  MX2X1    g27541(.A(new_n29972_), .B(new_n29892_), .S0(new_n4117_), .Y(new_n29978_));
  XOR2X1   g27542(.A(pi0561), .B(new_n4117_), .Y(new_n29979_));
  NAND2X1  g27543(.A(new_n29979_), .B(new_n29966_), .Y(new_n29980_));
  OAI21X1  g27544(.A0(new_n29980_), .A1(new_n3578_), .B0(pi0522), .Y(new_n29981_));
  AOI21X1  g27545(.A0(new_n29978_), .A1(new_n3578_), .B0(new_n29981_), .Y(new_n29982_));
  OR2X1    g27546(.A(new_n29982_), .B(pi0543), .Y(new_n29983_));
  INVX1    g27547(.A(pi0522), .Y(new_n29984_));
  AOI21X1  g27548(.A0(new_n29976_), .A1(pi0238), .B0(new_n29984_), .Y(new_n29985_));
  AND2X1   g27549(.A(new_n29978_), .B(pi0238), .Y(new_n29986_));
  OAI21X1  g27550(.A0(new_n29980_), .A1(pi0238), .B0(new_n29984_), .Y(new_n29987_));
  OAI21X1  g27551(.A0(new_n29987_), .A1(new_n29986_), .B0(pi0543), .Y(new_n29988_));
  OAI22X1  g27552(.A0(new_n29988_), .A1(new_n29985_), .B0(new_n29983_), .B1(new_n29977_), .Y(new_n29989_));
  AOI21X1  g27553(.A0(new_n29989_), .A1(new_n22718_), .B0(new_n22797_), .Y(new_n29990_));
  XOR2X1   g27554(.A(pi0492), .B(pi0240), .Y(new_n29991_));
  XOR2X1   g27555(.A(pi0490), .B(pi0241), .Y(new_n29992_));
  AOI21X1  g27556(.A0(new_n29516_), .A1(pi0234), .B0(new_n29573_), .Y(new_n29993_));
  XOR2X1   g27557(.A(pi0484), .B(pi0249), .Y(new_n29994_));
  XOR2X1   g27558(.A(pi0546), .B(pi0246), .Y(new_n29995_));
  XOR2X1   g27559(.A(pi0548), .B(pi0248), .Y(new_n29996_));
  NOR4X1   g27560(.A(new_n29996_), .B(new_n29995_), .C(new_n29994_), .D(new_n29993_), .Y(new_n29997_));
  OAI21X1  g27561(.A0(new_n29517_), .A1(pi0544), .B0(new_n29997_), .Y(new_n29998_));
  NOR3X1   g27562(.A(new_n29998_), .B(new_n29992_), .C(new_n29991_), .Y(new_n29999_));
  AOI21X1  g27563(.A0(new_n29999_), .A1(pi0494), .B0(pi0239), .Y(new_n30000_));
  AOI21X1  g27564(.A0(new_n29999_), .A1(new_n29502_), .B0(new_n3253_), .Y(new_n30001_));
  NOR2X1   g27565(.A(new_n30001_), .B(new_n30000_), .Y(new_n30002_));
  AOI21X1  g27566(.A0(new_n30002_), .A1(pi0483), .B0(new_n4894_), .Y(new_n30003_));
  INVX1    g27567(.A(pi0483), .Y(new_n30004_));
  AOI21X1  g27568(.A0(new_n30002_), .A1(new_n30004_), .B0(pi0242), .Y(new_n30005_));
  NOR2X1   g27569(.A(new_n30005_), .B(new_n30003_), .Y(new_n30006_));
  AOI21X1  g27570(.A0(new_n30006_), .A1(pi0495), .B0(new_n3392_), .Y(new_n30007_));
  INVX1    g27571(.A(pi0495), .Y(new_n30008_));
  AOI21X1  g27572(.A0(new_n30006_), .A1(new_n30008_), .B0(pi0235), .Y(new_n30009_));
  XOR2X1   g27573(.A(pi0493), .B(pi0244), .Y(new_n30010_));
  NOR3X1   g27574(.A(new_n30010_), .B(new_n30009_), .C(new_n30007_), .Y(new_n30011_));
  AOI21X1  g27575(.A0(new_n30011_), .A1(pi0545), .B0(new_n4550_), .Y(new_n30012_));
  INVX1    g27576(.A(pi0545), .Y(new_n30013_));
  AOI21X1  g27577(.A0(new_n30011_), .A1(new_n30013_), .B0(pi0245), .Y(new_n30014_));
  NOR2X1   g27578(.A(new_n30014_), .B(new_n30012_), .Y(new_n30015_));
  AOI21X1  g27579(.A0(new_n30015_), .A1(pi0547), .B0(new_n4117_), .Y(new_n30016_));
  INVX1    g27580(.A(new_n30016_), .Y(new_n30017_));
  INVX1    g27581(.A(pi0571), .Y(new_n30018_));
  NOR2X1   g27582(.A(new_n29756_), .B(new_n29547_), .Y(new_n30019_));
  NOR2X1   g27583(.A(new_n29528_), .B(pi0523), .Y(new_n30020_));
  XOR2X1   g27584(.A(pi0528), .B(new_n29717_), .Y(new_n30021_));
  XOR2X1   g27585(.A(pi0526), .B(new_n29757_), .Y(new_n30022_));
  XOR2X1   g27586(.A(pi0576), .B(new_n29726_), .Y(new_n30023_));
  NAND3X1  g27587(.A(new_n30023_), .B(new_n30022_), .C(new_n30021_), .Y(new_n30024_));
  OR4X1    g27588(.A(new_n30024_), .B(new_n30020_), .C(new_n30019_), .D(new_n30018_), .Y(new_n30025_));
  OR4X1    g27589(.A(new_n30024_), .B(new_n30020_), .C(new_n30019_), .D(pi0571), .Y(new_n30026_));
  MX2X1    g27590(.A(new_n30026_), .B(new_n30025_), .S0(pi0241), .Y(new_n30027_));
  NOR2X1   g27591(.A(new_n30027_), .B(pi0530), .Y(new_n30028_));
  NOR2X1   g27592(.A(new_n30028_), .B(pi0240), .Y(new_n30029_));
  INVX1    g27593(.A(pi0530), .Y(new_n30030_));
  NOR2X1   g27594(.A(new_n30027_), .B(new_n30030_), .Y(new_n30031_));
  NOR2X1   g27595(.A(new_n30031_), .B(new_n29753_), .Y(new_n30032_));
  XOR2X1   g27596(.A(pi0524), .B(new_n3253_), .Y(new_n30033_));
  XOR2X1   g27597(.A(pi0573), .B(pi0242), .Y(new_n30034_));
  NOR4X1   g27598(.A(new_n30034_), .B(new_n30033_), .C(new_n30032_), .D(new_n30029_), .Y(new_n30035_));
  XOR2X1   g27599(.A(pi0575), .B(new_n3392_), .Y(new_n30036_));
  AND2X1   g27600(.A(new_n30036_), .B(new_n30035_), .Y(new_n30037_));
  AOI21X1  g27601(.A0(new_n30037_), .A1(pi0572), .B0(new_n4697_), .Y(new_n30038_));
  AOI21X1  g27602(.A0(new_n30028_), .A1(pi0492), .B0(pi0240), .Y(new_n30039_));
  AND2X1   g27603(.A(new_n29998_), .B(new_n29729_), .Y(new_n30040_));
  AOI22X1  g27604(.A0(new_n30040_), .A1(new_n30026_), .B0(new_n30025_), .B1(pi0241), .Y(new_n30041_));
  AND2X1   g27605(.A(new_n29998_), .B(pi0241), .Y(new_n30042_));
  AOI22X1  g27606(.A0(new_n30042_), .A1(new_n30025_), .B0(new_n30026_), .B1(new_n29729_), .Y(new_n30043_));
  MX2X1    g27607(.A(new_n30041_), .B(new_n30043_), .S0(pi0490), .Y(new_n30044_));
  NOR2X1   g27608(.A(new_n29998_), .B(new_n29992_), .Y(new_n30045_));
  INVX1    g27609(.A(new_n30045_), .Y(new_n30046_));
  AOI21X1  g27610(.A0(new_n30046_), .A1(pi0530), .B0(pi0492), .Y(new_n30047_));
  OAI21X1  g27611(.A0(new_n30044_), .A1(pi0530), .B0(new_n30047_), .Y(new_n30048_));
  INVX1    g27612(.A(pi0492), .Y(new_n30049_));
  AOI21X1  g27613(.A0(new_n30031_), .A1(new_n30049_), .B0(new_n29753_), .Y(new_n30050_));
  AOI21X1  g27614(.A0(new_n30046_), .A1(new_n30030_), .B0(new_n30049_), .Y(new_n30051_));
  OAI21X1  g27615(.A0(new_n30044_), .A1(new_n30030_), .B0(new_n30051_), .Y(new_n30052_));
  AOI22X1  g27616(.A0(new_n30052_), .A1(new_n30050_), .B0(new_n30048_), .B1(new_n30039_), .Y(new_n30053_));
  OR2X1    g27617(.A(new_n30032_), .B(new_n30029_), .Y(new_n30054_));
  OAI21X1  g27618(.A0(new_n30054_), .A1(new_n29502_), .B0(pi0239), .Y(new_n30055_));
  AOI21X1  g27619(.A0(new_n30053_), .A1(new_n29502_), .B0(new_n30055_), .Y(new_n30056_));
  OAI21X1  g27620(.A0(new_n30056_), .A1(new_n30000_), .B0(new_n29551_), .Y(new_n30057_));
  OAI21X1  g27621(.A0(new_n30054_), .A1(pi0494), .B0(new_n3253_), .Y(new_n30058_));
  AOI21X1  g27622(.A0(new_n30053_), .A1(pi0494), .B0(new_n30058_), .Y(new_n30059_));
  OAI21X1  g27623(.A0(new_n30059_), .A1(new_n30001_), .B0(pi0524), .Y(new_n30060_));
  NAND3X1  g27624(.A(new_n30060_), .B(new_n30057_), .C(new_n30004_), .Y(new_n30061_));
  NOR3X1   g27625(.A(new_n30033_), .B(new_n30032_), .C(new_n30029_), .Y(new_n30062_));
  AOI21X1  g27626(.A0(new_n30062_), .A1(pi0483), .B0(pi0242), .Y(new_n30063_));
  AOI21X1  g27627(.A0(new_n30063_), .A1(new_n30061_), .B0(new_n30003_), .Y(new_n30064_));
  NAND3X1  g27628(.A(new_n30060_), .B(new_n30057_), .C(pi0483), .Y(new_n30065_));
  AOI21X1  g27629(.A0(new_n30062_), .A1(new_n30004_), .B0(new_n4894_), .Y(new_n30066_));
  AOI21X1  g27630(.A0(new_n30066_), .A1(new_n30065_), .B0(new_n30005_), .Y(new_n30067_));
  MX2X1    g27631(.A(new_n30064_), .B(new_n30067_), .S0(pi0573), .Y(new_n30068_));
  INVX1    g27632(.A(new_n30035_), .Y(new_n30069_));
  OAI21X1  g27633(.A0(new_n30069_), .A1(new_n30008_), .B0(new_n3392_), .Y(new_n30070_));
  AOI21X1  g27634(.A0(new_n30068_), .A1(new_n30008_), .B0(new_n30070_), .Y(new_n30071_));
  OR2X1    g27635(.A(new_n30071_), .B(new_n30007_), .Y(new_n30072_));
  OAI21X1  g27636(.A0(new_n30069_), .A1(pi0495), .B0(pi0235), .Y(new_n30073_));
  AOI21X1  g27637(.A0(new_n30068_), .A1(pi0495), .B0(new_n30073_), .Y(new_n30074_));
  OR2X1    g27638(.A(new_n30074_), .B(new_n30009_), .Y(new_n30075_));
  MX2X1    g27639(.A(new_n30072_), .B(new_n30075_), .S0(pi0575), .Y(new_n30076_));
  OR2X1    g27640(.A(new_n30076_), .B(pi0572), .Y(new_n30077_));
  NOR2X1   g27641(.A(new_n30009_), .B(new_n30007_), .Y(new_n30078_));
  AOI21X1  g27642(.A0(new_n30078_), .A1(pi0572), .B0(pi0244), .Y(new_n30079_));
  AOI21X1  g27643(.A0(new_n30079_), .A1(new_n30077_), .B0(new_n30038_), .Y(new_n30080_));
  INVX1    g27644(.A(pi0572), .Y(new_n30081_));
  AOI21X1  g27645(.A0(new_n30037_), .A1(new_n30081_), .B0(pi0244), .Y(new_n30082_));
  OR2X1    g27646(.A(new_n30076_), .B(new_n30081_), .Y(new_n30083_));
  AOI21X1  g27647(.A0(new_n30078_), .A1(new_n30081_), .B0(new_n4697_), .Y(new_n30084_));
  AOI21X1  g27648(.A0(new_n30084_), .A1(new_n30083_), .B0(new_n30082_), .Y(new_n30085_));
  MX2X1    g27649(.A(new_n30080_), .B(new_n30085_), .S0(pi0493), .Y(new_n30086_));
  OR2X1    g27650(.A(new_n30082_), .B(new_n30038_), .Y(new_n30087_));
  OAI21X1  g27651(.A0(new_n30087_), .A1(new_n30013_), .B0(new_n4550_), .Y(new_n30088_));
  AOI21X1  g27652(.A0(new_n30086_), .A1(new_n30013_), .B0(new_n30088_), .Y(new_n30089_));
  OR2X1    g27653(.A(new_n30089_), .B(new_n30012_), .Y(new_n30090_));
  OAI21X1  g27654(.A0(new_n30087_), .A1(pi0545), .B0(pi0245), .Y(new_n30091_));
  AOI21X1  g27655(.A0(new_n30086_), .A1(pi0545), .B0(new_n30091_), .Y(new_n30092_));
  OR2X1    g27656(.A(new_n30092_), .B(new_n30014_), .Y(new_n30093_));
  MX2X1    g27657(.A(new_n30090_), .B(new_n30093_), .S0(pi0525), .Y(new_n30094_));
  XOR2X1   g27658(.A(pi0525), .B(pi0245), .Y(new_n30095_));
  NOR3X1   g27659(.A(new_n30095_), .B(new_n30082_), .C(new_n30038_), .Y(new_n30096_));
  AOI21X1  g27660(.A0(new_n30096_), .A1(pi0547), .B0(pi0247), .Y(new_n30097_));
  OAI21X1  g27661(.A0(new_n30094_), .A1(pi0547), .B0(new_n30097_), .Y(new_n30098_));
  AOI21X1  g27662(.A0(new_n30098_), .A1(new_n30017_), .B0(pi0527), .Y(new_n30099_));
  NOR3X1   g27663(.A(new_n30014_), .B(new_n30012_), .C(pi0547), .Y(new_n30100_));
  INVX1    g27664(.A(pi0547), .Y(new_n30101_));
  AOI21X1  g27665(.A0(new_n30096_), .A1(new_n30101_), .B0(new_n4117_), .Y(new_n30102_));
  OAI21X1  g27666(.A0(new_n30094_), .A1(new_n30101_), .B0(new_n30102_), .Y(new_n30103_));
  OAI21X1  g27667(.A0(new_n30100_), .A1(pi0247), .B0(new_n30103_), .Y(new_n30104_));
  AOI21X1  g27668(.A0(new_n30104_), .A1(pi0527), .B0(new_n30099_), .Y(new_n30105_));
  AOI21X1  g27669(.A0(new_n30105_), .A1(new_n3578_), .B0(pi0529), .Y(new_n30106_));
  NOR3X1   g27670(.A(new_n30014_), .B(new_n30012_), .C(new_n30101_), .Y(new_n30107_));
  MX2X1    g27671(.A(new_n30100_), .B(new_n30107_), .S0(pi0247), .Y(new_n30108_));
  XOR2X1   g27672(.A(pi0527), .B(pi0247), .Y(new_n30109_));
  OR4X1    g27673(.A(new_n30109_), .B(new_n30095_), .C(new_n30082_), .D(new_n30038_), .Y(new_n30110_));
  OAI21X1  g27674(.A0(new_n30110_), .A1(new_n3578_), .B0(pi0529), .Y(new_n30111_));
  AOI21X1  g27675(.A0(new_n30108_), .A1(new_n3578_), .B0(new_n30111_), .Y(new_n30112_));
  NOR3X1   g27676(.A(new_n30112_), .B(new_n30106_), .C(pi0491), .Y(new_n30113_));
  INVX1    g27677(.A(pi0491), .Y(new_n30114_));
  INVX1    g27678(.A(pi0529), .Y(new_n30115_));
  AOI21X1  g27679(.A0(new_n30105_), .A1(pi0238), .B0(new_n30115_), .Y(new_n30116_));
  OAI21X1  g27680(.A0(new_n30110_), .A1(pi0238), .B0(new_n30115_), .Y(new_n30117_));
  AOI21X1  g27681(.A0(new_n30108_), .A1(pi0238), .B0(new_n30117_), .Y(new_n30118_));
  NOR3X1   g27682(.A(new_n30118_), .B(new_n30116_), .C(new_n30114_), .Y(new_n30119_));
  OAI21X1  g27683(.A0(new_n30119_), .A1(new_n30113_), .B0(pi0233), .Y(new_n30120_));
  INVX1    g27684(.A(pi0489), .Y(new_n30121_));
  INVX1    g27685(.A(pi0485), .Y(new_n30122_));
  AOI21X1  g27686(.A0(new_n29516_), .A1(pi0234), .B0(new_n30122_), .Y(new_n30123_));
  AOI21X1  g27687(.A0(new_n29516_), .A1(new_n2990_), .B0(pi0485), .Y(new_n30124_));
  XOR2X1   g27688(.A(pi0555), .B(new_n29717_), .Y(new_n30125_));
  XOR2X1   g27689(.A(pi0553), .B(new_n29729_), .Y(new_n30126_));
  XOR2X1   g27690(.A(pi0551), .B(pi0240), .Y(new_n30127_));
  XOR2X1   g27691(.A(pi0554), .B(pi0248), .Y(new_n30128_));
  XOR2X1   g27692(.A(pi0563), .B(pi0246), .Y(new_n30129_));
  NOR3X1   g27693(.A(new_n30129_), .B(new_n30128_), .C(new_n30127_), .Y(new_n30130_));
  NAND3X1  g27694(.A(new_n30130_), .B(new_n30126_), .C(new_n30125_), .Y(new_n30131_));
  NOR4X1   g27695(.A(new_n30131_), .B(new_n30124_), .C(new_n30123_), .D(new_n29582_), .Y(new_n30132_));
  INVX1    g27696(.A(new_n30132_), .Y(new_n30133_));
  OR4X1    g27697(.A(new_n30131_), .B(new_n30124_), .C(new_n30123_), .D(pi0550), .Y(new_n30134_));
  AND2X1   g27698(.A(new_n30134_), .B(pi0239), .Y(new_n30135_));
  AOI21X1  g27699(.A0(new_n30133_), .A1(new_n3253_), .B0(new_n30135_), .Y(new_n30136_));
  AOI21X1  g27700(.A0(new_n30136_), .A1(new_n30121_), .B0(pi0242), .Y(new_n30137_));
  AOI21X1  g27701(.A0(new_n30136_), .A1(pi0489), .B0(new_n4894_), .Y(new_n30138_));
  NOR2X1   g27702(.A(new_n30138_), .B(new_n30137_), .Y(new_n30139_));
  AOI21X1  g27703(.A0(new_n30139_), .A1(pi0549), .B0(new_n3392_), .Y(new_n30140_));
  INVX1    g27704(.A(pi0549), .Y(new_n30141_));
  AOI21X1  g27705(.A0(new_n30139_), .A1(new_n30141_), .B0(pi0235), .Y(new_n30142_));
  NOR2X1   g27706(.A(new_n30142_), .B(new_n30140_), .Y(new_n30143_));
  AOI21X1  g27707(.A0(new_n30143_), .A1(pi0486), .B0(new_n4697_), .Y(new_n30144_));
  INVX1    g27708(.A(pi0486), .Y(new_n30145_));
  AOI21X1  g27709(.A0(new_n30143_), .A1(new_n30145_), .B0(pi0244), .Y(new_n30146_));
  XOR2X1   g27710(.A(pi0580), .B(pi0245), .Y(new_n30147_));
  NOR3X1   g27711(.A(new_n30147_), .B(new_n30146_), .C(new_n30144_), .Y(new_n30148_));
  AOI21X1  g27712(.A0(new_n30148_), .A1(pi0552), .B0(new_n4117_), .Y(new_n30149_));
  INVX1    g27713(.A(pi0552), .Y(new_n30150_));
  NOR2X1   g27714(.A(pi0556), .B(pi0242), .Y(new_n30151_));
  AND2X1   g27715(.A(pi0556), .B(pi0242), .Y(new_n30152_));
  NOR2X1   g27716(.A(new_n29756_), .B(new_n29668_), .Y(new_n30153_));
  NOR2X1   g27717(.A(new_n29528_), .B(pi0570), .Y(new_n30154_));
  XOR2X1   g27718(.A(pi0562), .B(pi0241), .Y(new_n30155_));
  AOI22X1  g27719(.A0(pi0564), .A1(new_n29757_), .B0(pi0482), .B1(new_n29717_), .Y(new_n30156_));
  OAI21X1  g27720(.A0(pi0482), .A1(new_n29717_), .B0(new_n30156_), .Y(new_n30157_));
  OR4X1    g27721(.A(new_n30157_), .B(new_n30155_), .C(new_n30154_), .D(new_n30153_), .Y(new_n30158_));
  XOR2X1   g27722(.A(pi0565), .B(new_n29726_), .Y(new_n30159_));
  INVX1    g27723(.A(new_n30159_), .Y(new_n30160_));
  XOR2X1   g27724(.A(pi0560), .B(pi0240), .Y(new_n30161_));
  NOR2X1   g27725(.A(pi0564), .B(new_n29757_), .Y(new_n30162_));
  NOR4X1   g27726(.A(new_n30162_), .B(new_n30161_), .C(new_n30160_), .D(new_n30158_), .Y(new_n30163_));
  OAI21X1  g27727(.A0(pi0564), .A1(new_n29757_), .B0(pi0560), .Y(new_n30164_));
  NOR3X1   g27728(.A(new_n30164_), .B(new_n30160_), .C(new_n30158_), .Y(new_n30165_));
  MX2X1    g27729(.A(new_n30165_), .B(new_n30163_), .S0(new_n29753_), .Y(new_n30166_));
  XOR2X1   g27730(.A(pi0569), .B(pi0239), .Y(new_n30167_));
  AND2X1   g27731(.A(new_n30167_), .B(new_n30166_), .Y(new_n30168_));
  OAI21X1  g27732(.A0(new_n30152_), .A1(new_n30151_), .B0(new_n30168_), .Y(new_n30169_));
  XOR2X1   g27733(.A(pi0531), .B(pi0235), .Y(new_n30170_));
  NOR2X1   g27734(.A(new_n30170_), .B(new_n30169_), .Y(new_n30171_));
  XOR2X1   g27735(.A(pi0566), .B(new_n4697_), .Y(new_n30172_));
  AND2X1   g27736(.A(new_n30172_), .B(new_n30171_), .Y(new_n30173_));
  AOI21X1  g27737(.A0(new_n30173_), .A1(pi0568), .B0(new_n4550_), .Y(new_n30174_));
  INVX1    g27738(.A(new_n30174_), .Y(new_n30175_));
  AOI21X1  g27739(.A0(new_n30134_), .A1(pi0239), .B0(new_n29666_), .Y(new_n30176_));
  INVX1    g27740(.A(new_n30136_), .Y(new_n30177_));
  NAND3X1  g27741(.A(new_n30163_), .B(new_n29666_), .C(pi0239), .Y(new_n30178_));
  NAND2X1  g27742(.A(new_n30178_), .B(new_n30177_), .Y(new_n30179_));
  AOI21X1  g27743(.A0(new_n30176_), .A1(new_n30166_), .B0(new_n30179_), .Y(new_n30180_));
  AND2X1   g27744(.A(new_n30180_), .B(new_n30121_), .Y(new_n30181_));
  AOI21X1  g27745(.A0(new_n30167_), .A1(new_n30166_), .B0(new_n30121_), .Y(new_n30182_));
  OR2X1    g27746(.A(new_n30182_), .B(pi0556), .Y(new_n30183_));
  OAI22X1  g27747(.A0(new_n30183_), .A1(new_n30181_), .B0(new_n30151_), .B1(new_n30137_), .Y(new_n30184_));
  AND2X1   g27748(.A(new_n30180_), .B(pi0489), .Y(new_n30185_));
  OAI21X1  g27749(.A0(new_n30168_), .A1(pi0489), .B0(pi0556), .Y(new_n30186_));
  OAI22X1  g27750(.A0(new_n30186_), .A1(new_n30185_), .B0(new_n30152_), .B1(new_n30138_), .Y(new_n30187_));
  NAND3X1  g27751(.A(new_n30187_), .B(new_n30184_), .C(new_n30141_), .Y(new_n30188_));
  INVX1    g27752(.A(new_n30169_), .Y(new_n30189_));
  AOI21X1  g27753(.A0(new_n30189_), .A1(pi0549), .B0(pi0235), .Y(new_n30190_));
  AOI21X1  g27754(.A0(new_n30190_), .A1(new_n30188_), .B0(new_n30140_), .Y(new_n30191_));
  NAND3X1  g27755(.A(new_n30187_), .B(new_n30184_), .C(pi0549), .Y(new_n30192_));
  AOI21X1  g27756(.A0(new_n30189_), .A1(new_n30141_), .B0(new_n3392_), .Y(new_n30193_));
  AOI21X1  g27757(.A0(new_n30193_), .A1(new_n30192_), .B0(new_n30142_), .Y(new_n30194_));
  MX2X1    g27758(.A(new_n30191_), .B(new_n30194_), .S0(pi0531), .Y(new_n30195_));
  INVX1    g27759(.A(new_n30171_), .Y(new_n30196_));
  OAI21X1  g27760(.A0(new_n30196_), .A1(new_n30145_), .B0(new_n4697_), .Y(new_n30197_));
  AOI21X1  g27761(.A0(new_n30195_), .A1(new_n30145_), .B0(new_n30197_), .Y(new_n30198_));
  OR2X1    g27762(.A(new_n30198_), .B(new_n30144_), .Y(new_n30199_));
  OAI21X1  g27763(.A0(new_n30196_), .A1(pi0486), .B0(pi0244), .Y(new_n30200_));
  AOI21X1  g27764(.A0(new_n30195_), .A1(pi0486), .B0(new_n30200_), .Y(new_n30201_));
  OR2X1    g27765(.A(new_n30201_), .B(new_n30146_), .Y(new_n30202_));
  MX2X1    g27766(.A(new_n30199_), .B(new_n30202_), .S0(pi0566), .Y(new_n30203_));
  NOR2X1   g27767(.A(new_n30146_), .B(new_n30144_), .Y(new_n30204_));
  AOI21X1  g27768(.A0(new_n30204_), .A1(pi0568), .B0(pi0245), .Y(new_n30205_));
  OAI21X1  g27769(.A0(new_n30203_), .A1(pi0568), .B0(new_n30205_), .Y(new_n30206_));
  AOI21X1  g27770(.A0(new_n30206_), .A1(new_n30175_), .B0(pi0580), .Y(new_n30207_));
  INVX1    g27771(.A(pi0568), .Y(new_n30208_));
  NAND3X1  g27772(.A(new_n30172_), .B(new_n30171_), .C(new_n30208_), .Y(new_n30209_));
  AND2X1   g27773(.A(new_n30209_), .B(new_n4550_), .Y(new_n30210_));
  INVX1    g27774(.A(new_n30210_), .Y(new_n30211_));
  AOI21X1  g27775(.A0(new_n30204_), .A1(new_n30208_), .B0(new_n4550_), .Y(new_n30212_));
  OAI21X1  g27776(.A0(new_n30203_), .A1(new_n30208_), .B0(new_n30212_), .Y(new_n30213_));
  NAND2X1  g27777(.A(new_n30213_), .B(new_n30211_), .Y(new_n30214_));
  AOI21X1  g27778(.A0(new_n30214_), .A1(pi0580), .B0(new_n30207_), .Y(new_n30215_));
  NOR2X1   g27779(.A(new_n30210_), .B(new_n30174_), .Y(new_n30216_));
  INVX1    g27780(.A(new_n30216_), .Y(new_n30217_));
  OAI21X1  g27781(.A0(new_n30217_), .A1(new_n30150_), .B0(new_n4117_), .Y(new_n30218_));
  AOI21X1  g27782(.A0(new_n30215_), .A1(new_n30150_), .B0(new_n30218_), .Y(new_n30219_));
  NOR2X1   g27783(.A(new_n30219_), .B(new_n30149_), .Y(new_n30220_));
  AOI21X1  g27784(.A0(new_n30148_), .A1(new_n30150_), .B0(pi0247), .Y(new_n30221_));
  OAI21X1  g27785(.A0(new_n30217_), .A1(pi0552), .B0(pi0247), .Y(new_n30222_));
  AOI21X1  g27786(.A0(new_n30215_), .A1(pi0552), .B0(new_n30222_), .Y(new_n30223_));
  NOR2X1   g27787(.A(new_n30223_), .B(new_n30221_), .Y(new_n30224_));
  MX2X1    g27788(.A(new_n30220_), .B(new_n30224_), .S0(pi0532), .Y(new_n30225_));
  AOI21X1  g27789(.A0(new_n30225_), .A1(new_n3578_), .B0(pi0577), .Y(new_n30226_));
  INVX1    g27790(.A(pi0498), .Y(new_n30227_));
  NOR3X1   g27791(.A(new_n30221_), .B(new_n30149_), .C(new_n3578_), .Y(new_n30228_));
  XOR2X1   g27792(.A(pi0532), .B(new_n4117_), .Y(new_n30229_));
  NAND2X1  g27793(.A(new_n30229_), .B(new_n30216_), .Y(new_n30230_));
  OAI21X1  g27794(.A0(new_n30230_), .A1(pi0238), .B0(pi0577), .Y(new_n30231_));
  OAI21X1  g27795(.A0(new_n30231_), .A1(new_n30228_), .B0(new_n30227_), .Y(new_n30232_));
  INVX1    g27796(.A(pi0577), .Y(new_n30233_));
  AOI21X1  g27797(.A0(new_n30225_), .A1(pi0238), .B0(new_n30233_), .Y(new_n30234_));
  NOR3X1   g27798(.A(new_n30221_), .B(new_n30149_), .C(pi0238), .Y(new_n30235_));
  OAI21X1  g27799(.A0(new_n30230_), .A1(new_n3578_), .B0(new_n30233_), .Y(new_n30236_));
  OAI21X1  g27800(.A0(new_n30236_), .A1(new_n30235_), .B0(pi0498), .Y(new_n30237_));
  OAI22X1  g27801(.A0(new_n30237_), .A1(new_n30234_), .B0(new_n30232_), .B1(new_n30226_), .Y(new_n30238_));
  AOI21X1  g27802(.A0(new_n30238_), .A1(new_n22718_), .B0(pi0237), .Y(new_n30239_));
  AOI22X1  g27803(.A0(new_n30239_), .A1(new_n30120_), .B0(new_n29990_), .B1(new_n29867_), .Y(po0750));
  NOR4X1   g27804(.A(new_n29358_), .B(pi0806), .C(new_n29357_), .D(new_n29356_), .Y(new_n30241_));
  OR4X1    g27805(.A(new_n29358_), .B(pi0806), .C(new_n29357_), .D(pi0332), .Y(new_n30242_));
  OR2X1    g27806(.A(new_n29356_), .B(pi0332), .Y(new_n30243_));
  AOI21X1  g27807(.A0(new_n30243_), .A1(new_n30242_), .B0(new_n30241_), .Y(po0751));
  NAND3X1  g27808(.A(pi0600), .B(pi0597), .C(pi0594), .Y(new_n30245_));
  INVX1    g27809(.A(new_n30245_), .Y(new_n30246_));
  INVX1    g27810(.A(pi0806), .Y(new_n30247_));
  AND2X1   g27811(.A(new_n30247_), .B(pi0605), .Y(new_n30248_));
  NAND3X1  g27812(.A(new_n30248_), .B(new_n30246_), .C(pi0601), .Y(new_n30249_));
  OAI21X1  g27813(.A0(new_n30249_), .A1(new_n29341_), .B0(new_n2445_), .Y(new_n30250_));
  AOI21X1  g27814(.A0(new_n30249_), .A1(new_n29341_), .B0(new_n30250_), .Y(po0752));
  AND2X1   g27815(.A(pi0596), .B(new_n2445_), .Y(new_n30252_));
  NAND4X1  g27816(.A(pi0600), .B(pi0597), .C(pi0595), .D(pi0594), .Y(new_n30253_));
  NOR4X1   g27817(.A(new_n30253_), .B(new_n29358_), .C(pi0806), .D(pi0332), .Y(new_n30254_));
  MX2X1    g27818(.A(new_n30252_), .B(new_n29345_), .S0(new_n30254_), .Y(po0753));
  OR2X1    g27819(.A(new_n30241_), .B(pi0597), .Y(new_n30256_));
  AOI21X1  g27820(.A0(new_n30241_), .A1(pi0597), .B0(pi0332), .Y(new_n30257_));
  AND2X1   g27821(.A(new_n30257_), .B(new_n30256_), .Y(po0754));
  INVX1    g27822(.A(pi0598), .Y(new_n30259_));
  NOR4X1   g27823(.A(new_n5118_), .B(new_n14590_), .C(pi0882), .D(pi0057), .Y(new_n30260_));
  NAND3X1  g27824(.A(new_n5028_), .B(pi0780), .C(pi0740), .Y(new_n30261_));
  OAI21X1  g27825(.A0(new_n30260_), .A1(new_n30259_), .B0(new_n30261_), .Y(po0755));
  NAND2X1  g27826(.A(new_n30254_), .B(pi0596), .Y(new_n30263_));
  AND2X1   g27827(.A(pi0599), .B(new_n2445_), .Y(new_n30264_));
  MX2X1    g27828(.A(new_n29346_), .B(new_n30264_), .S0(new_n30263_), .Y(po0756));
  NOR3X1   g27829(.A(new_n29358_), .B(pi0806), .C(pi0332), .Y(new_n30266_));
  AND2X1   g27830(.A(pi0600), .B(new_n2445_), .Y(new_n30267_));
  MX2X1    g27831(.A(new_n30267_), .B(new_n29357_), .S0(new_n30266_), .Y(po0757));
  NOR2X1   g27832(.A(pi0989), .B(pi0806), .Y(new_n30269_));
  OAI21X1  g27833(.A0(new_n30247_), .A1(pi0601), .B0(new_n2445_), .Y(new_n30270_));
  NOR2X1   g27834(.A(new_n30270_), .B(new_n30269_), .Y(po0758));
  NOR3X1   g27835(.A(new_n12869_), .B(new_n12499_), .C(new_n24954_), .Y(new_n30272_));
  AOI21X1  g27836(.A0(pi1160), .A1(pi0715), .B0(new_n12897_), .Y(new_n30273_));
  OAI21X1  g27837(.A0(pi1160), .A1(pi0715), .B0(new_n30273_), .Y(new_n30274_));
  NAND4X1  g27838(.A(new_n30274_), .B(new_n30272_), .C(new_n14286_), .D(new_n13570_), .Y(new_n30275_));
  OAI22X1  g27839(.A0(new_n30275_), .A1(new_n13624_), .B0(new_n5293_), .B1(pi0230), .Y(po0759));
  INVX1    g27840(.A(pi1061), .Y(new_n30277_));
  INVX1    g27841(.A(pi0980), .Y(new_n30278_));
  AND2X1   g27842(.A(pi1038), .B(new_n30278_), .Y(new_n30279_));
  NAND4X1  g27843(.A(new_n30279_), .B(new_n30277_), .C(pi1060), .D(pi0952), .Y(new_n30280_));
  NOR2X1   g27844(.A(new_n30280_), .B(new_n12898_), .Y(po0897));
  NOR2X1   g27845(.A(po0897), .B(pi0603), .Y(new_n30282_));
  INVX1    g27846(.A(pi0966), .Y(new_n30283_));
  OR2X1    g27847(.A(pi1100), .B(new_n12898_), .Y(new_n30284_));
  OAI21X1  g27848(.A0(new_n30284_), .A1(new_n30280_), .B0(new_n30283_), .Y(new_n30285_));
  OAI21X1  g27849(.A0(pi0872), .A1(pi0871), .B0(pi0966), .Y(new_n30286_));
  OAI21X1  g27850(.A0(new_n30285_), .A1(new_n30282_), .B0(new_n30286_), .Y(po0760));
  NAND2X1  g27851(.A(new_n11993_), .B(pi0823), .Y(new_n30288_));
  NAND3X1  g27852(.A(pi0983), .B(pi0907), .C(new_n2953_), .Y(new_n30289_));
  NAND3X1  g27853(.A(new_n30289_), .B(new_n30288_), .C(pi0604), .Y(new_n30290_));
  OAI21X1  g27854(.A0(new_n30288_), .A1(pi0779), .B0(new_n30290_), .Y(po0761));
  AOI21X1  g27855(.A0(new_n30247_), .A1(new_n2445_), .B0(pi0605), .Y(new_n30292_));
  NOR3X1   g27856(.A(new_n30292_), .B(new_n30248_), .C(pi0332), .Y(po0762));
  MX2X1    g27857(.A(pi0606), .B(pi1104), .S0(po0897), .Y(new_n30294_));
  MX2X1    g27858(.A(new_n30294_), .B(pi0837), .S0(pi0966), .Y(po0763));
  INVX1    g27859(.A(po0897), .Y(new_n30296_));
  OAI21X1  g27860(.A0(new_n30296_), .A1(pi1107), .B0(new_n30283_), .Y(new_n30297_));
  AOI21X1  g27861(.A0(new_n30296_), .A1(new_n23127_), .B0(new_n30297_), .Y(po0764));
  OAI21X1  g27862(.A0(new_n30296_), .A1(pi1116), .B0(new_n30283_), .Y(new_n30299_));
  AOI21X1  g27863(.A0(new_n30296_), .A1(new_n12584_), .B0(new_n30299_), .Y(po0765));
  OAI21X1  g27864(.A0(new_n30296_), .A1(pi1118), .B0(new_n30283_), .Y(new_n30301_));
  AOI21X1  g27865(.A0(new_n30296_), .A1(new_n12590_), .B0(new_n30301_), .Y(po0766));
  NOR2X1   g27866(.A(po0897), .B(pi0610), .Y(new_n30303_));
  NOR3X1   g27867(.A(new_n30280_), .B(pi1113), .C(new_n12898_), .Y(new_n30304_));
  NOR3X1   g27868(.A(new_n30304_), .B(new_n30303_), .C(pi0966), .Y(po0767));
  NOR2X1   g27869(.A(po0897), .B(pi0611), .Y(new_n30306_));
  NOR3X1   g27870(.A(new_n30280_), .B(pi1114), .C(new_n12898_), .Y(new_n30307_));
  NOR3X1   g27871(.A(new_n30307_), .B(new_n30306_), .C(pi0966), .Y(po0768));
  OAI21X1  g27872(.A0(new_n30296_), .A1(pi1111), .B0(new_n30283_), .Y(new_n30309_));
  AOI21X1  g27873(.A0(new_n30296_), .A1(new_n23526_), .B0(new_n30309_), .Y(po0769));
  NOR2X1   g27874(.A(po0897), .B(pi0613), .Y(new_n30311_));
  NOR3X1   g27875(.A(new_n30280_), .B(pi1115), .C(new_n12898_), .Y(new_n30312_));
  NOR3X1   g27876(.A(new_n30312_), .B(new_n30311_), .C(pi0966), .Y(po0770));
  INVX1    g27877(.A(pi0871), .Y(new_n30314_));
  NOR2X1   g27878(.A(po0897), .B(pi0614), .Y(new_n30315_));
  OAI21X1  g27879(.A0(new_n30296_), .A1(pi1102), .B0(new_n30283_), .Y(new_n30316_));
  OAI22X1  g27880(.A0(new_n30316_), .A1(new_n30315_), .B0(new_n30283_), .B1(new_n30314_), .Y(po0771));
  NOR4X1   g27881(.A(new_n5118_), .B(new_n5297_), .C(pi0882), .D(pi0057), .Y(new_n30318_));
  NAND3X1  g27882(.A(new_n5030_), .B(pi0797), .C(pi0779), .Y(new_n30319_));
  OAI21X1  g27883(.A0(new_n30318_), .A1(pi0615), .B0(new_n30319_), .Y(po0772));
  INVX1    g27884(.A(pi0872), .Y(new_n30321_));
  NOR2X1   g27885(.A(po0897), .B(pi0616), .Y(new_n30322_));
  OAI21X1  g27886(.A0(new_n30296_), .A1(pi1101), .B0(new_n30283_), .Y(new_n30323_));
  OAI22X1  g27887(.A0(new_n30323_), .A1(new_n30322_), .B0(new_n30283_), .B1(new_n30321_), .Y(po0773));
  MX2X1    g27888(.A(pi0617), .B(pi1105), .S0(po0897), .Y(new_n30325_));
  MX2X1    g27889(.A(new_n30325_), .B(pi0850), .S0(pi0966), .Y(po0774));
  OAI21X1  g27890(.A0(new_n30296_), .A1(pi1117), .B0(new_n30283_), .Y(new_n30327_));
  AOI21X1  g27891(.A0(new_n30296_), .A1(new_n12614_), .B0(new_n30327_), .Y(po0775));
  OAI21X1  g27892(.A0(new_n30296_), .A1(pi1122), .B0(new_n30283_), .Y(new_n30329_));
  AOI21X1  g27893(.A0(new_n30296_), .A1(new_n12637_), .B0(new_n30329_), .Y(po0776));
  NOR2X1   g27894(.A(po0897), .B(pi0620), .Y(new_n30331_));
  NOR3X1   g27895(.A(new_n30280_), .B(pi1112), .C(new_n12898_), .Y(new_n30332_));
  NOR3X1   g27896(.A(new_n30332_), .B(new_n30331_), .C(pi0966), .Y(po0777));
  OAI21X1  g27897(.A0(new_n30296_), .A1(pi1108), .B0(new_n30283_), .Y(new_n30334_));
  AOI21X1  g27898(.A0(new_n30296_), .A1(new_n12092_), .B0(new_n30334_), .Y(po0778));
  OAI21X1  g27899(.A0(new_n30296_), .A1(pi1109), .B0(new_n30283_), .Y(new_n30336_));
  AOI21X1  g27900(.A0(new_n30296_), .A1(new_n23196_), .B0(new_n30336_), .Y(po0779));
  OAI21X1  g27901(.A0(new_n30296_), .A1(pi1106), .B0(new_n30283_), .Y(new_n30338_));
  AOI21X1  g27902(.A0(new_n30296_), .A1(new_n22925_), .B0(new_n30338_), .Y(po0780));
  NAND2X1  g27903(.A(new_n12125_), .B(pi0831), .Y(new_n30340_));
  NAND3X1  g27904(.A(pi0983), .B(pi0947), .C(new_n2953_), .Y(new_n30341_));
  NAND3X1  g27905(.A(new_n30341_), .B(new_n30340_), .C(pi0624), .Y(new_n30342_));
  OAI21X1  g27906(.A0(new_n30340_), .A1(pi0780), .B0(new_n30342_), .Y(po0781));
  INVX1    g27907(.A(pi1054), .Y(new_n30344_));
  NAND3X1  g27908(.A(pi1088), .B(pi1066), .C(new_n30344_), .Y(new_n30345_));
  NOR4X1   g27909(.A(new_n30345_), .B(pi0973), .C(pi0953), .D(new_n12898_), .Y(po0954));
  INVX1    g27910(.A(po0954), .Y(new_n30347_));
  INVX1    g27911(.A(pi0962), .Y(new_n30348_));
  OAI21X1  g27912(.A0(new_n30347_), .A1(pi1116), .B0(new_n30348_), .Y(new_n30349_));
  AOI21X1  g27913(.A0(new_n30347_), .A1(new_n12493_), .B0(new_n30349_), .Y(po0782));
  OAI21X1  g27914(.A0(new_n30296_), .A1(pi1121), .B0(new_n30283_), .Y(new_n30351_));
  AOI21X1  g27915(.A0(new_n30296_), .A1(new_n12664_), .B0(new_n30351_), .Y(po0783));
  OAI21X1  g27916(.A0(new_n30347_), .A1(pi1117), .B0(new_n30348_), .Y(new_n30353_));
  AOI21X1  g27917(.A0(new_n30347_), .A1(new_n12622_), .B0(new_n30353_), .Y(po0784));
  OAI21X1  g27918(.A0(new_n30347_), .A1(pi1119), .B0(new_n30348_), .Y(new_n30355_));
  AOI21X1  g27919(.A0(new_n30347_), .A1(new_n12683_), .B0(new_n30355_), .Y(po0785));
  OAI21X1  g27920(.A0(new_n30296_), .A1(pi1119), .B0(new_n30283_), .Y(new_n30357_));
  AOI21X1  g27921(.A0(new_n30296_), .A1(new_n12689_), .B0(new_n30357_), .Y(po0786));
  OAI21X1  g27922(.A0(new_n30296_), .A1(pi1120), .B0(new_n30283_), .Y(new_n30359_));
  AOI21X1  g27923(.A0(new_n30296_), .A1(new_n12723_), .B0(new_n30359_), .Y(po0787));
  INVX1    g27924(.A(pi1113), .Y(new_n30361_));
  INVX1    g27925(.A(pi0631), .Y(new_n30362_));
  OAI21X1  g27926(.A0(po0954), .A1(new_n30362_), .B0(new_n30348_), .Y(new_n30363_));
  AOI21X1  g27927(.A0(po0954), .A1(new_n30361_), .B0(new_n30363_), .Y(po0788));
  INVX1    g27928(.A(pi1115), .Y(new_n30365_));
  INVX1    g27929(.A(pi0632), .Y(new_n30366_));
  OAI21X1  g27930(.A0(po0954), .A1(new_n30366_), .B0(new_n30348_), .Y(new_n30367_));
  AOI21X1  g27931(.A0(po0954), .A1(new_n30365_), .B0(new_n30367_), .Y(po0789));
  OAI21X1  g27932(.A0(new_n30296_), .A1(pi1110), .B0(new_n30283_), .Y(new_n30369_));
  AOI21X1  g27933(.A0(new_n30296_), .A1(new_n21917_), .B0(new_n30369_), .Y(po0790));
  OAI21X1  g27934(.A0(new_n30347_), .A1(pi1110), .B0(new_n30348_), .Y(new_n30371_));
  AOI21X1  g27935(.A0(new_n30347_), .A1(new_n22072_), .B0(new_n30371_), .Y(po0791));
  INVX1    g27936(.A(pi1112), .Y(new_n30373_));
  INVX1    g27937(.A(pi0635), .Y(new_n30374_));
  OAI21X1  g27938(.A0(po0954), .A1(new_n30374_), .B0(new_n30348_), .Y(new_n30375_));
  AOI21X1  g27939(.A0(po0954), .A1(new_n30373_), .B0(new_n30375_), .Y(po0792));
  NOR2X1   g27940(.A(po0897), .B(pi0636), .Y(new_n30377_));
  NOR3X1   g27941(.A(new_n30280_), .B(pi1127), .C(new_n12898_), .Y(new_n30378_));
  NOR3X1   g27942(.A(new_n30378_), .B(new_n30377_), .C(pi0966), .Y(po0793));
  OAI21X1  g27943(.A0(new_n30347_), .A1(pi1105), .B0(new_n30348_), .Y(new_n30380_));
  AOI21X1  g27944(.A0(new_n30347_), .A1(new_n22270_), .B0(new_n30380_), .Y(po0794));
  OAI21X1  g27945(.A0(new_n30347_), .A1(pi1107), .B0(new_n30348_), .Y(new_n30382_));
  AOI21X1  g27946(.A0(new_n30347_), .A1(new_n23116_), .B0(new_n30382_), .Y(po0795));
  OAI21X1  g27947(.A0(new_n30347_), .A1(pi1109), .B0(new_n30348_), .Y(new_n30384_));
  AOI21X1  g27948(.A0(new_n30347_), .A1(new_n23151_), .B0(new_n30384_), .Y(po0796));
  NOR2X1   g27949(.A(po0897), .B(pi0640), .Y(new_n30386_));
  NOR3X1   g27950(.A(new_n30280_), .B(pi1128), .C(new_n12898_), .Y(new_n30387_));
  NOR3X1   g27951(.A(new_n30387_), .B(new_n30386_), .C(pi0966), .Y(po0797));
  OAI21X1  g27952(.A0(new_n30347_), .A1(pi1121), .B0(new_n30348_), .Y(new_n30389_));
  AOI21X1  g27953(.A0(new_n30347_), .A1(new_n12672_), .B0(new_n30389_), .Y(po0798));
  OAI21X1  g27954(.A0(new_n30296_), .A1(pi1103), .B0(new_n30283_), .Y(new_n30391_));
  AOI21X1  g27955(.A0(new_n30296_), .A1(new_n11968_), .B0(new_n30391_), .Y(po0799));
  OAI21X1  g27956(.A0(new_n30347_), .A1(pi1104), .B0(new_n30348_), .Y(new_n30393_));
  AOI21X1  g27957(.A0(new_n30347_), .A1(new_n22461_), .B0(new_n30393_), .Y(po0800));
  OAI21X1  g27958(.A0(new_n30296_), .A1(pi1123), .B0(new_n30283_), .Y(new_n30395_));
  AOI21X1  g27959(.A0(new_n30296_), .A1(new_n12743_), .B0(new_n30395_), .Y(po0801));
  NOR2X1   g27960(.A(po0897), .B(pi0645), .Y(new_n30397_));
  NOR3X1   g27961(.A(new_n30280_), .B(pi1125), .C(new_n12898_), .Y(new_n30398_));
  NOR3X1   g27962(.A(new_n30398_), .B(new_n30397_), .C(pi0966), .Y(po0802));
  INVX1    g27963(.A(pi1114), .Y(new_n30400_));
  INVX1    g27964(.A(pi0646), .Y(new_n30401_));
  OAI21X1  g27965(.A0(po0954), .A1(new_n30401_), .B0(new_n30348_), .Y(new_n30402_));
  AOI21X1  g27966(.A0(po0954), .A1(new_n30400_), .B0(new_n30402_), .Y(po0803));
  OAI21X1  g27967(.A0(new_n30347_), .A1(pi1120), .B0(new_n30348_), .Y(new_n30404_));
  AOI21X1  g27968(.A0(new_n30347_), .A1(new_n12705_), .B0(new_n30404_), .Y(po0804));
  OAI21X1  g27969(.A0(new_n30347_), .A1(pi1122), .B0(new_n30348_), .Y(new_n30406_));
  AOI21X1  g27970(.A0(new_n30347_), .A1(new_n12645_), .B0(new_n30406_), .Y(po0805));
  INVX1    g27971(.A(pi1126), .Y(new_n30408_));
  INVX1    g27972(.A(pi0649), .Y(new_n30409_));
  OAI21X1  g27973(.A0(po0954), .A1(new_n30409_), .B0(new_n30348_), .Y(new_n30410_));
  AOI21X1  g27974(.A0(po0954), .A1(new_n30408_), .B0(new_n30410_), .Y(po0806));
  INVX1    g27975(.A(pi1127), .Y(new_n30412_));
  INVX1    g27976(.A(pi0650), .Y(new_n30413_));
  OAI21X1  g27977(.A0(po0954), .A1(new_n30413_), .B0(new_n30348_), .Y(new_n30414_));
  AOI21X1  g27978(.A0(po0954), .A1(new_n30412_), .B0(new_n30414_), .Y(po0807));
  NOR2X1   g27979(.A(po0897), .B(pi0651), .Y(new_n30416_));
  NOR3X1   g27980(.A(new_n30280_), .B(pi1130), .C(new_n12898_), .Y(new_n30417_));
  NOR3X1   g27981(.A(new_n30417_), .B(new_n30416_), .C(pi0966), .Y(po0808));
  NOR2X1   g27982(.A(po0897), .B(pi0652), .Y(new_n30419_));
  NOR3X1   g27983(.A(new_n30280_), .B(pi1131), .C(new_n12898_), .Y(new_n30420_));
  NOR3X1   g27984(.A(new_n30420_), .B(new_n30419_), .C(pi0966), .Y(po0809));
  NOR2X1   g27985(.A(po0897), .B(pi0653), .Y(new_n30422_));
  NOR3X1   g27986(.A(new_n30280_), .B(pi1129), .C(new_n12898_), .Y(new_n30423_));
  NOR3X1   g27987(.A(new_n30423_), .B(new_n30422_), .C(pi0966), .Y(po0810));
  INVX1    g27988(.A(pi1130), .Y(new_n30425_));
  INVX1    g27989(.A(pi0654), .Y(new_n30426_));
  OAI21X1  g27990(.A0(po0954), .A1(new_n30426_), .B0(new_n30348_), .Y(new_n30427_));
  AOI21X1  g27991(.A0(po0954), .A1(new_n30425_), .B0(new_n30427_), .Y(po0811));
  INVX1    g27992(.A(pi1124), .Y(new_n30429_));
  INVX1    g27993(.A(pi0655), .Y(new_n30430_));
  OAI21X1  g27994(.A0(po0954), .A1(new_n30430_), .B0(new_n30348_), .Y(new_n30431_));
  AOI21X1  g27995(.A0(po0954), .A1(new_n30429_), .B0(new_n30431_), .Y(po0812));
  NOR2X1   g27996(.A(po0897), .B(pi0656), .Y(new_n30433_));
  NOR3X1   g27997(.A(new_n30280_), .B(pi1126), .C(new_n12898_), .Y(new_n30434_));
  NOR3X1   g27998(.A(new_n30434_), .B(new_n30433_), .C(pi0966), .Y(po0813));
  INVX1    g27999(.A(pi1131), .Y(new_n30436_));
  INVX1    g28000(.A(pi0657), .Y(new_n30437_));
  OAI21X1  g28001(.A0(po0954), .A1(new_n30437_), .B0(new_n30348_), .Y(new_n30438_));
  AOI21X1  g28002(.A0(po0954), .A1(new_n30436_), .B0(new_n30438_), .Y(po0814));
  NOR2X1   g28003(.A(po0897), .B(pi0658), .Y(new_n30440_));
  NOR3X1   g28004(.A(new_n30280_), .B(pi1124), .C(new_n12898_), .Y(new_n30441_));
  NOR3X1   g28005(.A(new_n30441_), .B(new_n30440_), .C(pi0966), .Y(po0815));
  INVX1    g28006(.A(pi0265), .Y(new_n30443_));
  INVX1    g28007(.A(pi0264), .Y(new_n30444_));
  INVX1    g28008(.A(pi0280), .Y(new_n30445_));
  AND2X1   g28009(.A(pi0992), .B(pi0266), .Y(new_n30446_));
  AND2X1   g28010(.A(new_n30446_), .B(new_n30445_), .Y(new_n30447_));
  INVX1    g28011(.A(new_n30447_), .Y(new_n30448_));
  OR2X1    g28012(.A(pi0277), .B(pi0270), .Y(new_n30449_));
  OR2X1    g28013(.A(new_n30449_), .B(pi0282), .Y(new_n30450_));
  NOR4X1   g28014(.A(new_n30450_), .B(new_n30448_), .C(pi0281), .D(pi0269), .Y(new_n30451_));
  AND2X1   g28015(.A(new_n30451_), .B(new_n30444_), .Y(new_n30452_));
  AND2X1   g28016(.A(new_n30452_), .B(new_n30443_), .Y(new_n30453_));
  XOR2X1   g28017(.A(new_n30453_), .B(new_n3360_), .Y(po0816));
  OAI21X1  g28018(.A0(new_n30347_), .A1(pi1118), .B0(new_n30348_), .Y(new_n30455_));
  AOI21X1  g28019(.A0(new_n30347_), .A1(new_n12596_), .B0(new_n30455_), .Y(po0817));
  OAI21X1  g28020(.A0(new_n30347_), .A1(pi1101), .B0(new_n30348_), .Y(new_n30457_));
  AOI21X1  g28021(.A0(new_n30347_), .A1(new_n11976_), .B0(new_n30457_), .Y(po0818));
  OAI21X1  g28022(.A0(new_n30347_), .A1(pi1102), .B0(new_n30348_), .Y(new_n30459_));
  AOI21X1  g28023(.A0(new_n30347_), .A1(new_n11977_), .B0(new_n30459_), .Y(po0819));
  NOR2X1   g28024(.A(pi0257), .B(pi0199), .Y(new_n30461_));
  OAI22X1  g28025(.A0(pi1065), .A1(new_n7941_), .B0(pi0224), .B1(pi0223), .Y(new_n30462_));
  NOR2X1   g28026(.A(new_n30462_), .B(new_n30461_), .Y(new_n30463_));
  AND2X1   g28027(.A(pi0592), .B(new_n6074_), .Y(new_n30464_));
  NOR3X1   g28028(.A(pi0592), .B(new_n6074_), .C(new_n6169_), .Y(new_n30465_));
  AOI21X1  g28029(.A0(new_n30464_), .A1(pi0365), .B0(new_n30465_), .Y(new_n30466_));
  NOR3X1   g28030(.A(pi0592), .B(pi0591), .C(new_n6168_), .Y(new_n30467_));
  AOI21X1  g28031(.A0(new_n30467_), .A1(pi0323), .B0(pi0588), .Y(new_n30468_));
  OAI21X1  g28032(.A0(new_n30466_), .A1(pi0590), .B0(new_n30468_), .Y(new_n30469_));
  NOR2X1   g28033(.A(pi0224), .B(pi0223), .Y(new_n30470_));
  INVX1    g28034(.A(new_n30470_), .Y(new_n30471_));
  NOR3X1   g28035(.A(pi0592), .B(pi0591), .C(pi0590), .Y(new_n30472_));
  AOI21X1  g28036(.A0(new_n30472_), .A1(pi0464), .B0(new_n9028_), .Y(new_n30473_));
  NOR2X1   g28037(.A(new_n30473_), .B(new_n30471_), .Y(new_n30474_));
  AOI21X1  g28038(.A0(new_n30474_), .A1(new_n30469_), .B0(new_n30463_), .Y(new_n30475_));
  NOR3X1   g28039(.A(pi1138), .B(pi1137), .C(pi1134), .Y(new_n30476_));
  INVX1    g28040(.A(new_n30476_), .Y(new_n30477_));
  AOI21X1  g28041(.A0(pi1136), .A1(new_n22072_), .B0(new_n28313_), .Y(new_n30478_));
  OAI21X1  g28042(.A0(pi1136), .A1(pi0784), .B0(new_n30478_), .Y(new_n30479_));
  AOI21X1  g28043(.A0(pi1136), .A1(new_n21917_), .B0(pi1135), .Y(new_n30480_));
  OAI21X1  g28044(.A0(pi1136), .A1(pi0815), .B0(new_n30480_), .Y(new_n30481_));
  AOI21X1  g28045(.A0(new_n30481_), .A1(new_n30479_), .B0(new_n30477_), .Y(new_n30482_));
  NOR2X1   g28046(.A(pi1138), .B(pi1137), .Y(new_n30483_));
  AOI21X1  g28047(.A0(new_n30483_), .A1(pi1135), .B0(new_n28946_), .Y(new_n30484_));
  AND2X1   g28048(.A(new_n30484_), .B(new_n14977_), .Y(new_n30485_));
  AND2X1   g28049(.A(new_n30483_), .B(pi1134), .Y(new_n30486_));
  OAI21X1  g28050(.A0(pi1136), .A1(new_n28313_), .B0(new_n30486_), .Y(new_n30487_));
  OAI22X1  g28051(.A0(pi1136), .A1(pi0855), .B0(new_n28313_), .B1(pi0700), .Y(new_n30488_));
  NOR3X1   g28052(.A(new_n30488_), .B(new_n30487_), .C(new_n30485_), .Y(new_n30489_));
  OAI21X1  g28053(.A0(new_n30489_), .A1(new_n30482_), .B0(new_n10265_), .Y(new_n30490_));
  OAI21X1  g28054(.A0(new_n30475_), .A1(new_n10265_), .B0(new_n30490_), .Y(po0820));
  INVX1    g28055(.A(new_n30467_), .Y(new_n30492_));
  AND2X1   g28056(.A(pi0591), .B(new_n6168_), .Y(new_n30493_));
  AOI21X1  g28057(.A0(pi0592), .A1(new_n6168_), .B0(pi0588), .Y(new_n30494_));
  INVX1    g28058(.A(new_n30494_), .Y(new_n30495_));
  AOI21X1  g28059(.A0(new_n30493_), .A1(pi0404), .B0(new_n30495_), .Y(new_n30496_));
  AOI21X1  g28060(.A0(new_n6074_), .A1(pi0380), .B0(new_n6120_), .Y(new_n30497_));
  OAI22X1  g28061(.A0(new_n30497_), .A1(new_n30496_), .B0(new_n30492_), .B1(new_n6039_), .Y(new_n30498_));
  AOI21X1  g28062(.A0(new_n30472_), .A1(pi0429), .B0(new_n9028_), .Y(new_n30499_));
  NOR2X1   g28063(.A(new_n30499_), .B(new_n30471_), .Y(new_n30500_));
  OR2X1    g28064(.A(pi0292), .B(pi0199), .Y(new_n30501_));
  INVX1    g28065(.A(pi1084), .Y(new_n30502_));
  AOI21X1  g28066(.A0(new_n30502_), .A1(pi0199), .B0(new_n30470_), .Y(new_n30503_));
  AOI22X1  g28067(.A0(new_n30503_), .A1(new_n30501_), .B0(new_n30500_), .B1(new_n30498_), .Y(new_n30504_));
  AOI21X1  g28068(.A0(pi1135), .A1(pi0662), .B0(new_n28946_), .Y(new_n30505_));
  OAI21X1  g28069(.A0(pi1135), .A1(new_n12051_), .B0(new_n30505_), .Y(new_n30506_));
  INVX1    g28070(.A(pi0811), .Y(new_n30507_));
  AOI21X1  g28071(.A0(pi1135), .A1(pi0785), .B0(pi1136), .Y(new_n30508_));
  OAI21X1  g28072(.A0(pi1135), .A1(new_n30507_), .B0(new_n30508_), .Y(new_n30509_));
  AOI21X1  g28073(.A0(new_n30509_), .A1(new_n30506_), .B0(pi1134), .Y(new_n30510_));
  OAI21X1  g28074(.A0(new_n28313_), .A1(pi0727), .B0(pi1136), .Y(new_n30511_));
  AOI21X1  g28075(.A0(new_n28313_), .A1(new_n15465_), .B0(new_n30511_), .Y(new_n30512_));
  NOR2X1   g28076(.A(pi1136), .B(pi1135), .Y(new_n30513_));
  INVX1    g28077(.A(new_n30513_), .Y(new_n30514_));
  OAI21X1  g28078(.A0(new_n30514_), .A1(new_n30321_), .B0(pi1134), .Y(new_n30515_));
  NOR3X1   g28079(.A(new_n6748_), .B(pi1138), .C(pi1137), .Y(new_n30516_));
  OAI21X1  g28080(.A0(new_n30515_), .A1(new_n30512_), .B0(new_n30516_), .Y(new_n30517_));
  OAI22X1  g28081(.A0(new_n30517_), .A1(new_n30510_), .B0(new_n30504_), .B1(new_n10265_), .Y(po0821));
  OAI21X1  g28082(.A0(new_n30347_), .A1(pi1108), .B0(new_n30348_), .Y(new_n30519_));
  AOI21X1  g28083(.A0(new_n30347_), .A1(new_n12255_), .B0(new_n30519_), .Y(po0822));
  AOI21X1  g28084(.A0(pi1135), .A1(new_n23116_), .B0(new_n28946_), .Y(new_n30521_));
  OAI21X1  g28085(.A0(pi1135), .A1(pi0607), .B0(new_n30521_), .Y(new_n30522_));
  AOI21X1  g28086(.A0(new_n28313_), .A1(pi0799), .B0(pi1136), .Y(new_n30523_));
  OAI21X1  g28087(.A0(new_n28313_), .A1(pi0790), .B0(new_n30523_), .Y(new_n30524_));
  AOI21X1  g28088(.A0(new_n30524_), .A1(new_n30522_), .B0(new_n30477_), .Y(new_n30525_));
  AND2X1   g28089(.A(new_n30484_), .B(new_n15641_), .Y(new_n30526_));
  OAI22X1  g28090(.A0(pi1136), .A1(pi0873), .B0(new_n28313_), .B1(pi0691), .Y(new_n30527_));
  NOR3X1   g28091(.A(new_n30527_), .B(new_n30526_), .C(new_n30487_), .Y(new_n30528_));
  OAI21X1  g28092(.A0(new_n30528_), .A1(new_n30525_), .B0(new_n10265_), .Y(new_n30529_));
  OR2X1    g28093(.A(pi0297), .B(pi0199), .Y(new_n30530_));
  AOI21X1  g28094(.A0(new_n28053_), .A1(pi0199), .B0(new_n30470_), .Y(new_n30531_));
  AOI21X1  g28095(.A0(new_n30493_), .A1(pi0456), .B0(new_n30495_), .Y(new_n30532_));
  AOI21X1  g28096(.A0(new_n6074_), .A1(pi0337), .B0(new_n6120_), .Y(new_n30533_));
  OAI22X1  g28097(.A0(new_n30533_), .A1(new_n30532_), .B0(new_n30492_), .B1(new_n6642_), .Y(new_n30534_));
  AOI21X1  g28098(.A0(new_n30472_), .A1(pi0443), .B0(new_n9028_), .Y(new_n30535_));
  NOR2X1   g28099(.A(new_n30535_), .B(new_n30471_), .Y(new_n30536_));
  AOI22X1  g28100(.A0(new_n30536_), .A1(new_n30534_), .B0(new_n30531_), .B1(new_n30530_), .Y(new_n30537_));
  OAI21X1  g28101(.A0(new_n30537_), .A1(new_n10265_), .B0(new_n30529_), .Y(po0823));
  AOI21X1  g28102(.A0(new_n30493_), .A1(pi0319), .B0(new_n30495_), .Y(new_n30539_));
  AOI21X1  g28103(.A0(new_n6074_), .A1(pi0338), .B0(new_n6120_), .Y(new_n30540_));
  OAI22X1  g28104(.A0(new_n30540_), .A1(new_n30539_), .B0(new_n30492_), .B1(new_n6038_), .Y(new_n30541_));
  AOI21X1  g28105(.A0(new_n30472_), .A1(pi0444), .B0(new_n9028_), .Y(new_n30542_));
  NOR2X1   g28106(.A(new_n30542_), .B(new_n30471_), .Y(new_n30543_));
  NOR2X1   g28107(.A(pi0294), .B(pi0199), .Y(new_n30544_));
  OAI22X1  g28108(.A0(pi1072), .A1(new_n7941_), .B0(pi0224), .B1(pi0223), .Y(new_n30545_));
  NOR2X1   g28109(.A(new_n30545_), .B(new_n30544_), .Y(new_n30546_));
  AOI21X1  g28110(.A0(new_n30543_), .A1(new_n30541_), .B0(new_n30546_), .Y(new_n30547_));
  AOI21X1  g28111(.A0(pi1136), .A1(pi0681), .B0(new_n28313_), .Y(new_n30548_));
  OAI21X1  g28112(.A0(pi1136), .A1(new_n11884_), .B0(new_n30548_), .Y(new_n30549_));
  AOI21X1  g28113(.A0(pi1136), .A1(pi0642), .B0(pi1135), .Y(new_n30550_));
  OAI21X1  g28114(.A0(pi1136), .A1(pi0809), .B0(new_n30550_), .Y(new_n30551_));
  AOI21X1  g28115(.A0(new_n30551_), .A1(new_n30549_), .B0(pi1134), .Y(new_n30552_));
  OAI21X1  g28116(.A0(new_n28313_), .A1(pi0699), .B0(pi1136), .Y(new_n30553_));
  AOI21X1  g28117(.A0(new_n28313_), .A1(new_n15495_), .B0(new_n30553_), .Y(new_n30554_));
  OAI21X1  g28118(.A0(new_n30514_), .A1(new_n30314_), .B0(pi1134), .Y(new_n30555_));
  OAI21X1  g28119(.A0(new_n30555_), .A1(new_n30554_), .B0(new_n30516_), .Y(new_n30556_));
  OAI22X1  g28120(.A0(new_n30556_), .A1(new_n30552_), .B0(new_n30547_), .B1(new_n10265_), .Y(po0824));
  AOI21X1  g28121(.A0(pi1135), .A1(new_n5029_), .B0(new_n28946_), .Y(new_n30558_));
  OAI21X1  g28122(.A0(pi1135), .A1(pi0603), .B0(new_n30558_), .Y(new_n30559_));
  AOI21X1  g28123(.A0(pi1135), .A1(new_n11889_), .B0(pi1136), .Y(new_n30560_));
  OAI21X1  g28124(.A0(pi1135), .A1(pi0981), .B0(new_n30560_), .Y(new_n30561_));
  AOI21X1  g28125(.A0(new_n30561_), .A1(new_n30559_), .B0(new_n30477_), .Y(new_n30562_));
  AND2X1   g28126(.A(new_n30484_), .B(new_n14908_), .Y(new_n30563_));
  OAI22X1  g28127(.A0(pi1136), .A1(pi0837), .B0(new_n28313_), .B1(pi0696), .Y(new_n30564_));
  NOR3X1   g28128(.A(new_n30564_), .B(new_n30563_), .C(new_n30487_), .Y(new_n30565_));
  OAI21X1  g28129(.A0(new_n30565_), .A1(new_n30562_), .B0(new_n10265_), .Y(new_n30566_));
  OR2X1    g28130(.A(pi0291), .B(pi0199), .Y(new_n30567_));
  INVX1    g28131(.A(pi1049), .Y(new_n30568_));
  AOI21X1  g28132(.A0(new_n30568_), .A1(pi0199), .B0(new_n30470_), .Y(new_n30569_));
  INVX1    g28133(.A(pi0342), .Y(new_n30570_));
  AOI21X1  g28134(.A0(new_n30493_), .A1(pi0390), .B0(new_n30495_), .Y(new_n30571_));
  AOI21X1  g28135(.A0(new_n6074_), .A1(pi0363), .B0(new_n6120_), .Y(new_n30572_));
  OAI22X1  g28136(.A0(new_n30572_), .A1(new_n30571_), .B0(new_n30492_), .B1(new_n30570_), .Y(new_n30573_));
  AOI21X1  g28137(.A0(new_n30472_), .A1(pi0414), .B0(new_n9028_), .Y(new_n30574_));
  NOR2X1   g28138(.A(new_n30574_), .B(new_n30471_), .Y(new_n30575_));
  AOI22X1  g28139(.A0(new_n30575_), .A1(new_n30573_), .B0(new_n30569_), .B1(new_n30567_), .Y(new_n30576_));
  OAI21X1  g28140(.A0(new_n30576_), .A1(new_n10265_), .B0(new_n30566_), .Y(po0825));
  INVX1    g28141(.A(pi1125), .Y(new_n30578_));
  INVX1    g28142(.A(pi0669), .Y(new_n30579_));
  OAI21X1  g28143(.A0(po0954), .A1(new_n30579_), .B0(new_n30348_), .Y(new_n30580_));
  AOI21X1  g28144(.A0(po0954), .A1(new_n30578_), .B0(new_n30580_), .Y(po0826));
  NOR2X1   g28145(.A(pi0258), .B(pi0199), .Y(new_n30582_));
  OAI22X1  g28146(.A0(pi1062), .A1(new_n7941_), .B0(pi0224), .B1(pi0223), .Y(new_n30583_));
  NOR2X1   g28147(.A(new_n30583_), .B(new_n30582_), .Y(new_n30584_));
  NOR3X1   g28148(.A(pi0592), .B(new_n6074_), .C(new_n6231_), .Y(new_n30585_));
  AOI21X1  g28149(.A0(new_n30464_), .A1(pi0364), .B0(new_n30585_), .Y(new_n30586_));
  AOI21X1  g28150(.A0(new_n30467_), .A1(pi0343), .B0(pi0588), .Y(new_n30587_));
  OAI21X1  g28151(.A0(new_n30586_), .A1(pi0590), .B0(new_n30587_), .Y(new_n30588_));
  AOI21X1  g28152(.A0(new_n30472_), .A1(pi0415), .B0(new_n9028_), .Y(new_n30589_));
  NOR2X1   g28153(.A(new_n30589_), .B(new_n30471_), .Y(new_n30590_));
  AOI21X1  g28154(.A0(new_n30590_), .A1(new_n30588_), .B0(new_n30584_), .Y(new_n30591_));
  AND2X1   g28155(.A(new_n30484_), .B(pi0745), .Y(new_n30592_));
  OAI22X1  g28156(.A0(pi1136), .A1(pi0852), .B0(new_n28313_), .B1(new_n14886_), .Y(new_n30593_));
  NOR3X1   g28157(.A(new_n30593_), .B(new_n30592_), .C(new_n30487_), .Y(new_n30594_));
  INVX1    g28158(.A(new_n30483_), .Y(new_n30595_));
  AND2X1   g28159(.A(pi1135), .B(pi0695), .Y(new_n30596_));
  OAI21X1  g28160(.A0(pi1135), .A1(pi0612), .B0(new_n4755_), .Y(new_n30597_));
  NOR4X1   g28161(.A(new_n30597_), .B(new_n30596_), .C(new_n30595_), .D(new_n28946_), .Y(new_n30598_));
  OAI21X1  g28162(.A0(new_n30598_), .A1(new_n30594_), .B0(new_n10265_), .Y(new_n30599_));
  OAI21X1  g28163(.A0(new_n30591_), .A1(new_n10265_), .B0(new_n30599_), .Y(po0827));
  NOR2X1   g28164(.A(pi0261), .B(pi0199), .Y(new_n30601_));
  OAI22X1  g28165(.A0(pi1040), .A1(new_n7941_), .B0(pi0224), .B1(pi0223), .Y(new_n30602_));
  NOR2X1   g28166(.A(new_n30602_), .B(new_n30601_), .Y(new_n30603_));
  NOR3X1   g28167(.A(pi0592), .B(new_n6074_), .C(new_n6172_), .Y(new_n30604_));
  AOI21X1  g28168(.A0(new_n30464_), .A1(pi0447), .B0(new_n30604_), .Y(new_n30605_));
  AOI21X1  g28169(.A0(new_n30467_), .A1(pi0327), .B0(pi0588), .Y(new_n30606_));
  OAI21X1  g28170(.A0(new_n30605_), .A1(pi0590), .B0(new_n30606_), .Y(new_n30607_));
  AOI21X1  g28171(.A0(new_n30472_), .A1(pi0453), .B0(new_n9028_), .Y(new_n30608_));
  NOR2X1   g28172(.A(new_n30608_), .B(new_n30471_), .Y(new_n30609_));
  AOI21X1  g28173(.A0(new_n30609_), .A1(new_n30607_), .B0(new_n30603_), .Y(new_n30610_));
  AND2X1   g28174(.A(new_n30484_), .B(pi0741), .Y(new_n30611_));
  OAI22X1  g28175(.A0(pi1136), .A1(pi0865), .B0(new_n28313_), .B1(new_n15092_), .Y(new_n30612_));
  NOR3X1   g28176(.A(new_n30612_), .B(new_n30611_), .C(new_n30487_), .Y(new_n30613_));
  AND2X1   g28177(.A(pi1135), .B(pi0646), .Y(new_n30614_));
  OAI21X1  g28178(.A0(pi1135), .A1(pi0611), .B0(new_n4755_), .Y(new_n30615_));
  NOR4X1   g28179(.A(new_n30615_), .B(new_n30614_), .C(new_n30595_), .D(new_n28946_), .Y(new_n30616_));
  OAI21X1  g28180(.A0(new_n30616_), .A1(new_n30613_), .B0(new_n10265_), .Y(new_n30617_));
  OAI21X1  g28181(.A0(new_n30610_), .A1(new_n10265_), .B0(new_n30617_), .Y(po0828));
  AOI21X1  g28182(.A0(pi1135), .A1(new_n11976_), .B0(new_n28946_), .Y(new_n30619_));
  OAI21X1  g28183(.A0(pi1135), .A1(pi0616), .B0(new_n30619_), .Y(new_n30620_));
  AOI21X1  g28184(.A0(pi1135), .A1(new_n11887_), .B0(pi1136), .Y(new_n30621_));
  OAI21X1  g28185(.A0(pi1135), .A1(pi0808), .B0(new_n30621_), .Y(new_n30622_));
  AOI21X1  g28186(.A0(new_n30622_), .A1(new_n30620_), .B0(new_n30477_), .Y(new_n30623_));
  AND2X1   g28187(.A(new_n30484_), .B(new_n13973_), .Y(new_n30624_));
  OAI22X1  g28188(.A0(pi1136), .A1(pi0850), .B0(new_n28313_), .B1(pi0736), .Y(new_n30625_));
  NOR3X1   g28189(.A(new_n30625_), .B(new_n30624_), .C(new_n30487_), .Y(new_n30626_));
  OAI21X1  g28190(.A0(new_n30626_), .A1(new_n30623_), .B0(new_n10265_), .Y(new_n30627_));
  NOR2X1   g28191(.A(pi0290), .B(pi0199), .Y(new_n30628_));
  OAI22X1  g28192(.A0(pi1048), .A1(new_n7941_), .B0(pi0224), .B1(pi0223), .Y(new_n30629_));
  NOR2X1   g28193(.A(new_n30629_), .B(new_n30628_), .Y(new_n30630_));
  INVX1    g28194(.A(pi0320), .Y(new_n30631_));
  AOI21X1  g28195(.A0(new_n30493_), .A1(pi0397), .B0(new_n30495_), .Y(new_n30632_));
  AOI21X1  g28196(.A0(new_n6074_), .A1(pi0372), .B0(new_n6120_), .Y(new_n30633_));
  OAI22X1  g28197(.A0(new_n30633_), .A1(new_n30632_), .B0(new_n30492_), .B1(new_n30631_), .Y(new_n30634_));
  AOI21X1  g28198(.A0(new_n30472_), .A1(pi0422), .B0(new_n9028_), .Y(new_n30635_));
  NOR2X1   g28199(.A(new_n30635_), .B(new_n30471_), .Y(new_n30636_));
  AOI21X1  g28200(.A0(new_n30636_), .A1(new_n30634_), .B0(new_n30630_), .Y(new_n30637_));
  OAI21X1  g28201(.A0(new_n30637_), .A1(new_n10265_), .B0(new_n30627_), .Y(po0829));
  AOI21X1  g28202(.A0(pi1135), .A1(new_n22270_), .B0(new_n28946_), .Y(new_n30639_));
  OAI21X1  g28203(.A0(pi1135), .A1(pi0617), .B0(new_n30639_), .Y(new_n30640_));
  AOI21X1  g28204(.A0(new_n28313_), .A1(pi0814), .B0(pi1136), .Y(new_n30641_));
  OAI21X1  g28205(.A0(new_n28313_), .A1(pi0788), .B0(new_n30641_), .Y(new_n30642_));
  AOI21X1  g28206(.A0(new_n30642_), .A1(new_n30640_), .B0(new_n30477_), .Y(new_n30643_));
  AND2X1   g28207(.A(new_n30484_), .B(new_n12911_), .Y(new_n30644_));
  OAI22X1  g28208(.A0(pi1136), .A1(pi0866), .B0(new_n28313_), .B1(pi0706), .Y(new_n30645_));
  NOR3X1   g28209(.A(new_n30645_), .B(new_n30644_), .C(new_n30487_), .Y(new_n30646_));
  OAI21X1  g28210(.A0(new_n30646_), .A1(new_n30643_), .B0(new_n10265_), .Y(new_n30647_));
  OR2X1    g28211(.A(pi0295), .B(pi0199), .Y(new_n30648_));
  AOI21X1  g28212(.A0(new_n27695_), .A1(pi0199), .B0(new_n30470_), .Y(new_n30649_));
  AOI21X1  g28213(.A0(new_n30493_), .A1(pi0411), .B0(new_n30495_), .Y(new_n30650_));
  AOI21X1  g28214(.A0(new_n6074_), .A1(pi0387), .B0(new_n6120_), .Y(new_n30651_));
  OAI22X1  g28215(.A0(new_n30651_), .A1(new_n30650_), .B0(new_n30492_), .B1(new_n6024_), .Y(new_n30652_));
  AOI21X1  g28216(.A0(new_n30472_), .A1(pi0435), .B0(new_n9028_), .Y(new_n30653_));
  NOR2X1   g28217(.A(new_n30653_), .B(new_n30471_), .Y(new_n30654_));
  AOI22X1  g28218(.A0(new_n30654_), .A1(new_n30652_), .B0(new_n30649_), .B1(new_n30648_), .Y(new_n30655_));
  OAI21X1  g28219(.A0(new_n30655_), .A1(new_n10265_), .B0(new_n30647_), .Y(po0830));
  NOR2X1   g28220(.A(pi0256), .B(pi0199), .Y(new_n30657_));
  OAI22X1  g28221(.A0(pi1070), .A1(new_n7941_), .B0(pi0224), .B1(pi0223), .Y(new_n30658_));
  NOR2X1   g28222(.A(new_n30658_), .B(new_n30657_), .Y(new_n30659_));
  AND2X1   g28223(.A(pi0591), .B(pi0463), .Y(new_n30660_));
  AOI22X1  g28224(.A0(new_n30660_), .A1(new_n6120_), .B0(new_n30464_), .B1(pi0336), .Y(new_n30661_));
  AOI21X1  g28225(.A0(new_n30467_), .A1(pi0362), .B0(pi0588), .Y(new_n30662_));
  OAI21X1  g28226(.A0(new_n30661_), .A1(pi0590), .B0(new_n30662_), .Y(new_n30663_));
  AOI21X1  g28227(.A0(new_n30472_), .A1(pi0437), .B0(new_n9028_), .Y(new_n30664_));
  NOR2X1   g28228(.A(new_n30664_), .B(new_n30471_), .Y(new_n30665_));
  AOI21X1  g28229(.A0(new_n30665_), .A1(new_n30663_), .B0(new_n30659_), .Y(new_n30666_));
  AOI21X1  g28230(.A0(pi1135), .A1(pi0639), .B0(new_n28946_), .Y(new_n30667_));
  OAI21X1  g28231(.A0(pi1135), .A1(new_n23196_), .B0(new_n30667_), .Y(new_n30668_));
  AOI21X1  g28232(.A0(pi1135), .A1(pi0783), .B0(pi1136), .Y(new_n30669_));
  OAI21X1  g28233(.A0(pi1135), .A1(new_n29342_), .B0(new_n30669_), .Y(new_n30670_));
  AOI21X1  g28234(.A0(new_n30670_), .A1(new_n30668_), .B0(pi1134), .Y(new_n30671_));
  OAI21X1  g28235(.A0(new_n28313_), .A1(pi0735), .B0(pi1136), .Y(new_n30672_));
  AOI21X1  g28236(.A0(new_n28313_), .A1(new_n13220_), .B0(new_n30672_), .Y(new_n30673_));
  AND2X1   g28237(.A(new_n30513_), .B(pi0859), .Y(new_n30674_));
  OR2X1    g28238(.A(new_n30674_), .B(new_n4755_), .Y(new_n30675_));
  OAI21X1  g28239(.A0(new_n30675_), .A1(new_n30673_), .B0(new_n30516_), .Y(new_n30676_));
  OAI22X1  g28240(.A0(new_n30676_), .A1(new_n30671_), .B0(new_n30666_), .B1(new_n10265_), .Y(po0831));
  INVX1    g28241(.A(new_n30486_), .Y(new_n30678_));
  OR2X1    g28242(.A(pi1135), .B(pi0748), .Y(new_n30679_));
  AOI21X1  g28243(.A0(pi1135), .A1(new_n21514_), .B0(new_n28946_), .Y(new_n30680_));
  AOI22X1  g28244(.A0(new_n30680_), .A1(new_n30679_), .B0(new_n30513_), .B1(pi0876), .Y(new_n30681_));
  AND2X1   g28245(.A(new_n30484_), .B(new_n22925_), .Y(new_n30682_));
  NOR3X1   g28246(.A(pi1136), .B(new_n28313_), .C(new_n11886_), .Y(new_n30683_));
  OAI21X1  g28247(.A0(new_n28313_), .A1(pi0710), .B0(pi1136), .Y(new_n30684_));
  OAI21X1  g28248(.A0(pi1135), .A1(pi0803), .B0(new_n30684_), .Y(new_n30685_));
  OAI21X1  g28249(.A0(new_n30685_), .A1(new_n30683_), .B0(new_n30476_), .Y(new_n30686_));
  OAI22X1  g28250(.A0(new_n30686_), .A1(new_n30682_), .B0(new_n30681_), .B1(new_n30678_), .Y(new_n30687_));
  AOI21X1  g28251(.A0(new_n28057_), .A1(pi0199), .B0(new_n30470_), .Y(new_n30688_));
  OAI21X1  g28252(.A0(pi0296), .A1(pi0199), .B0(new_n30688_), .Y(new_n30689_));
  NAND3X1  g28253(.A(pi0591), .B(new_n6168_), .C(pi0412), .Y(new_n30690_));
  NAND2X1  g28254(.A(new_n30690_), .B(new_n30494_), .Y(new_n30691_));
  INVX1    g28255(.A(pi0388), .Y(new_n30692_));
  OAI21X1  g28256(.A0(pi0591), .A1(new_n30692_), .B0(pi0592), .Y(new_n30693_));
  AOI22X1  g28257(.A0(new_n30693_), .A1(new_n30691_), .B0(new_n30467_), .B1(pi0455), .Y(new_n30694_));
  AOI21X1  g28258(.A0(new_n30472_), .A1(pi0436), .B0(new_n9028_), .Y(new_n30695_));
  OR2X1    g28259(.A(new_n30695_), .B(new_n30471_), .Y(new_n30696_));
  OAI21X1  g28260(.A0(new_n30696_), .A1(new_n30694_), .B0(new_n30689_), .Y(new_n30697_));
  MX2X1    g28261(.A(new_n30697_), .B(new_n30687_), .S0(new_n10265_), .Y(po0832));
  AOI21X1  g28262(.A0(pi1135), .A1(new_n22461_), .B0(new_n28946_), .Y(new_n30699_));
  OAI21X1  g28263(.A0(pi1135), .A1(pi0606), .B0(new_n30699_), .Y(new_n30700_));
  AOI21X1  g28264(.A0(new_n28313_), .A1(pi0812), .B0(pi1136), .Y(new_n30701_));
  OAI21X1  g28265(.A0(new_n28313_), .A1(pi0787), .B0(new_n30701_), .Y(new_n30702_));
  AOI21X1  g28266(.A0(new_n30702_), .A1(new_n30700_), .B0(new_n30477_), .Y(new_n30703_));
  AND2X1   g28267(.A(new_n30484_), .B(new_n15545_), .Y(new_n30704_));
  OAI22X1  g28268(.A0(pi1136), .A1(pi0881), .B0(new_n28313_), .B1(pi0729), .Y(new_n30705_));
  NOR3X1   g28269(.A(new_n30705_), .B(new_n30704_), .C(new_n30487_), .Y(new_n30706_));
  OAI21X1  g28270(.A0(new_n30706_), .A1(new_n30703_), .B0(new_n10265_), .Y(new_n30707_));
  NOR2X1   g28271(.A(pi0293), .B(pi0199), .Y(new_n30708_));
  OAI22X1  g28272(.A0(pi1059), .A1(new_n7941_), .B0(pi0224), .B1(pi0223), .Y(new_n30709_));
  NOR2X1   g28273(.A(new_n30709_), .B(new_n30708_), .Y(new_n30710_));
  AOI21X1  g28274(.A0(new_n30493_), .A1(pi0410), .B0(new_n30495_), .Y(new_n30711_));
  AOI21X1  g28275(.A0(new_n6074_), .A1(pi0386), .B0(new_n6120_), .Y(new_n30712_));
  OAI22X1  g28276(.A0(new_n30712_), .A1(new_n30711_), .B0(new_n30492_), .B1(new_n6029_), .Y(new_n30713_));
  AOI21X1  g28277(.A0(new_n30472_), .A1(pi0434), .B0(new_n9028_), .Y(new_n30714_));
  NOR2X1   g28278(.A(new_n30714_), .B(new_n30471_), .Y(new_n30715_));
  AOI21X1  g28279(.A0(new_n30715_), .A1(new_n30713_), .B0(new_n30710_), .Y(new_n30716_));
  OAI21X1  g28280(.A0(new_n30716_), .A1(new_n10265_), .B0(new_n30707_), .Y(po0833));
  NOR2X1   g28281(.A(pi0259), .B(pi0199), .Y(new_n30718_));
  OAI22X1  g28282(.A0(pi1069), .A1(new_n7941_), .B0(pi0224), .B1(pi0223), .Y(new_n30719_));
  NOR2X1   g28283(.A(new_n30719_), .B(new_n30718_), .Y(new_n30720_));
  NOR3X1   g28284(.A(pi0592), .B(new_n6074_), .C(new_n6237_), .Y(new_n30721_));
  AOI21X1  g28285(.A0(new_n30464_), .A1(pi0366), .B0(new_n30721_), .Y(new_n30722_));
  AOI21X1  g28286(.A0(new_n30467_), .A1(pi0344), .B0(pi0588), .Y(new_n30723_));
  OAI21X1  g28287(.A0(new_n30722_), .A1(pi0590), .B0(new_n30723_), .Y(new_n30724_));
  AOI21X1  g28288(.A0(new_n30472_), .A1(pi0416), .B0(new_n9028_), .Y(new_n30725_));
  NOR2X1   g28289(.A(new_n30725_), .B(new_n30471_), .Y(new_n30726_));
  AOI21X1  g28290(.A0(new_n30726_), .A1(new_n30724_), .B0(new_n30720_), .Y(new_n30727_));
  AND2X1   g28291(.A(new_n30484_), .B(pi0742), .Y(new_n30728_));
  OAI22X1  g28292(.A0(pi1136), .A1(pi0870), .B0(new_n28313_), .B1(new_n16615_), .Y(new_n30729_));
  NOR3X1   g28293(.A(new_n30729_), .B(new_n30728_), .C(new_n30487_), .Y(new_n30730_));
  AND2X1   g28294(.A(pi1135), .B(pi0635), .Y(new_n30731_));
  OAI21X1  g28295(.A0(pi1135), .A1(pi0620), .B0(new_n4755_), .Y(new_n30732_));
  NOR4X1   g28296(.A(new_n30732_), .B(new_n30731_), .C(new_n30595_), .D(new_n28946_), .Y(new_n30733_));
  OAI21X1  g28297(.A0(new_n30733_), .A1(new_n30730_), .B0(new_n10265_), .Y(new_n30734_));
  OAI21X1  g28298(.A0(new_n30727_), .A1(new_n10265_), .B0(new_n30734_), .Y(po0834));
  NOR2X1   g28299(.A(pi0260), .B(pi0199), .Y(new_n30736_));
  OAI22X1  g28300(.A0(pi1067), .A1(new_n7941_), .B0(pi0224), .B1(pi0223), .Y(new_n30737_));
  NOR2X1   g28301(.A(new_n30737_), .B(new_n30736_), .Y(new_n30738_));
  NOR3X1   g28302(.A(pi0592), .B(new_n6074_), .C(new_n6170_), .Y(new_n30739_));
  AOI21X1  g28303(.A0(new_n30464_), .A1(pi0368), .B0(new_n30739_), .Y(new_n30740_));
  AOI21X1  g28304(.A0(new_n30467_), .A1(pi0346), .B0(pi0588), .Y(new_n30741_));
  OAI21X1  g28305(.A0(new_n30740_), .A1(pi0590), .B0(new_n30741_), .Y(new_n30742_));
  AOI21X1  g28306(.A0(new_n30472_), .A1(pi0418), .B0(new_n9028_), .Y(new_n30743_));
  NOR2X1   g28307(.A(new_n30743_), .B(new_n30471_), .Y(new_n30744_));
  AOI21X1  g28308(.A0(new_n30744_), .A1(new_n30742_), .B0(new_n30738_), .Y(new_n30745_));
  AND2X1   g28309(.A(new_n30484_), .B(pi0760), .Y(new_n30746_));
  OAI22X1  g28310(.A0(pi1136), .A1(pi0856), .B0(new_n28313_), .B1(new_n15112_), .Y(new_n30747_));
  NOR3X1   g28311(.A(new_n30747_), .B(new_n30746_), .C(new_n30487_), .Y(new_n30748_));
  AND2X1   g28312(.A(pi1135), .B(pi0632), .Y(new_n30749_));
  OAI21X1  g28313(.A0(pi1135), .A1(pi0613), .B0(new_n4755_), .Y(new_n30750_));
  NOR4X1   g28314(.A(new_n30750_), .B(new_n30749_), .C(new_n30595_), .D(new_n28946_), .Y(new_n30751_));
  OAI21X1  g28315(.A0(new_n30751_), .A1(new_n30748_), .B0(new_n10265_), .Y(new_n30752_));
  OAI21X1  g28316(.A0(new_n30745_), .A1(new_n10265_), .B0(new_n30752_), .Y(po0835));
  NOR2X1   g28317(.A(pi0255), .B(pi0199), .Y(new_n30754_));
  OAI22X1  g28318(.A0(pi1036), .A1(new_n7941_), .B0(pi0224), .B1(pi0223), .Y(new_n30755_));
  NOR2X1   g28319(.A(new_n30755_), .B(new_n30754_), .Y(new_n30756_));
  AND2X1   g28320(.A(pi0591), .B(pi0413), .Y(new_n30757_));
  AOI22X1  g28321(.A0(new_n30757_), .A1(new_n6120_), .B0(new_n30464_), .B1(pi0389), .Y(new_n30758_));
  AOI21X1  g28322(.A0(new_n30467_), .A1(pi0450), .B0(pi0588), .Y(new_n30759_));
  OAI21X1  g28323(.A0(new_n30758_), .A1(pi0590), .B0(new_n30759_), .Y(new_n30760_));
  AOI21X1  g28324(.A0(new_n30472_), .A1(pi0438), .B0(new_n9028_), .Y(new_n30761_));
  NOR2X1   g28325(.A(new_n30761_), .B(new_n30471_), .Y(new_n30762_));
  AOI21X1  g28326(.A0(new_n30762_), .A1(new_n30760_), .B0(new_n30756_), .Y(new_n30763_));
  AOI21X1  g28327(.A0(pi1136), .A1(new_n12255_), .B0(new_n28313_), .Y(new_n30764_));
  OAI21X1  g28328(.A0(pi1136), .A1(pi0791), .B0(new_n30764_), .Y(new_n30765_));
  AOI21X1  g28329(.A0(pi1136), .A1(new_n12092_), .B0(pi1135), .Y(new_n30766_));
  OAI21X1  g28330(.A0(pi1136), .A1(pi0810), .B0(new_n30766_), .Y(new_n30767_));
  AOI21X1  g28331(.A0(new_n30767_), .A1(new_n30765_), .B0(new_n30477_), .Y(new_n30768_));
  AND2X1   g28332(.A(new_n30484_), .B(new_n15697_), .Y(new_n30769_));
  OAI22X1  g28333(.A0(pi1136), .A1(pi0874), .B0(new_n28313_), .B1(pi0690), .Y(new_n30770_));
  NOR3X1   g28334(.A(new_n30770_), .B(new_n30769_), .C(new_n30487_), .Y(new_n30771_));
  OAI21X1  g28335(.A0(new_n30771_), .A1(new_n30768_), .B0(new_n10265_), .Y(new_n30772_));
  OAI21X1  g28336(.A0(new_n30763_), .A1(new_n10265_), .B0(new_n30772_), .Y(po0836));
  OAI21X1  g28337(.A0(new_n30347_), .A1(pi1100), .B0(new_n30348_), .Y(new_n30774_));
  AOI21X1  g28338(.A0(new_n30347_), .A1(new_n5029_), .B0(new_n30774_), .Y(po0837));
  OAI21X1  g28339(.A0(new_n30347_), .A1(pi1103), .B0(new_n30348_), .Y(new_n30776_));
  AOI21X1  g28340(.A0(new_n30347_), .A1(new_n11949_), .B0(new_n30776_), .Y(po0838));
  NOR2X1   g28341(.A(pi0251), .B(pi0199), .Y(new_n30778_));
  OAI22X1  g28342(.A0(pi1039), .A1(new_n7941_), .B0(pi0224), .B1(pi0223), .Y(new_n30779_));
  NOR2X1   g28343(.A(new_n30779_), .B(new_n30778_), .Y(new_n30780_));
  NOR3X1   g28344(.A(pi0592), .B(new_n6074_), .C(new_n6171_), .Y(new_n30781_));
  AOI21X1  g28345(.A0(new_n30464_), .A1(pi0367), .B0(new_n30781_), .Y(new_n30782_));
  AOI21X1  g28346(.A0(new_n30467_), .A1(pi0345), .B0(pi0588), .Y(new_n30783_));
  OAI21X1  g28347(.A0(new_n30782_), .A1(pi0590), .B0(new_n30783_), .Y(new_n30784_));
  AOI21X1  g28348(.A0(new_n30472_), .A1(pi0417), .B0(new_n9028_), .Y(new_n30785_));
  NOR2X1   g28349(.A(new_n30785_), .B(new_n30471_), .Y(new_n30786_));
  AOI21X1  g28350(.A0(new_n30786_), .A1(new_n30784_), .B0(new_n30780_), .Y(new_n30787_));
  AND2X1   g28351(.A(new_n30484_), .B(pi0757), .Y(new_n30788_));
  OAI22X1  g28352(.A0(pi1136), .A1(pi0848), .B0(new_n28313_), .B1(new_n16855_), .Y(new_n30789_));
  NOR3X1   g28353(.A(new_n30789_), .B(new_n30788_), .C(new_n30487_), .Y(new_n30790_));
  AND2X1   g28354(.A(pi1135), .B(pi0631), .Y(new_n30791_));
  OAI21X1  g28355(.A0(pi1135), .A1(pi0610), .B0(new_n4755_), .Y(new_n30792_));
  NOR4X1   g28356(.A(new_n30792_), .B(new_n30791_), .C(new_n30595_), .D(new_n28946_), .Y(new_n30793_));
  OAI21X1  g28357(.A0(new_n30793_), .A1(new_n30790_), .B0(new_n10265_), .Y(new_n30794_));
  OAI21X1  g28358(.A0(new_n30787_), .A1(new_n10265_), .B0(new_n30794_), .Y(po0839));
  INVX1    g28359(.A(pi0953), .Y(new_n30796_));
  NOR4X1   g28360(.A(new_n30345_), .B(pi0973), .C(new_n30796_), .D(new_n12898_), .Y(po0980));
  INVX1    g28361(.A(pi0684), .Y(new_n30798_));
  OAI21X1  g28362(.A0(po0980), .A1(new_n30798_), .B0(new_n30348_), .Y(new_n30799_));
  AOI21X1  g28363(.A0(po0980), .A1(new_n30425_), .B0(new_n30799_), .Y(po0841));
  INVX1    g28364(.A(new_n28055_), .Y(new_n30801_));
  AND2X1   g28365(.A(pi0592), .B(new_n6168_), .Y(new_n30802_));
  AND2X1   g28366(.A(new_n6120_), .B(pi0590), .Y(new_n30803_));
  AOI22X1  g28367(.A0(new_n30803_), .A1(pi0357), .B0(new_n30802_), .B1(pi0382), .Y(new_n30804_));
  OR4X1    g28368(.A(pi0592), .B(new_n6074_), .C(pi0590), .D(new_n6203_), .Y(new_n30805_));
  OAI21X1  g28369(.A0(new_n30804_), .A1(pi0591), .B0(new_n30805_), .Y(new_n30806_));
  OR2X1    g28370(.A(pi0592), .B(pi0591), .Y(new_n30807_));
  NOR4X1   g28371(.A(new_n30807_), .B(pi0590), .C(new_n9028_), .D(new_n6582_), .Y(new_n30808_));
  AOI21X1  g28372(.A0(new_n30806_), .A1(new_n9028_), .B0(new_n30808_), .Y(new_n30809_));
  OAI22X1  g28373(.A0(pi1076), .A1(new_n7941_), .B0(pi0224), .B1(pi0223), .Y(new_n30810_));
  OAI22X1  g28374(.A0(new_n30810_), .A1(new_n30801_), .B0(new_n30809_), .B1(new_n30471_), .Y(new_n30811_));
  NAND2X1  g28375(.A(new_n28313_), .B(pi0744), .Y(new_n30812_));
  AOI21X1  g28376(.A0(pi1135), .A1(pi0728), .B0(new_n28946_), .Y(new_n30813_));
  AOI22X1  g28377(.A0(new_n30813_), .A1(new_n30812_), .B0(new_n30513_), .B1(pi0860), .Y(new_n30814_));
  OAI21X1  g28378(.A0(new_n30483_), .A1(new_n28946_), .B0(new_n4755_), .Y(new_n30815_));
  OR2X1    g28379(.A(pi1135), .B(pi0652), .Y(new_n30816_));
  AOI21X1  g28380(.A0(pi1135), .A1(pi0657), .B0(new_n28946_), .Y(new_n30817_));
  AND2X1   g28381(.A(new_n30483_), .B(pi0813), .Y(new_n30818_));
  AOI22X1  g28382(.A0(new_n30818_), .A1(new_n30513_), .B0(new_n30817_), .B1(new_n30816_), .Y(new_n30819_));
  OAI22X1  g28383(.A0(new_n30819_), .A1(new_n30815_), .B0(new_n30814_), .B1(new_n30678_), .Y(new_n30820_));
  MX2X1    g28384(.A(new_n30820_), .B(new_n30811_), .S0(new_n6748_), .Y(po0842));
  OAI21X1  g28385(.A0(po0980), .A1(new_n16855_), .B0(new_n30348_), .Y(new_n30822_));
  AOI21X1  g28386(.A0(po0980), .A1(new_n30361_), .B0(new_n30822_), .Y(po0843));
  INVX1    g28387(.A(po0980), .Y(new_n30824_));
  OAI21X1  g28388(.A0(new_n30824_), .A1(pi1127), .B0(new_n30348_), .Y(new_n30825_));
  AOI21X1  g28389(.A0(new_n30824_), .A1(new_n13680_), .B0(new_n30825_), .Y(po0844));
  OAI21X1  g28390(.A0(po0980), .A1(new_n15112_), .B0(new_n30348_), .Y(new_n30827_));
  AOI21X1  g28391(.A0(po0980), .A1(new_n30365_), .B0(new_n30827_), .Y(po0845));
  AOI22X1  g28392(.A0(new_n30803_), .A1(pi0351), .B0(new_n30802_), .B1(pi0376), .Y(new_n30829_));
  NAND4X1  g28393(.A(new_n6120_), .B(pi0591), .C(new_n6168_), .D(pi0401), .Y(new_n30830_));
  OAI21X1  g28394(.A0(new_n30829_), .A1(pi0591), .B0(new_n30830_), .Y(new_n30831_));
  NOR4X1   g28395(.A(new_n30807_), .B(pi0590), .C(new_n9028_), .D(new_n6585_), .Y(new_n30832_));
  AOI21X1  g28396(.A0(new_n30831_), .A1(new_n9028_), .B0(new_n30832_), .Y(new_n30833_));
  NOR2X1   g28397(.A(new_n28043_), .B(pi0199), .Y(new_n30834_));
  OAI22X1  g28398(.A0(pi1079), .A1(new_n7941_), .B0(pi0224), .B1(pi0223), .Y(new_n30835_));
  OAI22X1  g28399(.A0(new_n30835_), .A1(new_n30834_), .B0(new_n30833_), .B1(new_n30471_), .Y(new_n30836_));
  OR2X1    g28400(.A(pi1135), .B(pi0658), .Y(new_n30837_));
  AOI21X1  g28401(.A0(pi1135), .A1(pi0655), .B0(new_n28946_), .Y(new_n30838_));
  AOI22X1  g28402(.A0(new_n30838_), .A1(new_n30837_), .B0(new_n30513_), .B1(pi0798), .Y(new_n30839_));
  AND2X1   g28403(.A(new_n30484_), .B(pi0752), .Y(new_n30840_));
  OAI22X1  g28404(.A0(pi1136), .A1(pi0843), .B0(new_n28313_), .B1(pi0703), .Y(new_n30841_));
  OR2X1    g28405(.A(new_n30841_), .B(new_n30487_), .Y(new_n30842_));
  OAI22X1  g28406(.A0(new_n30842_), .A1(new_n30840_), .B0(new_n30839_), .B1(new_n30477_), .Y(new_n30843_));
  MX2X1    g28407(.A(new_n30843_), .B(new_n30836_), .S0(new_n6748_), .Y(po0846));
  OAI21X1  g28408(.A0(new_n30824_), .A1(pi1108), .B0(new_n30348_), .Y(new_n30845_));
  AOI21X1  g28409(.A0(new_n30824_), .A1(new_n15732_), .B0(new_n30845_), .Y(po0847));
  OAI21X1  g28410(.A0(new_n30824_), .A1(pi1107), .B0(new_n30348_), .Y(new_n30847_));
  AOI21X1  g28411(.A0(new_n30824_), .A1(new_n15681_), .B0(new_n30847_), .Y(po0848));
  NAND3X1  g28412(.A(new_n6120_), .B(pi0590), .C(pi0352), .Y(new_n30849_));
  NAND3X1  g28413(.A(pi0592), .B(new_n6168_), .C(pi0317), .Y(new_n30850_));
  AOI21X1  g28414(.A0(new_n30850_), .A1(new_n30849_), .B0(pi0591), .Y(new_n30851_));
  AND2X1   g28415(.A(new_n6120_), .B(pi0402), .Y(new_n30852_));
  AOI21X1  g28416(.A0(new_n30852_), .A1(new_n30493_), .B0(new_n30851_), .Y(new_n30853_));
  OR4X1    g28417(.A(new_n30807_), .B(pi0590), .C(new_n9028_), .D(new_n6527_), .Y(new_n30854_));
  OAI21X1  g28418(.A0(new_n30853_), .A1(pi0588), .B0(new_n30854_), .Y(new_n30855_));
  NOR2X1   g28419(.A(new_n28047_), .B(pi0199), .Y(new_n30856_));
  OAI22X1  g28420(.A0(pi1078), .A1(new_n7941_), .B0(pi0224), .B1(pi0223), .Y(new_n30857_));
  NOR2X1   g28421(.A(new_n30857_), .B(new_n30856_), .Y(new_n30858_));
  AOI21X1  g28422(.A0(new_n30855_), .A1(new_n30470_), .B0(new_n30858_), .Y(new_n30859_));
  AOI21X1  g28423(.A0(new_n28313_), .A1(pi0770), .B0(new_n28946_), .Y(new_n30860_));
  OAI21X1  g28424(.A0(new_n28313_), .A1(pi0726), .B0(new_n30860_), .Y(new_n30861_));
  AOI21X1  g28425(.A0(new_n30513_), .A1(pi0844), .B0(new_n4755_), .Y(new_n30862_));
  AND2X1   g28426(.A(new_n30862_), .B(new_n30861_), .Y(new_n30863_));
  OR2X1    g28427(.A(pi1135), .B(pi0656), .Y(new_n30864_));
  AOI21X1  g28428(.A0(pi1135), .A1(pi0649), .B0(new_n28946_), .Y(new_n30865_));
  INVX1    g28429(.A(pi0801), .Y(new_n30866_));
  OAI21X1  g28430(.A0(new_n30514_), .A1(new_n30866_), .B0(new_n4755_), .Y(new_n30867_));
  AOI21X1  g28431(.A0(new_n30865_), .A1(new_n30864_), .B0(new_n30867_), .Y(new_n30868_));
  OR4X1    g28432(.A(new_n30868_), .B(new_n30863_), .C(new_n30595_), .D(new_n6748_), .Y(new_n30869_));
  OAI21X1  g28433(.A0(new_n30859_), .A1(new_n10265_), .B0(new_n30869_), .Y(po0849));
  INVX1    g28434(.A(pi1129), .Y(new_n30871_));
  INVX1    g28435(.A(pi0693), .Y(new_n30872_));
  OAI21X1  g28436(.A0(po0954), .A1(new_n30872_), .B0(new_n30348_), .Y(new_n30873_));
  AOI21X1  g28437(.A0(po0954), .A1(new_n30871_), .B0(new_n30873_), .Y(po0850));
  INVX1    g28438(.A(pi1128), .Y(new_n30875_));
  INVX1    g28439(.A(pi0694), .Y(new_n30876_));
  OAI21X1  g28440(.A0(po0980), .A1(new_n30876_), .B0(new_n30348_), .Y(new_n30877_));
  AOI21X1  g28441(.A0(po0980), .A1(new_n30875_), .B0(new_n30877_), .Y(po0851));
  INVX1    g28442(.A(pi1111), .Y(new_n30879_));
  OAI21X1  g28443(.A0(po0954), .A1(new_n23523_), .B0(new_n30348_), .Y(new_n30880_));
  AOI21X1  g28444(.A0(po0954), .A1(new_n30879_), .B0(new_n30880_), .Y(po0852));
  OAI21X1  g28445(.A0(new_n30824_), .A1(pi1100), .B0(new_n30348_), .Y(new_n30882_));
  AOI21X1  g28446(.A0(new_n30824_), .A1(new_n14944_), .B0(new_n30882_), .Y(po0853));
  INVX1    g28447(.A(pi0697), .Y(new_n30884_));
  OAI21X1  g28448(.A0(po0980), .A1(new_n30884_), .B0(new_n30348_), .Y(new_n30885_));
  AOI21X1  g28449(.A0(po0980), .A1(new_n30871_), .B0(new_n30885_), .Y(po0854));
  INVX1    g28450(.A(pi1116), .Y(new_n30887_));
  OAI21X1  g28451(.A0(po0980), .A1(new_n14306_), .B0(new_n30348_), .Y(new_n30888_));
  AOI21X1  g28452(.A0(po0980), .A1(new_n30887_), .B0(new_n30888_), .Y(po0855));
  OAI21X1  g28453(.A0(new_n30824_), .A1(pi1103), .B0(new_n30348_), .Y(new_n30890_));
  AOI21X1  g28454(.A0(new_n30824_), .A1(new_n15535_), .B0(new_n30890_), .Y(po0856));
  OAI21X1  g28455(.A0(new_n30824_), .A1(pi1110), .B0(new_n30348_), .Y(new_n30892_));
  AOI21X1  g28456(.A0(new_n30824_), .A1(new_n15022_), .B0(new_n30892_), .Y(po0857));
  INVX1    g28457(.A(pi1123), .Y(new_n30894_));
  OAI21X1  g28458(.A0(po0980), .A1(new_n14840_), .B0(new_n30348_), .Y(new_n30895_));
  AOI21X1  g28459(.A0(po0980), .A1(new_n30894_), .B0(new_n30895_), .Y(po0858));
  INVX1    g28460(.A(pi1117), .Y(new_n30897_));
  OAI21X1  g28461(.A0(po0980), .A1(new_n15160_), .B0(new_n30348_), .Y(new_n30898_));
  AOI21X1  g28462(.A0(po0980), .A1(new_n30897_), .B0(new_n30898_), .Y(po0859));
  OAI21X1  g28463(.A0(new_n30824_), .A1(pi1124), .B0(new_n30348_), .Y(new_n30900_));
  AOI21X1  g28464(.A0(new_n30824_), .A1(new_n15364_), .B0(new_n30900_), .Y(po0860));
  OAI21X1  g28465(.A0(po0980), .A1(new_n16615_), .B0(new_n30348_), .Y(new_n30902_));
  AOI21X1  g28466(.A0(po0980), .A1(new_n30373_), .B0(new_n30902_), .Y(po0861));
  OAI21X1  g28467(.A0(new_n30824_), .A1(pi1125), .B0(new_n30348_), .Y(new_n30904_));
  AOI21X1  g28468(.A0(new_n30824_), .A1(new_n15470_), .B0(new_n30904_), .Y(po0862));
  OAI21X1  g28469(.A0(new_n30824_), .A1(pi1105), .B0(new_n30348_), .Y(new_n30906_));
  AOI21X1  g28470(.A0(new_n30824_), .A1(new_n12934_), .B0(new_n30906_), .Y(po0863));
  INVX1    g28471(.A(new_n30464_), .Y(new_n30908_));
  NAND3X1  g28472(.A(new_n6120_), .B(pi0591), .C(pi0395), .Y(new_n30909_));
  OAI21X1  g28473(.A0(new_n30908_), .A1(new_n6081_), .B0(new_n30909_), .Y(new_n30910_));
  AOI22X1  g28474(.A0(new_n30910_), .A1(new_n6168_), .B0(new_n30467_), .B1(pi0347), .Y(new_n30911_));
  NOR3X1   g28475(.A(pi0588), .B(pi0224), .C(pi0223), .Y(new_n30912_));
  INVX1    g28476(.A(new_n30912_), .Y(new_n30913_));
  MX2X1    g28477(.A(pi0304), .B(pi1048), .S0(pi0200), .Y(new_n30914_));
  OR2X1    g28478(.A(new_n30914_), .B(pi0199), .Y(new_n30915_));
  INVX1    g28479(.A(pi1055), .Y(new_n30916_));
  AOI21X1  g28480(.A0(new_n30916_), .A1(pi0199), .B0(new_n30470_), .Y(new_n30917_));
  AND2X1   g28481(.A(new_n30472_), .B(new_n30470_), .Y(new_n30918_));
  AND2X1   g28482(.A(pi0588), .B(pi0420), .Y(new_n30919_));
  AOI22X1  g28483(.A0(new_n30919_), .A1(new_n30918_), .B0(new_n30917_), .B1(new_n30915_), .Y(new_n30920_));
  OAI21X1  g28484(.A0(new_n30913_), .A1(new_n30911_), .B0(new_n30920_), .Y(new_n30921_));
  AND2X1   g28485(.A(new_n30483_), .B(pi1136), .Y(new_n30922_));
  INVX1    g28486(.A(new_n30922_), .Y(new_n30923_));
  AOI21X1  g28487(.A0(new_n28313_), .A1(new_n12614_), .B0(pi1134), .Y(new_n30924_));
  OAI21X1  g28488(.A0(new_n28313_), .A1(pi0627), .B0(new_n30924_), .Y(new_n30925_));
  AND2X1   g28489(.A(new_n30484_), .B(pi0753), .Y(new_n30926_));
  OAI22X1  g28490(.A0(pi1136), .A1(pi0847), .B0(new_n28313_), .B1(new_n15160_), .Y(new_n30927_));
  OR2X1    g28491(.A(new_n30927_), .B(new_n30487_), .Y(new_n30928_));
  OAI22X1  g28492(.A0(new_n30928_), .A1(new_n30926_), .B0(new_n30925_), .B1(new_n30923_), .Y(new_n30929_));
  MX2X1    g28493(.A(new_n30929_), .B(new_n30921_), .S0(new_n6748_), .Y(po0864));
  NAND4X1  g28494(.A(new_n30470_), .B(pi0592), .C(new_n6074_), .D(pi0442), .Y(new_n30931_));
  NAND4X1  g28495(.A(new_n30470_), .B(new_n6120_), .C(pi0591), .D(pi0328), .Y(new_n30932_));
  AOI21X1  g28496(.A0(new_n30932_), .A1(new_n30931_), .B0(pi0590), .Y(new_n30933_));
  NOR3X1   g28497(.A(new_n30492_), .B(new_n30471_), .C(new_n6008_), .Y(new_n30934_));
  OAI21X1  g28498(.A0(new_n30934_), .A1(new_n30933_), .B0(new_n9028_), .Y(new_n30935_));
  INVX1    g28499(.A(pi0305), .Y(new_n30936_));
  MX2X1    g28500(.A(new_n30502_), .B(new_n30936_), .S0(new_n8009_), .Y(new_n30937_));
  OAI22X1  g28501(.A0(pi1058), .A1(new_n7941_), .B0(pi0224), .B1(pi0223), .Y(new_n30938_));
  AOI21X1  g28502(.A0(new_n30937_), .A1(new_n7941_), .B0(new_n30938_), .Y(new_n30939_));
  INVX1    g28503(.A(pi0459), .Y(new_n30940_));
  OR4X1    g28504(.A(pi0592), .B(pi0591), .C(pi0224), .D(pi0223), .Y(new_n30941_));
  NOR4X1   g28505(.A(new_n30941_), .B(pi0590), .C(new_n9028_), .D(new_n30940_), .Y(new_n30942_));
  NOR3X1   g28506(.A(new_n30942_), .B(new_n30939_), .C(new_n10265_), .Y(new_n30943_));
  NAND2X1  g28507(.A(new_n30484_), .B(pi0754), .Y(new_n30944_));
  AOI21X1  g28508(.A0(new_n28946_), .A1(pi1135), .B0(new_n30595_), .Y(new_n30945_));
  OAI21X1  g28509(.A0(pi1136), .A1(pi0857), .B0(pi1134), .Y(new_n30946_));
  AOI21X1  g28510(.A0(pi1135), .A1(pi0709), .B0(new_n30946_), .Y(new_n30947_));
  NAND3X1  g28511(.A(new_n30947_), .B(new_n30945_), .C(new_n30944_), .Y(new_n30948_));
  OAI21X1  g28512(.A0(new_n28313_), .A1(pi0660), .B0(new_n4755_), .Y(new_n30949_));
  AOI21X1  g28513(.A0(new_n28313_), .A1(new_n12590_), .B0(new_n30949_), .Y(new_n30950_));
  AOI21X1  g28514(.A0(new_n30950_), .A1(new_n30922_), .B0(new_n6748_), .Y(new_n30951_));
  AOI22X1  g28515(.A0(new_n30951_), .A1(new_n30948_), .B0(new_n30943_), .B1(new_n30935_), .Y(po0865));
  INVX1    g28516(.A(pi1118), .Y(new_n30953_));
  OAI21X1  g28517(.A0(po0980), .A1(new_n15191_), .B0(new_n30348_), .Y(new_n30954_));
  AOI21X1  g28518(.A0(po0980), .A1(new_n30953_), .B0(new_n30954_), .Y(po0866));
  OAI21X1  g28519(.A0(new_n30347_), .A1(pi1106), .B0(new_n30348_), .Y(new_n30956_));
  AOI21X1  g28520(.A0(new_n30347_), .A1(new_n22840_), .B0(new_n30956_), .Y(po0867));
  NAND3X1  g28521(.A(new_n6120_), .B(pi0591), .C(pi0398), .Y(new_n30958_));
  OAI21X1  g28522(.A0(new_n30908_), .A1(new_n6079_), .B0(new_n30958_), .Y(new_n30959_));
  AOI22X1  g28523(.A0(new_n30959_), .A1(new_n6168_), .B0(new_n30467_), .B1(pi0348), .Y(new_n30960_));
  MX2X1    g28524(.A(pi0306), .B(pi1059), .S0(pi0200), .Y(new_n30961_));
  OR2X1    g28525(.A(new_n30961_), .B(pi0199), .Y(new_n30962_));
  INVX1    g28526(.A(pi1087), .Y(new_n30963_));
  AOI21X1  g28527(.A0(new_n30963_), .A1(pi0199), .B0(new_n30470_), .Y(new_n30964_));
  AND2X1   g28528(.A(pi0588), .B(pi0423), .Y(new_n30965_));
  AOI22X1  g28529(.A0(new_n30965_), .A1(new_n30918_), .B0(new_n30964_), .B1(new_n30962_), .Y(new_n30966_));
  OAI21X1  g28530(.A0(new_n30960_), .A1(new_n30913_), .B0(new_n30966_), .Y(new_n30967_));
  AOI21X1  g28531(.A0(new_n28313_), .A1(new_n12723_), .B0(pi1134), .Y(new_n30968_));
  OAI21X1  g28532(.A0(new_n28313_), .A1(pi0647), .B0(new_n30968_), .Y(new_n30969_));
  AND2X1   g28533(.A(new_n30484_), .B(pi0755), .Y(new_n30970_));
  OAI22X1  g28534(.A0(pi1136), .A1(pi0858), .B0(new_n28313_), .B1(new_n14788_), .Y(new_n30971_));
  OR2X1    g28535(.A(new_n30971_), .B(new_n30487_), .Y(new_n30972_));
  OAI22X1  g28536(.A0(new_n30972_), .A1(new_n30970_), .B0(new_n30969_), .B1(new_n30923_), .Y(new_n30973_));
  MX2X1    g28537(.A(new_n30973_), .B(new_n30967_), .S0(new_n6748_), .Y(po0868));
  NAND2X1  g28538(.A(new_n30484_), .B(pi0751), .Y(new_n30975_));
  OAI21X1  g28539(.A0(pi1136), .A1(pi0842), .B0(pi1134), .Y(new_n30976_));
  AOI21X1  g28540(.A0(pi1135), .A1(pi0701), .B0(new_n30976_), .Y(new_n30977_));
  AND2X1   g28541(.A(new_n30977_), .B(new_n30945_), .Y(new_n30978_));
  OAI21X1  g28542(.A0(pi1135), .A1(pi0644), .B0(new_n4755_), .Y(new_n30979_));
  AOI21X1  g28543(.A0(pi1135), .A1(new_n12739_), .B0(new_n30979_), .Y(new_n30980_));
  AOI22X1  g28544(.A0(new_n30980_), .A1(new_n30922_), .B0(new_n30978_), .B1(new_n30975_), .Y(new_n30981_));
  NOR3X1   g28545(.A(pi0592), .B(new_n6074_), .C(new_n6177_), .Y(new_n30982_));
  AOI21X1  g28546(.A0(new_n30464_), .A1(pi0374), .B0(new_n30982_), .Y(new_n30983_));
  OAI22X1  g28547(.A0(new_n30983_), .A1(pi0590), .B0(new_n30492_), .B1(new_n6019_), .Y(new_n30984_));
  NAND3X1  g28548(.A(new_n6168_), .B(pi0588), .C(pi0425), .Y(new_n30985_));
  OAI21X1  g28549(.A0(new_n30985_), .A1(new_n30807_), .B0(new_n30470_), .Y(new_n30986_));
  AOI21X1  g28550(.A0(new_n30984_), .A1(new_n9028_), .B0(new_n30986_), .Y(new_n30987_));
  AND2X1   g28551(.A(new_n8130_), .B(pi0298), .Y(new_n30988_));
  NAND3X1  g28552(.A(pi1044), .B(pi0200), .C(new_n7941_), .Y(new_n30989_));
  AOI21X1  g28553(.A0(pi1035), .A1(pi0199), .B0(new_n30470_), .Y(new_n30990_));
  NAND2X1  g28554(.A(new_n30990_), .B(new_n30989_), .Y(new_n30991_));
  OAI21X1  g28555(.A0(new_n30991_), .A1(new_n30988_), .B0(new_n6748_), .Y(new_n30992_));
  OAI22X1  g28556(.A0(new_n30992_), .A1(new_n30987_), .B0(new_n30981_), .B1(new_n6748_), .Y(po0869));
  NAND3X1  g28557(.A(new_n6120_), .B(pi0591), .C(pi0396), .Y(new_n30994_));
  OAI21X1  g28558(.A0(new_n30908_), .A1(new_n6080_), .B0(new_n30994_), .Y(new_n30995_));
  AOI22X1  g28559(.A0(new_n30995_), .A1(new_n6168_), .B0(new_n30467_), .B1(pi0322), .Y(new_n30996_));
  MX2X1    g28560(.A(pi0309), .B(pi1072), .S0(pi0200), .Y(new_n30997_));
  OR2X1    g28561(.A(new_n30997_), .B(pi0199), .Y(new_n30998_));
  INVX1    g28562(.A(pi1051), .Y(new_n30999_));
  AOI21X1  g28563(.A0(new_n30999_), .A1(pi0199), .B0(new_n30470_), .Y(new_n31000_));
  AND2X1   g28564(.A(pi0588), .B(pi0421), .Y(new_n31001_));
  AOI22X1  g28565(.A0(new_n31001_), .A1(new_n30918_), .B0(new_n31000_), .B1(new_n30998_), .Y(new_n31002_));
  OAI21X1  g28566(.A0(new_n30996_), .A1(new_n30913_), .B0(new_n31002_), .Y(new_n31003_));
  AOI21X1  g28567(.A0(new_n28313_), .A1(new_n12689_), .B0(pi1134), .Y(new_n31004_));
  OAI21X1  g28568(.A0(new_n28313_), .A1(pi0628), .B0(new_n31004_), .Y(new_n31005_));
  AND2X1   g28569(.A(new_n30484_), .B(pi0756), .Y(new_n31006_));
  OAI22X1  g28570(.A0(pi1136), .A1(pi0854), .B0(new_n28313_), .B1(new_n15209_), .Y(new_n31007_));
  OR2X1    g28571(.A(new_n31007_), .B(new_n30487_), .Y(new_n31008_));
  OAI22X1  g28572(.A0(new_n31008_), .A1(new_n31006_), .B0(new_n31005_), .B1(new_n30923_), .Y(new_n31009_));
  MX2X1    g28573(.A(new_n31009_), .B(new_n31003_), .S0(new_n6748_), .Y(po0870));
  INVX1    g28574(.A(new_n27697_), .Y(new_n31011_));
  AOI22X1  g28575(.A0(new_n30803_), .A1(pi0461), .B0(new_n30802_), .B1(pi0439), .Y(new_n31012_));
  NAND4X1  g28576(.A(new_n6120_), .B(pi0591), .C(new_n6168_), .D(pi0326), .Y(new_n31013_));
  OAI21X1  g28577(.A0(new_n31012_), .A1(pi0591), .B0(new_n31013_), .Y(new_n31014_));
  NOR4X1   g28578(.A(new_n30807_), .B(pi0590), .C(new_n9028_), .D(new_n6523_), .Y(new_n31015_));
  AOI21X1  g28579(.A0(new_n31014_), .A1(new_n9028_), .B0(new_n31015_), .Y(new_n31016_));
  OAI22X1  g28580(.A0(pi1057), .A1(new_n7941_), .B0(pi0224), .B1(pi0223), .Y(new_n31017_));
  OAI22X1  g28581(.A0(new_n31017_), .A1(new_n31011_), .B0(new_n31016_), .B1(new_n30471_), .Y(new_n31018_));
  NAND2X1  g28582(.A(new_n28313_), .B(pi0762), .Y(new_n31019_));
  AOI21X1  g28583(.A0(pi1135), .A1(pi0697), .B0(new_n28946_), .Y(new_n31020_));
  AOI22X1  g28584(.A0(new_n31020_), .A1(new_n31019_), .B0(new_n30513_), .B1(pi0867), .Y(new_n31021_));
  OR2X1    g28585(.A(pi1135), .B(pi0653), .Y(new_n31022_));
  AOI21X1  g28586(.A0(pi1135), .A1(pi0693), .B0(new_n28946_), .Y(new_n31023_));
  AND2X1   g28587(.A(new_n30483_), .B(pi0816), .Y(new_n31024_));
  AOI22X1  g28588(.A0(new_n31024_), .A1(new_n30513_), .B0(new_n31023_), .B1(new_n31022_), .Y(new_n31025_));
  OAI22X1  g28589(.A0(new_n31025_), .A1(new_n30815_), .B0(new_n31021_), .B1(new_n30678_), .Y(new_n31026_));
  MX2X1    g28590(.A(new_n31026_), .B(new_n31018_), .S0(new_n6748_), .Y(po0871));
  OAI21X1  g28591(.A0(new_n30347_), .A1(pi1123), .B0(new_n30348_), .Y(new_n31028_));
  AOI21X1  g28592(.A0(new_n30347_), .A1(new_n12739_), .B0(new_n31028_), .Y(po0872));
  NAND4X1  g28593(.A(new_n30470_), .B(pi0592), .C(new_n6074_), .D(pi0440), .Y(new_n31030_));
  NAND4X1  g28594(.A(new_n30470_), .B(new_n6120_), .C(pi0591), .D(pi0329), .Y(new_n31031_));
  AOI21X1  g28595(.A0(new_n31031_), .A1(new_n31030_), .B0(pi0590), .Y(new_n31032_));
  AND2X1   g28596(.A(new_n30470_), .B(pi0349), .Y(new_n31033_));
  AND2X1   g28597(.A(new_n31033_), .B(new_n30467_), .Y(new_n31034_));
  OAI21X1  g28598(.A0(new_n31034_), .A1(new_n31032_), .B0(new_n9028_), .Y(new_n31035_));
  INVX1    g28599(.A(pi0307), .Y(new_n31036_));
  MX2X1    g28600(.A(new_n27695_), .B(new_n31036_), .S0(new_n8009_), .Y(new_n31037_));
  OAI22X1  g28601(.A0(pi1043), .A1(new_n7941_), .B0(pi0224), .B1(pi0223), .Y(new_n31038_));
  AOI21X1  g28602(.A0(new_n31037_), .A1(new_n7941_), .B0(new_n31038_), .Y(new_n31039_));
  INVX1    g28603(.A(pi0454), .Y(new_n31040_));
  NOR4X1   g28604(.A(new_n30941_), .B(pi0590), .C(new_n9028_), .D(new_n31040_), .Y(new_n31041_));
  NOR3X1   g28605(.A(new_n31041_), .B(new_n31039_), .C(new_n10265_), .Y(new_n31042_));
  NAND2X1  g28606(.A(new_n30484_), .B(pi0761), .Y(new_n31043_));
  OAI21X1  g28607(.A0(pi1136), .A1(pi0845), .B0(pi1134), .Y(new_n31044_));
  AOI21X1  g28608(.A0(pi1135), .A1(pi0738), .B0(new_n31044_), .Y(new_n31045_));
  NAND3X1  g28609(.A(new_n31045_), .B(new_n31043_), .C(new_n30945_), .Y(new_n31046_));
  OAI21X1  g28610(.A0(new_n28313_), .A1(pi0641), .B0(new_n4755_), .Y(new_n31047_));
  AOI21X1  g28611(.A0(new_n28313_), .A1(new_n12664_), .B0(new_n31047_), .Y(new_n31048_));
  AOI21X1  g28612(.A0(new_n31048_), .A1(new_n30922_), .B0(new_n6748_), .Y(new_n31049_));
  AOI22X1  g28613(.A0(new_n31049_), .A1(new_n31046_), .B0(new_n31042_), .B1(new_n31035_), .Y(po0873));
  NAND2X1  g28614(.A(pi0591), .B(pi0318), .Y(new_n31051_));
  OAI22X1  g28615(.A0(new_n31051_), .A1(pi0592), .B0(new_n6108_), .B1(pi0591), .Y(new_n31052_));
  AOI22X1  g28616(.A0(new_n31052_), .A1(new_n6168_), .B0(new_n30467_), .B1(pi0462), .Y(new_n31053_));
  OR2X1    g28617(.A(new_n28045_), .B(pi0199), .Y(new_n31054_));
  INVX1    g28618(.A(pi1074), .Y(new_n31055_));
  AOI21X1  g28619(.A0(new_n31055_), .A1(pi0199), .B0(new_n30470_), .Y(new_n31056_));
  AND2X1   g28620(.A(pi0588), .B(pi0448), .Y(new_n31057_));
  AOI22X1  g28621(.A0(new_n31057_), .A1(new_n30918_), .B0(new_n31056_), .B1(new_n31054_), .Y(new_n31058_));
  OAI21X1  g28622(.A0(new_n31053_), .A1(new_n30913_), .B0(new_n31058_), .Y(new_n31059_));
  AND2X1   g28623(.A(new_n30484_), .B(pi0768), .Y(new_n31060_));
  OAI21X1  g28624(.A0(pi1136), .A1(pi0839), .B0(pi1134), .Y(new_n31061_));
  AOI21X1  g28625(.A0(pi1135), .A1(new_n15470_), .B0(new_n31061_), .Y(new_n31062_));
  NAND2X1  g28626(.A(new_n31062_), .B(new_n30945_), .Y(new_n31063_));
  OR2X1    g28627(.A(pi1135), .B(pi0645), .Y(new_n31064_));
  AOI21X1  g28628(.A0(pi1135), .A1(pi0669), .B0(new_n28946_), .Y(new_n31065_));
  AOI22X1  g28629(.A0(new_n31065_), .A1(new_n31064_), .B0(new_n30513_), .B1(pi0800), .Y(new_n31066_));
  OAI22X1  g28630(.A0(new_n31066_), .A1(new_n30477_), .B0(new_n31063_), .B1(new_n31060_), .Y(new_n31067_));
  MX2X1    g28631(.A(new_n31067_), .B(new_n31059_), .S0(new_n6748_), .Y(po0874));
  NAND4X1  g28632(.A(new_n30470_), .B(pi0592), .C(new_n6074_), .D(pi0369), .Y(new_n31069_));
  NAND4X1  g28633(.A(new_n30470_), .B(new_n6120_), .C(pi0591), .D(pi0394), .Y(new_n31070_));
  AOI21X1  g28634(.A0(new_n31070_), .A1(new_n31069_), .B0(pi0590), .Y(new_n31071_));
  NOR3X1   g28635(.A(new_n30492_), .B(new_n30471_), .C(new_n6012_), .Y(new_n31072_));
  OAI21X1  g28636(.A0(new_n31072_), .A1(new_n31071_), .B0(new_n9028_), .Y(new_n31073_));
  INVX1    g28637(.A(pi0303), .Y(new_n31074_));
  MX2X1    g28638(.A(new_n30568_), .B(new_n31074_), .S0(new_n8009_), .Y(new_n31075_));
  OAI22X1  g28639(.A0(pi1080), .A1(new_n7941_), .B0(pi0224), .B1(pi0223), .Y(new_n31076_));
  AOI21X1  g28640(.A0(new_n31075_), .A1(new_n7941_), .B0(new_n31076_), .Y(new_n31077_));
  INVX1    g28641(.A(pi0419), .Y(new_n31078_));
  NOR4X1   g28642(.A(new_n30941_), .B(pi0590), .C(new_n9028_), .D(new_n31078_), .Y(new_n31079_));
  NOR3X1   g28643(.A(new_n31079_), .B(new_n31077_), .C(new_n10265_), .Y(new_n31080_));
  NAND2X1  g28644(.A(new_n30484_), .B(pi0767), .Y(new_n31081_));
  OAI21X1  g28645(.A0(pi1136), .A1(pi0853), .B0(pi1134), .Y(new_n31082_));
  AOI21X1  g28646(.A0(pi1135), .A1(pi0698), .B0(new_n31082_), .Y(new_n31083_));
  NAND3X1  g28647(.A(new_n31083_), .B(new_n31081_), .C(new_n30945_), .Y(new_n31084_));
  OAI21X1  g28648(.A0(new_n28313_), .A1(pi0625), .B0(new_n4755_), .Y(new_n31085_));
  AOI21X1  g28649(.A0(new_n28313_), .A1(new_n12584_), .B0(new_n31085_), .Y(new_n31086_));
  AOI21X1  g28650(.A0(new_n31086_), .A1(new_n30922_), .B0(new_n6748_), .Y(new_n31087_));
  AOI22X1  g28651(.A0(new_n31087_), .A1(new_n31084_), .B0(new_n31080_), .B1(new_n31073_), .Y(po0875));
  NAND3X1  g28652(.A(new_n6120_), .B(pi0591), .C(pi0325), .Y(new_n31089_));
  OAI21X1  g28653(.A0(new_n30908_), .A1(new_n6113_), .B0(new_n31089_), .Y(new_n31090_));
  AOI22X1  g28654(.A0(new_n31090_), .A1(new_n6168_), .B0(new_n30467_), .B1(pi0353), .Y(new_n31091_));
  OR2X1    g28655(.A(new_n28049_), .B(pi0199), .Y(new_n31092_));
  INVX1    g28656(.A(pi1063), .Y(new_n31093_));
  AOI21X1  g28657(.A0(new_n31093_), .A1(pi0199), .B0(new_n30470_), .Y(new_n31094_));
  AND2X1   g28658(.A(pi0588), .B(pi0451), .Y(new_n31095_));
  AOI22X1  g28659(.A0(new_n31095_), .A1(new_n30918_), .B0(new_n31094_), .B1(new_n31092_), .Y(new_n31096_));
  OAI21X1  g28660(.A0(new_n31091_), .A1(new_n30913_), .B0(new_n31096_), .Y(new_n31097_));
  AND2X1   g28661(.A(new_n30484_), .B(pi0774), .Y(new_n31098_));
  OAI21X1  g28662(.A0(pi1136), .A1(pi0868), .B0(pi1134), .Y(new_n31099_));
  AOI21X1  g28663(.A0(pi1135), .A1(new_n13680_), .B0(new_n31099_), .Y(new_n31100_));
  NAND2X1  g28664(.A(new_n31100_), .B(new_n30945_), .Y(new_n31101_));
  OR2X1    g28665(.A(pi1135), .B(pi0636), .Y(new_n31102_));
  AOI21X1  g28666(.A0(pi1135), .A1(pi0650), .B0(new_n28946_), .Y(new_n31103_));
  AOI22X1  g28667(.A0(new_n31103_), .A1(new_n31102_), .B0(new_n30513_), .B1(pi0807), .Y(new_n31104_));
  OAI22X1  g28668(.A0(new_n31104_), .A1(new_n30477_), .B0(new_n31101_), .B1(new_n31098_), .Y(new_n31105_));
  MX2X1    g28669(.A(new_n31105_), .B(new_n31097_), .S0(new_n6748_), .Y(po0876));
  INVX1    g28670(.A(new_n28059_), .Y(new_n31107_));
  AOI22X1  g28671(.A0(new_n30803_), .A1(pi0356), .B0(new_n30802_), .B1(pi0381), .Y(new_n31108_));
  NAND4X1  g28672(.A(new_n6120_), .B(pi0591), .C(new_n6168_), .D(pi0405), .Y(new_n31109_));
  OAI21X1  g28673(.A0(new_n31108_), .A1(pi0591), .B0(new_n31109_), .Y(new_n31110_));
  NOR4X1   g28674(.A(new_n30807_), .B(pi0590), .C(new_n9028_), .D(new_n6589_), .Y(new_n31111_));
  AOI21X1  g28675(.A0(new_n31110_), .A1(new_n9028_), .B0(new_n31111_), .Y(new_n31112_));
  OAI22X1  g28676(.A0(pi1081), .A1(new_n7941_), .B0(pi0224), .B1(pi0223), .Y(new_n31113_));
  OAI22X1  g28677(.A0(new_n31113_), .A1(new_n31107_), .B0(new_n31112_), .B1(new_n30471_), .Y(new_n31114_));
  NAND2X1  g28678(.A(new_n28313_), .B(pi0750), .Y(new_n31115_));
  AOI21X1  g28679(.A0(pi1135), .A1(pi0684), .B0(new_n28946_), .Y(new_n31116_));
  AOI22X1  g28680(.A0(new_n31116_), .A1(new_n31115_), .B0(new_n30513_), .B1(pi0880), .Y(new_n31117_));
  OR2X1    g28681(.A(pi1135), .B(pi0651), .Y(new_n31118_));
  AOI21X1  g28682(.A0(pi1135), .A1(pi0654), .B0(new_n28946_), .Y(new_n31119_));
  AND2X1   g28683(.A(new_n30483_), .B(pi0794), .Y(new_n31120_));
  AOI22X1  g28684(.A0(new_n31120_), .A1(new_n30513_), .B0(new_n31119_), .B1(new_n31118_), .Y(new_n31121_));
  OAI22X1  g28685(.A0(new_n31121_), .A1(new_n30815_), .B0(new_n31117_), .B1(new_n30678_), .Y(new_n31122_));
  MX2X1    g28686(.A(new_n31122_), .B(new_n31114_), .S0(new_n6748_), .Y(po0877));
  INVX1    g28687(.A(pi0795), .Y(new_n31124_));
  INVX1    g28688(.A(pi0775), .Y(new_n31125_));
  INVX1    g28689(.A(pi0721), .Y(new_n31126_));
  INVX1    g28690(.A(pi0747), .Y(new_n31127_));
  INVX1    g28691(.A(pi0769), .Y(new_n31128_));
  INVX1    g28692(.A(pi0773), .Y(new_n31129_));
  NOR4X1   g28693(.A(new_n31129_), .B(new_n31128_), .C(new_n31127_), .D(new_n31126_), .Y(new_n31130_));
  AND2X1   g28694(.A(pi0773), .B(pi0747), .Y(new_n31131_));
  AOI21X1  g28695(.A0(new_n31131_), .A1(pi0769), .B0(pi0721), .Y(new_n31132_));
  NOR3X1   g28696(.A(new_n31132_), .B(new_n31130_), .C(new_n31125_), .Y(new_n31133_));
  INVX1    g28697(.A(pi0813), .Y(new_n31134_));
  XOR2X1   g28698(.A(pi0801), .B(pi0773), .Y(new_n31135_));
  XOR2X1   g28699(.A(pi0800), .B(pi0771), .Y(new_n31136_));
  XOR2X1   g28700(.A(pi0794), .B(pi0769), .Y(new_n31137_));
  INVX1    g28701(.A(pi0807), .Y(new_n31138_));
  XOR2X1   g28702(.A(pi0798), .B(pi0765), .Y(new_n31139_));
  NOR3X1   g28703(.A(new_n31139_), .B(new_n31138_), .C(new_n31127_), .Y(new_n31140_));
  OR2X1    g28704(.A(pi0807), .B(pi0747), .Y(new_n31141_));
  NOR2X1   g28705(.A(new_n31141_), .B(new_n31139_), .Y(new_n31142_));
  NOR2X1   g28706(.A(new_n31142_), .B(new_n31140_), .Y(new_n31143_));
  OR4X1    g28707(.A(new_n31143_), .B(new_n31137_), .C(new_n31136_), .D(new_n31135_), .Y(new_n31144_));
  NOR3X1   g28708(.A(new_n31144_), .B(new_n31134_), .C(new_n31126_), .Y(new_n31145_));
  NOR3X1   g28709(.A(new_n31139_), .B(new_n31136_), .C(new_n31138_), .Y(new_n31146_));
  INVX1    g28710(.A(pi0794), .Y(new_n31147_));
  NOR4X1   g28711(.A(pi0813), .B(new_n30866_), .C(new_n31147_), .D(pi0721), .Y(new_n31148_));
  AND2X1   g28712(.A(new_n31148_), .B(new_n31146_), .Y(new_n31149_));
  OAI21X1  g28713(.A0(new_n31149_), .A1(new_n31145_), .B0(pi0816), .Y(new_n31150_));
  AOI21X1  g28714(.A0(new_n31150_), .A1(new_n31133_), .B0(new_n31124_), .Y(new_n31151_));
  INVX1    g28715(.A(pi0945), .Y(new_n31152_));
  AND2X1   g28716(.A(pi0988), .B(new_n31152_), .Y(new_n31153_));
  AND2X1   g28717(.A(new_n31153_), .B(pi0731), .Y(new_n31154_));
  AND2X1   g28718(.A(new_n31125_), .B(pi0721), .Y(new_n31155_));
  OAI21X1  g28719(.A0(new_n31155_), .A1(new_n31133_), .B0(new_n31154_), .Y(new_n31156_));
  XOR2X1   g28720(.A(pi0816), .B(pi0775), .Y(new_n31157_));
  OR4X1    g28721(.A(new_n31157_), .B(new_n31144_), .C(new_n31134_), .D(new_n31126_), .Y(new_n31158_));
  XOR2X1   g28722(.A(pi0795), .B(pi0731), .Y(new_n31159_));
  OR2X1    g28723(.A(new_n31159_), .B(new_n31158_), .Y(new_n31160_));
  AOI21X1  g28724(.A0(new_n31153_), .A1(pi0731), .B0(new_n31126_), .Y(new_n31161_));
  AOI22X1  g28725(.A0(new_n31161_), .A1(new_n31160_), .B0(new_n31158_), .B1(new_n31155_), .Y(new_n31162_));
  OAI21X1  g28726(.A0(new_n31156_), .A1(new_n31151_), .B0(new_n31162_), .Y(po0878));
  INVX1    g28727(.A(new_n30516_), .Y(new_n31164_));
  AND2X1   g28728(.A(pi0591), .B(pi0403), .Y(new_n31165_));
  AOI22X1  g28729(.A0(new_n31165_), .A1(new_n6120_), .B0(new_n30464_), .B1(pi0379), .Y(new_n31166_));
  OAI22X1  g28730(.A0(new_n31166_), .A1(pi0590), .B0(new_n30492_), .B1(new_n9116_), .Y(new_n31167_));
  NOR2X1   g28731(.A(new_n28051_), .B(pi0199), .Y(new_n31168_));
  OAI22X1  g28732(.A0(pi1045), .A1(new_n7941_), .B0(pi0224), .B1(pi0223), .Y(new_n31169_));
  NAND4X1  g28733(.A(new_n30472_), .B(new_n30470_), .C(pi0588), .D(pi0428), .Y(new_n31170_));
  OAI21X1  g28734(.A0(new_n31169_), .A1(new_n31168_), .B0(new_n31170_), .Y(new_n31171_));
  AOI21X1  g28735(.A0(new_n31167_), .A1(new_n30912_), .B0(new_n31171_), .Y(new_n31172_));
  NOR2X1   g28736(.A(pi1134), .B(pi0795), .Y(new_n31173_));
  OAI21X1  g28737(.A0(new_n4755_), .A1(pi0851), .B0(new_n28946_), .Y(new_n31174_));
  NOR2X1   g28738(.A(pi1134), .B(pi0640), .Y(new_n31175_));
  AND2X1   g28739(.A(pi1134), .B(pi0776), .Y(new_n31176_));
  OR2X1    g28740(.A(new_n31176_), .B(new_n28946_), .Y(new_n31177_));
  OAI22X1  g28741(.A0(new_n31177_), .A1(new_n31175_), .B0(new_n31174_), .B1(new_n31173_), .Y(new_n31178_));
  INVX1    g28742(.A(pi0732), .Y(new_n31179_));
  AND2X1   g28743(.A(pi1136), .B(pi1135), .Y(new_n31180_));
  OAI21X1  g28744(.A0(pi1134), .A1(new_n31179_), .B0(new_n31180_), .Y(new_n31181_));
  AOI21X1  g28745(.A0(pi1134), .A1(pi0694), .B0(new_n31181_), .Y(new_n31182_));
  AOI21X1  g28746(.A0(new_n31178_), .A1(new_n28313_), .B0(new_n31182_), .Y(new_n31183_));
  OAI22X1  g28747(.A0(new_n31183_), .A1(new_n31164_), .B0(new_n31172_), .B1(new_n10265_), .Y(po0879));
  OAI21X1  g28748(.A0(po0980), .A1(new_n14886_), .B0(new_n30348_), .Y(new_n31185_));
  AOI21X1  g28749(.A0(po0980), .A1(new_n30879_), .B0(new_n31185_), .Y(po0880));
  OAI21X1  g28750(.A0(po0980), .A1(new_n15092_), .B0(new_n30348_), .Y(new_n31187_));
  AOI21X1  g28751(.A0(po0980), .A1(new_n30400_), .B0(new_n31187_), .Y(po0881));
  INVX1    g28752(.A(pi1120), .Y(new_n31189_));
  OAI21X1  g28753(.A0(po0980), .A1(new_n14788_), .B0(new_n30348_), .Y(new_n31190_));
  AOI21X1  g28754(.A0(po0980), .A1(new_n31189_), .B0(new_n31190_), .Y(po0882));
  OAI21X1  g28755(.A0(new_n30824_), .A1(pi1126), .B0(new_n30348_), .Y(new_n31192_));
  AOI21X1  g28756(.A0(new_n30824_), .A1(new_n14637_), .B0(new_n31192_), .Y(po0883));
  OAI21X1  g28757(.A0(new_n30824_), .A1(pi1102), .B0(new_n30348_), .Y(new_n31194_));
  AOI21X1  g28758(.A0(new_n30824_), .A1(new_n15428_), .B0(new_n31194_), .Y(po0884));
  INVX1    g28759(.A(pi0728), .Y(new_n31196_));
  OAI21X1  g28760(.A0(po0980), .A1(new_n31196_), .B0(new_n30348_), .Y(new_n31197_));
  AOI21X1  g28761(.A0(po0980), .A1(new_n30436_), .B0(new_n31197_), .Y(po0885));
  OAI21X1  g28762(.A0(new_n30824_), .A1(pi1104), .B0(new_n30348_), .Y(new_n31199_));
  AOI21X1  g28763(.A0(new_n30824_), .A1(new_n15585_), .B0(new_n31199_), .Y(po0886));
  OAI21X1  g28764(.A0(new_n30824_), .A1(pi1106), .B0(new_n30348_), .Y(new_n31201_));
  AOI21X1  g28765(.A0(new_n30824_), .A1(new_n21514_), .B0(new_n31201_), .Y(po0887));
  INVX1    g28766(.A(new_n31131_), .Y(new_n31203_));
  XOR2X1   g28767(.A(pi0813), .B(pi0721), .Y(new_n31204_));
  OR4X1    g28768(.A(new_n31204_), .B(new_n31157_), .C(new_n31144_), .D(new_n31124_), .Y(new_n31205_));
  NAND2X1  g28769(.A(new_n31205_), .B(new_n31203_), .Y(new_n31206_));
  AND2X1   g28770(.A(new_n31205_), .B(pi0731), .Y(new_n31207_));
  INVX1    g28771(.A(new_n31207_), .Y(new_n31208_));
  OR2X1    g28772(.A(new_n31204_), .B(new_n31157_), .Y(new_n31209_));
  NOR4X1   g28773(.A(new_n31209_), .B(new_n31137_), .C(new_n30866_), .D(pi0795), .Y(new_n31210_));
  AOI21X1  g28774(.A0(new_n31210_), .A1(new_n31146_), .B0(new_n31203_), .Y(new_n31211_));
  OAI21X1  g28775(.A0(new_n31211_), .A1(pi0731), .B0(new_n31153_), .Y(new_n31212_));
  AOI22X1  g28776(.A0(new_n31212_), .A1(new_n31208_), .B0(new_n31206_), .B1(new_n31154_), .Y(po0888));
  OAI21X1  g28777(.A0(po0954), .A1(new_n31179_), .B0(new_n30348_), .Y(new_n31214_));
  AOI21X1  g28778(.A0(po0954), .A1(new_n30875_), .B0(new_n31214_), .Y(po0889));
  NAND4X1  g28779(.A(new_n30470_), .B(pi0592), .C(new_n6074_), .D(pi0375), .Y(new_n31216_));
  NAND4X1  g28780(.A(new_n30470_), .B(new_n6120_), .C(pi0591), .D(pi0399), .Y(new_n31217_));
  AOI21X1  g28781(.A0(new_n31217_), .A1(new_n31216_), .B0(pi0590), .Y(new_n31218_));
  AND2X1   g28782(.A(new_n30470_), .B(pi0316), .Y(new_n31219_));
  AND2X1   g28783(.A(new_n31219_), .B(new_n30467_), .Y(new_n31220_));
  OAI21X1  g28784(.A0(new_n31220_), .A1(new_n31218_), .B0(new_n9028_), .Y(new_n31221_));
  INVX1    g28785(.A(pi0308), .Y(new_n31222_));
  MX2X1    g28786(.A(new_n28057_), .B(new_n31222_), .S0(new_n8009_), .Y(new_n31223_));
  OAI22X1  g28787(.A0(pi1047), .A1(new_n7941_), .B0(pi0224), .B1(pi0223), .Y(new_n31224_));
  AOI21X1  g28788(.A0(new_n31223_), .A1(new_n7941_), .B0(new_n31224_), .Y(new_n31225_));
  INVX1    g28789(.A(pi0424), .Y(new_n31226_));
  NOR4X1   g28790(.A(new_n30941_), .B(pi0590), .C(new_n9028_), .D(new_n31226_), .Y(new_n31227_));
  NOR3X1   g28791(.A(new_n31227_), .B(new_n31225_), .C(new_n10265_), .Y(new_n31228_));
  NAND2X1  g28792(.A(new_n30484_), .B(pi0777), .Y(new_n31229_));
  OAI21X1  g28793(.A0(pi1136), .A1(pi0838), .B0(pi1134), .Y(new_n31230_));
  AOI21X1  g28794(.A0(pi1135), .A1(pi0737), .B0(new_n31230_), .Y(new_n31231_));
  NAND3X1  g28795(.A(new_n31231_), .B(new_n31229_), .C(new_n30945_), .Y(new_n31232_));
  OAI21X1  g28796(.A0(new_n28313_), .A1(pi0648), .B0(new_n4755_), .Y(new_n31233_));
  AOI21X1  g28797(.A0(new_n28313_), .A1(new_n12637_), .B0(new_n31233_), .Y(new_n31234_));
  AOI21X1  g28798(.A0(new_n31234_), .A1(new_n30922_), .B0(new_n6748_), .Y(new_n31235_));
  AOI22X1  g28799(.A0(new_n31235_), .A1(new_n31232_), .B0(new_n31228_), .B1(new_n31221_), .Y(po0890));
  INVX1    g28800(.A(pi1119), .Y(new_n31237_));
  OAI21X1  g28801(.A0(po0980), .A1(new_n15209_), .B0(new_n30348_), .Y(new_n31238_));
  AOI21X1  g28802(.A0(po0980), .A1(new_n31237_), .B0(new_n31238_), .Y(po0891));
  OAI21X1  g28803(.A0(new_n30824_), .A1(pi1109), .B0(new_n30348_), .Y(new_n31240_));
  AOI21X1  g28804(.A0(new_n30824_), .A1(new_n13294_), .B0(new_n31240_), .Y(po0892));
  OAI21X1  g28805(.A0(new_n30824_), .A1(pi1101), .B0(new_n30348_), .Y(new_n31242_));
  AOI21X1  g28806(.A0(new_n30824_), .A1(new_n13969_), .B0(new_n31242_), .Y(po0893));
  INVX1    g28807(.A(pi1122), .Y(new_n31244_));
  OAI21X1  g28808(.A0(po0980), .A1(new_n15335_), .B0(new_n30348_), .Y(new_n31245_));
  AOI21X1  g28809(.A0(po0980), .A1(new_n31244_), .B0(new_n31245_), .Y(po0894));
  INVX1    g28810(.A(pi1121), .Y(new_n31247_));
  OAI21X1  g28811(.A0(po0980), .A1(new_n12565_), .B0(new_n30348_), .Y(new_n31248_));
  AOI21X1  g28812(.A0(po0980), .A1(new_n31247_), .B0(new_n31248_), .Y(po0895));
  AND2X1   g28813(.A(new_n30279_), .B(pi1060), .Y(new_n31250_));
  INVX1    g28814(.A(new_n31250_), .Y(new_n31251_));
  NOR4X1   g28815(.A(new_n31251_), .B(pi1061), .C(pi0952), .D(new_n12898_), .Y(po0988));
  AND2X1   g28816(.A(po0988), .B(pi1108), .Y(new_n31253_));
  OAI21X1  g28817(.A0(po0988), .A1(new_n15697_), .B0(new_n30283_), .Y(new_n31254_));
  OR2X1    g28818(.A(new_n31254_), .B(new_n31253_), .Y(po0896));
  AOI21X1  g28819(.A0(po0988), .A1(pi1114), .B0(pi0966), .Y(new_n31256_));
  OAI21X1  g28820(.A0(po0988), .A1(pi0741), .B0(new_n31256_), .Y(po0898));
  AOI21X1  g28821(.A0(po0988), .A1(pi1112), .B0(pi0966), .Y(new_n31258_));
  OAI21X1  g28822(.A0(po0988), .A1(pi0742), .B0(new_n31258_), .Y(po0899));
  AND2X1   g28823(.A(po0988), .B(pi1109), .Y(new_n31260_));
  OAI21X1  g28824(.A0(po0988), .A1(new_n13220_), .B0(new_n30283_), .Y(new_n31261_));
  OR2X1    g28825(.A(new_n31261_), .B(new_n31260_), .Y(po0900));
  AOI21X1  g28826(.A0(po0988), .A1(pi1131), .B0(pi0966), .Y(new_n31263_));
  OAI21X1  g28827(.A0(po0988), .A1(pi0744), .B0(new_n31263_), .Y(po0901));
  AOI21X1  g28828(.A0(po0988), .A1(pi1111), .B0(pi0966), .Y(new_n31265_));
  OAI21X1  g28829(.A0(po0988), .A1(pi0745), .B0(new_n31265_), .Y(po0902));
  AND2X1   g28830(.A(po0988), .B(pi1104), .Y(new_n31267_));
  OAI21X1  g28831(.A0(po0988), .A1(new_n15545_), .B0(new_n30283_), .Y(new_n31268_));
  OR2X1    g28832(.A(new_n31268_), .B(new_n31267_), .Y(po0903));
  NOR3X1   g28833(.A(new_n31141_), .B(new_n31139_), .C(new_n30866_), .Y(new_n31270_));
  AND2X1   g28834(.A(new_n31153_), .B(pi0773), .Y(new_n31271_));
  NOR4X1   g28835(.A(new_n31271_), .B(new_n31139_), .C(new_n31135_), .D(new_n31138_), .Y(new_n31272_));
  NOR4X1   g28836(.A(new_n31209_), .B(new_n31159_), .C(new_n31137_), .D(new_n31136_), .Y(new_n31273_));
  OAI21X1  g28837(.A0(new_n31272_), .A1(new_n31270_), .B0(new_n31273_), .Y(new_n31274_));
  AOI21X1  g28838(.A0(new_n31153_), .A1(pi0773), .B0(pi0747), .Y(new_n31275_));
  AOI21X1  g28839(.A0(new_n31153_), .A1(new_n31131_), .B0(new_n31275_), .Y(new_n31276_));
  AND2X1   g28840(.A(new_n31276_), .B(new_n31274_), .Y(po0904));
  AND2X1   g28841(.A(po0988), .B(pi1106), .Y(new_n31278_));
  OAI21X1  g28842(.A0(po0988), .A1(new_n15595_), .B0(new_n30283_), .Y(new_n31279_));
  OR2X1    g28843(.A(new_n31279_), .B(new_n31278_), .Y(po0905));
  AND2X1   g28844(.A(po0988), .B(pi1105), .Y(new_n31281_));
  OAI21X1  g28845(.A0(po0988), .A1(new_n12911_), .B0(new_n30283_), .Y(new_n31282_));
  OR2X1    g28846(.A(new_n31282_), .B(new_n31281_), .Y(po0906));
  AOI21X1  g28847(.A0(po0988), .A1(pi1130), .B0(pi0966), .Y(new_n31284_));
  OAI21X1  g28848(.A0(po0988), .A1(pi0750), .B0(new_n31284_), .Y(po0907));
  AOI21X1  g28849(.A0(po0988), .A1(pi1123), .B0(pi0966), .Y(new_n31286_));
  OAI21X1  g28850(.A0(po0988), .A1(pi0751), .B0(new_n31286_), .Y(po0908));
  AOI21X1  g28851(.A0(po0988), .A1(pi1124), .B0(pi0966), .Y(new_n31288_));
  OAI21X1  g28852(.A0(po0988), .A1(pi0752), .B0(new_n31288_), .Y(po0909));
  AOI21X1  g28853(.A0(po0988), .A1(pi1117), .B0(pi0966), .Y(new_n31290_));
  OAI21X1  g28854(.A0(po0988), .A1(pi0753), .B0(new_n31290_), .Y(po0910));
  AOI21X1  g28855(.A0(po0988), .A1(pi1118), .B0(pi0966), .Y(new_n31292_));
  OAI21X1  g28856(.A0(po0988), .A1(pi0754), .B0(new_n31292_), .Y(po0911));
  AOI21X1  g28857(.A0(po0988), .A1(pi1120), .B0(pi0966), .Y(new_n31294_));
  OAI21X1  g28858(.A0(po0988), .A1(pi0755), .B0(new_n31294_), .Y(po0912));
  AOI21X1  g28859(.A0(po0988), .A1(pi1119), .B0(pi0966), .Y(new_n31296_));
  OAI21X1  g28860(.A0(po0988), .A1(pi0756), .B0(new_n31296_), .Y(po0913));
  AOI21X1  g28861(.A0(po0988), .A1(pi1113), .B0(pi0966), .Y(new_n31298_));
  OAI21X1  g28862(.A0(po0988), .A1(pi0757), .B0(new_n31298_), .Y(po0914));
  AND2X1   g28863(.A(po0988), .B(pi1101), .Y(new_n31300_));
  OAI21X1  g28864(.A0(po0988), .A1(new_n13973_), .B0(new_n30283_), .Y(new_n31301_));
  OR2X1    g28865(.A(new_n31301_), .B(new_n31300_), .Y(po0915));
  NOR2X1   g28866(.A(po0988), .B(pi0759), .Y(new_n31303_));
  NOR4X1   g28867(.A(new_n30284_), .B(new_n31251_), .C(pi1061), .D(pi0952), .Y(new_n31304_));
  OAI21X1  g28868(.A0(new_n31304_), .A1(new_n31303_), .B0(new_n30283_), .Y(po0916));
  AOI21X1  g28869(.A0(po0988), .A1(pi1115), .B0(pi0966), .Y(new_n31306_));
  OAI21X1  g28870(.A0(po0988), .A1(pi0760), .B0(new_n31306_), .Y(po0917));
  AOI21X1  g28871(.A0(po0988), .A1(pi1121), .B0(pi0966), .Y(new_n31308_));
  OAI21X1  g28872(.A0(po0988), .A1(pi0761), .B0(new_n31308_), .Y(po0918));
  AOI21X1  g28873(.A0(po0988), .A1(pi1129), .B0(pi0966), .Y(new_n31310_));
  OAI21X1  g28874(.A0(po0988), .A1(pi0762), .B0(new_n31310_), .Y(po0919));
  INVX1    g28875(.A(pi1103), .Y(new_n31312_));
  INVX1    g28876(.A(po0988), .Y(new_n31313_));
  AOI21X1  g28877(.A0(new_n31313_), .A1(pi0763), .B0(pi0966), .Y(new_n31314_));
  OAI21X1  g28878(.A0(new_n31313_), .A1(new_n31312_), .B0(new_n31314_), .Y(po0920));
  INVX1    g28879(.A(pi1107), .Y(new_n31316_));
  AOI21X1  g28880(.A0(new_n31313_), .A1(pi0764), .B0(pi0966), .Y(new_n31317_));
  OAI21X1  g28881(.A0(new_n31313_), .A1(new_n31316_), .B0(new_n31317_), .Y(po0921));
  NOR3X1   g28882(.A(new_n31204_), .B(new_n31159_), .C(new_n31157_), .Y(new_n31319_));
  INVX1    g28883(.A(new_n31319_), .Y(new_n31320_));
  NOR2X1   g28884(.A(new_n31320_), .B(new_n31144_), .Y(po0978));
  INVX1    g28885(.A(po0978), .Y(new_n31322_));
  AOI21X1  g28886(.A0(new_n31322_), .A1(pi0765), .B0(new_n31152_), .Y(new_n31323_));
  INVX1    g28887(.A(pi0765), .Y(new_n31324_));
  AOI21X1  g28888(.A0(new_n31134_), .A1(new_n31126_), .B0(new_n31145_), .Y(new_n31325_));
  OR2X1    g28889(.A(pi0816), .B(pi0775), .Y(new_n31326_));
  AND2X1   g28890(.A(pi0801), .B(pi0773), .Y(new_n31327_));
  NOR3X1   g28891(.A(new_n31143_), .B(new_n31137_), .C(new_n31136_), .Y(new_n31328_));
  AOI21X1  g28892(.A0(pi0800), .A1(pi0771), .B0(pi0765), .Y(new_n31329_));
  OAI21X1  g28893(.A0(new_n31147_), .A1(new_n31128_), .B0(new_n31329_), .Y(new_n31330_));
  NOR2X1   g28894(.A(new_n31330_), .B(new_n31140_), .Y(new_n31331_));
  NOR3X1   g28895(.A(new_n31331_), .B(pi0801), .C(pi0773), .Y(new_n31332_));
  OAI21X1  g28896(.A0(new_n31332_), .A1(new_n31327_), .B0(new_n31328_), .Y(new_n31333_));
  AOI21X1  g28897(.A0(new_n31333_), .A1(new_n31126_), .B0(new_n31326_), .Y(new_n31334_));
  INVX1    g28898(.A(new_n31334_), .Y(new_n31335_));
  AND2X1   g28899(.A(pi0816), .B(pi0775), .Y(new_n31336_));
  NOR2X1   g28900(.A(new_n31204_), .B(new_n31144_), .Y(new_n31337_));
  AOI21X1  g28901(.A0(new_n31337_), .A1(new_n31336_), .B0(pi0765), .Y(new_n31338_));
  OAI21X1  g28902(.A0(new_n31335_), .A1(new_n31325_), .B0(new_n31338_), .Y(new_n31339_));
  AOI21X1  g28903(.A0(new_n31339_), .A1(new_n31124_), .B0(pi0731), .Y(new_n31340_));
  NOR3X1   g28904(.A(new_n31339_), .B(pi0795), .C(pi0731), .Y(new_n31341_));
  OAI22X1  g28905(.A0(new_n31341_), .A1(new_n31324_), .B0(new_n31340_), .B1(new_n31207_), .Y(new_n31342_));
  AOI21X1  g28906(.A0(new_n31342_), .A1(new_n31152_), .B0(new_n31323_), .Y(po0922));
  INVX1    g28907(.A(pi1110), .Y(new_n31344_));
  AOI21X1  g28908(.A0(new_n31313_), .A1(pi0766), .B0(pi0966), .Y(new_n31345_));
  OAI21X1  g28909(.A0(new_n31313_), .A1(new_n31344_), .B0(new_n31345_), .Y(po0923));
  AOI21X1  g28910(.A0(po0988), .A1(pi1116), .B0(pi0966), .Y(new_n31347_));
  OAI21X1  g28911(.A0(po0988), .A1(pi0767), .B0(new_n31347_), .Y(po0924));
  AOI21X1  g28912(.A0(po0988), .A1(pi1125), .B0(pi0966), .Y(new_n31349_));
  OAI21X1  g28913(.A0(po0988), .A1(pi0768), .B0(new_n31349_), .Y(po0925));
  INVX1    g28914(.A(new_n31336_), .Y(new_n31351_));
  NOR3X1   g28915(.A(new_n31204_), .B(new_n31351_), .C(new_n31144_), .Y(new_n31352_));
  OR4X1    g28916(.A(new_n31209_), .B(new_n31136_), .C(new_n31135_), .D(new_n31147_), .Y(new_n31353_));
  NOR3X1   g28917(.A(new_n31353_), .B(new_n31143_), .C(pi0775), .Y(new_n31354_));
  OAI21X1  g28918(.A0(new_n31354_), .A1(new_n31352_), .B0(pi0795), .Y(new_n31355_));
  NAND3X1  g28919(.A(pi0775), .B(pi0773), .C(pi0747), .Y(new_n31356_));
  XOR2X1   g28920(.A(new_n31356_), .B(new_n31128_), .Y(new_n31357_));
  NAND3X1  g28921(.A(new_n31357_), .B(new_n31355_), .C(new_n31154_), .Y(new_n31358_));
  NOR3X1   g28922(.A(new_n31353_), .B(new_n31159_), .C(new_n31143_), .Y(new_n31359_));
  OR2X1    g28923(.A(new_n31154_), .B(new_n31128_), .Y(new_n31360_));
  OAI21X1  g28924(.A0(new_n31360_), .A1(new_n31359_), .B0(new_n31358_), .Y(po0926));
  AOI21X1  g28925(.A0(po0988), .A1(pi1126), .B0(pi0966), .Y(new_n31362_));
  OAI21X1  g28926(.A0(po0988), .A1(pi0770), .B0(new_n31362_), .Y(po0927));
  INVX1    g28927(.A(new_n31337_), .Y(new_n31364_));
  NOR2X1   g28928(.A(pi0795), .B(pi0731), .Y(new_n31365_));
  OAI21X1  g28929(.A0(new_n31334_), .A1(new_n31336_), .B0(new_n31365_), .Y(new_n31366_));
  NAND2X1  g28930(.A(pi0795), .B(pi0731), .Y(new_n31367_));
  NOR2X1   g28931(.A(new_n31367_), .B(new_n31157_), .Y(new_n31368_));
  INVX1    g28932(.A(new_n31368_), .Y(new_n31369_));
  AOI21X1  g28933(.A0(new_n31369_), .A1(new_n31366_), .B0(new_n31364_), .Y(po0963));
  NAND2X1  g28934(.A(pi0987), .B(new_n31152_), .Y(new_n31371_));
  NAND3X1  g28935(.A(new_n31322_), .B(pi0945), .C(pi0771), .Y(new_n31372_));
  OAI21X1  g28936(.A0(new_n31371_), .A1(po0963), .B0(new_n31372_), .Y(po0928));
  AND2X1   g28937(.A(po0988), .B(pi1102), .Y(new_n31374_));
  OAI21X1  g28938(.A0(po0988), .A1(new_n15465_), .B0(new_n30283_), .Y(new_n31375_));
  OR2X1    g28939(.A(new_n31375_), .B(new_n31374_), .Y(po0929));
  NAND3X1  g28940(.A(po0963), .B(new_n31328_), .C(new_n30866_), .Y(new_n31377_));
  NAND2X1  g28941(.A(new_n31377_), .B(new_n31153_), .Y(new_n31378_));
  NOR2X1   g28942(.A(new_n31319_), .B(new_n30866_), .Y(new_n31379_));
  OAI21X1  g28943(.A0(new_n31379_), .A1(new_n31144_), .B0(pi0773), .Y(new_n31380_));
  AOI21X1  g28944(.A0(new_n31380_), .A1(new_n31378_), .B0(new_n31271_), .Y(po0930));
  AOI21X1  g28945(.A0(po0988), .A1(pi1127), .B0(pi0966), .Y(new_n31382_));
  OAI21X1  g28946(.A0(po0988), .A1(pi0774), .B0(new_n31382_), .Y(po0931));
  AND2X1   g28947(.A(new_n31152_), .B(pi0731), .Y(new_n31384_));
  NAND4X1  g28948(.A(pi0773), .B(pi0771), .C(pi0765), .D(pi0747), .Y(new_n31385_));
  INVX1    g28949(.A(pi0800), .Y(new_n31386_));
  OR4X1    g28950(.A(pi0816), .B(new_n30866_), .C(new_n31386_), .D(new_n31124_), .Y(new_n31387_));
  NOR4X1   g28951(.A(new_n31387_), .B(new_n31204_), .C(new_n31143_), .D(new_n31137_), .Y(new_n31388_));
  OAI21X1  g28952(.A0(new_n31388_), .A1(new_n31385_), .B0(new_n31125_), .Y(new_n31389_));
  AOI22X1  g28953(.A0(new_n31389_), .A1(new_n31384_), .B0(new_n31322_), .B1(pi0775), .Y(new_n31390_));
  NAND3X1  g28954(.A(new_n31152_), .B(pi0775), .C(pi0731), .Y(new_n31391_));
  AOI21X1  g28955(.A0(new_n31385_), .A1(new_n31205_), .B0(new_n31391_), .Y(new_n31392_));
  NOR2X1   g28956(.A(new_n31392_), .B(new_n31390_), .Y(po0932));
  AOI21X1  g28957(.A0(po0988), .A1(pi1128), .B0(pi0966), .Y(new_n31394_));
  OAI21X1  g28958(.A0(po0988), .A1(pi0776), .B0(new_n31394_), .Y(po0933));
  AOI21X1  g28959(.A0(po0988), .A1(pi1122), .B0(pi0966), .Y(new_n31396_));
  OAI21X1  g28960(.A0(po0988), .A1(pi0777), .B0(new_n31396_), .Y(po0934));
  INVX1    g28961(.A(pi0968), .Y(new_n31398_));
  AND2X1   g28962(.A(pi0956), .B(pi0832), .Y(new_n31399_));
  NOR2X1   g28963(.A(pi1083), .B(pi1046), .Y(new_n31400_));
  NAND4X1  g28964(.A(new_n31400_), .B(new_n31399_), .C(pi1085), .D(new_n31398_), .Y(new_n31401_));
  MX2X1    g28965(.A(pi1100), .B(pi0778), .S0(new_n31401_), .Y(po0935));
  OR4X1    g28966(.A(new_n22606_), .B(pi0882), .C(pi0059), .D(pi0057), .Y(new_n31403_));
  OAI21X1  g28967(.A0(new_n31403_), .A1(new_n5297_), .B0(pi0779), .Y(po0936));
  OAI21X1  g28968(.A0(new_n31403_), .A1(new_n14590_), .B0(pi0780), .Y(po0937));
  MX2X1    g28969(.A(pi1101), .B(pi0781), .S0(new_n31401_), .Y(po0938));
  AOI22X1  g28970(.A0(new_n5244_), .A1(new_n5035_), .B0(pi0983), .B1(new_n2953_), .Y(new_n31407_));
  NAND2X1  g28971(.A(new_n31407_), .B(new_n31403_), .Y(po0939));
  MX2X1    g28972(.A(pi1109), .B(pi0783), .S0(new_n31401_), .Y(po0940));
  MX2X1    g28973(.A(pi1110), .B(pi0784), .S0(new_n31401_), .Y(po0941));
  MX2X1    g28974(.A(pi1102), .B(pi0785), .S0(new_n31401_), .Y(po0942));
  MX2X1    g28975(.A(new_n7704_), .B(new_n5787_), .S0(po1110), .Y(po0943));
  MX2X1    g28976(.A(pi1104), .B(pi0787), .S0(new_n31401_), .Y(po0944));
  MX2X1    g28977(.A(pi1105), .B(pi0788), .S0(new_n31401_), .Y(po0945));
  MX2X1    g28978(.A(pi1106), .B(pi0789), .S0(new_n31401_), .Y(po0946));
  MX2X1    g28979(.A(pi1107), .B(pi0790), .S0(new_n31401_), .Y(po0947));
  MX2X1    g28980(.A(pi1108), .B(pi0791), .S0(new_n31401_), .Y(po0948));
  MX2X1    g28981(.A(pi1103), .B(pi0792), .S0(new_n31401_), .Y(po0949));
  NAND4X1  g28982(.A(new_n31400_), .B(new_n31399_), .C(pi1085), .D(pi0968), .Y(new_n31419_));
  MX2X1    g28983(.A(pi1130), .B(pi0794), .S0(new_n31419_), .Y(po0951));
  MX2X1    g28984(.A(pi1128), .B(pi0795), .S0(new_n31419_), .Y(po0952));
  INVX1    g28985(.A(pi0281), .Y(new_n31422_));
  NAND2X1  g28986(.A(pi0279), .B(pi0278), .Y(new_n31423_));
  NOR4X1   g28987(.A(new_n31423_), .B(pi0280), .C(pi0269), .D(new_n4505_), .Y(new_n31424_));
  NAND2X1  g28988(.A(new_n31424_), .B(new_n31422_), .Y(new_n31425_));
  NOR2X1   g28989(.A(new_n31425_), .B(new_n30450_), .Y(new_n31426_));
  XOR2X1   g28990(.A(new_n31426_), .B(new_n30444_), .Y(po0953));
  MX2X1    g28991(.A(pi1124), .B(pi0798), .S0(new_n31419_), .Y(po0955));
  INVX1    g28992(.A(pi0799), .Y(new_n31429_));
  MX2X1    g28993(.A(pi1107), .B(new_n31429_), .S0(new_n31419_), .Y(po0956));
  MX2X1    g28994(.A(pi1125), .B(pi0800), .S0(new_n31419_), .Y(po0957));
  MX2X1    g28995(.A(pi1126), .B(pi0801), .S0(new_n31419_), .Y(po0958));
  AND2X1   g28996(.A(new_n30453_), .B(new_n3360_), .Y(po0959));
  INVX1    g28997(.A(pi0803), .Y(new_n31434_));
  MX2X1    g28998(.A(pi1106), .B(new_n31434_), .S0(new_n31419_), .Y(po0960));
  MX2X1    g28999(.A(pi1109), .B(pi0804), .S0(new_n31419_), .Y(po0961));
  NOR4X1   g29000(.A(new_n30448_), .B(pi0282), .C(pi0281), .D(pi0269), .Y(new_n31437_));
  XOR2X1   g29001(.A(new_n31437_), .B(new_n28613_), .Y(po0962));
  MX2X1    g29002(.A(pi1127), .B(pi0807), .S0(new_n31419_), .Y(po0964));
  MX2X1    g29003(.A(pi1101), .B(pi0808), .S0(new_n31419_), .Y(po0965));
  INVX1    g29004(.A(pi0809), .Y(new_n31441_));
  MX2X1    g29005(.A(pi1103), .B(new_n31441_), .S0(new_n31419_), .Y(po0966));
  MX2X1    g29006(.A(pi1108), .B(pi0810), .S0(new_n31419_), .Y(po0967));
  MX2X1    g29007(.A(pi1102), .B(pi0811), .S0(new_n31419_), .Y(po0968));
  INVX1    g29008(.A(pi0812), .Y(new_n31445_));
  MX2X1    g29009(.A(pi1104), .B(new_n31445_), .S0(new_n31419_), .Y(po0969));
  MX2X1    g29010(.A(pi1131), .B(pi0813), .S0(new_n31419_), .Y(po0970));
  INVX1    g29011(.A(pi0814), .Y(new_n31448_));
  MX2X1    g29012(.A(pi1105), .B(new_n31448_), .S0(new_n31419_), .Y(po0971));
  MX2X1    g29013(.A(pi1110), .B(pi0815), .S0(new_n31419_), .Y(po0972));
  MX2X1    g29014(.A(pi1129), .B(pi0816), .S0(new_n31419_), .Y(po0973));
  XOR2X1   g29015(.A(new_n30448_), .B(pi0269), .Y(po0974));
  OAI21X1  g29016(.A0(new_n10309_), .A1(new_n10265_), .B0(new_n10168_), .Y(po0975));
  XOR2X1   g29017(.A(new_n30452_), .B(new_n30443_), .Y(po0976));
  NAND2X1  g29018(.A(new_n31437_), .B(new_n28613_), .Y(new_n31455_));
  AOI21X1  g29019(.A0(new_n31455_), .A1(pi0277), .B0(new_n30451_), .Y(po0977));
  NOR2X1   g29020(.A(pi0893), .B(pi0811), .Y(po0979));
  OAI22X1  g29021(.A0(new_n7607_), .A1(pi0982), .B0(new_n10265_), .B1(new_n5983_), .Y(new_n31458_));
  AND2X1   g29022(.A(new_n31458_), .B(new_n2783_), .Y(po0981));
  INVX1    g29023(.A(pi0825), .Y(po1147));
  AND2X1   g29024(.A(new_n3008_), .B(pi0123), .Y(new_n31461_));
  AOI22X1  g29025(.A0(new_n3008_), .A1(pi0123), .B0(new_n30436_), .B1(new_n30412_), .Y(new_n31462_));
  AOI21X1  g29026(.A0(new_n31461_), .A1(po1147), .B0(new_n31462_), .Y(new_n31463_));
  NOR3X1   g29027(.A(new_n31461_), .B(new_n30436_), .C(new_n30412_), .Y(new_n31464_));
  OR2X1    g29028(.A(new_n31464_), .B(new_n31463_), .Y(new_n31465_));
  XOR2X1   g29029(.A(pi1130), .B(new_n30429_), .Y(new_n31466_));
  XOR2X1   g29030(.A(pi1129), .B(pi1128), .Y(new_n31467_));
  XOR2X1   g29031(.A(pi1126), .B(pi1125), .Y(new_n31468_));
  XOR2X1   g29032(.A(new_n31468_), .B(new_n31467_), .Y(new_n31469_));
  XOR2X1   g29033(.A(new_n31469_), .B(new_n31466_), .Y(new_n31470_));
  AOI21X1  g29034(.A0(new_n31461_), .A1(pi0825), .B0(new_n31462_), .Y(new_n31471_));
  NOR3X1   g29035(.A(new_n31471_), .B(new_n31470_), .C(new_n31464_), .Y(new_n31472_));
  AOI21X1  g29036(.A0(new_n31470_), .A1(new_n31465_), .B0(new_n31472_), .Y(po0982));
  INVX1    g29037(.A(pi0826), .Y(po1148));
  AOI22X1  g29038(.A0(new_n3008_), .A1(pi0123), .B0(new_n30894_), .B1(new_n31244_), .Y(new_n31475_));
  AOI21X1  g29039(.A0(new_n31461_), .A1(po1148), .B0(new_n31475_), .Y(new_n31476_));
  NOR3X1   g29040(.A(new_n31461_), .B(new_n30894_), .C(new_n31244_), .Y(new_n31477_));
  OR2X1    g29041(.A(new_n31477_), .B(new_n31476_), .Y(new_n31478_));
  XOR2X1   g29042(.A(pi1119), .B(new_n30953_), .Y(new_n31479_));
  XOR2X1   g29043(.A(pi1121), .B(pi1120), .Y(new_n31480_));
  XOR2X1   g29044(.A(pi1117), .B(pi1116), .Y(new_n31481_));
  XOR2X1   g29045(.A(new_n31481_), .B(new_n31480_), .Y(new_n31482_));
  XOR2X1   g29046(.A(new_n31482_), .B(new_n31479_), .Y(new_n31483_));
  AOI21X1  g29047(.A0(new_n31461_), .A1(pi0826), .B0(new_n31475_), .Y(new_n31484_));
  NOR3X1   g29048(.A(new_n31484_), .B(new_n31483_), .C(new_n31477_), .Y(new_n31485_));
  AOI21X1  g29049(.A0(new_n31483_), .A1(new_n31478_), .B0(new_n31485_), .Y(po0983));
  INVX1    g29050(.A(pi0827), .Y(po1178));
  INVX1    g29051(.A(pi1100), .Y(new_n31488_));
  AOI22X1  g29052(.A0(new_n3008_), .A1(pi0123), .B0(new_n31316_), .B1(new_n31488_), .Y(new_n31489_));
  AOI21X1  g29053(.A0(new_n31461_), .A1(po1178), .B0(new_n31489_), .Y(new_n31490_));
  NOR3X1   g29054(.A(new_n31461_), .B(new_n31316_), .C(new_n31488_), .Y(new_n31491_));
  OR2X1    g29055(.A(new_n31491_), .B(new_n31490_), .Y(new_n31492_));
  XOR2X1   g29056(.A(pi1105), .B(new_n31312_), .Y(new_n31493_));
  XOR2X1   g29057(.A(pi1102), .B(pi1101), .Y(new_n31494_));
  XOR2X1   g29058(.A(pi1106), .B(pi1104), .Y(new_n31495_));
  XOR2X1   g29059(.A(new_n31495_), .B(new_n31494_), .Y(new_n31496_));
  XOR2X1   g29060(.A(new_n31496_), .B(new_n31493_), .Y(new_n31497_));
  AOI21X1  g29061(.A0(new_n31461_), .A1(pi0827), .B0(new_n31489_), .Y(new_n31498_));
  NOR3X1   g29062(.A(new_n31498_), .B(new_n31497_), .C(new_n31491_), .Y(new_n31499_));
  AOI21X1  g29063(.A0(new_n31497_), .A1(new_n31492_), .B0(new_n31499_), .Y(po0984));
  INVX1    g29064(.A(pi0828), .Y(po1182));
  AOI22X1  g29065(.A0(new_n3008_), .A1(pi0123), .B0(new_n30365_), .B1(new_n30400_), .Y(new_n31502_));
  AOI21X1  g29066(.A0(new_n31461_), .A1(po1182), .B0(new_n31502_), .Y(new_n31503_));
  NOR3X1   g29067(.A(new_n31461_), .B(new_n30365_), .C(new_n30400_), .Y(new_n31504_));
  OR2X1    g29068(.A(new_n31504_), .B(new_n31503_), .Y(new_n31505_));
  XOR2X1   g29069(.A(pi1111), .B(new_n31344_), .Y(new_n31506_));
  XOR2X1   g29070(.A(pi1113), .B(pi1112), .Y(new_n31507_));
  XOR2X1   g29071(.A(pi1109), .B(pi1108), .Y(new_n31508_));
  XOR2X1   g29072(.A(new_n31508_), .B(new_n31507_), .Y(new_n31509_));
  XOR2X1   g29073(.A(new_n31509_), .B(new_n31506_), .Y(new_n31510_));
  AOI21X1  g29074(.A0(new_n31461_), .A1(pi0828), .B0(new_n31502_), .Y(new_n31511_));
  NOR3X1   g29075(.A(new_n31511_), .B(new_n31510_), .C(new_n31504_), .Y(new_n31512_));
  AOI21X1  g29076(.A0(new_n31510_), .A1(new_n31505_), .B0(new_n31512_), .Y(po0985));
  NAND2X1  g29077(.A(new_n6748_), .B(new_n2781_), .Y(new_n31514_));
  AOI21X1  g29078(.A0(new_n31514_), .A1(pi0951), .B0(new_n2755_), .Y(po0986));
  XOR2X1   g29079(.A(new_n31424_), .B(new_n31422_), .Y(po0987));
  NAND3X1  g29080(.A(pi1162), .B(pi1091), .C(new_n12898_), .Y(new_n31517_));
  NOR4X1   g29081(.A(new_n31517_), .B(new_n2740_), .C(pi1163), .D(new_n6751_), .Y(po0989));
  OAI22X1  g29082(.A0(new_n11923_), .A1(new_n2755_), .B0(new_n2739_), .B1(new_n2721_), .Y(po0990));
  AND2X1   g29083(.A(new_n2739_), .B(pi0946), .Y(po0991));
  INVX1    g29084(.A(pi0282), .Y(new_n31521_));
  NOR3X1   g29085(.A(new_n30448_), .B(pi0281), .C(pi0269), .Y(new_n31522_));
  XOR2X1   g29086(.A(new_n31522_), .B(new_n31521_), .Y(po0992));
  MX2X1    g29087(.A(pi1049), .B(pi0837), .S0(pi0955), .Y(po0993));
  MX2X1    g29088(.A(pi1047), .B(pi0838), .S0(pi0955), .Y(po0994));
  MX2X1    g29089(.A(pi1074), .B(pi0839), .S0(pi0955), .Y(po0995));
  MX2X1    g29090(.A(pi0840), .B(pi1196), .S0(new_n2739_), .Y(po0996));
  NOR3X1   g29091(.A(new_n6819_), .B(pi0034), .C(pi0033), .Y(po0997));
  MX2X1    g29092(.A(pi1035), .B(pi0842), .S0(pi0955), .Y(po0998));
  MX2X1    g29093(.A(pi1079), .B(pi0843), .S0(pi0955), .Y(po0999));
  MX2X1    g29094(.A(pi1078), .B(pi0844), .S0(pi0955), .Y(po1000));
  MX2X1    g29095(.A(pi1043), .B(pi0845), .S0(pi0955), .Y(po1001));
  MX2X1    g29096(.A(pi0846), .B(pi1134), .S0(new_n28069_), .Y(po1002));
  MX2X1    g29097(.A(pi1055), .B(pi0847), .S0(pi0955), .Y(po1003));
  MX2X1    g29098(.A(pi1039), .B(pi0848), .S0(pi0955), .Y(po1004));
  MX2X1    g29099(.A(pi0849), .B(pi1198), .S0(new_n2739_), .Y(po1005));
  MX2X1    g29100(.A(pi1048), .B(pi0850), .S0(pi0955), .Y(po1006));
  MX2X1    g29101(.A(pi1045), .B(pi0851), .S0(pi0955), .Y(po1007));
  MX2X1    g29102(.A(pi1062), .B(pi0852), .S0(pi0955), .Y(po1008));
  MX2X1    g29103(.A(pi1080), .B(pi0853), .S0(pi0955), .Y(po1009));
  MX2X1    g29104(.A(pi1051), .B(pi0854), .S0(pi0955), .Y(po1010));
  MX2X1    g29105(.A(pi1065), .B(pi0855), .S0(pi0955), .Y(po1011));
  MX2X1    g29106(.A(pi1067), .B(pi0856), .S0(pi0955), .Y(po1012));
  MX2X1    g29107(.A(pi1058), .B(pi0857), .S0(pi0955), .Y(po1013));
  MX2X1    g29108(.A(pi1087), .B(pi0858), .S0(pi0955), .Y(po1014));
  MX2X1    g29109(.A(pi1070), .B(pi0859), .S0(pi0955), .Y(po1015));
  MX2X1    g29110(.A(pi1076), .B(pi0860), .S0(pi0955), .Y(po1016));
  MX2X1    g29111(.A(new_n3847_), .B(new_n3744_), .S0(new_n2756_), .Y(new_n31548_));
  NOR2X1   g29112(.A(pi1141), .B(pi0123), .Y(new_n31549_));
  OAI21X1  g29113(.A0(pi0861), .A1(new_n28068_), .B0(pi0228), .Y(new_n31550_));
  OAI22X1  g29114(.A0(new_n31550_), .A1(new_n31549_), .B0(new_n31548_), .B1(pi0228), .Y(po1017));
  MX2X1    g29115(.A(pi0862), .B(pi1139), .S0(new_n28069_), .Y(po1018));
  MX2X1    g29116(.A(pi0863), .B(pi1199), .S0(new_n2739_), .Y(po1019));
  MX2X1    g29117(.A(pi0864), .B(pi1197), .S0(new_n2739_), .Y(po1020));
  MX2X1    g29118(.A(pi1040), .B(pi0865), .S0(pi0955), .Y(po1021));
  MX2X1    g29119(.A(pi1053), .B(pi0866), .S0(pi0955), .Y(po1022));
  MX2X1    g29120(.A(pi1057), .B(pi0867), .S0(pi0955), .Y(po1023));
  MX2X1    g29121(.A(pi1063), .B(pi0868), .S0(pi0955), .Y(po1024));
  MX2X1    g29122(.A(new_n3988_), .B(new_n3887_), .S0(new_n2756_), .Y(new_n31559_));
  NOR2X1   g29123(.A(pi1140), .B(pi0123), .Y(new_n31560_));
  OAI21X1  g29124(.A0(pi0869), .A1(new_n28068_), .B0(pi0228), .Y(new_n31561_));
  OAI22X1  g29125(.A0(new_n31561_), .A1(new_n31560_), .B0(new_n31559_), .B1(pi0228), .Y(po1025));
  MX2X1    g29126(.A(pi1069), .B(pi0870), .S0(pi0955), .Y(po1026));
  MX2X1    g29127(.A(pi1072), .B(pi0871), .S0(pi0955), .Y(po1027));
  MX2X1    g29128(.A(pi1084), .B(pi0872), .S0(pi0955), .Y(po1028));
  MX2X1    g29129(.A(pi1044), .B(pi0873), .S0(pi0955), .Y(po1029));
  MX2X1    g29130(.A(pi1036), .B(pi0874), .S0(pi0955), .Y(po1030));
  MX2X1    g29131(.A(new_n28946_), .B(new_n4460_), .S0(new_n2756_), .Y(new_n31568_));
  OR2X1    g29132(.A(new_n28946_), .B(pi0123), .Y(new_n31569_));
  AOI21X1  g29133(.A0(pi0875), .A1(pi0123), .B0(new_n3013_), .Y(new_n31570_));
  AOI22X1  g29134(.A0(new_n31570_), .A1(new_n31569_), .B0(new_n31568_), .B1(new_n3013_), .Y(po1031));
  MX2X1    g29135(.A(pi1037), .B(pi0876), .S0(pi0955), .Y(po1032));
  MX2X1    g29136(.A(new_n4281_), .B(new_n4180_), .S0(new_n2756_), .Y(new_n31573_));
  NOR2X1   g29137(.A(pi1138), .B(pi0123), .Y(new_n31574_));
  OAI21X1  g29138(.A0(pi0877), .A1(new_n28068_), .B0(pi0228), .Y(new_n31575_));
  OAI22X1  g29139(.A0(new_n31575_), .A1(new_n31574_), .B0(new_n31573_), .B1(pi0228), .Y(po1033));
  MX2X1    g29140(.A(new_n4422_), .B(new_n4321_), .S0(new_n2756_), .Y(new_n31577_));
  NOR2X1   g29141(.A(pi1137), .B(pi0123), .Y(new_n31578_));
  OAI21X1  g29142(.A0(pi0878), .A1(new_n28068_), .B0(pi0228), .Y(new_n31579_));
  OAI22X1  g29143(.A0(new_n31579_), .A1(new_n31578_), .B0(new_n31577_), .B1(pi0228), .Y(po1034));
  MX2X1    g29144(.A(new_n28313_), .B(new_n4609_), .S0(new_n2756_), .Y(new_n31581_));
  NOR2X1   g29145(.A(pi1135), .B(pi0123), .Y(new_n31582_));
  OAI21X1  g29146(.A0(pi0879), .A1(new_n28068_), .B0(pi0228), .Y(new_n31583_));
  OAI22X1  g29147(.A0(new_n31583_), .A1(new_n31582_), .B0(new_n31581_), .B1(pi0228), .Y(po1035));
  MX2X1    g29148(.A(pi1081), .B(pi0880), .S0(pi0955), .Y(po1036));
  MX2X1    g29149(.A(pi1059), .B(pi0881), .S0(pi0955), .Y(po1037));
  INVX1    g29150(.A(pi0883), .Y(po1163));
  MX2X1    g29151(.A(pi1107), .B(po1163), .S0(new_n31461_), .Y(po1039));
  INVX1    g29152(.A(pi0884), .Y(po1180));
  MX2X1    g29153(.A(pi1124), .B(po1180), .S0(new_n31461_), .Y(po1040));
  INVX1    g29154(.A(pi0885), .Y(po1172));
  MX2X1    g29155(.A(pi1125), .B(po1172), .S0(new_n31461_), .Y(po1041));
  INVX1    g29156(.A(pi0886), .Y(po1166));
  MX2X1    g29157(.A(pi1109), .B(po1166), .S0(new_n31461_), .Y(po1042));
  INVX1    g29158(.A(pi0887), .Y(po1179));
  MX2X1    g29159(.A(pi1100), .B(po1179), .S0(new_n31461_), .Y(po1043));
  INVX1    g29160(.A(pi0888), .Y(po1164));
  MX2X1    g29161(.A(pi1120), .B(po1164), .S0(new_n31461_), .Y(po1044));
  INVX1    g29162(.A(pi0889), .Y(po1170));
  MX2X1    g29163(.A(pi1103), .B(po1170), .S0(new_n31461_), .Y(po1045));
  INVX1    g29164(.A(pi0890), .Y(po1153));
  MX2X1    g29165(.A(pi1126), .B(po1153), .S0(new_n31461_), .Y(po1046));
  INVX1    g29166(.A(pi0891), .Y(po1160));
  MX2X1    g29167(.A(pi1116), .B(po1160), .S0(new_n31461_), .Y(po1047));
  INVX1    g29168(.A(pi0892), .Y(po1183));
  MX2X1    g29169(.A(pi1101), .B(po1183), .S0(new_n31461_), .Y(po1048));
  INVX1    g29170(.A(pi0894), .Y(po1150));
  MX2X1    g29171(.A(pi1119), .B(po1150), .S0(new_n31461_), .Y(po1050));
  INVX1    g29172(.A(pi0895), .Y(po1168));
  MX2X1    g29173(.A(pi1113), .B(po1168), .S0(new_n31461_), .Y(po1051));
  INVX1    g29174(.A(pi0896), .Y(po1156));
  MX2X1    g29175(.A(pi1118), .B(po1156), .S0(new_n31461_), .Y(po1052));
  INVX1    g29176(.A(pi0898), .Y(po1176));
  MX2X1    g29177(.A(pi1129), .B(po1176), .S0(new_n31461_), .Y(po1054));
  INVX1    g29178(.A(pi0899), .Y(po1174));
  MX2X1    g29179(.A(pi1115), .B(po1174), .S0(new_n31461_), .Y(po1055));
  INVX1    g29180(.A(pi0900), .Y(po1171));
  MX2X1    g29181(.A(pi1110), .B(po1171), .S0(new_n31461_), .Y(po1056));
  INVX1    g29182(.A(pi0902), .Y(po1161));
  MX2X1    g29183(.A(pi1111), .B(po1161), .S0(new_n31461_), .Y(po1058));
  INVX1    g29184(.A(pi0903), .Y(po1162));
  MX2X1    g29185(.A(pi1121), .B(po1162), .S0(new_n31461_), .Y(po1059));
  INVX1    g29186(.A(pi0904), .Y(po1173));
  MX2X1    g29187(.A(pi1127), .B(po1173), .S0(new_n31461_), .Y(po1060));
  INVX1    g29188(.A(pi0905), .Y(po1151));
  MX2X1    g29189(.A(pi1131), .B(po1151), .S0(new_n31461_), .Y(po1061));
  INVX1    g29190(.A(pi0906), .Y(po1155));
  MX2X1    g29191(.A(pi1128), .B(po1155), .S0(new_n31461_), .Y(po1062));
  INVX1    g29192(.A(pi0782), .Y(new_n31629_));
  AOI21X1  g29193(.A0(pi0979), .A1(new_n30259_), .B0(new_n31629_), .Y(new_n31630_));
  OAI21X1  g29194(.A0(pi0979), .A1(pi0624), .B0(new_n31630_), .Y(new_n31631_));
  INVX1    g29195(.A(pi0615), .Y(new_n31632_));
  MX2X1    g29196(.A(new_n31632_), .B(pi0604), .S0(new_n5035_), .Y(new_n31633_));
  MX2X1    g29197(.A(new_n31633_), .B(pi0907), .S0(new_n31629_), .Y(new_n31634_));
  AND2X1   g29198(.A(new_n31634_), .B(new_n31631_), .Y(po1063));
  INVX1    g29199(.A(pi0908), .Y(po1159));
  MX2X1    g29200(.A(pi1122), .B(po1159), .S0(new_n31461_), .Y(po1064));
  INVX1    g29201(.A(pi0909), .Y(po1157));
  MX2X1    g29202(.A(pi1105), .B(po1157), .S0(new_n31461_), .Y(po1065));
  INVX1    g29203(.A(pi0910), .Y(po1181));
  MX2X1    g29204(.A(pi1117), .B(po1181), .S0(new_n31461_), .Y(po1066));
  INVX1    g29205(.A(pi0911), .Y(po1158));
  MX2X1    g29206(.A(pi1130), .B(po1158), .S0(new_n31461_), .Y(po1067));
  INVX1    g29207(.A(pi0912), .Y(po1167));
  MX2X1    g29208(.A(pi1114), .B(po1167), .S0(new_n31461_), .Y(po1068));
  INVX1    g29209(.A(pi0913), .Y(po1149));
  MX2X1    g29210(.A(pi1106), .B(po1149), .S0(new_n31461_), .Y(po1069));
  XOR2X1   g29211(.A(new_n30446_), .B(new_n30445_), .Y(po1070));
  INVX1    g29212(.A(pi0915), .Y(po1146));
  MX2X1    g29213(.A(pi1108), .B(po1146), .S0(new_n31461_), .Y(po1071));
  INVX1    g29214(.A(pi0916), .Y(po1169));
  MX2X1    g29215(.A(pi1123), .B(po1169), .S0(new_n31461_), .Y(po1072));
  INVX1    g29216(.A(pi0917), .Y(po1177));
  MX2X1    g29217(.A(pi1112), .B(po1177), .S0(new_n31461_), .Y(po1073));
  INVX1    g29218(.A(pi0918), .Y(po1175));
  MX2X1    g29219(.A(pi1104), .B(po1175), .S0(new_n31461_), .Y(po1074));
  INVX1    g29220(.A(pi0919), .Y(po1165));
  MX2X1    g29221(.A(pi1102), .B(po1165), .S0(new_n31461_), .Y(po1075));
  MX2X1    g29222(.A(pi0920), .B(pi1139), .S0(pi1093), .Y(po1076));
  MX2X1    g29223(.A(pi0921), .B(pi1140), .S0(pi1093), .Y(po1077));
  MX2X1    g29224(.A(pi0922), .B(pi1152), .S0(pi1093), .Y(po1078));
  MX2X1    g29225(.A(pi0923), .B(pi1154), .S0(pi1093), .Y(po1079));
  INVX1    g29226(.A(pi0311), .Y(new_n31663_));
  NOR4X1   g29227(.A(pi0312), .B(new_n31663_), .C(new_n29116_), .D(pi0300), .Y(po1080));
  MX2X1    g29228(.A(pi0925), .B(pi1155), .S0(pi1093), .Y(po1081));
  MX2X1    g29229(.A(pi0926), .B(pi1157), .S0(pi1093), .Y(po1082));
  MX2X1    g29230(.A(pi0927), .B(pi1145), .S0(pi1093), .Y(po1083));
  MX2X1    g29231(.A(pi0928), .B(pi1136), .S0(pi1093), .Y(po1084));
  MX2X1    g29232(.A(pi0929), .B(pi1144), .S0(pi1093), .Y(po1085));
  MX2X1    g29233(.A(pi0930), .B(pi1134), .S0(pi1093), .Y(po1086));
  MX2X1    g29234(.A(pi0931), .B(pi1150), .S0(pi1093), .Y(po1087));
  MX2X1    g29235(.A(pi0932), .B(pi1142), .S0(pi1093), .Y(po1088));
  MX2X1    g29236(.A(pi0933), .B(pi1137), .S0(pi1093), .Y(po1089));
  MX2X1    g29237(.A(pi0934), .B(pi1147), .S0(pi1093), .Y(po1090));
  MX2X1    g29238(.A(pi0935), .B(pi1141), .S0(pi1093), .Y(po1091));
  MX2X1    g29239(.A(pi0936), .B(pi1149), .S0(pi1093), .Y(po1092));
  MX2X1    g29240(.A(pi0937), .B(pi1148), .S0(pi1093), .Y(po1093));
  MX2X1    g29241(.A(pi0938), .B(pi1135), .S0(pi1093), .Y(po1094));
  MX2X1    g29242(.A(pi0939), .B(pi1146), .S0(pi1093), .Y(po1095));
  MX2X1    g29243(.A(pi0940), .B(pi1138), .S0(pi1093), .Y(po1096));
  MX2X1    g29244(.A(pi0941), .B(pi1153), .S0(pi1093), .Y(po1097));
  MX2X1    g29245(.A(pi0942), .B(pi1156), .S0(pi1093), .Y(po1098));
  MX2X1    g29246(.A(pi0943), .B(pi1151), .S0(pi1093), .Y(po1099));
  MX2X1    g29247(.A(pi0944), .B(pi1143), .S0(pi1093), .Y(po1100));
  AND2X1   g29248(.A(new_n2739_), .B(pi0230), .Y(po1102));
  OAI21X1  g29249(.A0(new_n14590_), .A1(pi0782), .B0(new_n31631_), .Y(po1103));
  XOR2X1   g29250(.A(pi0992), .B(pi0266), .Y(po1104));
  MX2X1    g29251(.A(pi0949), .B(new_n29164_), .S0(po1110), .Y(po1105));
  NOR3X1   g29252(.A(new_n5982_), .B(new_n2755_), .C(new_n5258_), .Y(po1107));
  OAI21X1  g29253(.A0(new_n2755_), .A1(new_n2780_), .B0(new_n6750_), .Y(po1112));
  AND2X1   g29254(.A(pi0960), .B(new_n31629_), .Y(po1115));
  AND2X1   g29255(.A(pi0961), .B(new_n24954_), .Y(po1116));
  AND2X1   g29256(.A(pi0963), .B(new_n31629_), .Y(po1118));
  AND2X1   g29257(.A(pi0967), .B(new_n24954_), .Y(po1122));
  AND2X1   g29258(.A(pi0969), .B(new_n24954_), .Y(po1124));
  AND2X1   g29259(.A(pi0970), .B(new_n31629_), .Y(po1125));
  AND2X1   g29260(.A(pi0971), .B(new_n24954_), .Y(po1126));
  AND2X1   g29261(.A(pi0972), .B(new_n31629_), .Y(po1127));
  AND2X1   g29262(.A(pi0974), .B(new_n24954_), .Y(po1128));
  AND2X1   g29263(.A(pi0975), .B(new_n31629_), .Y(po1129));
  AND2X1   g29264(.A(pi0977), .B(new_n24954_), .Y(po1131));
  AND2X1   g29265(.A(pi0978), .B(new_n31629_), .Y(po1132));
  OR2X1    g29266(.A(new_n31632_), .B(pi0598), .Y(po1133));
  AND2X1   g29267(.A(pi1092), .B(pi0824), .Y(po1135));
  OR2X1    g29268(.A(pi0624), .B(pi0604), .Y(po1137));
  ONE      g29269(.Y(po0166));
  BUFX1    g29270(.A(pi0668), .Y(po0000));
  BUFX1    g29271(.A(pi0672), .Y(po0001));
  BUFX1    g29272(.A(pi0664), .Y(po0002));
  BUFX1    g29273(.A(pi0667), .Y(po0003));
  BUFX1    g29274(.A(pi0676), .Y(po0004));
  BUFX1    g29275(.A(pi0673), .Y(po0005));
  BUFX1    g29276(.A(pi0675), .Y(po0006));
  BUFX1    g29277(.A(pi0666), .Y(po0007));
  BUFX1    g29278(.A(pi0679), .Y(po0008));
  BUFX1    g29279(.A(pi0674), .Y(po0009));
  BUFX1    g29280(.A(pi0663), .Y(po0010));
  BUFX1    g29281(.A(pi0670), .Y(po0011));
  BUFX1    g29282(.A(pi0677), .Y(po0012));
  BUFX1    g29283(.A(pi0682), .Y(po0013));
  BUFX1    g29284(.A(pi0671), .Y(po0014));
  BUFX1    g29285(.A(pi0678), .Y(po0015));
  BUFX1    g29286(.A(pi0718), .Y(po0016));
  BUFX1    g29287(.A(pi0707), .Y(po0017));
  BUFX1    g29288(.A(pi0708), .Y(po0018));
  BUFX1    g29289(.A(pi0713), .Y(po0019));
  BUFX1    g29290(.A(pi0711), .Y(po0020));
  BUFX1    g29291(.A(pi0716), .Y(po0021));
  BUFX1    g29292(.A(pi0733), .Y(po0022));
  BUFX1    g29293(.A(pi0712), .Y(po0023));
  BUFX1    g29294(.A(pi0689), .Y(po0024));
  BUFX1    g29295(.A(pi0717), .Y(po0025));
  BUFX1    g29296(.A(pi0692), .Y(po0026));
  BUFX1    g29297(.A(pi0719), .Y(po0027));
  BUFX1    g29298(.A(pi0722), .Y(po0028));
  BUFX1    g29299(.A(pi0714), .Y(po0029));
  BUFX1    g29300(.A(pi0720), .Y(po0030));
  BUFX1    g29301(.A(pi0685), .Y(po0031));
  BUFX1    g29302(.A(pi0837), .Y(po0032));
  BUFX1    g29303(.A(pi0850), .Y(po0033));
  BUFX1    g29304(.A(pi0872), .Y(po0034));
  BUFX1    g29305(.A(pi0871), .Y(po0035));
  BUFX1    g29306(.A(pi0881), .Y(po0036));
  BUFX1    g29307(.A(pi0866), .Y(po0037));
  BUFX1    g29308(.A(pi0876), .Y(po0038));
  BUFX1    g29309(.A(pi0873), .Y(po0039));
  BUFX1    g29310(.A(pi0874), .Y(po0040));
  BUFX1    g29311(.A(pi0859), .Y(po0041));
  BUFX1    g29312(.A(pi0855), .Y(po0042));
  BUFX1    g29313(.A(pi0852), .Y(po0043));
  BUFX1    g29314(.A(pi0870), .Y(po0044));
  BUFX1    g29315(.A(pi0848), .Y(po0045));
  BUFX1    g29316(.A(pi0865), .Y(po0046));
  BUFX1    g29317(.A(pi0856), .Y(po0047));
  BUFX1    g29318(.A(pi0853), .Y(po0048));
  BUFX1    g29319(.A(pi0847), .Y(po0049));
  BUFX1    g29320(.A(pi0857), .Y(po0050));
  BUFX1    g29321(.A(pi0854), .Y(po0051));
  BUFX1    g29322(.A(pi0858), .Y(po0052));
  BUFX1    g29323(.A(pi0845), .Y(po0053));
  BUFX1    g29324(.A(pi0838), .Y(po0054));
  BUFX1    g29325(.A(pi0842), .Y(po0055));
  BUFX1    g29326(.A(pi0843), .Y(po0056));
  BUFX1    g29327(.A(pi0839), .Y(po0057));
  BUFX1    g29328(.A(pi0844), .Y(po0058));
  BUFX1    g29329(.A(pi0868), .Y(po0059));
  BUFX1    g29330(.A(pi0851), .Y(po0060));
  BUFX1    g29331(.A(pi0867), .Y(po0061));
  BUFX1    g29332(.A(pi0880), .Y(po0062));
  BUFX1    g29333(.A(pi0860), .Y(po0063));
  BUFX1    g29334(.A(pi1030), .Y(po0064));
  BUFX1    g29335(.A(pi1034), .Y(po0065));
  BUFX1    g29336(.A(pi1015), .Y(po0066));
  BUFX1    g29337(.A(pi1020), .Y(po0067));
  BUFX1    g29338(.A(pi1025), .Y(po0068));
  BUFX1    g29339(.A(pi1005), .Y(po0069));
  BUFX1    g29340(.A(pi0996), .Y(po0070));
  BUFX1    g29341(.A(pi1012), .Y(po0071));
  BUFX1    g29342(.A(pi0993), .Y(po0072));
  BUFX1    g29343(.A(pi1016), .Y(po0073));
  BUFX1    g29344(.A(pi1021), .Y(po0074));
  BUFX1    g29345(.A(pi1010), .Y(po0075));
  BUFX1    g29346(.A(pi1027), .Y(po0076));
  BUFX1    g29347(.A(pi1018), .Y(po0077));
  BUFX1    g29348(.A(pi1017), .Y(po0078));
  BUFX1    g29349(.A(pi1024), .Y(po0079));
  BUFX1    g29350(.A(pi1009), .Y(po0080));
  BUFX1    g29351(.A(pi1032), .Y(po0081));
  BUFX1    g29352(.A(pi1003), .Y(po0082));
  BUFX1    g29353(.A(pi0997), .Y(po0083));
  BUFX1    g29354(.A(pi1013), .Y(po0084));
  BUFX1    g29355(.A(pi1011), .Y(po0085));
  BUFX1    g29356(.A(pi1008), .Y(po0086));
  BUFX1    g29357(.A(pi1019), .Y(po0087));
  BUFX1    g29358(.A(pi1031), .Y(po0088));
  BUFX1    g29359(.A(pi1022), .Y(po0089));
  BUFX1    g29360(.A(pi1000), .Y(po0090));
  BUFX1    g29361(.A(pi1023), .Y(po0091));
  BUFX1    g29362(.A(pi1002), .Y(po0092));
  BUFX1    g29363(.A(pi1026), .Y(po0093));
  BUFX1    g29364(.A(pi1006), .Y(po0094));
  BUFX1    g29365(.A(pi0998), .Y(po0095));
  BUFX1    g29366(.A(pi0031), .Y(po0096));
  BUFX1    g29367(.A(pi0080), .Y(po0097));
  BUFX1    g29368(.A(pi0893), .Y(po0098));
  BUFX1    g29369(.A(pi0467), .Y(po0099));
  BUFX1    g29370(.A(pi0078), .Y(po0100));
  BUFX1    g29371(.A(pi0112), .Y(po0101));
  BUFX1    g29372(.A(pi0013), .Y(po0102));
  BUFX1    g29373(.A(pi0025), .Y(po0103));
  BUFX1    g29374(.A(pi0226), .Y(po0104));
  BUFX1    g29375(.A(pi0127), .Y(po0105));
  BUFX1    g29376(.A(pi0822), .Y(po0106));
  BUFX1    g29377(.A(pi0808), .Y(po0107));
  BUFX1    g29378(.A(pi0227), .Y(po0108));
  BUFX1    g29379(.A(pi0477), .Y(po0109));
  BUFX1    g29380(.A(pi0834), .Y(po0110));
  BUFX1    g29381(.A(pi0229), .Y(po0111));
  BUFX1    g29382(.A(pi0012), .Y(po0112));
  BUFX1    g29383(.A(pi0011), .Y(po0113));
  BUFX1    g29384(.A(pi0010), .Y(po0114));
  BUFX1    g29385(.A(pi0009), .Y(po0115));
  BUFX1    g29386(.A(pi0008), .Y(po0116));
  BUFX1    g29387(.A(pi0007), .Y(po0117));
  BUFX1    g29388(.A(pi0006), .Y(po0118));
  BUFX1    g29389(.A(pi0005), .Y(po0119));
  BUFX1    g29390(.A(pi0004), .Y(po0120));
  BUFX1    g29391(.A(pi0003), .Y(po0121));
  BUFX1    g29392(.A(pi0000), .Y(po0122));
  BUFX1    g29393(.A(pi0002), .Y(po0123));
  BUFX1    g29394(.A(pi0001), .Y(po0124));
  BUFX1    g29395(.A(pi0310), .Y(po0125));
  BUFX1    g29396(.A(pi0302), .Y(po0126));
  BUFX1    g29397(.A(pi0475), .Y(po0127));
  BUFX1    g29398(.A(pi0474), .Y(po0128));
  BUFX1    g29399(.A(pi0466), .Y(po0129));
  BUFX1    g29400(.A(pi0473), .Y(po0130));
  BUFX1    g29401(.A(pi0471), .Y(po0131));
  BUFX1    g29402(.A(pi0472), .Y(po0132));
  BUFX1    g29403(.A(pi0470), .Y(po0133));
  BUFX1    g29404(.A(pi0469), .Y(po0134));
  BUFX1    g29405(.A(pi0465), .Y(po0135));
  BUFX1    g29406(.A(pi1028), .Y(po0136));
  BUFX1    g29407(.A(pi1033), .Y(po0137));
  BUFX1    g29408(.A(pi0995), .Y(po0138));
  BUFX1    g29409(.A(pi0994), .Y(po0139));
  BUFX1    g29410(.A(pi0028), .Y(po0140));
  BUFX1    g29411(.A(pi0027), .Y(po0141));
  BUFX1    g29412(.A(pi0026), .Y(po0142));
  BUFX1    g29413(.A(pi0029), .Y(po0143));
  BUFX1    g29414(.A(pi0015), .Y(po0144));
  BUFX1    g29415(.A(pi0014), .Y(po0145));
  BUFX1    g29416(.A(pi0021), .Y(po0146));
  BUFX1    g29417(.A(pi0020), .Y(po0147));
  BUFX1    g29418(.A(pi0019), .Y(po0148));
  BUFX1    g29419(.A(pi0018), .Y(po0149));
  BUFX1    g29420(.A(pi0017), .Y(po0150));
  BUFX1    g29421(.A(pi0016), .Y(po0151));
  BUFX1    g29422(.A(pi1096), .Y(po0152));
  BUFX1    g29423(.A(pi0228), .Y(po0168));
  BUFX1    g29424(.A(pi0022), .Y(po0169));
  BUFX1    g29425(.A(pi1089), .Y(po0179));
  BUFX1    g29426(.A(pi0023), .Y(po0180));
  MX2X1    g29427(.A(new_n5114_), .B(new_n4986_), .S0(pi0057), .Y(po0181));
  BUFX1    g29428(.A(pi0037), .Y(po0188));
  BUFX1    g29429(.A(pi0117), .Y(po0263));
  BUFX1    g29430(.A(pi0131), .Y(po0285));
  BUFX1    g29431(.A(pi0232), .Y(po0386));
  BUFX1    g29432(.A(pi0236), .Y(po0388));
  BUFX1    g29433(.A(pi0583), .Y(po0636));
  BUFX1    g29434(.A(pi0067), .Y(po1053));
  BUFX1    g29435(.A(pi1134), .Y(po1108));
  BUFX1    g29436(.A(pi0964), .Y(po1109));
  BUFX1    g29437(.A(pi0965), .Y(po1111));
  BUFX1    g29438(.A(pi0991), .Y(po1113));
  BUFX1    g29439(.A(pi0985), .Y(po1114));
  BUFX1    g29440(.A(pi1014), .Y(po1117));
  BUFX1    g29441(.A(pi1029), .Y(po1119));
  BUFX1    g29442(.A(pi1004), .Y(po1120));
  BUFX1    g29443(.A(pi1007), .Y(po1121));
  BUFX1    g29444(.A(pi1135), .Y(po1123));
  BUFX1    g29445(.A(pi1064), .Y(po1134));
  BUFX1    g29446(.A(pi0299), .Y(po1136));
  BUFX1    g29447(.A(pi1075), .Y(po1138));
  BUFX1    g29448(.A(pi1052), .Y(po1139));
  BUFX1    g29449(.A(pi0771), .Y(po1140));
  BUFX1    g29450(.A(pi0765), .Y(po1141));
  BUFX1    g29451(.A(pi0605), .Y(po1142));
  BUFX1    g29452(.A(pi0601), .Y(po1143));
  BUFX1    g29453(.A(pi0278), .Y(po1144));
  BUFX1    g29454(.A(pi0279), .Y(po1145));
  BUFX1    g29455(.A(pi1095), .Y(po1152));
  BUFX1    g29456(.A(pi1094), .Y(po1154));
  BUFX1    g29457(.A(pi1187), .Y(po1184));
  BUFX1    g29458(.A(pi1172), .Y(po1185));
  BUFX1    g29459(.A(pi1170), .Y(po1186));
  BUFX1    g29460(.A(pi1138), .Y(po1187));
  BUFX1    g29461(.A(pi1177), .Y(po1188));
  BUFX1    g29462(.A(pi1178), .Y(po1189));
  BUFX1    g29463(.A(pi0863), .Y(po1190));
  BUFX1    g29464(.A(pi1203), .Y(po1191));
  BUFX1    g29465(.A(pi1185), .Y(po1192));
  BUFX1    g29466(.A(pi1171), .Y(po1193));
  BUFX1    g29467(.A(pi1192), .Y(po1194));
  BUFX1    g29468(.A(pi1137), .Y(po1195));
  BUFX1    g29469(.A(pi1186), .Y(po1196));
  BUFX1    g29470(.A(pi1165), .Y(po1197));
  BUFX1    g29471(.A(pi1164), .Y(po1198));
  BUFX1    g29472(.A(pi1098), .Y(po1199));
  BUFX1    g29473(.A(pi1183), .Y(po1200));
  BUFX1    g29474(.A(pi0230), .Y(po1201));
  BUFX1    g29475(.A(pi1169), .Y(po1202));
  BUFX1    g29476(.A(pi1136), .Y(po1203));
  BUFX1    g29477(.A(pi1181), .Y(po1204));
  BUFX1    g29478(.A(pi0849), .Y(po1205));
  BUFX1    g29479(.A(pi1193), .Y(po1206));
  BUFX1    g29480(.A(pi1182), .Y(po1207));
  BUFX1    g29481(.A(pi1168), .Y(po1208));
  BUFX1    g29482(.A(pi1175), .Y(po1209));
  BUFX1    g29483(.A(pi1191), .Y(po1210));
  BUFX1    g29484(.A(pi1099), .Y(po1211));
  BUFX1    g29485(.A(pi1174), .Y(po1212));
  BUFX1    g29486(.A(pi1179), .Y(po1213));
  BUFX1    g29487(.A(pi1202), .Y(po1214));
  BUFX1    g29488(.A(pi1176), .Y(po1215));
  BUFX1    g29489(.A(pi1173), .Y(po1216));
  BUFX1    g29490(.A(pi1201), .Y(po1217));
  BUFX1    g29491(.A(pi1167), .Y(po1218));
  BUFX1    g29492(.A(pi0840), .Y(po1219));
  BUFX1    g29493(.A(pi1189), .Y(po1220));
  BUFX1    g29494(.A(pi1195), .Y(po1221));
  BUFX1    g29495(.A(pi0864), .Y(po1222));
  BUFX1    g29496(.A(pi1190), .Y(po1223));
  BUFX1    g29497(.A(pi1188), .Y(po1224));
  BUFX1    g29498(.A(pi1180), .Y(po1225));
  BUFX1    g29499(.A(pi1194), .Y(po1226));
  BUFX1    g29500(.A(pi1097), .Y(po1227));
  BUFX1    g29501(.A(pi1166), .Y(po1228));
  BUFX1    g29502(.A(pi1200), .Y(po1229));
  BUFX1    g29503(.A(pi1184), .Y(po1230));
endmodule


