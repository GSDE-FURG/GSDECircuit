// Benchmark "top" written by ABC on Mon Sep 21 03:36:50 2020

module top ( 
    \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] , \a[24] ,
    \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] , \a[32] ,
    \a[33] , \a[34] , \a[35] , \a[36] , \a[37] , \a[38] , \a[39] , \a[40] ,
    \a[41] , \a[42] , \a[43] , \a[44] , \a[45] , \a[46] , \a[47] , \a[48] ,
    \a[49] , \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] , \a[56] ,
    \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] , \a[64] ,
    \a[65] , \a[66] , \a[67] , \a[68] , \a[69] , \a[70] , \a[71] , \a[72] ,
    \a[73] , \a[74] , \a[75] , \a[76] , \a[77] , \a[78] , \a[79] , \a[80] ,
    \a[81] , \a[82] , \a[83] , \a[84] , \a[85] , \a[86] , \a[87] , \a[88] ,
    \a[89] , \a[90] , \a[91] , \a[92] , \a[93] , \a[94] , \a[95] , \a[96] ,
    \a[97] , \a[98] , \a[99] , \a[100] , \a[101] , \a[102] , \a[103] ,
    \a[104] , \a[105] , \a[106] , \a[107] , \a[108] , \a[109] , \a[110] ,
    \a[111] , \a[112] , \a[113] , \a[114] , \a[115] , \a[116] , \a[117] ,
    \a[118] , \a[119] , \a[120] , \a[121] , \a[122] , \a[123] , \a[124] ,
    \a[125] , \a[126] , \a[127] , \shift[0] , \shift[1] , \shift[2] ,
    \shift[3] , \shift[4] , \shift[5] , \shift[6] ,
    \result[0] , \result[1] , \result[2] , \result[3] , \result[4] ,
    \result[5] , \result[6] , \result[7] , \result[8] , \result[9] ,
    \result[10] , \result[11] , \result[12] , \result[13] , \result[14] ,
    \result[15] , \result[16] , \result[17] , \result[18] , \result[19] ,
    \result[20] , \result[21] , \result[22] , \result[23] , \result[24] ,
    \result[25] , \result[26] , \result[27] , \result[28] , \result[29] ,
    \result[30] , \result[31] , \result[32] , \result[33] , \result[34] ,
    \result[35] , \result[36] , \result[37] , \result[38] , \result[39] ,
    \result[40] , \result[41] , \result[42] , \result[43] , \result[44] ,
    \result[45] , \result[46] , \result[47] , \result[48] , \result[49] ,
    \result[50] , \result[51] , \result[52] , \result[53] , \result[54] ,
    \result[55] , \result[56] , \result[57] , \result[58] , \result[59] ,
    \result[60] , \result[61] , \result[62] , \result[63] , \result[64] ,
    \result[65] , \result[66] , \result[67] , \result[68] , \result[69] ,
    \result[70] , \result[71] , \result[72] , \result[73] , \result[74] ,
    \result[75] , \result[76] , \result[77] , \result[78] , \result[79] ,
    \result[80] , \result[81] , \result[82] , \result[83] , \result[84] ,
    \result[85] , \result[86] , \result[87] , \result[88] , \result[89] ,
    \result[90] , \result[91] , \result[92] , \result[93] , \result[94] ,
    \result[95] , \result[96] , \result[97] , \result[98] , \result[99] ,
    \result[100] , \result[101] , \result[102] , \result[103] ,
    \result[104] , \result[105] , \result[106] , \result[107] ,
    \result[108] , \result[109] , \result[110] , \result[111] ,
    \result[112] , \result[113] , \result[114] , \result[115] ,
    \result[116] , \result[117] , \result[118] , \result[119] ,
    \result[120] , \result[121] , \result[122] , \result[123] ,
    \result[124] , \result[125] , \result[126] , \result[127]   );
  input  \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] ,
    \a[8] , \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] ,
    \a[32] , \a[33] , \a[34] , \a[35] , \a[36] , \a[37] , \a[38] , \a[39] ,
    \a[40] , \a[41] , \a[42] , \a[43] , \a[44] , \a[45] , \a[46] , \a[47] ,
    \a[48] , \a[49] , \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] ,
    \a[56] , \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] ,
    \a[64] , \a[65] , \a[66] , \a[67] , \a[68] , \a[69] , \a[70] , \a[71] ,
    \a[72] , \a[73] , \a[74] , \a[75] , \a[76] , \a[77] , \a[78] , \a[79] ,
    \a[80] , \a[81] , \a[82] , \a[83] , \a[84] , \a[85] , \a[86] , \a[87] ,
    \a[88] , \a[89] , \a[90] , \a[91] , \a[92] , \a[93] , \a[94] , \a[95] ,
    \a[96] , \a[97] , \a[98] , \a[99] , \a[100] , \a[101] , \a[102] ,
    \a[103] , \a[104] , \a[105] , \a[106] , \a[107] , \a[108] , \a[109] ,
    \a[110] , \a[111] , \a[112] , \a[113] , \a[114] , \a[115] , \a[116] ,
    \a[117] , \a[118] , \a[119] , \a[120] , \a[121] , \a[122] , \a[123] ,
    \a[124] , \a[125] , \a[126] , \a[127] , \shift[0] , \shift[1] ,
    \shift[2] , \shift[3] , \shift[4] , \shift[5] , \shift[6] ;
  output \result[0] , \result[1] , \result[2] , \result[3] , \result[4] ,
    \result[5] , \result[6] , \result[7] , \result[8] , \result[9] ,
    \result[10] , \result[11] , \result[12] , \result[13] , \result[14] ,
    \result[15] , \result[16] , \result[17] , \result[18] , \result[19] ,
    \result[20] , \result[21] , \result[22] , \result[23] , \result[24] ,
    \result[25] , \result[26] , \result[27] , \result[28] , \result[29] ,
    \result[30] , \result[31] , \result[32] , \result[33] , \result[34] ,
    \result[35] , \result[36] , \result[37] , \result[38] , \result[39] ,
    \result[40] , \result[41] , \result[42] , \result[43] , \result[44] ,
    \result[45] , \result[46] , \result[47] , \result[48] , \result[49] ,
    \result[50] , \result[51] , \result[52] , \result[53] , \result[54] ,
    \result[55] , \result[56] , \result[57] , \result[58] , \result[59] ,
    \result[60] , \result[61] , \result[62] , \result[63] , \result[64] ,
    \result[65] , \result[66] , \result[67] , \result[68] , \result[69] ,
    \result[70] , \result[71] , \result[72] , \result[73] , \result[74] ,
    \result[75] , \result[76] , \result[77] , \result[78] , \result[79] ,
    \result[80] , \result[81] , \result[82] , \result[83] , \result[84] ,
    \result[85] , \result[86] , \result[87] , \result[88] , \result[89] ,
    \result[90] , \result[91] , \result[92] , \result[93] , \result[94] ,
    \result[95] , \result[96] , \result[97] , \result[98] , \result[99] ,
    \result[100] , \result[101] , \result[102] , \result[103] ,
    \result[104] , \result[105] , \result[106] , \result[107] ,
    \result[108] , \result[109] , \result[110] , \result[111] ,
    \result[112] , \result[113] , \result[114] , \result[115] ,
    \result[116] , \result[117] , \result[118] , \result[119] ,
    \result[120] , \result[121] , \result[122] , \result[123] ,
    \result[124] , \result[125] , \result[126] , \result[127] ;
  wire new_n264_, new_n265_, new_n266_, new_n267_, new_n268_, new_n269_,
    new_n270_, new_n271_, new_n272_, new_n273_, new_n274_, new_n275_,
    new_n276_, new_n277_, new_n278_, new_n279_, new_n280_, new_n281_,
    new_n282_, new_n283_, new_n284_, new_n285_, new_n286_, new_n287_,
    new_n288_, new_n289_, new_n290_, new_n291_, new_n292_, new_n293_,
    new_n294_, new_n295_, new_n296_, new_n297_, new_n298_, new_n299_,
    new_n300_, new_n301_, new_n302_, new_n303_, new_n304_, new_n305_,
    new_n306_, new_n307_, new_n308_, new_n309_, new_n310_, new_n311_,
    new_n312_, new_n313_, new_n314_, new_n315_, new_n316_, new_n317_,
    new_n318_, new_n319_, new_n320_, new_n321_, new_n322_, new_n323_,
    new_n324_, new_n325_, new_n326_, new_n327_, new_n328_, new_n329_,
    new_n330_, new_n331_, new_n332_, new_n333_, new_n334_, new_n335_,
    new_n336_, new_n337_, new_n338_, new_n339_, new_n340_, new_n341_,
    new_n342_, new_n343_, new_n344_, new_n345_, new_n346_, new_n347_,
    new_n348_, new_n349_, new_n350_, new_n351_, new_n352_, new_n353_,
    new_n354_, new_n355_, new_n356_, new_n357_, new_n358_, new_n359_,
    new_n360_, new_n361_, new_n362_, new_n363_, new_n364_, new_n365_,
    new_n366_, new_n367_, new_n368_, new_n369_, new_n370_, new_n371_,
    new_n372_, new_n373_, new_n374_, new_n375_, new_n376_, new_n377_,
    new_n378_, new_n379_, new_n380_, new_n381_, new_n382_, new_n383_,
    new_n384_, new_n385_, new_n386_, new_n387_, new_n388_, new_n389_,
    new_n390_, new_n391_, new_n392_, new_n393_, new_n394_, new_n395_,
    new_n396_, new_n397_, new_n398_, new_n399_, new_n400_, new_n401_,
    new_n402_, new_n403_, new_n404_, new_n405_, new_n406_, new_n407_,
    new_n408_, new_n409_, new_n410_, new_n411_, new_n412_, new_n413_,
    new_n414_, new_n415_, new_n416_, new_n417_, new_n418_, new_n419_,
    new_n420_, new_n421_, new_n422_, new_n423_, new_n424_, new_n425_,
    new_n426_, new_n427_, new_n428_, new_n429_, new_n430_, new_n431_,
    new_n432_, new_n433_, new_n434_, new_n435_, new_n436_, new_n437_,
    new_n438_, new_n439_, new_n440_, new_n441_, new_n442_, new_n443_,
    new_n444_, new_n445_, new_n446_, new_n447_, new_n448_, new_n449_,
    new_n450_, new_n451_, new_n452_, new_n453_, new_n454_, new_n455_,
    new_n456_, new_n457_, new_n458_, new_n459_, new_n460_, new_n461_,
    new_n462_, new_n463_, new_n464_, new_n465_, new_n466_, new_n467_,
    new_n468_, new_n469_, new_n470_, new_n471_, new_n472_, new_n473_,
    new_n474_, new_n475_, new_n476_, new_n477_, new_n478_, new_n479_,
    new_n480_, new_n481_, new_n482_, new_n483_, new_n484_, new_n485_,
    new_n486_, new_n487_, new_n488_, new_n489_, new_n490_, new_n491_,
    new_n492_, new_n493_, new_n494_, new_n495_, new_n496_, new_n497_,
    new_n498_, new_n499_, new_n500_, new_n501_, new_n502_, new_n503_,
    new_n504_, new_n505_, new_n506_, new_n507_, new_n508_, new_n509_,
    new_n510_, new_n511_, new_n512_, new_n513_, new_n514_, new_n515_,
    new_n516_, new_n517_, new_n518_, new_n519_, new_n520_, new_n521_,
    new_n522_, new_n523_, new_n524_, new_n525_, new_n526_, new_n527_,
    new_n528_, new_n529_, new_n530_, new_n531_, new_n532_, new_n533_,
    new_n534_, new_n535_, new_n536_, new_n537_, new_n538_, new_n539_,
    new_n540_, new_n541_, new_n542_, new_n543_, new_n544_, new_n545_,
    new_n546_, new_n547_, new_n548_, new_n549_, new_n550_, new_n551_,
    new_n552_, new_n553_, new_n554_, new_n555_, new_n556_, new_n557_,
    new_n558_, new_n559_, new_n560_, new_n561_, new_n562_, new_n563_,
    new_n564_, new_n565_, new_n566_, new_n567_, new_n568_, new_n569_,
    new_n570_, new_n571_, new_n572_, new_n573_, new_n574_, new_n575_,
    new_n576_, new_n577_, new_n578_, new_n579_, new_n580_, new_n581_,
    new_n582_, new_n583_, new_n584_, new_n585_, new_n586_, new_n587_,
    new_n588_, new_n589_, new_n590_, new_n592_, new_n593_, new_n594_,
    new_n595_, new_n596_, new_n597_, new_n598_, new_n599_, new_n600_,
    new_n601_, new_n602_, new_n603_, new_n604_, new_n605_, new_n606_,
    new_n607_, new_n608_, new_n609_, new_n610_, new_n611_, new_n612_,
    new_n613_, new_n614_, new_n615_, new_n616_, new_n617_, new_n618_,
    new_n619_, new_n620_, new_n621_, new_n622_, new_n623_, new_n624_,
    new_n625_, new_n626_, new_n627_, new_n628_, new_n629_, new_n630_,
    new_n631_, new_n632_, new_n633_, new_n634_, new_n635_, new_n636_,
    new_n637_, new_n638_, new_n639_, new_n640_, new_n641_, new_n642_,
    new_n643_, new_n644_, new_n645_, new_n646_, new_n647_, new_n648_,
    new_n649_, new_n650_, new_n651_, new_n652_, new_n653_, new_n654_,
    new_n655_, new_n656_, new_n657_, new_n658_, new_n659_, new_n660_,
    new_n661_, new_n662_, new_n663_, new_n664_, new_n665_, new_n666_,
    new_n667_, new_n668_, new_n669_, new_n670_, new_n671_, new_n672_,
    new_n673_, new_n674_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n687_, new_n688_, new_n689_, new_n690_,
    new_n691_, new_n692_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n927_, new_n928_, new_n929_, new_n930_, new_n931_,
    new_n932_, new_n933_, new_n934_, new_n935_, new_n936_, new_n937_,
    new_n938_, new_n939_, new_n940_, new_n941_, new_n942_, new_n943_,
    new_n944_, new_n945_, new_n946_, new_n947_, new_n948_, new_n949_,
    new_n950_, new_n951_, new_n952_, new_n953_, new_n954_, new_n955_,
    new_n956_, new_n957_, new_n958_, new_n959_, new_n960_, new_n961_,
    new_n962_, new_n963_, new_n964_, new_n966_, new_n967_, new_n968_,
    new_n969_, new_n970_, new_n971_, new_n972_, new_n973_, new_n974_,
    new_n975_, new_n976_, new_n977_, new_n978_, new_n979_, new_n980_,
    new_n981_, new_n982_, new_n983_, new_n984_, new_n985_, new_n986_,
    new_n987_, new_n988_, new_n989_, new_n990_, new_n991_, new_n992_,
    new_n993_, new_n994_, new_n995_, new_n996_, new_n997_, new_n998_,
    new_n999_, new_n1000_, new_n1001_, new_n1002_, new_n1003_, new_n1004_,
    new_n1005_, new_n1006_, new_n1007_, new_n1008_, new_n1009_, new_n1010_,
    new_n1011_, new_n1012_, new_n1013_, new_n1014_, new_n1015_, new_n1016_,
    new_n1017_, new_n1018_, new_n1019_, new_n1020_, new_n1021_, new_n1022_,
    new_n1023_, new_n1024_, new_n1025_, new_n1026_, new_n1027_, new_n1028_,
    new_n1029_, new_n1030_, new_n1031_, new_n1032_, new_n1033_, new_n1034_,
    new_n1035_, new_n1036_, new_n1037_, new_n1038_, new_n1039_, new_n1040_,
    new_n1041_, new_n1042_, new_n1043_, new_n1044_, new_n1045_, new_n1046_,
    new_n1047_, new_n1048_, new_n1049_, new_n1050_, new_n1051_, new_n1052_,
    new_n1053_, new_n1054_, new_n1055_, new_n1056_, new_n1057_, new_n1058_,
    new_n1059_, new_n1060_, new_n1061_, new_n1062_, new_n1063_, new_n1064_,
    new_n1065_, new_n1066_, new_n1067_, new_n1068_, new_n1069_, new_n1070_,
    new_n1071_, new_n1072_, new_n1073_, new_n1074_, new_n1075_, new_n1076_,
    new_n1077_, new_n1078_, new_n1079_, new_n1080_, new_n1081_, new_n1082_,
    new_n1083_, new_n1084_, new_n1085_, new_n1086_, new_n1087_, new_n1088_,
    new_n1089_, new_n1090_, new_n1091_, new_n1092_, new_n1093_, new_n1094_,
    new_n1095_, new_n1096_, new_n1097_, new_n1098_, new_n1099_, new_n1100_,
    new_n1101_, new_n1102_, new_n1103_, new_n1104_, new_n1105_, new_n1106_,
    new_n1107_, new_n1108_, new_n1109_, new_n1110_, new_n1111_, new_n1112_,
    new_n1113_, new_n1114_, new_n1115_, new_n1116_, new_n1117_, new_n1118_,
    new_n1119_, new_n1120_, new_n1121_, new_n1122_, new_n1123_, new_n1124_,
    new_n1125_, new_n1126_, new_n1127_, new_n1128_, new_n1129_, new_n1130_,
    new_n1131_, new_n1132_, new_n1133_, new_n1134_, new_n1135_, new_n1136_,
    new_n1137_, new_n1138_, new_n1139_, new_n1140_, new_n1141_, new_n1142_,
    new_n1143_, new_n1144_, new_n1145_, new_n1146_, new_n1147_, new_n1148_,
    new_n1149_, new_n1150_, new_n1151_, new_n1153_, new_n1154_, new_n1155_,
    new_n1156_, new_n1157_, new_n1158_, new_n1159_, new_n1160_, new_n1161_,
    new_n1162_, new_n1163_, new_n1164_, new_n1165_, new_n1166_, new_n1167_,
    new_n1168_, new_n1169_, new_n1170_, new_n1171_, new_n1172_, new_n1173_,
    new_n1174_, new_n1175_, new_n1176_, new_n1177_, new_n1178_, new_n1180_,
    new_n1181_, new_n1182_, new_n1183_, new_n1184_, new_n1185_, new_n1186_,
    new_n1187_, new_n1188_, new_n1189_, new_n1190_, new_n1191_, new_n1192_,
    new_n1193_, new_n1194_, new_n1195_, new_n1196_, new_n1197_, new_n1198_,
    new_n1199_, new_n1200_, new_n1201_, new_n1202_, new_n1203_, new_n1204_,
    new_n1205_, new_n1207_, new_n1208_, new_n1209_, new_n1210_, new_n1211_,
    new_n1212_, new_n1213_, new_n1214_, new_n1215_, new_n1216_, new_n1217_,
    new_n1218_, new_n1219_, new_n1220_, new_n1221_, new_n1222_, new_n1223_,
    new_n1224_, new_n1225_, new_n1226_, new_n1227_, new_n1228_, new_n1229_,
    new_n1230_, new_n1231_, new_n1232_, new_n1234_, new_n1235_, new_n1236_,
    new_n1237_, new_n1238_, new_n1239_, new_n1240_, new_n1241_, new_n1242_,
    new_n1243_, new_n1244_, new_n1245_, new_n1246_, new_n1247_, new_n1248_,
    new_n1249_, new_n1250_, new_n1251_, new_n1252_, new_n1253_, new_n1254_,
    new_n1255_, new_n1256_, new_n1257_, new_n1258_, new_n1259_, new_n1261_,
    new_n1262_, new_n1263_, new_n1264_, new_n1265_, new_n1266_, new_n1267_,
    new_n1268_, new_n1269_, new_n1270_, new_n1271_, new_n1272_, new_n1273_,
    new_n1274_, new_n1275_, new_n1276_, new_n1277_, new_n1278_, new_n1279_,
    new_n1280_, new_n1281_, new_n1282_, new_n1283_, new_n1284_, new_n1285_,
    new_n1286_, new_n1288_, new_n1289_, new_n1290_, new_n1291_, new_n1292_,
    new_n1293_, new_n1294_, new_n1295_, new_n1296_, new_n1297_, new_n1298_,
    new_n1299_, new_n1300_, new_n1301_, new_n1302_, new_n1303_, new_n1304_,
    new_n1305_, new_n1306_, new_n1307_, new_n1308_, new_n1309_, new_n1310_,
    new_n1311_, new_n1312_, new_n1313_, new_n1315_, new_n1316_, new_n1317_,
    new_n1318_, new_n1319_, new_n1320_, new_n1321_, new_n1322_, new_n1323_,
    new_n1324_, new_n1325_, new_n1326_, new_n1327_, new_n1328_, new_n1329_,
    new_n1330_, new_n1331_, new_n1332_, new_n1333_, new_n1334_, new_n1335_,
    new_n1336_, new_n1337_, new_n1338_, new_n1339_, new_n1340_, new_n1342_,
    new_n1343_, new_n1344_, new_n1345_, new_n1346_, new_n1347_, new_n1348_,
    new_n1349_, new_n1350_, new_n1351_, new_n1352_, new_n1353_, new_n1354_,
    new_n1355_, new_n1356_, new_n1357_, new_n1358_, new_n1359_, new_n1360_,
    new_n1361_, new_n1362_, new_n1363_, new_n1364_, new_n1365_, new_n1366_,
    new_n1367_, new_n1369_, new_n1370_, new_n1371_, new_n1372_, new_n1373_,
    new_n1374_, new_n1375_, new_n1376_, new_n1377_, new_n1378_, new_n1379_,
    new_n1380_, new_n1381_, new_n1382_, new_n1383_, new_n1384_, new_n1385_,
    new_n1386_, new_n1387_, new_n1388_, new_n1389_, new_n1390_, new_n1391_,
    new_n1392_, new_n1393_, new_n1394_, new_n1396_, new_n1397_, new_n1398_,
    new_n1399_, new_n1400_, new_n1401_, new_n1402_, new_n1403_, new_n1404_,
    new_n1405_, new_n1406_, new_n1407_, new_n1408_, new_n1409_, new_n1410_,
    new_n1411_, new_n1412_, new_n1413_, new_n1414_, new_n1415_, new_n1416_,
    new_n1417_, new_n1418_, new_n1419_, new_n1420_, new_n1421_, new_n1423_,
    new_n1424_, new_n1425_, new_n1426_, new_n1427_, new_n1428_, new_n1429_,
    new_n1430_, new_n1431_, new_n1432_, new_n1433_, new_n1434_, new_n1435_,
    new_n1436_, new_n1437_, new_n1438_, new_n1439_, new_n1440_, new_n1441_,
    new_n1442_, new_n1443_, new_n1444_, new_n1445_, new_n1446_, new_n1447_,
    new_n1448_, new_n1450_, new_n1451_, new_n1452_, new_n1453_, new_n1454_,
    new_n1455_, new_n1456_, new_n1457_, new_n1458_, new_n1459_, new_n1460_,
    new_n1461_, new_n1462_, new_n1463_, new_n1464_, new_n1465_, new_n1466_,
    new_n1467_, new_n1468_, new_n1469_, new_n1470_, new_n1471_, new_n1472_,
    new_n1473_, new_n1474_, new_n1475_, new_n1477_, new_n1478_, new_n1479_,
    new_n1480_, new_n1481_, new_n1482_, new_n1483_, new_n1484_, new_n1485_,
    new_n1486_, new_n1488_, new_n1489_, new_n1490_, new_n1491_, new_n1492_,
    new_n1493_, new_n1494_, new_n1495_, new_n1496_, new_n1497_, new_n1499_,
    new_n1500_, new_n1501_, new_n1502_, new_n1503_, new_n1504_, new_n1505_,
    new_n1506_, new_n1507_, new_n1508_, new_n1510_, new_n1511_, new_n1512_,
    new_n1513_, new_n1514_, new_n1515_, new_n1516_, new_n1517_, new_n1518_,
    new_n1519_, new_n1521_, new_n1522_, new_n1523_, new_n1524_, new_n1525_,
    new_n1526_, new_n1527_, new_n1528_, new_n1529_, new_n1530_, new_n1532_,
    new_n1533_, new_n1534_, new_n1535_, new_n1536_, new_n1537_, new_n1538_,
    new_n1539_, new_n1540_, new_n1541_, new_n1543_, new_n1544_, new_n1545_,
    new_n1546_, new_n1547_, new_n1548_, new_n1549_, new_n1550_, new_n1551_,
    new_n1552_, new_n1554_, new_n1555_, new_n1556_, new_n1557_, new_n1558_,
    new_n1559_, new_n1560_, new_n1561_, new_n1562_, new_n1563_, new_n1565_,
    new_n1566_, new_n1567_, new_n1568_, new_n1569_, new_n1570_, new_n1571_,
    new_n1572_, new_n1573_, new_n1574_, new_n1576_, new_n1577_, new_n1578_,
    new_n1579_, new_n1580_, new_n1581_, new_n1582_, new_n1583_, new_n1584_,
    new_n1585_, new_n1587_, new_n1588_, new_n1589_, new_n1590_, new_n1591_,
    new_n1592_, new_n1593_, new_n1594_, new_n1595_, new_n1596_, new_n1598_,
    new_n1599_, new_n1600_, new_n1601_, new_n1602_, new_n1603_, new_n1604_,
    new_n1605_, new_n1606_, new_n1607_, new_n1609_, new_n1610_, new_n1611_,
    new_n1612_, new_n1613_, new_n1614_, new_n1615_, new_n1616_, new_n1617_,
    new_n1618_, new_n1620_, new_n1621_, new_n1622_, new_n1623_, new_n1624_,
    new_n1625_, new_n1626_, new_n1627_, new_n1628_, new_n1629_, new_n1631_,
    new_n1632_, new_n1633_, new_n1634_, new_n1635_, new_n1636_, new_n1637_,
    new_n1638_, new_n1639_, new_n1640_, new_n1642_, new_n1643_, new_n1644_,
    new_n1645_, new_n1646_, new_n1647_, new_n1648_, new_n1649_, new_n1650_,
    new_n1651_, new_n1653_, new_n1654_, new_n1655_, new_n1656_, new_n1657_,
    new_n1658_, new_n1659_, new_n1660_, new_n1661_, new_n1662_, new_n1664_,
    new_n1665_, new_n1666_, new_n1667_, new_n1668_, new_n1669_, new_n1670_,
    new_n1671_, new_n1672_, new_n1673_, new_n1675_, new_n1676_, new_n1677_,
    new_n1678_, new_n1679_, new_n1680_, new_n1681_, new_n1682_, new_n1683_,
    new_n1684_, new_n1686_, new_n1687_, new_n1688_, new_n1689_, new_n1690_,
    new_n1691_, new_n1692_, new_n1693_, new_n1694_, new_n1695_, new_n1697_,
    new_n1698_, new_n1699_, new_n1700_, new_n1701_, new_n1702_, new_n1703_,
    new_n1704_, new_n1705_, new_n1706_, new_n1708_, new_n1709_, new_n1710_,
    new_n1711_, new_n1712_, new_n1713_, new_n1714_, new_n1715_, new_n1716_,
    new_n1717_, new_n1719_, new_n1720_, new_n1721_, new_n1722_, new_n1723_,
    new_n1724_, new_n1725_, new_n1726_, new_n1727_, new_n1728_, new_n1730_,
    new_n1731_, new_n1732_, new_n1733_, new_n1734_, new_n1735_, new_n1736_,
    new_n1737_, new_n1738_, new_n1739_, new_n1741_, new_n1742_, new_n1743_,
    new_n1744_, new_n1745_, new_n1746_, new_n1747_, new_n1748_, new_n1749_,
    new_n1750_, new_n1752_, new_n1753_, new_n1754_, new_n1755_, new_n1756_,
    new_n1757_, new_n1758_, new_n1759_, new_n1760_, new_n1761_, new_n1763_,
    new_n1764_, new_n1765_, new_n1766_, new_n1767_, new_n1768_, new_n1769_,
    new_n1770_, new_n1771_, new_n1772_, new_n1774_, new_n1775_, new_n1776_,
    new_n1777_, new_n1778_, new_n1779_, new_n1780_, new_n1781_, new_n1782_,
    new_n1783_, new_n1785_, new_n1786_, new_n1787_, new_n1788_, new_n1789_,
    new_n1790_, new_n1791_, new_n1792_, new_n1793_, new_n1794_, new_n1796_,
    new_n1797_, new_n1798_, new_n1799_, new_n1800_, new_n1801_, new_n1802_,
    new_n1803_, new_n1804_, new_n1805_, new_n1807_, new_n1808_, new_n1809_,
    new_n1810_, new_n1811_, new_n1812_, new_n1813_, new_n1814_, new_n1815_,
    new_n1816_, new_n1818_, new_n1819_, new_n1820_, new_n1821_, new_n1822_,
    new_n1823_, new_n1824_, new_n1825_, new_n1826_, new_n1827_, new_n1829_,
    new_n1830_, new_n1831_, new_n1832_, new_n1833_, new_n1834_, new_n1835_,
    new_n1836_, new_n1837_, new_n1838_, new_n1840_, new_n1841_, new_n1842_,
    new_n1843_, new_n1844_, new_n1845_, new_n1846_, new_n1847_, new_n1848_,
    new_n1849_, new_n1851_, new_n1852_, new_n1853_, new_n1854_, new_n1855_,
    new_n1856_, new_n1857_, new_n1858_, new_n1859_, new_n1860_, new_n1862_,
    new_n1863_, new_n1864_, new_n1865_, new_n1866_, new_n1867_, new_n1868_,
    new_n1869_, new_n1870_, new_n1871_, new_n1873_, new_n1874_, new_n1875_,
    new_n1876_, new_n1877_, new_n1878_, new_n1879_, new_n1880_, new_n1881_,
    new_n1882_, new_n1884_, new_n1885_, new_n1886_, new_n1887_, new_n1888_,
    new_n1889_, new_n1890_, new_n1891_, new_n1892_, new_n1893_, new_n1895_,
    new_n1896_, new_n1897_, new_n1898_, new_n1899_, new_n1900_, new_n1901_,
    new_n1902_, new_n1903_, new_n1904_, new_n1906_, new_n1907_, new_n1908_,
    new_n1909_, new_n1910_, new_n1911_, new_n1912_, new_n1913_, new_n1914_,
    new_n1915_, new_n1917_, new_n1918_, new_n1919_, new_n1920_, new_n1921_,
    new_n1922_, new_n1923_, new_n1924_, new_n1925_, new_n1926_, new_n1928_,
    new_n1929_, new_n1930_, new_n1931_, new_n1932_, new_n1933_, new_n1934_,
    new_n1935_, new_n1936_, new_n1937_, new_n1939_, new_n1940_, new_n1941_,
    new_n1942_, new_n1943_, new_n1944_, new_n1945_, new_n1946_, new_n1947_,
    new_n1948_, new_n1950_, new_n1951_, new_n1952_, new_n1953_, new_n1954_,
    new_n1955_, new_n1956_, new_n1957_, new_n1958_, new_n1959_, new_n1961_,
    new_n1962_, new_n1963_, new_n1964_, new_n1965_, new_n1966_, new_n1967_,
    new_n1968_, new_n1969_, new_n1970_, new_n1972_, new_n1973_, new_n1974_,
    new_n1975_, new_n1976_, new_n1977_, new_n1978_, new_n1979_, new_n1980_,
    new_n1981_, new_n1983_, new_n1984_, new_n1985_, new_n1986_, new_n1987_,
    new_n1988_, new_n1989_, new_n1990_, new_n1991_, new_n1992_, new_n1994_,
    new_n1995_, new_n1996_, new_n1997_, new_n1998_, new_n1999_, new_n2000_,
    new_n2001_, new_n2002_, new_n2003_;
  INVX1    g0000(.A(\shift[6] ), .Y(new_n264_));
  INVX1    g0001(.A(\a[77] ), .Y(new_n265_));
  INVX1    g0002(.A(\shift[0] ), .Y(new_n266_));
  INVX1    g0003(.A(\shift[1] ), .Y(new_n267_));
  NOR3X1   g0004(.A(new_n267_), .B(new_n266_), .C(new_n265_), .Y(new_n268_));
  INVX1    g0005(.A(\a[78] ), .Y(new_n269_));
  NOR3X1   g0006(.A(new_n267_), .B(\shift[0] ), .C(new_n269_), .Y(new_n270_));
  INVX1    g0007(.A(\a[80] ), .Y(new_n271_));
  NOR3X1   g0008(.A(\shift[1] ), .B(\shift[0] ), .C(new_n271_), .Y(new_n272_));
  INVX1    g0009(.A(\a[79] ), .Y(new_n273_));
  NOR3X1   g0010(.A(\shift[1] ), .B(new_n266_), .C(new_n273_), .Y(new_n274_));
  OR4X1    g0011(.A(new_n274_), .B(new_n272_), .C(new_n270_), .D(new_n268_), .Y(new_n275_));
  NOR2X1   g0012(.A(\shift[3] ), .B(\shift[2] ), .Y(new_n276_));
  INVX1    g0013(.A(\a[73] ), .Y(new_n277_));
  NOR3X1   g0014(.A(new_n267_), .B(new_n266_), .C(new_n277_), .Y(new_n278_));
  INVX1    g0015(.A(\a[74] ), .Y(new_n279_));
  NOR3X1   g0016(.A(new_n267_), .B(\shift[0] ), .C(new_n279_), .Y(new_n280_));
  INVX1    g0017(.A(\a[76] ), .Y(new_n281_));
  NOR3X1   g0018(.A(\shift[1] ), .B(\shift[0] ), .C(new_n281_), .Y(new_n282_));
  INVX1    g0019(.A(\a[75] ), .Y(new_n283_));
  NOR3X1   g0020(.A(\shift[1] ), .B(new_n266_), .C(new_n283_), .Y(new_n284_));
  OR4X1    g0021(.A(new_n284_), .B(new_n282_), .C(new_n280_), .D(new_n278_), .Y(new_n285_));
  INVX1    g0022(.A(\shift[2] ), .Y(new_n286_));
  NOR2X1   g0023(.A(\shift[3] ), .B(new_n286_), .Y(new_n287_));
  AOI22X1  g0024(.A0(new_n287_), .A1(new_n285_), .B0(new_n276_), .B1(new_n275_), .Y(new_n288_));
  INVX1    g0025(.A(\a[65] ), .Y(new_n289_));
  NOR3X1   g0026(.A(new_n267_), .B(new_n266_), .C(new_n289_), .Y(new_n290_));
  INVX1    g0027(.A(\a[66] ), .Y(new_n291_));
  NOR3X1   g0028(.A(new_n267_), .B(\shift[0] ), .C(new_n291_), .Y(new_n292_));
  INVX1    g0029(.A(\a[68] ), .Y(new_n293_));
  NOR3X1   g0030(.A(\shift[1] ), .B(\shift[0] ), .C(new_n293_), .Y(new_n294_));
  INVX1    g0031(.A(\a[67] ), .Y(new_n295_));
  NOR3X1   g0032(.A(\shift[1] ), .B(new_n266_), .C(new_n295_), .Y(new_n296_));
  OR4X1    g0033(.A(new_n296_), .B(new_n294_), .C(new_n292_), .D(new_n290_), .Y(new_n297_));
  AND2X1   g0034(.A(\shift[3] ), .B(\shift[2] ), .Y(new_n298_));
  INVX1    g0035(.A(\a[69] ), .Y(new_n299_));
  NOR3X1   g0036(.A(new_n267_), .B(new_n266_), .C(new_n299_), .Y(new_n300_));
  INVX1    g0037(.A(\a[70] ), .Y(new_n301_));
  NOR3X1   g0038(.A(new_n267_), .B(\shift[0] ), .C(new_n301_), .Y(new_n302_));
  INVX1    g0039(.A(\a[72] ), .Y(new_n303_));
  NOR3X1   g0040(.A(\shift[1] ), .B(\shift[0] ), .C(new_n303_), .Y(new_n304_));
  INVX1    g0041(.A(\a[71] ), .Y(new_n305_));
  NOR3X1   g0042(.A(\shift[1] ), .B(new_n266_), .C(new_n305_), .Y(new_n306_));
  OR4X1    g0043(.A(new_n306_), .B(new_n304_), .C(new_n302_), .D(new_n300_), .Y(new_n307_));
  AND2X1   g0044(.A(\shift[3] ), .B(new_n286_), .Y(new_n308_));
  AOI22X1  g0045(.A0(new_n308_), .A1(new_n307_), .B0(new_n298_), .B1(new_n297_), .Y(new_n309_));
  NAND2X1  g0046(.A(\shift[5] ), .B(\shift[4] ), .Y(new_n310_));
  AOI21X1  g0047(.A0(new_n309_), .A1(new_n288_), .B0(new_n310_), .Y(new_n311_));
  INVX1    g0048(.A(\a[93] ), .Y(new_n312_));
  NOR3X1   g0049(.A(new_n267_), .B(new_n266_), .C(new_n312_), .Y(new_n313_));
  INVX1    g0050(.A(\a[94] ), .Y(new_n314_));
  NOR3X1   g0051(.A(new_n267_), .B(\shift[0] ), .C(new_n314_), .Y(new_n315_));
  INVX1    g0052(.A(\a[96] ), .Y(new_n316_));
  NOR3X1   g0053(.A(\shift[1] ), .B(\shift[0] ), .C(new_n316_), .Y(new_n317_));
  INVX1    g0054(.A(\a[95] ), .Y(new_n318_));
  NOR3X1   g0055(.A(\shift[1] ), .B(new_n266_), .C(new_n318_), .Y(new_n319_));
  OR4X1    g0056(.A(new_n319_), .B(new_n317_), .C(new_n315_), .D(new_n313_), .Y(new_n320_));
  INVX1    g0057(.A(\a[89] ), .Y(new_n321_));
  NOR3X1   g0058(.A(new_n267_), .B(new_n266_), .C(new_n321_), .Y(new_n322_));
  INVX1    g0059(.A(\a[90] ), .Y(new_n323_));
  NOR3X1   g0060(.A(new_n267_), .B(\shift[0] ), .C(new_n323_), .Y(new_n324_));
  INVX1    g0061(.A(\a[92] ), .Y(new_n325_));
  NOR3X1   g0062(.A(\shift[1] ), .B(\shift[0] ), .C(new_n325_), .Y(new_n326_));
  INVX1    g0063(.A(\a[91] ), .Y(new_n327_));
  NOR3X1   g0064(.A(\shift[1] ), .B(new_n266_), .C(new_n327_), .Y(new_n328_));
  OR4X1    g0065(.A(new_n328_), .B(new_n326_), .C(new_n324_), .D(new_n322_), .Y(new_n329_));
  AOI22X1  g0066(.A0(new_n329_), .A1(new_n287_), .B0(new_n320_), .B1(new_n276_), .Y(new_n330_));
  INVX1    g0067(.A(\a[81] ), .Y(new_n331_));
  NOR3X1   g0068(.A(new_n267_), .B(new_n266_), .C(new_n331_), .Y(new_n332_));
  INVX1    g0069(.A(\a[82] ), .Y(new_n333_));
  NOR3X1   g0070(.A(new_n267_), .B(\shift[0] ), .C(new_n333_), .Y(new_n334_));
  INVX1    g0071(.A(\a[84] ), .Y(new_n335_));
  NOR3X1   g0072(.A(\shift[1] ), .B(\shift[0] ), .C(new_n335_), .Y(new_n336_));
  INVX1    g0073(.A(\a[83] ), .Y(new_n337_));
  NOR3X1   g0074(.A(\shift[1] ), .B(new_n266_), .C(new_n337_), .Y(new_n338_));
  OR4X1    g0075(.A(new_n338_), .B(new_n336_), .C(new_n334_), .D(new_n332_), .Y(new_n339_));
  INVX1    g0076(.A(\a[85] ), .Y(new_n340_));
  NOR3X1   g0077(.A(new_n267_), .B(new_n266_), .C(new_n340_), .Y(new_n341_));
  INVX1    g0078(.A(\a[86] ), .Y(new_n342_));
  NOR3X1   g0079(.A(new_n267_), .B(\shift[0] ), .C(new_n342_), .Y(new_n343_));
  INVX1    g0080(.A(\a[88] ), .Y(new_n344_));
  NOR3X1   g0081(.A(\shift[1] ), .B(\shift[0] ), .C(new_n344_), .Y(new_n345_));
  INVX1    g0082(.A(\a[87] ), .Y(new_n346_));
  NOR3X1   g0083(.A(\shift[1] ), .B(new_n266_), .C(new_n346_), .Y(new_n347_));
  OR4X1    g0084(.A(new_n347_), .B(new_n345_), .C(new_n343_), .D(new_n341_), .Y(new_n348_));
  AOI22X1  g0085(.A0(new_n348_), .A1(new_n308_), .B0(new_n339_), .B1(new_n298_), .Y(new_n349_));
  INVX1    g0086(.A(\shift[4] ), .Y(new_n350_));
  NAND2X1  g0087(.A(\shift[5] ), .B(new_n350_), .Y(new_n351_));
  AOI21X1  g0088(.A0(new_n349_), .A1(new_n330_), .B0(new_n351_), .Y(new_n352_));
  INVX1    g0089(.A(\a[125] ), .Y(new_n353_));
  NOR3X1   g0090(.A(new_n267_), .B(new_n266_), .C(new_n353_), .Y(new_n354_));
  INVX1    g0091(.A(\a[126] ), .Y(new_n355_));
  NOR3X1   g0092(.A(new_n267_), .B(\shift[0] ), .C(new_n355_), .Y(new_n356_));
  INVX1    g0093(.A(\a[0] ), .Y(new_n357_));
  NOR3X1   g0094(.A(\shift[1] ), .B(\shift[0] ), .C(new_n357_), .Y(new_n358_));
  INVX1    g0095(.A(\a[127] ), .Y(new_n359_));
  NOR3X1   g0096(.A(\shift[1] ), .B(new_n266_), .C(new_n359_), .Y(new_n360_));
  OR4X1    g0097(.A(new_n360_), .B(new_n358_), .C(new_n356_), .D(new_n354_), .Y(new_n361_));
  INVX1    g0098(.A(\a[121] ), .Y(new_n362_));
  NOR3X1   g0099(.A(new_n267_), .B(new_n266_), .C(new_n362_), .Y(new_n363_));
  INVX1    g0100(.A(\a[122] ), .Y(new_n364_));
  NOR3X1   g0101(.A(new_n267_), .B(\shift[0] ), .C(new_n364_), .Y(new_n365_));
  INVX1    g0102(.A(\a[124] ), .Y(new_n366_));
  NOR3X1   g0103(.A(\shift[1] ), .B(\shift[0] ), .C(new_n366_), .Y(new_n367_));
  INVX1    g0104(.A(\a[123] ), .Y(new_n368_));
  NOR3X1   g0105(.A(\shift[1] ), .B(new_n266_), .C(new_n368_), .Y(new_n369_));
  OR4X1    g0106(.A(new_n369_), .B(new_n367_), .C(new_n365_), .D(new_n363_), .Y(new_n370_));
  AOI22X1  g0107(.A0(new_n370_), .A1(new_n287_), .B0(new_n361_), .B1(new_n276_), .Y(new_n371_));
  INVX1    g0108(.A(\a[113] ), .Y(new_n372_));
  NOR3X1   g0109(.A(new_n267_), .B(new_n266_), .C(new_n372_), .Y(new_n373_));
  INVX1    g0110(.A(\a[114] ), .Y(new_n374_));
  NOR3X1   g0111(.A(new_n267_), .B(\shift[0] ), .C(new_n374_), .Y(new_n375_));
  INVX1    g0112(.A(\a[116] ), .Y(new_n376_));
  NOR3X1   g0113(.A(\shift[1] ), .B(\shift[0] ), .C(new_n376_), .Y(new_n377_));
  INVX1    g0114(.A(\a[115] ), .Y(new_n378_));
  NOR3X1   g0115(.A(\shift[1] ), .B(new_n266_), .C(new_n378_), .Y(new_n379_));
  OR4X1    g0116(.A(new_n379_), .B(new_n377_), .C(new_n375_), .D(new_n373_), .Y(new_n380_));
  INVX1    g0117(.A(\a[117] ), .Y(new_n381_));
  NOR3X1   g0118(.A(new_n267_), .B(new_n266_), .C(new_n381_), .Y(new_n382_));
  INVX1    g0119(.A(\a[118] ), .Y(new_n383_));
  NOR3X1   g0120(.A(new_n267_), .B(\shift[0] ), .C(new_n383_), .Y(new_n384_));
  INVX1    g0121(.A(\a[120] ), .Y(new_n385_));
  NOR3X1   g0122(.A(\shift[1] ), .B(\shift[0] ), .C(new_n385_), .Y(new_n386_));
  INVX1    g0123(.A(\a[119] ), .Y(new_n387_));
  NOR3X1   g0124(.A(\shift[1] ), .B(new_n266_), .C(new_n387_), .Y(new_n388_));
  OR4X1    g0125(.A(new_n388_), .B(new_n386_), .C(new_n384_), .D(new_n382_), .Y(new_n389_));
  AOI22X1  g0126(.A0(new_n389_), .A1(new_n308_), .B0(new_n380_), .B1(new_n298_), .Y(new_n390_));
  OR2X1    g0127(.A(\shift[5] ), .B(\shift[4] ), .Y(new_n391_));
  AOI21X1  g0128(.A0(new_n390_), .A1(new_n371_), .B0(new_n391_), .Y(new_n392_));
  INVX1    g0129(.A(\a[109] ), .Y(new_n393_));
  NOR3X1   g0130(.A(new_n267_), .B(new_n266_), .C(new_n393_), .Y(new_n394_));
  INVX1    g0131(.A(\a[110] ), .Y(new_n395_));
  NOR3X1   g0132(.A(new_n267_), .B(\shift[0] ), .C(new_n395_), .Y(new_n396_));
  INVX1    g0133(.A(\a[112] ), .Y(new_n397_));
  NOR3X1   g0134(.A(\shift[1] ), .B(\shift[0] ), .C(new_n397_), .Y(new_n398_));
  INVX1    g0135(.A(\a[111] ), .Y(new_n399_));
  NOR3X1   g0136(.A(\shift[1] ), .B(new_n266_), .C(new_n399_), .Y(new_n400_));
  OR4X1    g0137(.A(new_n400_), .B(new_n398_), .C(new_n396_), .D(new_n394_), .Y(new_n401_));
  INVX1    g0138(.A(\a[105] ), .Y(new_n402_));
  NOR3X1   g0139(.A(new_n267_), .B(new_n266_), .C(new_n402_), .Y(new_n403_));
  INVX1    g0140(.A(\a[106] ), .Y(new_n404_));
  NOR3X1   g0141(.A(new_n267_), .B(\shift[0] ), .C(new_n404_), .Y(new_n405_));
  INVX1    g0142(.A(\a[108] ), .Y(new_n406_));
  NOR3X1   g0143(.A(\shift[1] ), .B(\shift[0] ), .C(new_n406_), .Y(new_n407_));
  INVX1    g0144(.A(\a[107] ), .Y(new_n408_));
  NOR3X1   g0145(.A(\shift[1] ), .B(new_n266_), .C(new_n408_), .Y(new_n409_));
  OR4X1    g0146(.A(new_n409_), .B(new_n407_), .C(new_n405_), .D(new_n403_), .Y(new_n410_));
  AOI22X1  g0147(.A0(new_n410_), .A1(new_n287_), .B0(new_n401_), .B1(new_n276_), .Y(new_n411_));
  INVX1    g0148(.A(\a[97] ), .Y(new_n412_));
  NOR3X1   g0149(.A(new_n267_), .B(new_n266_), .C(new_n412_), .Y(new_n413_));
  INVX1    g0150(.A(\a[98] ), .Y(new_n414_));
  NOR3X1   g0151(.A(new_n267_), .B(\shift[0] ), .C(new_n414_), .Y(new_n415_));
  INVX1    g0152(.A(\a[100] ), .Y(new_n416_));
  NOR3X1   g0153(.A(\shift[1] ), .B(\shift[0] ), .C(new_n416_), .Y(new_n417_));
  INVX1    g0154(.A(\a[99] ), .Y(new_n418_));
  NOR3X1   g0155(.A(\shift[1] ), .B(new_n266_), .C(new_n418_), .Y(new_n419_));
  OR4X1    g0156(.A(new_n419_), .B(new_n417_), .C(new_n415_), .D(new_n413_), .Y(new_n420_));
  INVX1    g0157(.A(\a[101] ), .Y(new_n421_));
  NOR3X1   g0158(.A(new_n267_), .B(new_n266_), .C(new_n421_), .Y(new_n422_));
  INVX1    g0159(.A(\a[102] ), .Y(new_n423_));
  NOR3X1   g0160(.A(new_n267_), .B(\shift[0] ), .C(new_n423_), .Y(new_n424_));
  INVX1    g0161(.A(\a[104] ), .Y(new_n425_));
  NOR3X1   g0162(.A(\shift[1] ), .B(\shift[0] ), .C(new_n425_), .Y(new_n426_));
  INVX1    g0163(.A(\a[103] ), .Y(new_n427_));
  NOR3X1   g0164(.A(\shift[1] ), .B(new_n266_), .C(new_n427_), .Y(new_n428_));
  OR4X1    g0165(.A(new_n428_), .B(new_n426_), .C(new_n424_), .D(new_n422_), .Y(new_n429_));
  AOI22X1  g0166(.A0(new_n429_), .A1(new_n308_), .B0(new_n420_), .B1(new_n298_), .Y(new_n430_));
  OR2X1    g0167(.A(\shift[5] ), .B(new_n350_), .Y(new_n431_));
  AOI21X1  g0168(.A0(new_n430_), .A1(new_n411_), .B0(new_n431_), .Y(new_n432_));
  OR4X1    g0169(.A(new_n432_), .B(new_n392_), .C(new_n352_), .D(new_n311_), .Y(new_n433_));
  INVX1    g0170(.A(\a[13] ), .Y(new_n434_));
  NOR3X1   g0171(.A(new_n267_), .B(new_n266_), .C(new_n434_), .Y(new_n435_));
  INVX1    g0172(.A(\a[14] ), .Y(new_n436_));
  NOR3X1   g0173(.A(new_n267_), .B(\shift[0] ), .C(new_n436_), .Y(new_n437_));
  INVX1    g0174(.A(\a[16] ), .Y(new_n438_));
  NOR3X1   g0175(.A(\shift[1] ), .B(\shift[0] ), .C(new_n438_), .Y(new_n439_));
  INVX1    g0176(.A(\a[15] ), .Y(new_n440_));
  NOR3X1   g0177(.A(\shift[1] ), .B(new_n266_), .C(new_n440_), .Y(new_n441_));
  OR4X1    g0178(.A(new_n441_), .B(new_n439_), .C(new_n437_), .D(new_n435_), .Y(new_n442_));
  INVX1    g0179(.A(\a[9] ), .Y(new_n443_));
  NOR3X1   g0180(.A(new_n267_), .B(new_n266_), .C(new_n443_), .Y(new_n444_));
  INVX1    g0181(.A(\a[10] ), .Y(new_n445_));
  NOR3X1   g0182(.A(new_n267_), .B(\shift[0] ), .C(new_n445_), .Y(new_n446_));
  INVX1    g0183(.A(\a[12] ), .Y(new_n447_));
  NOR3X1   g0184(.A(\shift[1] ), .B(\shift[0] ), .C(new_n447_), .Y(new_n448_));
  INVX1    g0185(.A(\a[11] ), .Y(new_n449_));
  NOR3X1   g0186(.A(\shift[1] ), .B(new_n266_), .C(new_n449_), .Y(new_n450_));
  OR4X1    g0187(.A(new_n450_), .B(new_n448_), .C(new_n446_), .D(new_n444_), .Y(new_n451_));
  AOI22X1  g0188(.A0(new_n451_), .A1(new_n287_), .B0(new_n442_), .B1(new_n276_), .Y(new_n452_));
  INVX1    g0189(.A(\a[1] ), .Y(new_n453_));
  NOR3X1   g0190(.A(new_n267_), .B(new_n266_), .C(new_n453_), .Y(new_n454_));
  INVX1    g0191(.A(\a[2] ), .Y(new_n455_));
  NOR3X1   g0192(.A(new_n267_), .B(\shift[0] ), .C(new_n455_), .Y(new_n456_));
  INVX1    g0193(.A(\a[4] ), .Y(new_n457_));
  NOR3X1   g0194(.A(\shift[1] ), .B(\shift[0] ), .C(new_n457_), .Y(new_n458_));
  INVX1    g0195(.A(\a[3] ), .Y(new_n459_));
  NOR3X1   g0196(.A(\shift[1] ), .B(new_n266_), .C(new_n459_), .Y(new_n460_));
  OR4X1    g0197(.A(new_n460_), .B(new_n458_), .C(new_n456_), .D(new_n454_), .Y(new_n461_));
  INVX1    g0198(.A(\a[5] ), .Y(new_n462_));
  NOR3X1   g0199(.A(new_n267_), .B(new_n266_), .C(new_n462_), .Y(new_n463_));
  INVX1    g0200(.A(\a[6] ), .Y(new_n464_));
  NOR3X1   g0201(.A(new_n267_), .B(\shift[0] ), .C(new_n464_), .Y(new_n465_));
  INVX1    g0202(.A(\a[8] ), .Y(new_n466_));
  NOR3X1   g0203(.A(\shift[1] ), .B(\shift[0] ), .C(new_n466_), .Y(new_n467_));
  INVX1    g0204(.A(\a[7] ), .Y(new_n468_));
  NOR3X1   g0205(.A(\shift[1] ), .B(new_n266_), .C(new_n468_), .Y(new_n469_));
  OR4X1    g0206(.A(new_n469_), .B(new_n467_), .C(new_n465_), .D(new_n463_), .Y(new_n470_));
  AOI22X1  g0207(.A0(new_n470_), .A1(new_n308_), .B0(new_n461_), .B1(new_n298_), .Y(new_n471_));
  AOI21X1  g0208(.A0(new_n471_), .A1(new_n452_), .B0(new_n310_), .Y(new_n472_));
  INVX1    g0209(.A(\a[29] ), .Y(new_n473_));
  NOR3X1   g0210(.A(new_n267_), .B(new_n266_), .C(new_n473_), .Y(new_n474_));
  INVX1    g0211(.A(\a[30] ), .Y(new_n475_));
  NOR3X1   g0212(.A(new_n267_), .B(\shift[0] ), .C(new_n475_), .Y(new_n476_));
  INVX1    g0213(.A(\a[32] ), .Y(new_n477_));
  NOR3X1   g0214(.A(\shift[1] ), .B(\shift[0] ), .C(new_n477_), .Y(new_n478_));
  INVX1    g0215(.A(\a[31] ), .Y(new_n479_));
  NOR3X1   g0216(.A(\shift[1] ), .B(new_n266_), .C(new_n479_), .Y(new_n480_));
  OR4X1    g0217(.A(new_n480_), .B(new_n478_), .C(new_n476_), .D(new_n474_), .Y(new_n481_));
  INVX1    g0218(.A(\a[25] ), .Y(new_n482_));
  NOR3X1   g0219(.A(new_n267_), .B(new_n266_), .C(new_n482_), .Y(new_n483_));
  INVX1    g0220(.A(\a[26] ), .Y(new_n484_));
  NOR3X1   g0221(.A(new_n267_), .B(\shift[0] ), .C(new_n484_), .Y(new_n485_));
  INVX1    g0222(.A(\a[28] ), .Y(new_n486_));
  NOR3X1   g0223(.A(\shift[1] ), .B(\shift[0] ), .C(new_n486_), .Y(new_n487_));
  INVX1    g0224(.A(\a[27] ), .Y(new_n488_));
  NOR3X1   g0225(.A(\shift[1] ), .B(new_n266_), .C(new_n488_), .Y(new_n489_));
  OR4X1    g0226(.A(new_n489_), .B(new_n487_), .C(new_n485_), .D(new_n483_), .Y(new_n490_));
  AOI22X1  g0227(.A0(new_n490_), .A1(new_n287_), .B0(new_n481_), .B1(new_n276_), .Y(new_n491_));
  INVX1    g0228(.A(\a[17] ), .Y(new_n492_));
  NOR3X1   g0229(.A(new_n267_), .B(new_n266_), .C(new_n492_), .Y(new_n493_));
  INVX1    g0230(.A(\a[18] ), .Y(new_n494_));
  NOR3X1   g0231(.A(new_n267_), .B(\shift[0] ), .C(new_n494_), .Y(new_n495_));
  INVX1    g0232(.A(\a[20] ), .Y(new_n496_));
  NOR3X1   g0233(.A(\shift[1] ), .B(\shift[0] ), .C(new_n496_), .Y(new_n497_));
  INVX1    g0234(.A(\a[19] ), .Y(new_n498_));
  NOR3X1   g0235(.A(\shift[1] ), .B(new_n266_), .C(new_n498_), .Y(new_n499_));
  OR4X1    g0236(.A(new_n499_), .B(new_n497_), .C(new_n495_), .D(new_n493_), .Y(new_n500_));
  INVX1    g0237(.A(\a[21] ), .Y(new_n501_));
  NOR3X1   g0238(.A(new_n267_), .B(new_n266_), .C(new_n501_), .Y(new_n502_));
  INVX1    g0239(.A(\a[22] ), .Y(new_n503_));
  NOR3X1   g0240(.A(new_n267_), .B(\shift[0] ), .C(new_n503_), .Y(new_n504_));
  INVX1    g0241(.A(\a[24] ), .Y(new_n505_));
  NOR3X1   g0242(.A(\shift[1] ), .B(\shift[0] ), .C(new_n505_), .Y(new_n506_));
  INVX1    g0243(.A(\a[23] ), .Y(new_n507_));
  NOR3X1   g0244(.A(\shift[1] ), .B(new_n266_), .C(new_n507_), .Y(new_n508_));
  OR4X1    g0245(.A(new_n508_), .B(new_n506_), .C(new_n504_), .D(new_n502_), .Y(new_n509_));
  AOI22X1  g0246(.A0(new_n509_), .A1(new_n308_), .B0(new_n500_), .B1(new_n298_), .Y(new_n510_));
  AOI21X1  g0247(.A0(new_n510_), .A1(new_n491_), .B0(new_n351_), .Y(new_n511_));
  INVX1    g0248(.A(\a[61] ), .Y(new_n512_));
  NOR3X1   g0249(.A(new_n267_), .B(new_n266_), .C(new_n512_), .Y(new_n513_));
  INVX1    g0250(.A(\a[62] ), .Y(new_n514_));
  NOR3X1   g0251(.A(new_n267_), .B(\shift[0] ), .C(new_n514_), .Y(new_n515_));
  INVX1    g0252(.A(\a[64] ), .Y(new_n516_));
  NOR3X1   g0253(.A(\shift[1] ), .B(\shift[0] ), .C(new_n516_), .Y(new_n517_));
  INVX1    g0254(.A(\a[63] ), .Y(new_n518_));
  NOR3X1   g0255(.A(\shift[1] ), .B(new_n266_), .C(new_n518_), .Y(new_n519_));
  OR4X1    g0256(.A(new_n519_), .B(new_n517_), .C(new_n515_), .D(new_n513_), .Y(new_n520_));
  INVX1    g0257(.A(\a[57] ), .Y(new_n521_));
  NOR3X1   g0258(.A(new_n267_), .B(new_n266_), .C(new_n521_), .Y(new_n522_));
  INVX1    g0259(.A(\a[58] ), .Y(new_n523_));
  NOR3X1   g0260(.A(new_n267_), .B(\shift[0] ), .C(new_n523_), .Y(new_n524_));
  INVX1    g0261(.A(\a[60] ), .Y(new_n525_));
  NOR3X1   g0262(.A(\shift[1] ), .B(\shift[0] ), .C(new_n525_), .Y(new_n526_));
  INVX1    g0263(.A(\a[59] ), .Y(new_n527_));
  NOR3X1   g0264(.A(\shift[1] ), .B(new_n266_), .C(new_n527_), .Y(new_n528_));
  OR4X1    g0265(.A(new_n528_), .B(new_n526_), .C(new_n524_), .D(new_n522_), .Y(new_n529_));
  AOI22X1  g0266(.A0(new_n529_), .A1(new_n287_), .B0(new_n520_), .B1(new_n276_), .Y(new_n530_));
  INVX1    g0267(.A(\a[49] ), .Y(new_n531_));
  NOR3X1   g0268(.A(new_n267_), .B(new_n266_), .C(new_n531_), .Y(new_n532_));
  INVX1    g0269(.A(\a[50] ), .Y(new_n533_));
  NOR3X1   g0270(.A(new_n267_), .B(\shift[0] ), .C(new_n533_), .Y(new_n534_));
  INVX1    g0271(.A(\a[52] ), .Y(new_n535_));
  NOR3X1   g0272(.A(\shift[1] ), .B(\shift[0] ), .C(new_n535_), .Y(new_n536_));
  INVX1    g0273(.A(\a[51] ), .Y(new_n537_));
  NOR3X1   g0274(.A(\shift[1] ), .B(new_n266_), .C(new_n537_), .Y(new_n538_));
  OR4X1    g0275(.A(new_n538_), .B(new_n536_), .C(new_n534_), .D(new_n532_), .Y(new_n539_));
  INVX1    g0276(.A(\a[53] ), .Y(new_n540_));
  NOR3X1   g0277(.A(new_n267_), .B(new_n266_), .C(new_n540_), .Y(new_n541_));
  INVX1    g0278(.A(\a[54] ), .Y(new_n542_));
  NOR3X1   g0279(.A(new_n267_), .B(\shift[0] ), .C(new_n542_), .Y(new_n543_));
  INVX1    g0280(.A(\a[56] ), .Y(new_n544_));
  NOR3X1   g0281(.A(\shift[1] ), .B(\shift[0] ), .C(new_n544_), .Y(new_n545_));
  INVX1    g0282(.A(\a[55] ), .Y(new_n546_));
  NOR3X1   g0283(.A(\shift[1] ), .B(new_n266_), .C(new_n546_), .Y(new_n547_));
  OR4X1    g0284(.A(new_n547_), .B(new_n545_), .C(new_n543_), .D(new_n541_), .Y(new_n548_));
  AOI22X1  g0285(.A0(new_n548_), .A1(new_n308_), .B0(new_n539_), .B1(new_n298_), .Y(new_n549_));
  AOI21X1  g0286(.A0(new_n549_), .A1(new_n530_), .B0(new_n391_), .Y(new_n550_));
  INVX1    g0287(.A(\a[45] ), .Y(new_n551_));
  NOR3X1   g0288(.A(new_n267_), .B(new_n266_), .C(new_n551_), .Y(new_n552_));
  INVX1    g0289(.A(\a[46] ), .Y(new_n553_));
  NOR3X1   g0290(.A(new_n267_), .B(\shift[0] ), .C(new_n553_), .Y(new_n554_));
  INVX1    g0291(.A(\a[48] ), .Y(new_n555_));
  NOR3X1   g0292(.A(\shift[1] ), .B(\shift[0] ), .C(new_n555_), .Y(new_n556_));
  INVX1    g0293(.A(\a[47] ), .Y(new_n557_));
  NOR3X1   g0294(.A(\shift[1] ), .B(new_n266_), .C(new_n557_), .Y(new_n558_));
  OR4X1    g0295(.A(new_n558_), .B(new_n556_), .C(new_n554_), .D(new_n552_), .Y(new_n559_));
  INVX1    g0296(.A(\a[41] ), .Y(new_n560_));
  NOR3X1   g0297(.A(new_n267_), .B(new_n266_), .C(new_n560_), .Y(new_n561_));
  INVX1    g0298(.A(\a[42] ), .Y(new_n562_));
  NOR3X1   g0299(.A(new_n267_), .B(\shift[0] ), .C(new_n562_), .Y(new_n563_));
  INVX1    g0300(.A(\a[44] ), .Y(new_n564_));
  NOR3X1   g0301(.A(\shift[1] ), .B(\shift[0] ), .C(new_n564_), .Y(new_n565_));
  INVX1    g0302(.A(\a[43] ), .Y(new_n566_));
  NOR3X1   g0303(.A(\shift[1] ), .B(new_n266_), .C(new_n566_), .Y(new_n567_));
  OR4X1    g0304(.A(new_n567_), .B(new_n565_), .C(new_n563_), .D(new_n561_), .Y(new_n568_));
  AOI22X1  g0305(.A0(new_n568_), .A1(new_n287_), .B0(new_n559_), .B1(new_n276_), .Y(new_n569_));
  INVX1    g0306(.A(\a[33] ), .Y(new_n570_));
  NOR3X1   g0307(.A(new_n267_), .B(new_n266_), .C(new_n570_), .Y(new_n571_));
  INVX1    g0308(.A(\a[34] ), .Y(new_n572_));
  NOR3X1   g0309(.A(new_n267_), .B(\shift[0] ), .C(new_n572_), .Y(new_n573_));
  INVX1    g0310(.A(\a[36] ), .Y(new_n574_));
  NOR3X1   g0311(.A(\shift[1] ), .B(\shift[0] ), .C(new_n574_), .Y(new_n575_));
  INVX1    g0312(.A(\a[35] ), .Y(new_n576_));
  NOR3X1   g0313(.A(\shift[1] ), .B(new_n266_), .C(new_n576_), .Y(new_n577_));
  OR4X1    g0314(.A(new_n577_), .B(new_n575_), .C(new_n573_), .D(new_n571_), .Y(new_n578_));
  INVX1    g0315(.A(\a[40] ), .Y(new_n579_));
  NOR3X1   g0316(.A(\shift[1] ), .B(\shift[0] ), .C(new_n579_), .Y(new_n580_));
  INVX1    g0317(.A(\a[37] ), .Y(new_n581_));
  NOR3X1   g0318(.A(new_n267_), .B(new_n266_), .C(new_n581_), .Y(new_n582_));
  INVX1    g0319(.A(\a[39] ), .Y(new_n583_));
  NOR3X1   g0320(.A(\shift[1] ), .B(new_n266_), .C(new_n583_), .Y(new_n584_));
  INVX1    g0321(.A(\a[38] ), .Y(new_n585_));
  NOR3X1   g0322(.A(new_n267_), .B(\shift[0] ), .C(new_n585_), .Y(new_n586_));
  OR4X1    g0323(.A(new_n586_), .B(new_n584_), .C(new_n582_), .D(new_n580_), .Y(new_n587_));
  AOI22X1  g0324(.A0(new_n587_), .A1(new_n308_), .B0(new_n578_), .B1(new_n298_), .Y(new_n588_));
  AOI21X1  g0325(.A0(new_n588_), .A1(new_n569_), .B0(new_n431_), .Y(new_n589_));
  OR4X1    g0326(.A(new_n589_), .B(new_n550_), .C(new_n511_), .D(new_n472_), .Y(new_n590_));
  MX2X1    g0327(.A(new_n590_), .B(new_n433_), .S0(new_n264_), .Y(\result[0] ));
  NOR3X1   g0328(.A(\shift[1] ), .B(\shift[0] ), .C(new_n331_), .Y(new_n592_));
  NOR3X1   g0329(.A(new_n267_), .B(new_n266_), .C(new_n269_), .Y(new_n593_));
  NOR3X1   g0330(.A(\shift[1] ), .B(new_n266_), .C(new_n271_), .Y(new_n594_));
  NOR3X1   g0331(.A(new_n267_), .B(\shift[0] ), .C(new_n273_), .Y(new_n595_));
  OR4X1    g0332(.A(new_n595_), .B(new_n594_), .C(new_n593_), .D(new_n592_), .Y(new_n596_));
  NOR3X1   g0333(.A(\shift[1] ), .B(\shift[0] ), .C(new_n265_), .Y(new_n597_));
  NOR3X1   g0334(.A(new_n267_), .B(new_n266_), .C(new_n279_), .Y(new_n598_));
  NOR3X1   g0335(.A(\shift[1] ), .B(new_n266_), .C(new_n281_), .Y(new_n599_));
  NOR3X1   g0336(.A(new_n267_), .B(\shift[0] ), .C(new_n283_), .Y(new_n600_));
  OR4X1    g0337(.A(new_n600_), .B(new_n599_), .C(new_n598_), .D(new_n597_), .Y(new_n601_));
  AOI22X1  g0338(.A0(new_n601_), .A1(new_n287_), .B0(new_n596_), .B1(new_n276_), .Y(new_n602_));
  NOR3X1   g0339(.A(\shift[1] ), .B(\shift[0] ), .C(new_n299_), .Y(new_n603_));
  NOR3X1   g0340(.A(new_n267_), .B(new_n266_), .C(new_n291_), .Y(new_n604_));
  NOR3X1   g0341(.A(\shift[1] ), .B(new_n266_), .C(new_n293_), .Y(new_n605_));
  NOR3X1   g0342(.A(new_n267_), .B(\shift[0] ), .C(new_n295_), .Y(new_n606_));
  OR4X1    g0343(.A(new_n606_), .B(new_n605_), .C(new_n604_), .D(new_n603_), .Y(new_n607_));
  NOR3X1   g0344(.A(\shift[1] ), .B(\shift[0] ), .C(new_n277_), .Y(new_n608_));
  NOR3X1   g0345(.A(new_n267_), .B(new_n266_), .C(new_n301_), .Y(new_n609_));
  NOR3X1   g0346(.A(\shift[1] ), .B(new_n266_), .C(new_n303_), .Y(new_n610_));
  NOR3X1   g0347(.A(new_n267_), .B(\shift[0] ), .C(new_n305_), .Y(new_n611_));
  OR4X1    g0348(.A(new_n611_), .B(new_n610_), .C(new_n609_), .D(new_n608_), .Y(new_n612_));
  AOI22X1  g0349(.A0(new_n612_), .A1(new_n308_), .B0(new_n607_), .B1(new_n298_), .Y(new_n613_));
  AOI21X1  g0350(.A0(new_n613_), .A1(new_n602_), .B0(new_n310_), .Y(new_n614_));
  NOR3X1   g0351(.A(\shift[1] ), .B(\shift[0] ), .C(new_n412_), .Y(new_n615_));
  NOR3X1   g0352(.A(new_n267_), .B(new_n266_), .C(new_n314_), .Y(new_n616_));
  NOR3X1   g0353(.A(\shift[1] ), .B(new_n266_), .C(new_n316_), .Y(new_n617_));
  NOR3X1   g0354(.A(new_n267_), .B(\shift[0] ), .C(new_n318_), .Y(new_n618_));
  OR4X1    g0355(.A(new_n618_), .B(new_n617_), .C(new_n616_), .D(new_n615_), .Y(new_n619_));
  NOR3X1   g0356(.A(\shift[1] ), .B(\shift[0] ), .C(new_n312_), .Y(new_n620_));
  NOR3X1   g0357(.A(new_n267_), .B(new_n266_), .C(new_n323_), .Y(new_n621_));
  NOR3X1   g0358(.A(\shift[1] ), .B(new_n266_), .C(new_n325_), .Y(new_n622_));
  NOR3X1   g0359(.A(new_n267_), .B(\shift[0] ), .C(new_n327_), .Y(new_n623_));
  OR4X1    g0360(.A(new_n623_), .B(new_n622_), .C(new_n621_), .D(new_n620_), .Y(new_n624_));
  AOI22X1  g0361(.A0(new_n624_), .A1(new_n287_), .B0(new_n619_), .B1(new_n276_), .Y(new_n625_));
  NOR3X1   g0362(.A(\shift[1] ), .B(\shift[0] ), .C(new_n340_), .Y(new_n626_));
  NOR3X1   g0363(.A(new_n267_), .B(new_n266_), .C(new_n333_), .Y(new_n627_));
  NOR3X1   g0364(.A(\shift[1] ), .B(new_n266_), .C(new_n335_), .Y(new_n628_));
  NOR3X1   g0365(.A(new_n267_), .B(\shift[0] ), .C(new_n337_), .Y(new_n629_));
  OR4X1    g0366(.A(new_n629_), .B(new_n628_), .C(new_n627_), .D(new_n626_), .Y(new_n630_));
  NOR3X1   g0367(.A(\shift[1] ), .B(\shift[0] ), .C(new_n321_), .Y(new_n631_));
  NOR3X1   g0368(.A(new_n267_), .B(new_n266_), .C(new_n342_), .Y(new_n632_));
  NOR3X1   g0369(.A(\shift[1] ), .B(new_n266_), .C(new_n344_), .Y(new_n633_));
  NOR3X1   g0370(.A(new_n267_), .B(\shift[0] ), .C(new_n346_), .Y(new_n634_));
  OR4X1    g0371(.A(new_n634_), .B(new_n633_), .C(new_n632_), .D(new_n631_), .Y(new_n635_));
  AOI22X1  g0372(.A0(new_n635_), .A1(new_n308_), .B0(new_n630_), .B1(new_n298_), .Y(new_n636_));
  AOI21X1  g0373(.A0(new_n636_), .A1(new_n625_), .B0(new_n351_), .Y(new_n637_));
  NOR3X1   g0374(.A(\shift[1] ), .B(\shift[0] ), .C(new_n453_), .Y(new_n638_));
  NOR3X1   g0375(.A(new_n267_), .B(new_n266_), .C(new_n355_), .Y(new_n639_));
  NOR3X1   g0376(.A(\shift[1] ), .B(new_n266_), .C(new_n357_), .Y(new_n640_));
  NOR3X1   g0377(.A(new_n267_), .B(\shift[0] ), .C(new_n359_), .Y(new_n641_));
  OR4X1    g0378(.A(new_n641_), .B(new_n640_), .C(new_n639_), .D(new_n638_), .Y(new_n642_));
  NOR3X1   g0379(.A(\shift[1] ), .B(\shift[0] ), .C(new_n353_), .Y(new_n643_));
  NOR3X1   g0380(.A(new_n267_), .B(new_n266_), .C(new_n364_), .Y(new_n644_));
  NOR3X1   g0381(.A(\shift[1] ), .B(new_n266_), .C(new_n366_), .Y(new_n645_));
  NOR3X1   g0382(.A(new_n267_), .B(\shift[0] ), .C(new_n368_), .Y(new_n646_));
  OR4X1    g0383(.A(new_n646_), .B(new_n645_), .C(new_n644_), .D(new_n643_), .Y(new_n647_));
  AOI22X1  g0384(.A0(new_n647_), .A1(new_n287_), .B0(new_n642_), .B1(new_n276_), .Y(new_n648_));
  NOR3X1   g0385(.A(\shift[1] ), .B(\shift[0] ), .C(new_n381_), .Y(new_n649_));
  NOR3X1   g0386(.A(new_n267_), .B(new_n266_), .C(new_n374_), .Y(new_n650_));
  NOR3X1   g0387(.A(\shift[1] ), .B(new_n266_), .C(new_n376_), .Y(new_n651_));
  NOR3X1   g0388(.A(new_n267_), .B(\shift[0] ), .C(new_n378_), .Y(new_n652_));
  OR4X1    g0389(.A(new_n652_), .B(new_n651_), .C(new_n650_), .D(new_n649_), .Y(new_n653_));
  NOR3X1   g0390(.A(\shift[1] ), .B(\shift[0] ), .C(new_n362_), .Y(new_n654_));
  NOR3X1   g0391(.A(new_n267_), .B(new_n266_), .C(new_n383_), .Y(new_n655_));
  NOR3X1   g0392(.A(\shift[1] ), .B(new_n266_), .C(new_n385_), .Y(new_n656_));
  NOR3X1   g0393(.A(new_n267_), .B(\shift[0] ), .C(new_n387_), .Y(new_n657_));
  OR4X1    g0394(.A(new_n657_), .B(new_n656_), .C(new_n655_), .D(new_n654_), .Y(new_n658_));
  AOI22X1  g0395(.A0(new_n658_), .A1(new_n308_), .B0(new_n653_), .B1(new_n298_), .Y(new_n659_));
  AOI21X1  g0396(.A0(new_n659_), .A1(new_n648_), .B0(new_n391_), .Y(new_n660_));
  NOR3X1   g0397(.A(\shift[1] ), .B(\shift[0] ), .C(new_n372_), .Y(new_n661_));
  NOR3X1   g0398(.A(new_n267_), .B(new_n266_), .C(new_n395_), .Y(new_n662_));
  NOR3X1   g0399(.A(\shift[1] ), .B(new_n266_), .C(new_n397_), .Y(new_n663_));
  NOR3X1   g0400(.A(new_n267_), .B(\shift[0] ), .C(new_n399_), .Y(new_n664_));
  OR4X1    g0401(.A(new_n664_), .B(new_n663_), .C(new_n662_), .D(new_n661_), .Y(new_n665_));
  NOR3X1   g0402(.A(\shift[1] ), .B(\shift[0] ), .C(new_n393_), .Y(new_n666_));
  NOR3X1   g0403(.A(new_n267_), .B(new_n266_), .C(new_n404_), .Y(new_n667_));
  NOR3X1   g0404(.A(\shift[1] ), .B(new_n266_), .C(new_n406_), .Y(new_n668_));
  NOR3X1   g0405(.A(new_n267_), .B(\shift[0] ), .C(new_n408_), .Y(new_n669_));
  OR4X1    g0406(.A(new_n669_), .B(new_n668_), .C(new_n667_), .D(new_n666_), .Y(new_n670_));
  AOI22X1  g0407(.A0(new_n670_), .A1(new_n287_), .B0(new_n665_), .B1(new_n276_), .Y(new_n671_));
  NOR3X1   g0408(.A(\shift[1] ), .B(\shift[0] ), .C(new_n421_), .Y(new_n672_));
  NOR3X1   g0409(.A(new_n267_), .B(new_n266_), .C(new_n414_), .Y(new_n673_));
  NOR3X1   g0410(.A(\shift[1] ), .B(new_n266_), .C(new_n416_), .Y(new_n674_));
  NOR3X1   g0411(.A(new_n267_), .B(\shift[0] ), .C(new_n418_), .Y(new_n675_));
  OR4X1    g0412(.A(new_n675_), .B(new_n674_), .C(new_n673_), .D(new_n672_), .Y(new_n676_));
  NOR3X1   g0413(.A(\shift[1] ), .B(\shift[0] ), .C(new_n402_), .Y(new_n677_));
  NOR3X1   g0414(.A(new_n267_), .B(new_n266_), .C(new_n423_), .Y(new_n678_));
  NOR3X1   g0415(.A(\shift[1] ), .B(new_n266_), .C(new_n425_), .Y(new_n679_));
  NOR3X1   g0416(.A(new_n267_), .B(\shift[0] ), .C(new_n427_), .Y(new_n680_));
  OR4X1    g0417(.A(new_n680_), .B(new_n679_), .C(new_n678_), .D(new_n677_), .Y(new_n681_));
  AOI22X1  g0418(.A0(new_n681_), .A1(new_n308_), .B0(new_n676_), .B1(new_n298_), .Y(new_n682_));
  AOI21X1  g0419(.A0(new_n682_), .A1(new_n671_), .B0(new_n431_), .Y(new_n683_));
  OR4X1    g0420(.A(new_n683_), .B(new_n660_), .C(new_n637_), .D(new_n614_), .Y(new_n684_));
  NOR3X1   g0421(.A(\shift[1] ), .B(\shift[0] ), .C(new_n289_), .Y(new_n685_));
  NOR3X1   g0422(.A(new_n267_), .B(new_n266_), .C(new_n514_), .Y(new_n686_));
  NOR3X1   g0423(.A(\shift[1] ), .B(new_n266_), .C(new_n516_), .Y(new_n687_));
  NOR3X1   g0424(.A(new_n267_), .B(\shift[0] ), .C(new_n518_), .Y(new_n688_));
  OR4X1    g0425(.A(new_n688_), .B(new_n687_), .C(new_n686_), .D(new_n685_), .Y(new_n689_));
  NOR3X1   g0426(.A(\shift[1] ), .B(\shift[0] ), .C(new_n512_), .Y(new_n690_));
  NOR3X1   g0427(.A(new_n267_), .B(new_n266_), .C(new_n523_), .Y(new_n691_));
  NOR3X1   g0428(.A(\shift[1] ), .B(new_n266_), .C(new_n525_), .Y(new_n692_));
  NOR3X1   g0429(.A(new_n267_), .B(\shift[0] ), .C(new_n527_), .Y(new_n693_));
  OR4X1    g0430(.A(new_n693_), .B(new_n692_), .C(new_n691_), .D(new_n690_), .Y(new_n694_));
  AOI22X1  g0431(.A0(new_n694_), .A1(new_n287_), .B0(new_n689_), .B1(new_n276_), .Y(new_n695_));
  NOR3X1   g0432(.A(\shift[1] ), .B(\shift[0] ), .C(new_n540_), .Y(new_n696_));
  NOR3X1   g0433(.A(new_n267_), .B(new_n266_), .C(new_n533_), .Y(new_n697_));
  NOR3X1   g0434(.A(\shift[1] ), .B(new_n266_), .C(new_n535_), .Y(new_n698_));
  NOR3X1   g0435(.A(new_n267_), .B(\shift[0] ), .C(new_n537_), .Y(new_n699_));
  OR4X1    g0436(.A(new_n699_), .B(new_n698_), .C(new_n697_), .D(new_n696_), .Y(new_n700_));
  NOR3X1   g0437(.A(\shift[1] ), .B(\shift[0] ), .C(new_n521_), .Y(new_n701_));
  NOR3X1   g0438(.A(new_n267_), .B(new_n266_), .C(new_n542_), .Y(new_n702_));
  NOR3X1   g0439(.A(\shift[1] ), .B(new_n266_), .C(new_n544_), .Y(new_n703_));
  NOR3X1   g0440(.A(new_n267_), .B(\shift[0] ), .C(new_n546_), .Y(new_n704_));
  OR4X1    g0441(.A(new_n704_), .B(new_n703_), .C(new_n702_), .D(new_n701_), .Y(new_n705_));
  AOI22X1  g0442(.A0(new_n705_), .A1(new_n308_), .B0(new_n700_), .B1(new_n298_), .Y(new_n706_));
  AOI21X1  g0443(.A0(new_n706_), .A1(new_n695_), .B0(new_n391_), .Y(new_n707_));
  NOR3X1   g0444(.A(\shift[1] ), .B(\shift[0] ), .C(new_n492_), .Y(new_n708_));
  NOR3X1   g0445(.A(new_n267_), .B(new_n266_), .C(new_n436_), .Y(new_n709_));
  NOR3X1   g0446(.A(\shift[1] ), .B(new_n266_), .C(new_n438_), .Y(new_n710_));
  NOR3X1   g0447(.A(new_n267_), .B(\shift[0] ), .C(new_n440_), .Y(new_n711_));
  OR4X1    g0448(.A(new_n711_), .B(new_n710_), .C(new_n709_), .D(new_n708_), .Y(new_n712_));
  NOR3X1   g0449(.A(\shift[1] ), .B(\shift[0] ), .C(new_n434_), .Y(new_n713_));
  NOR3X1   g0450(.A(new_n267_), .B(new_n266_), .C(new_n445_), .Y(new_n714_));
  NOR3X1   g0451(.A(\shift[1] ), .B(new_n266_), .C(new_n447_), .Y(new_n715_));
  NOR3X1   g0452(.A(new_n267_), .B(\shift[0] ), .C(new_n449_), .Y(new_n716_));
  OR4X1    g0453(.A(new_n716_), .B(new_n715_), .C(new_n714_), .D(new_n713_), .Y(new_n717_));
  AOI22X1  g0454(.A0(new_n717_), .A1(new_n287_), .B0(new_n712_), .B1(new_n276_), .Y(new_n718_));
  NOR3X1   g0455(.A(\shift[1] ), .B(\shift[0] ), .C(new_n462_), .Y(new_n719_));
  NOR3X1   g0456(.A(new_n267_), .B(new_n266_), .C(new_n455_), .Y(new_n720_));
  NOR3X1   g0457(.A(\shift[1] ), .B(new_n266_), .C(new_n457_), .Y(new_n721_));
  NOR3X1   g0458(.A(new_n267_), .B(\shift[0] ), .C(new_n459_), .Y(new_n722_));
  OR4X1    g0459(.A(new_n722_), .B(new_n721_), .C(new_n720_), .D(new_n719_), .Y(new_n723_));
  NOR3X1   g0460(.A(\shift[1] ), .B(\shift[0] ), .C(new_n443_), .Y(new_n724_));
  NOR3X1   g0461(.A(new_n267_), .B(new_n266_), .C(new_n464_), .Y(new_n725_));
  NOR3X1   g0462(.A(\shift[1] ), .B(new_n266_), .C(new_n466_), .Y(new_n726_));
  NOR3X1   g0463(.A(new_n267_), .B(\shift[0] ), .C(new_n468_), .Y(new_n727_));
  OR4X1    g0464(.A(new_n727_), .B(new_n726_), .C(new_n725_), .D(new_n724_), .Y(new_n728_));
  AOI22X1  g0465(.A0(new_n728_), .A1(new_n308_), .B0(new_n723_), .B1(new_n298_), .Y(new_n729_));
  AOI21X1  g0466(.A0(new_n729_), .A1(new_n718_), .B0(new_n310_), .Y(new_n730_));
  NOR3X1   g0467(.A(\shift[1] ), .B(\shift[0] ), .C(new_n531_), .Y(new_n731_));
  NOR3X1   g0468(.A(new_n267_), .B(new_n266_), .C(new_n553_), .Y(new_n732_));
  NOR3X1   g0469(.A(\shift[1] ), .B(new_n266_), .C(new_n555_), .Y(new_n733_));
  NOR3X1   g0470(.A(new_n267_), .B(\shift[0] ), .C(new_n557_), .Y(new_n734_));
  OR4X1    g0471(.A(new_n734_), .B(new_n733_), .C(new_n732_), .D(new_n731_), .Y(new_n735_));
  NOR3X1   g0472(.A(new_n267_), .B(new_n266_), .C(new_n562_), .Y(new_n736_));
  NOR3X1   g0473(.A(new_n267_), .B(\shift[0] ), .C(new_n566_), .Y(new_n737_));
  NOR3X1   g0474(.A(\shift[1] ), .B(\shift[0] ), .C(new_n551_), .Y(new_n738_));
  NOR3X1   g0475(.A(\shift[1] ), .B(new_n266_), .C(new_n564_), .Y(new_n739_));
  OR4X1    g0476(.A(new_n739_), .B(new_n738_), .C(new_n737_), .D(new_n736_), .Y(new_n740_));
  AOI22X1  g0477(.A0(new_n740_), .A1(new_n287_), .B0(new_n735_), .B1(new_n276_), .Y(new_n741_));
  NOR3X1   g0478(.A(\shift[1] ), .B(\shift[0] ), .C(new_n581_), .Y(new_n742_));
  NOR3X1   g0479(.A(new_n267_), .B(new_n266_), .C(new_n572_), .Y(new_n743_));
  NOR3X1   g0480(.A(\shift[1] ), .B(new_n266_), .C(new_n574_), .Y(new_n744_));
  NOR3X1   g0481(.A(new_n267_), .B(\shift[0] ), .C(new_n576_), .Y(new_n745_));
  OR4X1    g0482(.A(new_n745_), .B(new_n744_), .C(new_n743_), .D(new_n742_), .Y(new_n746_));
  NOR3X1   g0483(.A(\shift[1] ), .B(\shift[0] ), .C(new_n560_), .Y(new_n747_));
  NOR3X1   g0484(.A(\shift[1] ), .B(new_n266_), .C(new_n579_), .Y(new_n748_));
  NOR3X1   g0485(.A(new_n267_), .B(\shift[0] ), .C(new_n583_), .Y(new_n749_));
  NOR3X1   g0486(.A(new_n267_), .B(new_n266_), .C(new_n585_), .Y(new_n750_));
  OR4X1    g0487(.A(new_n750_), .B(new_n749_), .C(new_n748_), .D(new_n747_), .Y(new_n751_));
  AOI22X1  g0488(.A0(new_n751_), .A1(new_n308_), .B0(new_n746_), .B1(new_n298_), .Y(new_n752_));
  AOI21X1  g0489(.A0(new_n752_), .A1(new_n741_), .B0(new_n431_), .Y(new_n753_));
  NOR3X1   g0490(.A(\shift[1] ), .B(\shift[0] ), .C(new_n570_), .Y(new_n754_));
  NOR3X1   g0491(.A(new_n267_), .B(new_n266_), .C(new_n475_), .Y(new_n755_));
  NOR3X1   g0492(.A(\shift[1] ), .B(new_n266_), .C(new_n477_), .Y(new_n756_));
  NOR3X1   g0493(.A(new_n267_), .B(\shift[0] ), .C(new_n479_), .Y(new_n757_));
  OR4X1    g0494(.A(new_n757_), .B(new_n756_), .C(new_n755_), .D(new_n754_), .Y(new_n758_));
  NOR3X1   g0495(.A(\shift[1] ), .B(\shift[0] ), .C(new_n473_), .Y(new_n759_));
  NOR3X1   g0496(.A(new_n267_), .B(new_n266_), .C(new_n484_), .Y(new_n760_));
  NOR3X1   g0497(.A(\shift[1] ), .B(new_n266_), .C(new_n486_), .Y(new_n761_));
  NOR3X1   g0498(.A(new_n267_), .B(\shift[0] ), .C(new_n488_), .Y(new_n762_));
  OR4X1    g0499(.A(new_n762_), .B(new_n761_), .C(new_n760_), .D(new_n759_), .Y(new_n763_));
  AOI22X1  g0500(.A0(new_n763_), .A1(new_n287_), .B0(new_n758_), .B1(new_n276_), .Y(new_n764_));
  NOR3X1   g0501(.A(\shift[1] ), .B(\shift[0] ), .C(new_n501_), .Y(new_n765_));
  NOR3X1   g0502(.A(new_n267_), .B(new_n266_), .C(new_n494_), .Y(new_n766_));
  NOR3X1   g0503(.A(\shift[1] ), .B(new_n266_), .C(new_n496_), .Y(new_n767_));
  NOR3X1   g0504(.A(new_n267_), .B(\shift[0] ), .C(new_n498_), .Y(new_n768_));
  OR4X1    g0505(.A(new_n768_), .B(new_n767_), .C(new_n766_), .D(new_n765_), .Y(new_n769_));
  NOR3X1   g0506(.A(\shift[1] ), .B(\shift[0] ), .C(new_n482_), .Y(new_n770_));
  NOR3X1   g0507(.A(new_n267_), .B(new_n266_), .C(new_n503_), .Y(new_n771_));
  NOR3X1   g0508(.A(\shift[1] ), .B(new_n266_), .C(new_n505_), .Y(new_n772_));
  NOR3X1   g0509(.A(new_n267_), .B(\shift[0] ), .C(new_n507_), .Y(new_n773_));
  OR4X1    g0510(.A(new_n773_), .B(new_n772_), .C(new_n771_), .D(new_n770_), .Y(new_n774_));
  AOI22X1  g0511(.A0(new_n774_), .A1(new_n308_), .B0(new_n769_), .B1(new_n298_), .Y(new_n775_));
  AOI21X1  g0512(.A0(new_n775_), .A1(new_n764_), .B0(new_n351_), .Y(new_n776_));
  OR4X1    g0513(.A(new_n776_), .B(new_n753_), .C(new_n730_), .D(new_n707_), .Y(new_n777_));
  MX2X1    g0514(.A(new_n777_), .B(new_n684_), .S0(new_n264_), .Y(\result[1] ));
  NOR3X1   g0515(.A(\shift[1] ), .B(new_n266_), .C(new_n331_), .Y(new_n779_));
  NOR3X1   g0516(.A(\shift[1] ), .B(\shift[0] ), .C(new_n333_), .Y(new_n780_));
  NOR3X1   g0517(.A(new_n267_), .B(\shift[0] ), .C(new_n271_), .Y(new_n781_));
  NOR3X1   g0518(.A(new_n267_), .B(new_n266_), .C(new_n273_), .Y(new_n782_));
  OR4X1    g0519(.A(new_n782_), .B(new_n781_), .C(new_n780_), .D(new_n779_), .Y(new_n783_));
  NOR3X1   g0520(.A(\shift[1] ), .B(new_n266_), .C(new_n265_), .Y(new_n784_));
  NOR3X1   g0521(.A(\shift[1] ), .B(\shift[0] ), .C(new_n269_), .Y(new_n785_));
  NOR3X1   g0522(.A(new_n267_), .B(\shift[0] ), .C(new_n281_), .Y(new_n786_));
  NOR3X1   g0523(.A(new_n267_), .B(new_n266_), .C(new_n283_), .Y(new_n787_));
  OR4X1    g0524(.A(new_n787_), .B(new_n786_), .C(new_n785_), .D(new_n784_), .Y(new_n788_));
  AOI22X1  g0525(.A0(new_n788_), .A1(new_n287_), .B0(new_n783_), .B1(new_n276_), .Y(new_n789_));
  NOR3X1   g0526(.A(\shift[1] ), .B(new_n266_), .C(new_n299_), .Y(new_n790_));
  NOR3X1   g0527(.A(\shift[1] ), .B(\shift[0] ), .C(new_n301_), .Y(new_n791_));
  NOR3X1   g0528(.A(new_n267_), .B(\shift[0] ), .C(new_n293_), .Y(new_n792_));
  NOR3X1   g0529(.A(new_n267_), .B(new_n266_), .C(new_n295_), .Y(new_n793_));
  OR4X1    g0530(.A(new_n793_), .B(new_n792_), .C(new_n791_), .D(new_n790_), .Y(new_n794_));
  NOR3X1   g0531(.A(\shift[1] ), .B(new_n266_), .C(new_n277_), .Y(new_n795_));
  NOR3X1   g0532(.A(\shift[1] ), .B(\shift[0] ), .C(new_n279_), .Y(new_n796_));
  NOR3X1   g0533(.A(new_n267_), .B(\shift[0] ), .C(new_n303_), .Y(new_n797_));
  NOR3X1   g0534(.A(new_n267_), .B(new_n266_), .C(new_n305_), .Y(new_n798_));
  OR4X1    g0535(.A(new_n798_), .B(new_n797_), .C(new_n796_), .D(new_n795_), .Y(new_n799_));
  AOI22X1  g0536(.A0(new_n799_), .A1(new_n308_), .B0(new_n794_), .B1(new_n298_), .Y(new_n800_));
  AOI21X1  g0537(.A0(new_n800_), .A1(new_n789_), .B0(new_n310_), .Y(new_n801_));
  NOR3X1   g0538(.A(\shift[1] ), .B(new_n266_), .C(new_n412_), .Y(new_n802_));
  NOR3X1   g0539(.A(\shift[1] ), .B(\shift[0] ), .C(new_n414_), .Y(new_n803_));
  NOR3X1   g0540(.A(new_n267_), .B(\shift[0] ), .C(new_n316_), .Y(new_n804_));
  NOR3X1   g0541(.A(new_n267_), .B(new_n266_), .C(new_n318_), .Y(new_n805_));
  OR4X1    g0542(.A(new_n805_), .B(new_n804_), .C(new_n803_), .D(new_n802_), .Y(new_n806_));
  NOR3X1   g0543(.A(\shift[1] ), .B(new_n266_), .C(new_n312_), .Y(new_n807_));
  NOR3X1   g0544(.A(\shift[1] ), .B(\shift[0] ), .C(new_n314_), .Y(new_n808_));
  NOR3X1   g0545(.A(new_n267_), .B(\shift[0] ), .C(new_n325_), .Y(new_n809_));
  NOR3X1   g0546(.A(new_n267_), .B(new_n266_), .C(new_n327_), .Y(new_n810_));
  OR4X1    g0547(.A(new_n810_), .B(new_n809_), .C(new_n808_), .D(new_n807_), .Y(new_n811_));
  AOI22X1  g0548(.A0(new_n811_), .A1(new_n287_), .B0(new_n806_), .B1(new_n276_), .Y(new_n812_));
  NOR3X1   g0549(.A(\shift[1] ), .B(new_n266_), .C(new_n340_), .Y(new_n813_));
  NOR3X1   g0550(.A(\shift[1] ), .B(\shift[0] ), .C(new_n342_), .Y(new_n814_));
  NOR3X1   g0551(.A(new_n267_), .B(\shift[0] ), .C(new_n335_), .Y(new_n815_));
  NOR3X1   g0552(.A(new_n267_), .B(new_n266_), .C(new_n337_), .Y(new_n816_));
  OR4X1    g0553(.A(new_n816_), .B(new_n815_), .C(new_n814_), .D(new_n813_), .Y(new_n817_));
  NOR3X1   g0554(.A(\shift[1] ), .B(new_n266_), .C(new_n321_), .Y(new_n818_));
  NOR3X1   g0555(.A(\shift[1] ), .B(\shift[0] ), .C(new_n323_), .Y(new_n819_));
  NOR3X1   g0556(.A(new_n267_), .B(\shift[0] ), .C(new_n344_), .Y(new_n820_));
  NOR3X1   g0557(.A(new_n267_), .B(new_n266_), .C(new_n346_), .Y(new_n821_));
  OR4X1    g0558(.A(new_n821_), .B(new_n820_), .C(new_n819_), .D(new_n818_), .Y(new_n822_));
  AOI22X1  g0559(.A0(new_n822_), .A1(new_n308_), .B0(new_n817_), .B1(new_n298_), .Y(new_n823_));
  AOI21X1  g0560(.A0(new_n823_), .A1(new_n812_), .B0(new_n351_), .Y(new_n824_));
  NOR3X1   g0561(.A(\shift[1] ), .B(new_n266_), .C(new_n453_), .Y(new_n825_));
  NOR3X1   g0562(.A(\shift[1] ), .B(\shift[0] ), .C(new_n455_), .Y(new_n826_));
  NOR3X1   g0563(.A(new_n267_), .B(\shift[0] ), .C(new_n357_), .Y(new_n827_));
  NOR3X1   g0564(.A(new_n267_), .B(new_n266_), .C(new_n359_), .Y(new_n828_));
  OR4X1    g0565(.A(new_n828_), .B(new_n827_), .C(new_n826_), .D(new_n825_), .Y(new_n829_));
  NOR3X1   g0566(.A(\shift[1] ), .B(new_n266_), .C(new_n353_), .Y(new_n830_));
  NOR3X1   g0567(.A(\shift[1] ), .B(\shift[0] ), .C(new_n355_), .Y(new_n831_));
  NOR3X1   g0568(.A(new_n267_), .B(\shift[0] ), .C(new_n366_), .Y(new_n832_));
  NOR3X1   g0569(.A(new_n267_), .B(new_n266_), .C(new_n368_), .Y(new_n833_));
  OR4X1    g0570(.A(new_n833_), .B(new_n832_), .C(new_n831_), .D(new_n830_), .Y(new_n834_));
  AOI22X1  g0571(.A0(new_n834_), .A1(new_n287_), .B0(new_n829_), .B1(new_n276_), .Y(new_n835_));
  NOR3X1   g0572(.A(\shift[1] ), .B(new_n266_), .C(new_n381_), .Y(new_n836_));
  NOR3X1   g0573(.A(\shift[1] ), .B(\shift[0] ), .C(new_n383_), .Y(new_n837_));
  NOR3X1   g0574(.A(new_n267_), .B(\shift[0] ), .C(new_n376_), .Y(new_n838_));
  NOR3X1   g0575(.A(new_n267_), .B(new_n266_), .C(new_n378_), .Y(new_n839_));
  OR4X1    g0576(.A(new_n839_), .B(new_n838_), .C(new_n837_), .D(new_n836_), .Y(new_n840_));
  NOR3X1   g0577(.A(\shift[1] ), .B(new_n266_), .C(new_n362_), .Y(new_n841_));
  NOR3X1   g0578(.A(\shift[1] ), .B(\shift[0] ), .C(new_n364_), .Y(new_n842_));
  NOR3X1   g0579(.A(new_n267_), .B(\shift[0] ), .C(new_n385_), .Y(new_n843_));
  NOR3X1   g0580(.A(new_n267_), .B(new_n266_), .C(new_n387_), .Y(new_n844_));
  OR4X1    g0581(.A(new_n844_), .B(new_n843_), .C(new_n842_), .D(new_n841_), .Y(new_n845_));
  AOI22X1  g0582(.A0(new_n845_), .A1(new_n308_), .B0(new_n840_), .B1(new_n298_), .Y(new_n846_));
  AOI21X1  g0583(.A0(new_n846_), .A1(new_n835_), .B0(new_n391_), .Y(new_n847_));
  NOR3X1   g0584(.A(\shift[1] ), .B(new_n266_), .C(new_n372_), .Y(new_n848_));
  NOR3X1   g0585(.A(\shift[1] ), .B(\shift[0] ), .C(new_n374_), .Y(new_n849_));
  NOR3X1   g0586(.A(new_n267_), .B(\shift[0] ), .C(new_n397_), .Y(new_n850_));
  NOR3X1   g0587(.A(new_n267_), .B(new_n266_), .C(new_n399_), .Y(new_n851_));
  OR4X1    g0588(.A(new_n851_), .B(new_n850_), .C(new_n849_), .D(new_n848_), .Y(new_n852_));
  NOR3X1   g0589(.A(\shift[1] ), .B(new_n266_), .C(new_n393_), .Y(new_n853_));
  NOR3X1   g0590(.A(\shift[1] ), .B(\shift[0] ), .C(new_n395_), .Y(new_n854_));
  NOR3X1   g0591(.A(new_n267_), .B(\shift[0] ), .C(new_n406_), .Y(new_n855_));
  NOR3X1   g0592(.A(new_n267_), .B(new_n266_), .C(new_n408_), .Y(new_n856_));
  OR4X1    g0593(.A(new_n856_), .B(new_n855_), .C(new_n854_), .D(new_n853_), .Y(new_n857_));
  AOI22X1  g0594(.A0(new_n857_), .A1(new_n287_), .B0(new_n852_), .B1(new_n276_), .Y(new_n858_));
  NOR3X1   g0595(.A(\shift[1] ), .B(new_n266_), .C(new_n421_), .Y(new_n859_));
  NOR3X1   g0596(.A(\shift[1] ), .B(\shift[0] ), .C(new_n423_), .Y(new_n860_));
  NOR3X1   g0597(.A(new_n267_), .B(\shift[0] ), .C(new_n416_), .Y(new_n861_));
  NOR3X1   g0598(.A(new_n267_), .B(new_n266_), .C(new_n418_), .Y(new_n862_));
  OR4X1    g0599(.A(new_n862_), .B(new_n861_), .C(new_n860_), .D(new_n859_), .Y(new_n863_));
  NOR3X1   g0600(.A(\shift[1] ), .B(new_n266_), .C(new_n402_), .Y(new_n864_));
  NOR3X1   g0601(.A(\shift[1] ), .B(\shift[0] ), .C(new_n404_), .Y(new_n865_));
  NOR3X1   g0602(.A(new_n267_), .B(\shift[0] ), .C(new_n425_), .Y(new_n866_));
  NOR3X1   g0603(.A(new_n267_), .B(new_n266_), .C(new_n427_), .Y(new_n867_));
  OR4X1    g0604(.A(new_n867_), .B(new_n866_), .C(new_n865_), .D(new_n864_), .Y(new_n868_));
  AOI22X1  g0605(.A0(new_n868_), .A1(new_n308_), .B0(new_n863_), .B1(new_n298_), .Y(new_n869_));
  AOI21X1  g0606(.A0(new_n869_), .A1(new_n858_), .B0(new_n431_), .Y(new_n870_));
  OR4X1    g0607(.A(new_n870_), .B(new_n847_), .C(new_n824_), .D(new_n801_), .Y(new_n871_));
  NOR3X1   g0608(.A(\shift[1] ), .B(new_n266_), .C(new_n289_), .Y(new_n872_));
  NOR3X1   g0609(.A(\shift[1] ), .B(\shift[0] ), .C(new_n291_), .Y(new_n873_));
  NOR3X1   g0610(.A(new_n267_), .B(\shift[0] ), .C(new_n516_), .Y(new_n874_));
  NOR3X1   g0611(.A(new_n267_), .B(new_n266_), .C(new_n518_), .Y(new_n875_));
  OR4X1    g0612(.A(new_n875_), .B(new_n874_), .C(new_n873_), .D(new_n872_), .Y(new_n876_));
  NOR3X1   g0613(.A(\shift[1] ), .B(new_n266_), .C(new_n512_), .Y(new_n877_));
  NOR3X1   g0614(.A(\shift[1] ), .B(\shift[0] ), .C(new_n514_), .Y(new_n878_));
  NOR3X1   g0615(.A(new_n267_), .B(\shift[0] ), .C(new_n525_), .Y(new_n879_));
  NOR3X1   g0616(.A(new_n267_), .B(new_n266_), .C(new_n527_), .Y(new_n880_));
  OR4X1    g0617(.A(new_n880_), .B(new_n879_), .C(new_n878_), .D(new_n877_), .Y(new_n881_));
  AOI22X1  g0618(.A0(new_n881_), .A1(new_n287_), .B0(new_n876_), .B1(new_n276_), .Y(new_n882_));
  NOR3X1   g0619(.A(\shift[1] ), .B(new_n266_), .C(new_n540_), .Y(new_n883_));
  NOR3X1   g0620(.A(\shift[1] ), .B(\shift[0] ), .C(new_n542_), .Y(new_n884_));
  NOR3X1   g0621(.A(new_n267_), .B(\shift[0] ), .C(new_n535_), .Y(new_n885_));
  NOR3X1   g0622(.A(new_n267_), .B(new_n266_), .C(new_n537_), .Y(new_n886_));
  OR4X1    g0623(.A(new_n886_), .B(new_n885_), .C(new_n884_), .D(new_n883_), .Y(new_n887_));
  NOR3X1   g0624(.A(\shift[1] ), .B(new_n266_), .C(new_n521_), .Y(new_n888_));
  NOR3X1   g0625(.A(\shift[1] ), .B(\shift[0] ), .C(new_n523_), .Y(new_n889_));
  NOR3X1   g0626(.A(new_n267_), .B(\shift[0] ), .C(new_n544_), .Y(new_n890_));
  NOR3X1   g0627(.A(new_n267_), .B(new_n266_), .C(new_n546_), .Y(new_n891_));
  OR4X1    g0628(.A(new_n891_), .B(new_n890_), .C(new_n889_), .D(new_n888_), .Y(new_n892_));
  AOI22X1  g0629(.A0(new_n892_), .A1(new_n308_), .B0(new_n887_), .B1(new_n298_), .Y(new_n893_));
  AOI21X1  g0630(.A0(new_n893_), .A1(new_n882_), .B0(new_n391_), .Y(new_n894_));
  NOR3X1   g0631(.A(\shift[1] ), .B(new_n266_), .C(new_n492_), .Y(new_n895_));
  NOR3X1   g0632(.A(\shift[1] ), .B(\shift[0] ), .C(new_n494_), .Y(new_n896_));
  NOR3X1   g0633(.A(new_n267_), .B(\shift[0] ), .C(new_n438_), .Y(new_n897_));
  NOR3X1   g0634(.A(new_n267_), .B(new_n266_), .C(new_n440_), .Y(new_n898_));
  OR4X1    g0635(.A(new_n898_), .B(new_n897_), .C(new_n896_), .D(new_n895_), .Y(new_n899_));
  NOR3X1   g0636(.A(\shift[1] ), .B(new_n266_), .C(new_n434_), .Y(new_n900_));
  NOR3X1   g0637(.A(\shift[1] ), .B(\shift[0] ), .C(new_n436_), .Y(new_n901_));
  NOR3X1   g0638(.A(new_n267_), .B(\shift[0] ), .C(new_n447_), .Y(new_n902_));
  NOR3X1   g0639(.A(new_n267_), .B(new_n266_), .C(new_n449_), .Y(new_n903_));
  OR4X1    g0640(.A(new_n903_), .B(new_n902_), .C(new_n901_), .D(new_n900_), .Y(new_n904_));
  AOI22X1  g0641(.A0(new_n904_), .A1(new_n287_), .B0(new_n899_), .B1(new_n276_), .Y(new_n905_));
  NOR3X1   g0642(.A(\shift[1] ), .B(new_n266_), .C(new_n462_), .Y(new_n906_));
  NOR3X1   g0643(.A(\shift[1] ), .B(\shift[0] ), .C(new_n464_), .Y(new_n907_));
  NOR3X1   g0644(.A(new_n267_), .B(\shift[0] ), .C(new_n457_), .Y(new_n908_));
  NOR3X1   g0645(.A(new_n267_), .B(new_n266_), .C(new_n459_), .Y(new_n909_));
  OR4X1    g0646(.A(new_n909_), .B(new_n908_), .C(new_n907_), .D(new_n906_), .Y(new_n910_));
  NOR3X1   g0647(.A(\shift[1] ), .B(new_n266_), .C(new_n443_), .Y(new_n911_));
  NOR3X1   g0648(.A(\shift[1] ), .B(\shift[0] ), .C(new_n445_), .Y(new_n912_));
  NOR3X1   g0649(.A(new_n267_), .B(\shift[0] ), .C(new_n466_), .Y(new_n913_));
  NOR3X1   g0650(.A(new_n267_), .B(new_n266_), .C(new_n468_), .Y(new_n914_));
  OR4X1    g0651(.A(new_n914_), .B(new_n913_), .C(new_n912_), .D(new_n911_), .Y(new_n915_));
  AOI22X1  g0652(.A0(new_n915_), .A1(new_n308_), .B0(new_n910_), .B1(new_n298_), .Y(new_n916_));
  AOI21X1  g0653(.A0(new_n916_), .A1(new_n905_), .B0(new_n310_), .Y(new_n917_));
  NOR3X1   g0654(.A(\shift[1] ), .B(new_n266_), .C(new_n531_), .Y(new_n918_));
  NOR3X1   g0655(.A(\shift[1] ), .B(\shift[0] ), .C(new_n533_), .Y(new_n919_));
  NOR3X1   g0656(.A(new_n267_), .B(\shift[0] ), .C(new_n555_), .Y(new_n920_));
  NOR3X1   g0657(.A(new_n267_), .B(new_n266_), .C(new_n557_), .Y(new_n921_));
  OR4X1    g0658(.A(new_n921_), .B(new_n920_), .C(new_n919_), .D(new_n918_), .Y(new_n922_));
  NOR3X1   g0659(.A(new_n267_), .B(new_n266_), .C(new_n566_), .Y(new_n923_));
  NOR3X1   g0660(.A(new_n267_), .B(\shift[0] ), .C(new_n564_), .Y(new_n924_));
  NOR3X1   g0661(.A(\shift[1] ), .B(\shift[0] ), .C(new_n553_), .Y(new_n925_));
  NOR3X1   g0662(.A(\shift[1] ), .B(new_n266_), .C(new_n551_), .Y(new_n926_));
  OR4X1    g0663(.A(new_n926_), .B(new_n925_), .C(new_n924_), .D(new_n923_), .Y(new_n927_));
  AOI22X1  g0664(.A0(new_n927_), .A1(new_n287_), .B0(new_n922_), .B1(new_n276_), .Y(new_n928_));
  NOR3X1   g0665(.A(\shift[1] ), .B(new_n266_), .C(new_n581_), .Y(new_n929_));
  NOR3X1   g0666(.A(\shift[1] ), .B(\shift[0] ), .C(new_n585_), .Y(new_n930_));
  NOR3X1   g0667(.A(new_n267_), .B(\shift[0] ), .C(new_n574_), .Y(new_n931_));
  NOR3X1   g0668(.A(new_n267_), .B(new_n266_), .C(new_n576_), .Y(new_n932_));
  OR4X1    g0669(.A(new_n932_), .B(new_n931_), .C(new_n930_), .D(new_n929_), .Y(new_n933_));
  NOR3X1   g0670(.A(\shift[1] ), .B(new_n266_), .C(new_n560_), .Y(new_n934_));
  NOR3X1   g0671(.A(\shift[1] ), .B(\shift[0] ), .C(new_n562_), .Y(new_n935_));
  NOR3X1   g0672(.A(new_n267_), .B(new_n266_), .C(new_n583_), .Y(new_n936_));
  NOR3X1   g0673(.A(new_n267_), .B(\shift[0] ), .C(new_n579_), .Y(new_n937_));
  OR4X1    g0674(.A(new_n937_), .B(new_n936_), .C(new_n935_), .D(new_n934_), .Y(new_n938_));
  AOI22X1  g0675(.A0(new_n938_), .A1(new_n308_), .B0(new_n933_), .B1(new_n298_), .Y(new_n939_));
  AOI21X1  g0676(.A0(new_n939_), .A1(new_n928_), .B0(new_n431_), .Y(new_n940_));
  NOR3X1   g0677(.A(\shift[1] ), .B(new_n266_), .C(new_n570_), .Y(new_n941_));
  NOR3X1   g0678(.A(\shift[1] ), .B(\shift[0] ), .C(new_n572_), .Y(new_n942_));
  NOR3X1   g0679(.A(new_n267_), .B(\shift[0] ), .C(new_n477_), .Y(new_n943_));
  NOR3X1   g0680(.A(new_n267_), .B(new_n266_), .C(new_n479_), .Y(new_n944_));
  OR4X1    g0681(.A(new_n944_), .B(new_n943_), .C(new_n942_), .D(new_n941_), .Y(new_n945_));
  NOR3X1   g0682(.A(\shift[1] ), .B(new_n266_), .C(new_n473_), .Y(new_n946_));
  NOR3X1   g0683(.A(\shift[1] ), .B(\shift[0] ), .C(new_n475_), .Y(new_n947_));
  NOR3X1   g0684(.A(new_n267_), .B(\shift[0] ), .C(new_n486_), .Y(new_n948_));
  NOR3X1   g0685(.A(new_n267_), .B(new_n266_), .C(new_n488_), .Y(new_n949_));
  OR4X1    g0686(.A(new_n949_), .B(new_n948_), .C(new_n947_), .D(new_n946_), .Y(new_n950_));
  AOI22X1  g0687(.A0(new_n950_), .A1(new_n287_), .B0(new_n945_), .B1(new_n276_), .Y(new_n951_));
  NOR3X1   g0688(.A(\shift[1] ), .B(new_n266_), .C(new_n501_), .Y(new_n952_));
  NOR3X1   g0689(.A(\shift[1] ), .B(\shift[0] ), .C(new_n503_), .Y(new_n953_));
  NOR3X1   g0690(.A(new_n267_), .B(\shift[0] ), .C(new_n496_), .Y(new_n954_));
  NOR3X1   g0691(.A(new_n267_), .B(new_n266_), .C(new_n498_), .Y(new_n955_));
  OR4X1    g0692(.A(new_n955_), .B(new_n954_), .C(new_n953_), .D(new_n952_), .Y(new_n956_));
  NOR3X1   g0693(.A(\shift[1] ), .B(new_n266_), .C(new_n482_), .Y(new_n957_));
  NOR3X1   g0694(.A(\shift[1] ), .B(\shift[0] ), .C(new_n484_), .Y(new_n958_));
  NOR3X1   g0695(.A(new_n267_), .B(\shift[0] ), .C(new_n505_), .Y(new_n959_));
  NOR3X1   g0696(.A(new_n267_), .B(new_n266_), .C(new_n507_), .Y(new_n960_));
  OR4X1    g0697(.A(new_n960_), .B(new_n959_), .C(new_n958_), .D(new_n957_), .Y(new_n961_));
  AOI22X1  g0698(.A0(new_n961_), .A1(new_n308_), .B0(new_n956_), .B1(new_n298_), .Y(new_n962_));
  AOI21X1  g0699(.A0(new_n962_), .A1(new_n951_), .B0(new_n351_), .Y(new_n963_));
  OR4X1    g0700(.A(new_n963_), .B(new_n940_), .C(new_n917_), .D(new_n894_), .Y(new_n964_));
  MX2X1    g0701(.A(new_n964_), .B(new_n871_), .S0(new_n264_), .Y(\result[2] ));
  NOR3X1   g0702(.A(new_n267_), .B(\shift[0] ), .C(new_n372_), .Y(new_n966_));
  NOR3X1   g0703(.A(\shift[1] ), .B(new_n266_), .C(new_n374_), .Y(new_n967_));
  NOR3X1   g0704(.A(new_n267_), .B(new_n266_), .C(new_n397_), .Y(new_n968_));
  NOR3X1   g0705(.A(\shift[1] ), .B(\shift[0] ), .C(new_n378_), .Y(new_n969_));
  OR4X1    g0706(.A(new_n969_), .B(new_n968_), .C(new_n967_), .D(new_n966_), .Y(new_n970_));
  NOR3X1   g0707(.A(new_n267_), .B(\shift[0] ), .C(new_n393_), .Y(new_n971_));
  NOR3X1   g0708(.A(\shift[1] ), .B(new_n266_), .C(new_n395_), .Y(new_n972_));
  NOR3X1   g0709(.A(new_n267_), .B(new_n266_), .C(new_n406_), .Y(new_n973_));
  NOR3X1   g0710(.A(\shift[1] ), .B(\shift[0] ), .C(new_n399_), .Y(new_n974_));
  OR4X1    g0711(.A(new_n974_), .B(new_n973_), .C(new_n972_), .D(new_n971_), .Y(new_n975_));
  AOI22X1  g0712(.A0(new_n975_), .A1(new_n287_), .B0(new_n970_), .B1(new_n276_), .Y(new_n976_));
  NOR3X1   g0713(.A(new_n267_), .B(\shift[0] ), .C(new_n421_), .Y(new_n977_));
  NOR3X1   g0714(.A(\shift[1] ), .B(new_n266_), .C(new_n423_), .Y(new_n978_));
  NOR3X1   g0715(.A(new_n267_), .B(new_n266_), .C(new_n416_), .Y(new_n979_));
  NOR3X1   g0716(.A(\shift[1] ), .B(\shift[0] ), .C(new_n427_), .Y(new_n980_));
  OR4X1    g0717(.A(new_n980_), .B(new_n979_), .C(new_n978_), .D(new_n977_), .Y(new_n981_));
  NOR3X1   g0718(.A(new_n267_), .B(\shift[0] ), .C(new_n402_), .Y(new_n982_));
  NOR3X1   g0719(.A(\shift[1] ), .B(new_n266_), .C(new_n404_), .Y(new_n983_));
  NOR3X1   g0720(.A(new_n267_), .B(new_n266_), .C(new_n425_), .Y(new_n984_));
  NOR3X1   g0721(.A(\shift[1] ), .B(\shift[0] ), .C(new_n408_), .Y(new_n985_));
  OR4X1    g0722(.A(new_n985_), .B(new_n984_), .C(new_n983_), .D(new_n982_), .Y(new_n986_));
  AOI22X1  g0723(.A0(new_n986_), .A1(new_n308_), .B0(new_n981_), .B1(new_n298_), .Y(new_n987_));
  AOI21X1  g0724(.A0(new_n987_), .A1(new_n976_), .B0(new_n431_), .Y(new_n988_));
  NOR3X1   g0725(.A(new_n267_), .B(\shift[0] ), .C(new_n412_), .Y(new_n989_));
  NOR3X1   g0726(.A(\shift[1] ), .B(new_n266_), .C(new_n414_), .Y(new_n990_));
  NOR3X1   g0727(.A(new_n267_), .B(new_n266_), .C(new_n316_), .Y(new_n991_));
  NOR3X1   g0728(.A(\shift[1] ), .B(\shift[0] ), .C(new_n418_), .Y(new_n992_));
  OR4X1    g0729(.A(new_n992_), .B(new_n991_), .C(new_n990_), .D(new_n989_), .Y(new_n993_));
  NOR3X1   g0730(.A(new_n267_), .B(\shift[0] ), .C(new_n312_), .Y(new_n994_));
  NOR3X1   g0731(.A(\shift[1] ), .B(new_n266_), .C(new_n314_), .Y(new_n995_));
  NOR3X1   g0732(.A(new_n267_), .B(new_n266_), .C(new_n325_), .Y(new_n996_));
  NOR3X1   g0733(.A(\shift[1] ), .B(\shift[0] ), .C(new_n318_), .Y(new_n997_));
  OR4X1    g0734(.A(new_n997_), .B(new_n996_), .C(new_n995_), .D(new_n994_), .Y(new_n998_));
  AOI22X1  g0735(.A0(new_n998_), .A1(new_n287_), .B0(new_n993_), .B1(new_n276_), .Y(new_n999_));
  NOR3X1   g0736(.A(new_n267_), .B(\shift[0] ), .C(new_n340_), .Y(new_n1000_));
  NOR3X1   g0737(.A(\shift[1] ), .B(new_n266_), .C(new_n342_), .Y(new_n1001_));
  NOR3X1   g0738(.A(new_n267_), .B(new_n266_), .C(new_n335_), .Y(new_n1002_));
  NOR3X1   g0739(.A(\shift[1] ), .B(\shift[0] ), .C(new_n346_), .Y(new_n1003_));
  OR4X1    g0740(.A(new_n1003_), .B(new_n1002_), .C(new_n1001_), .D(new_n1000_), .Y(new_n1004_));
  NOR3X1   g0741(.A(new_n267_), .B(\shift[0] ), .C(new_n321_), .Y(new_n1005_));
  NOR3X1   g0742(.A(\shift[1] ), .B(new_n266_), .C(new_n323_), .Y(new_n1006_));
  NOR3X1   g0743(.A(new_n267_), .B(new_n266_), .C(new_n344_), .Y(new_n1007_));
  NOR3X1   g0744(.A(\shift[1] ), .B(\shift[0] ), .C(new_n327_), .Y(new_n1008_));
  OR4X1    g0745(.A(new_n1008_), .B(new_n1007_), .C(new_n1006_), .D(new_n1005_), .Y(new_n1009_));
  AOI22X1  g0746(.A0(new_n1009_), .A1(new_n308_), .B0(new_n1004_), .B1(new_n298_), .Y(new_n1010_));
  AOI21X1  g0747(.A0(new_n1010_), .A1(new_n999_), .B0(new_n351_), .Y(new_n1011_));
  NOR3X1   g0748(.A(new_n267_), .B(\shift[0] ), .C(new_n453_), .Y(new_n1012_));
  NOR3X1   g0749(.A(\shift[1] ), .B(new_n266_), .C(new_n455_), .Y(new_n1013_));
  NOR3X1   g0750(.A(new_n267_), .B(new_n266_), .C(new_n357_), .Y(new_n1014_));
  NOR3X1   g0751(.A(\shift[1] ), .B(\shift[0] ), .C(new_n459_), .Y(new_n1015_));
  OR4X1    g0752(.A(new_n1015_), .B(new_n1014_), .C(new_n1013_), .D(new_n1012_), .Y(new_n1016_));
  NOR3X1   g0753(.A(new_n267_), .B(\shift[0] ), .C(new_n353_), .Y(new_n1017_));
  NOR3X1   g0754(.A(\shift[1] ), .B(new_n266_), .C(new_n355_), .Y(new_n1018_));
  NOR3X1   g0755(.A(new_n267_), .B(new_n266_), .C(new_n366_), .Y(new_n1019_));
  NOR3X1   g0756(.A(\shift[1] ), .B(\shift[0] ), .C(new_n359_), .Y(new_n1020_));
  OR4X1    g0757(.A(new_n1020_), .B(new_n1019_), .C(new_n1018_), .D(new_n1017_), .Y(new_n1021_));
  AOI22X1  g0758(.A0(new_n1021_), .A1(new_n287_), .B0(new_n1016_), .B1(new_n276_), .Y(new_n1022_));
  NOR3X1   g0759(.A(new_n267_), .B(\shift[0] ), .C(new_n381_), .Y(new_n1023_));
  NOR3X1   g0760(.A(\shift[1] ), .B(new_n266_), .C(new_n383_), .Y(new_n1024_));
  NOR3X1   g0761(.A(new_n267_), .B(new_n266_), .C(new_n376_), .Y(new_n1025_));
  NOR3X1   g0762(.A(\shift[1] ), .B(\shift[0] ), .C(new_n387_), .Y(new_n1026_));
  OR4X1    g0763(.A(new_n1026_), .B(new_n1025_), .C(new_n1024_), .D(new_n1023_), .Y(new_n1027_));
  NOR3X1   g0764(.A(new_n267_), .B(\shift[0] ), .C(new_n362_), .Y(new_n1028_));
  NOR3X1   g0765(.A(\shift[1] ), .B(new_n266_), .C(new_n364_), .Y(new_n1029_));
  NOR3X1   g0766(.A(new_n267_), .B(new_n266_), .C(new_n385_), .Y(new_n1030_));
  NOR3X1   g0767(.A(\shift[1] ), .B(\shift[0] ), .C(new_n368_), .Y(new_n1031_));
  OR4X1    g0768(.A(new_n1031_), .B(new_n1030_), .C(new_n1029_), .D(new_n1028_), .Y(new_n1032_));
  AOI22X1  g0769(.A0(new_n1032_), .A1(new_n308_), .B0(new_n1027_), .B1(new_n298_), .Y(new_n1033_));
  AOI21X1  g0770(.A0(new_n1033_), .A1(new_n1022_), .B0(new_n391_), .Y(new_n1034_));
  NOR3X1   g0771(.A(new_n267_), .B(\shift[0] ), .C(new_n331_), .Y(new_n1035_));
  NOR3X1   g0772(.A(\shift[1] ), .B(new_n266_), .C(new_n333_), .Y(new_n1036_));
  NOR3X1   g0773(.A(new_n267_), .B(new_n266_), .C(new_n271_), .Y(new_n1037_));
  NOR3X1   g0774(.A(\shift[1] ), .B(\shift[0] ), .C(new_n337_), .Y(new_n1038_));
  OR4X1    g0775(.A(new_n1038_), .B(new_n1037_), .C(new_n1036_), .D(new_n1035_), .Y(new_n1039_));
  NOR3X1   g0776(.A(new_n267_), .B(\shift[0] ), .C(new_n265_), .Y(new_n1040_));
  NOR3X1   g0777(.A(\shift[1] ), .B(new_n266_), .C(new_n269_), .Y(new_n1041_));
  NOR3X1   g0778(.A(new_n267_), .B(new_n266_), .C(new_n281_), .Y(new_n1042_));
  NOR3X1   g0779(.A(\shift[1] ), .B(\shift[0] ), .C(new_n273_), .Y(new_n1043_));
  OR4X1    g0780(.A(new_n1043_), .B(new_n1042_), .C(new_n1041_), .D(new_n1040_), .Y(new_n1044_));
  AOI22X1  g0781(.A0(new_n1044_), .A1(new_n287_), .B0(new_n1039_), .B1(new_n276_), .Y(new_n1045_));
  NOR3X1   g0782(.A(new_n267_), .B(\shift[0] ), .C(new_n299_), .Y(new_n1046_));
  NOR3X1   g0783(.A(\shift[1] ), .B(new_n266_), .C(new_n301_), .Y(new_n1047_));
  NOR3X1   g0784(.A(new_n267_), .B(new_n266_), .C(new_n293_), .Y(new_n1048_));
  NOR3X1   g0785(.A(\shift[1] ), .B(\shift[0] ), .C(new_n305_), .Y(new_n1049_));
  OR4X1    g0786(.A(new_n1049_), .B(new_n1048_), .C(new_n1047_), .D(new_n1046_), .Y(new_n1050_));
  NOR3X1   g0787(.A(new_n267_), .B(\shift[0] ), .C(new_n277_), .Y(new_n1051_));
  NOR3X1   g0788(.A(\shift[1] ), .B(new_n266_), .C(new_n279_), .Y(new_n1052_));
  NOR3X1   g0789(.A(new_n267_), .B(new_n266_), .C(new_n303_), .Y(new_n1053_));
  NOR3X1   g0790(.A(\shift[1] ), .B(\shift[0] ), .C(new_n283_), .Y(new_n1054_));
  OR4X1    g0791(.A(new_n1054_), .B(new_n1053_), .C(new_n1052_), .D(new_n1051_), .Y(new_n1055_));
  AOI22X1  g0792(.A0(new_n1055_), .A1(new_n308_), .B0(new_n1050_), .B1(new_n298_), .Y(new_n1056_));
  AOI21X1  g0793(.A0(new_n1056_), .A1(new_n1045_), .B0(new_n310_), .Y(new_n1057_));
  OR4X1    g0794(.A(new_n1057_), .B(new_n1034_), .C(new_n1011_), .D(new_n988_), .Y(new_n1058_));
  NOR3X1   g0795(.A(new_n267_), .B(\shift[0] ), .C(new_n289_), .Y(new_n1059_));
  NOR3X1   g0796(.A(\shift[1] ), .B(new_n266_), .C(new_n291_), .Y(new_n1060_));
  NOR3X1   g0797(.A(new_n267_), .B(new_n266_), .C(new_n516_), .Y(new_n1061_));
  NOR3X1   g0798(.A(\shift[1] ), .B(\shift[0] ), .C(new_n295_), .Y(new_n1062_));
  OR4X1    g0799(.A(new_n1062_), .B(new_n1061_), .C(new_n1060_), .D(new_n1059_), .Y(new_n1063_));
  NOR3X1   g0800(.A(new_n267_), .B(\shift[0] ), .C(new_n512_), .Y(new_n1064_));
  NOR3X1   g0801(.A(\shift[1] ), .B(new_n266_), .C(new_n514_), .Y(new_n1065_));
  NOR3X1   g0802(.A(new_n267_), .B(new_n266_), .C(new_n525_), .Y(new_n1066_));
  NOR3X1   g0803(.A(\shift[1] ), .B(\shift[0] ), .C(new_n518_), .Y(new_n1067_));
  OR4X1    g0804(.A(new_n1067_), .B(new_n1066_), .C(new_n1065_), .D(new_n1064_), .Y(new_n1068_));
  AOI22X1  g0805(.A0(new_n1068_), .A1(new_n287_), .B0(new_n1063_), .B1(new_n276_), .Y(new_n1069_));
  NOR3X1   g0806(.A(new_n267_), .B(\shift[0] ), .C(new_n540_), .Y(new_n1070_));
  NOR3X1   g0807(.A(\shift[1] ), .B(new_n266_), .C(new_n542_), .Y(new_n1071_));
  NOR3X1   g0808(.A(new_n267_), .B(new_n266_), .C(new_n535_), .Y(new_n1072_));
  NOR3X1   g0809(.A(\shift[1] ), .B(\shift[0] ), .C(new_n546_), .Y(new_n1073_));
  OR4X1    g0810(.A(new_n1073_), .B(new_n1072_), .C(new_n1071_), .D(new_n1070_), .Y(new_n1074_));
  NOR3X1   g0811(.A(new_n267_), .B(\shift[0] ), .C(new_n521_), .Y(new_n1075_));
  NOR3X1   g0812(.A(\shift[1] ), .B(new_n266_), .C(new_n523_), .Y(new_n1076_));
  NOR3X1   g0813(.A(new_n267_), .B(new_n266_), .C(new_n544_), .Y(new_n1077_));
  NOR3X1   g0814(.A(\shift[1] ), .B(\shift[0] ), .C(new_n527_), .Y(new_n1078_));
  OR4X1    g0815(.A(new_n1078_), .B(new_n1077_), .C(new_n1076_), .D(new_n1075_), .Y(new_n1079_));
  AOI22X1  g0816(.A0(new_n1079_), .A1(new_n308_), .B0(new_n1074_), .B1(new_n298_), .Y(new_n1080_));
  AOI21X1  g0817(.A0(new_n1080_), .A1(new_n1069_), .B0(new_n391_), .Y(new_n1081_));
  NOR3X1   g0818(.A(new_n267_), .B(\shift[0] ), .C(new_n531_), .Y(new_n1082_));
  NOR3X1   g0819(.A(\shift[1] ), .B(new_n266_), .C(new_n533_), .Y(new_n1083_));
  NOR3X1   g0820(.A(new_n267_), .B(new_n266_), .C(new_n555_), .Y(new_n1084_));
  NOR3X1   g0821(.A(\shift[1] ), .B(\shift[0] ), .C(new_n537_), .Y(new_n1085_));
  OR4X1    g0822(.A(new_n1085_), .B(new_n1084_), .C(new_n1083_), .D(new_n1082_), .Y(new_n1086_));
  NOR3X1   g0823(.A(new_n267_), .B(new_n266_), .C(new_n564_), .Y(new_n1087_));
  NOR3X1   g0824(.A(new_n267_), .B(\shift[0] ), .C(new_n551_), .Y(new_n1088_));
  NOR3X1   g0825(.A(\shift[1] ), .B(\shift[0] ), .C(new_n557_), .Y(new_n1089_));
  NOR3X1   g0826(.A(\shift[1] ), .B(new_n266_), .C(new_n553_), .Y(new_n1090_));
  OR4X1    g0827(.A(new_n1090_), .B(new_n1089_), .C(new_n1088_), .D(new_n1087_), .Y(new_n1091_));
  AOI22X1  g0828(.A0(new_n1091_), .A1(new_n287_), .B0(new_n1086_), .B1(new_n276_), .Y(new_n1092_));
  NOR3X1   g0829(.A(new_n267_), .B(\shift[0] ), .C(new_n581_), .Y(new_n1093_));
  NOR3X1   g0830(.A(\shift[1] ), .B(new_n266_), .C(new_n585_), .Y(new_n1094_));
  NOR3X1   g0831(.A(new_n267_), .B(new_n266_), .C(new_n574_), .Y(new_n1095_));
  NOR3X1   g0832(.A(\shift[1] ), .B(\shift[0] ), .C(new_n583_), .Y(new_n1096_));
  OR4X1    g0833(.A(new_n1096_), .B(new_n1095_), .C(new_n1094_), .D(new_n1093_), .Y(new_n1097_));
  NOR3X1   g0834(.A(new_n267_), .B(\shift[0] ), .C(new_n560_), .Y(new_n1098_));
  NOR3X1   g0835(.A(\shift[1] ), .B(new_n266_), .C(new_n562_), .Y(new_n1099_));
  NOR3X1   g0836(.A(new_n267_), .B(new_n266_), .C(new_n579_), .Y(new_n1100_));
  NOR3X1   g0837(.A(\shift[1] ), .B(\shift[0] ), .C(new_n566_), .Y(new_n1101_));
  OR4X1    g0838(.A(new_n1101_), .B(new_n1100_), .C(new_n1099_), .D(new_n1098_), .Y(new_n1102_));
  AOI22X1  g0839(.A0(new_n1102_), .A1(new_n308_), .B0(new_n1097_), .B1(new_n298_), .Y(new_n1103_));
  AOI21X1  g0840(.A0(new_n1103_), .A1(new_n1092_), .B0(new_n431_), .Y(new_n1104_));
  NOR3X1   g0841(.A(new_n267_), .B(\shift[0] ), .C(new_n492_), .Y(new_n1105_));
  NOR3X1   g0842(.A(\shift[1] ), .B(new_n266_), .C(new_n494_), .Y(new_n1106_));
  NOR3X1   g0843(.A(new_n267_), .B(new_n266_), .C(new_n438_), .Y(new_n1107_));
  NOR3X1   g0844(.A(\shift[1] ), .B(\shift[0] ), .C(new_n498_), .Y(new_n1108_));
  OR4X1    g0845(.A(new_n1108_), .B(new_n1107_), .C(new_n1106_), .D(new_n1105_), .Y(new_n1109_));
  NOR3X1   g0846(.A(new_n267_), .B(\shift[0] ), .C(new_n434_), .Y(new_n1110_));
  NOR3X1   g0847(.A(\shift[1] ), .B(new_n266_), .C(new_n436_), .Y(new_n1111_));
  NOR3X1   g0848(.A(new_n267_), .B(new_n266_), .C(new_n447_), .Y(new_n1112_));
  NOR3X1   g0849(.A(\shift[1] ), .B(\shift[0] ), .C(new_n440_), .Y(new_n1113_));
  OR4X1    g0850(.A(new_n1113_), .B(new_n1112_), .C(new_n1111_), .D(new_n1110_), .Y(new_n1114_));
  AOI22X1  g0851(.A0(new_n1114_), .A1(new_n287_), .B0(new_n1109_), .B1(new_n276_), .Y(new_n1115_));
  NOR3X1   g0852(.A(new_n267_), .B(\shift[0] ), .C(new_n462_), .Y(new_n1116_));
  NOR3X1   g0853(.A(\shift[1] ), .B(new_n266_), .C(new_n464_), .Y(new_n1117_));
  NOR3X1   g0854(.A(new_n267_), .B(new_n266_), .C(new_n457_), .Y(new_n1118_));
  NOR3X1   g0855(.A(\shift[1] ), .B(\shift[0] ), .C(new_n468_), .Y(new_n1119_));
  OR4X1    g0856(.A(new_n1119_), .B(new_n1118_), .C(new_n1117_), .D(new_n1116_), .Y(new_n1120_));
  NOR3X1   g0857(.A(new_n267_), .B(\shift[0] ), .C(new_n443_), .Y(new_n1121_));
  NOR3X1   g0858(.A(\shift[1] ), .B(new_n266_), .C(new_n445_), .Y(new_n1122_));
  NOR3X1   g0859(.A(new_n267_), .B(new_n266_), .C(new_n466_), .Y(new_n1123_));
  NOR3X1   g0860(.A(\shift[1] ), .B(\shift[0] ), .C(new_n449_), .Y(new_n1124_));
  OR4X1    g0861(.A(new_n1124_), .B(new_n1123_), .C(new_n1122_), .D(new_n1121_), .Y(new_n1125_));
  AOI22X1  g0862(.A0(new_n1125_), .A1(new_n308_), .B0(new_n1120_), .B1(new_n298_), .Y(new_n1126_));
  AOI21X1  g0863(.A0(new_n1126_), .A1(new_n1115_), .B0(new_n310_), .Y(new_n1127_));
  NOR3X1   g0864(.A(new_n267_), .B(\shift[0] ), .C(new_n570_), .Y(new_n1128_));
  NOR3X1   g0865(.A(\shift[1] ), .B(new_n266_), .C(new_n572_), .Y(new_n1129_));
  NOR3X1   g0866(.A(new_n267_), .B(new_n266_), .C(new_n477_), .Y(new_n1130_));
  NOR3X1   g0867(.A(\shift[1] ), .B(\shift[0] ), .C(new_n576_), .Y(new_n1131_));
  OR4X1    g0868(.A(new_n1131_), .B(new_n1130_), .C(new_n1129_), .D(new_n1128_), .Y(new_n1132_));
  NOR3X1   g0869(.A(new_n267_), .B(\shift[0] ), .C(new_n473_), .Y(new_n1133_));
  NOR3X1   g0870(.A(\shift[1] ), .B(new_n266_), .C(new_n475_), .Y(new_n1134_));
  NOR3X1   g0871(.A(new_n267_), .B(new_n266_), .C(new_n486_), .Y(new_n1135_));
  NOR3X1   g0872(.A(\shift[1] ), .B(\shift[0] ), .C(new_n479_), .Y(new_n1136_));
  OR4X1    g0873(.A(new_n1136_), .B(new_n1135_), .C(new_n1134_), .D(new_n1133_), .Y(new_n1137_));
  AOI22X1  g0874(.A0(new_n1137_), .A1(new_n287_), .B0(new_n1132_), .B1(new_n276_), .Y(new_n1138_));
  NOR3X1   g0875(.A(new_n267_), .B(\shift[0] ), .C(new_n501_), .Y(new_n1139_));
  NOR3X1   g0876(.A(\shift[1] ), .B(new_n266_), .C(new_n503_), .Y(new_n1140_));
  NOR3X1   g0877(.A(new_n267_), .B(new_n266_), .C(new_n496_), .Y(new_n1141_));
  NOR3X1   g0878(.A(\shift[1] ), .B(\shift[0] ), .C(new_n507_), .Y(new_n1142_));
  OR4X1    g0879(.A(new_n1142_), .B(new_n1141_), .C(new_n1140_), .D(new_n1139_), .Y(new_n1143_));
  NOR3X1   g0880(.A(new_n267_), .B(\shift[0] ), .C(new_n482_), .Y(new_n1144_));
  NOR3X1   g0881(.A(\shift[1] ), .B(new_n266_), .C(new_n484_), .Y(new_n1145_));
  NOR3X1   g0882(.A(new_n267_), .B(new_n266_), .C(new_n505_), .Y(new_n1146_));
  NOR3X1   g0883(.A(\shift[1] ), .B(\shift[0] ), .C(new_n488_), .Y(new_n1147_));
  OR4X1    g0884(.A(new_n1147_), .B(new_n1146_), .C(new_n1145_), .D(new_n1144_), .Y(new_n1148_));
  AOI22X1  g0885(.A0(new_n1148_), .A1(new_n308_), .B0(new_n1143_), .B1(new_n298_), .Y(new_n1149_));
  AOI21X1  g0886(.A0(new_n1149_), .A1(new_n1138_), .B0(new_n351_), .Y(new_n1150_));
  OR4X1    g0887(.A(new_n1150_), .B(new_n1127_), .C(new_n1104_), .D(new_n1081_), .Y(new_n1151_));
  MX2X1    g0888(.A(new_n1151_), .B(new_n1058_), .S0(new_n264_), .Y(\result[3] ));
  AOI22X1  g0889(.A0(new_n339_), .A1(new_n276_), .B0(new_n287_), .B1(new_n275_), .Y(new_n1153_));
  AOI22X1  g0890(.A0(new_n308_), .A1(new_n285_), .B0(new_n307_), .B1(new_n298_), .Y(new_n1154_));
  AOI21X1  g0891(.A0(new_n1154_), .A1(new_n1153_), .B0(new_n310_), .Y(new_n1155_));
  AOI22X1  g0892(.A0(new_n420_), .A1(new_n276_), .B0(new_n320_), .B1(new_n287_), .Y(new_n1156_));
  AOI22X1  g0893(.A0(new_n348_), .A1(new_n298_), .B0(new_n329_), .B1(new_n308_), .Y(new_n1157_));
  AOI21X1  g0894(.A0(new_n1157_), .A1(new_n1156_), .B0(new_n351_), .Y(new_n1158_));
  AOI22X1  g0895(.A0(new_n461_), .A1(new_n276_), .B0(new_n361_), .B1(new_n287_), .Y(new_n1159_));
  AOI22X1  g0896(.A0(new_n389_), .A1(new_n298_), .B0(new_n370_), .B1(new_n308_), .Y(new_n1160_));
  AOI21X1  g0897(.A0(new_n1160_), .A1(new_n1159_), .B0(new_n391_), .Y(new_n1161_));
  AOI22X1  g0898(.A0(new_n401_), .A1(new_n287_), .B0(new_n380_), .B1(new_n276_), .Y(new_n1162_));
  AOI22X1  g0899(.A0(new_n429_), .A1(new_n298_), .B0(new_n410_), .B1(new_n308_), .Y(new_n1163_));
  AOI21X1  g0900(.A0(new_n1163_), .A1(new_n1162_), .B0(new_n431_), .Y(new_n1164_));
  OR4X1    g0901(.A(new_n1164_), .B(new_n1161_), .C(new_n1158_), .D(new_n1155_), .Y(new_n1165_));
  AOI22X1  g0902(.A0(new_n559_), .A1(new_n287_), .B0(new_n539_), .B1(new_n276_), .Y(new_n1166_));
  AOI22X1  g0903(.A0(new_n587_), .A1(new_n298_), .B0(new_n568_), .B1(new_n308_), .Y(new_n1167_));
  AOI21X1  g0904(.A0(new_n1167_), .A1(new_n1166_), .B0(new_n431_), .Y(new_n1168_));
  AOI22X1  g0905(.A0(new_n520_), .A1(new_n287_), .B0(new_n297_), .B1(new_n276_), .Y(new_n1169_));
  AOI22X1  g0906(.A0(new_n548_), .A1(new_n298_), .B0(new_n529_), .B1(new_n308_), .Y(new_n1170_));
  AOI21X1  g0907(.A0(new_n1170_), .A1(new_n1169_), .B0(new_n391_), .Y(new_n1171_));
  AOI22X1  g0908(.A0(new_n578_), .A1(new_n276_), .B0(new_n481_), .B1(new_n287_), .Y(new_n1172_));
  AOI22X1  g0909(.A0(new_n509_), .A1(new_n298_), .B0(new_n490_), .B1(new_n308_), .Y(new_n1173_));
  AOI21X1  g0910(.A0(new_n1173_), .A1(new_n1172_), .B0(new_n351_), .Y(new_n1174_));
  AOI22X1  g0911(.A0(new_n500_), .A1(new_n276_), .B0(new_n442_), .B1(new_n287_), .Y(new_n1175_));
  AOI22X1  g0912(.A0(new_n470_), .A1(new_n298_), .B0(new_n451_), .B1(new_n308_), .Y(new_n1176_));
  AOI21X1  g0913(.A0(new_n1176_), .A1(new_n1175_), .B0(new_n310_), .Y(new_n1177_));
  OR4X1    g0914(.A(new_n1177_), .B(new_n1174_), .C(new_n1171_), .D(new_n1168_), .Y(new_n1178_));
  MX2X1    g0915(.A(new_n1178_), .B(new_n1165_), .S0(new_n264_), .Y(\result[4] ));
  AOI22X1  g0916(.A0(new_n630_), .A1(new_n276_), .B0(new_n596_), .B1(new_n287_), .Y(new_n1180_));
  AOI22X1  g0917(.A0(new_n612_), .A1(new_n298_), .B0(new_n601_), .B1(new_n308_), .Y(new_n1181_));
  AOI21X1  g0918(.A0(new_n1181_), .A1(new_n1180_), .B0(new_n310_), .Y(new_n1182_));
  AOI22X1  g0919(.A0(new_n676_), .A1(new_n276_), .B0(new_n619_), .B1(new_n287_), .Y(new_n1183_));
  AOI22X1  g0920(.A0(new_n635_), .A1(new_n298_), .B0(new_n624_), .B1(new_n308_), .Y(new_n1184_));
  AOI21X1  g0921(.A0(new_n1184_), .A1(new_n1183_), .B0(new_n351_), .Y(new_n1185_));
  AOI22X1  g0922(.A0(new_n723_), .A1(new_n276_), .B0(new_n642_), .B1(new_n287_), .Y(new_n1186_));
  AOI22X1  g0923(.A0(new_n658_), .A1(new_n298_), .B0(new_n647_), .B1(new_n308_), .Y(new_n1187_));
  AOI21X1  g0924(.A0(new_n1187_), .A1(new_n1186_), .B0(new_n391_), .Y(new_n1188_));
  AOI22X1  g0925(.A0(new_n665_), .A1(new_n287_), .B0(new_n653_), .B1(new_n276_), .Y(new_n1189_));
  AOI22X1  g0926(.A0(new_n681_), .A1(new_n298_), .B0(new_n670_), .B1(new_n308_), .Y(new_n1190_));
  AOI21X1  g0927(.A0(new_n1190_), .A1(new_n1189_), .B0(new_n431_), .Y(new_n1191_));
  OR4X1    g0928(.A(new_n1191_), .B(new_n1188_), .C(new_n1185_), .D(new_n1182_), .Y(new_n1192_));
  AOI22X1  g0929(.A0(new_n735_), .A1(new_n287_), .B0(new_n700_), .B1(new_n276_), .Y(new_n1193_));
  AOI22X1  g0930(.A0(new_n751_), .A1(new_n298_), .B0(new_n740_), .B1(new_n308_), .Y(new_n1194_));
  AOI21X1  g0931(.A0(new_n1194_), .A1(new_n1193_), .B0(new_n431_), .Y(new_n1195_));
  AOI22X1  g0932(.A0(new_n689_), .A1(new_n287_), .B0(new_n607_), .B1(new_n276_), .Y(new_n1196_));
  AOI22X1  g0933(.A0(new_n705_), .A1(new_n298_), .B0(new_n694_), .B1(new_n308_), .Y(new_n1197_));
  AOI21X1  g0934(.A0(new_n1197_), .A1(new_n1196_), .B0(new_n391_), .Y(new_n1198_));
  AOI22X1  g0935(.A0(new_n758_), .A1(new_n287_), .B0(new_n746_), .B1(new_n276_), .Y(new_n1199_));
  AOI22X1  g0936(.A0(new_n774_), .A1(new_n298_), .B0(new_n763_), .B1(new_n308_), .Y(new_n1200_));
  AOI21X1  g0937(.A0(new_n1200_), .A1(new_n1199_), .B0(new_n351_), .Y(new_n1201_));
  AOI22X1  g0938(.A0(new_n769_), .A1(new_n276_), .B0(new_n712_), .B1(new_n287_), .Y(new_n1202_));
  AOI22X1  g0939(.A0(new_n728_), .A1(new_n298_), .B0(new_n717_), .B1(new_n308_), .Y(new_n1203_));
  AOI21X1  g0940(.A0(new_n1203_), .A1(new_n1202_), .B0(new_n310_), .Y(new_n1204_));
  OR4X1    g0941(.A(new_n1204_), .B(new_n1201_), .C(new_n1198_), .D(new_n1195_), .Y(new_n1205_));
  MX2X1    g0942(.A(new_n1205_), .B(new_n1192_), .S0(new_n264_), .Y(\result[5] ));
  AOI22X1  g0943(.A0(new_n817_), .A1(new_n276_), .B0(new_n783_), .B1(new_n287_), .Y(new_n1207_));
  AOI22X1  g0944(.A0(new_n799_), .A1(new_n298_), .B0(new_n788_), .B1(new_n308_), .Y(new_n1208_));
  AOI21X1  g0945(.A0(new_n1208_), .A1(new_n1207_), .B0(new_n310_), .Y(new_n1209_));
  AOI22X1  g0946(.A0(new_n863_), .A1(new_n276_), .B0(new_n806_), .B1(new_n287_), .Y(new_n1210_));
  AOI22X1  g0947(.A0(new_n822_), .A1(new_n298_), .B0(new_n811_), .B1(new_n308_), .Y(new_n1211_));
  AOI21X1  g0948(.A0(new_n1211_), .A1(new_n1210_), .B0(new_n351_), .Y(new_n1212_));
  AOI22X1  g0949(.A0(new_n910_), .A1(new_n276_), .B0(new_n829_), .B1(new_n287_), .Y(new_n1213_));
  AOI22X1  g0950(.A0(new_n845_), .A1(new_n298_), .B0(new_n834_), .B1(new_n308_), .Y(new_n1214_));
  AOI21X1  g0951(.A0(new_n1214_), .A1(new_n1213_), .B0(new_n391_), .Y(new_n1215_));
  AOI22X1  g0952(.A0(new_n852_), .A1(new_n287_), .B0(new_n840_), .B1(new_n276_), .Y(new_n1216_));
  AOI22X1  g0953(.A0(new_n868_), .A1(new_n298_), .B0(new_n857_), .B1(new_n308_), .Y(new_n1217_));
  AOI21X1  g0954(.A0(new_n1217_), .A1(new_n1216_), .B0(new_n431_), .Y(new_n1218_));
  OR4X1    g0955(.A(new_n1218_), .B(new_n1215_), .C(new_n1212_), .D(new_n1209_), .Y(new_n1219_));
  AOI22X1  g0956(.A0(new_n922_), .A1(new_n287_), .B0(new_n887_), .B1(new_n276_), .Y(new_n1220_));
  AOI22X1  g0957(.A0(new_n938_), .A1(new_n298_), .B0(new_n927_), .B1(new_n308_), .Y(new_n1221_));
  AOI21X1  g0958(.A0(new_n1221_), .A1(new_n1220_), .B0(new_n431_), .Y(new_n1222_));
  AOI22X1  g0959(.A0(new_n876_), .A1(new_n287_), .B0(new_n794_), .B1(new_n276_), .Y(new_n1223_));
  AOI22X1  g0960(.A0(new_n892_), .A1(new_n298_), .B0(new_n881_), .B1(new_n308_), .Y(new_n1224_));
  AOI21X1  g0961(.A0(new_n1224_), .A1(new_n1223_), .B0(new_n391_), .Y(new_n1225_));
  AOI22X1  g0962(.A0(new_n945_), .A1(new_n287_), .B0(new_n933_), .B1(new_n276_), .Y(new_n1226_));
  AOI22X1  g0963(.A0(new_n961_), .A1(new_n298_), .B0(new_n950_), .B1(new_n308_), .Y(new_n1227_));
  AOI21X1  g0964(.A0(new_n1227_), .A1(new_n1226_), .B0(new_n351_), .Y(new_n1228_));
  AOI22X1  g0965(.A0(new_n956_), .A1(new_n276_), .B0(new_n899_), .B1(new_n287_), .Y(new_n1229_));
  AOI22X1  g0966(.A0(new_n915_), .A1(new_n298_), .B0(new_n904_), .B1(new_n308_), .Y(new_n1230_));
  AOI21X1  g0967(.A0(new_n1230_), .A1(new_n1229_), .B0(new_n310_), .Y(new_n1231_));
  OR4X1    g0968(.A(new_n1231_), .B(new_n1228_), .C(new_n1225_), .D(new_n1222_), .Y(new_n1232_));
  MX2X1    g0969(.A(new_n1232_), .B(new_n1219_), .S0(new_n264_), .Y(\result[6] ));
  AOI22X1  g0970(.A0(new_n1039_), .A1(new_n287_), .B0(new_n1004_), .B1(new_n276_), .Y(new_n1234_));
  AOI22X1  g0971(.A0(new_n1055_), .A1(new_n298_), .B0(new_n1044_), .B1(new_n308_), .Y(new_n1235_));
  AOI21X1  g0972(.A0(new_n1235_), .A1(new_n1234_), .B0(new_n310_), .Y(new_n1236_));
  AOI22X1  g0973(.A0(new_n993_), .A1(new_n287_), .B0(new_n981_), .B1(new_n276_), .Y(new_n1237_));
  AOI22X1  g0974(.A0(new_n1009_), .A1(new_n298_), .B0(new_n998_), .B1(new_n308_), .Y(new_n1238_));
  AOI21X1  g0975(.A0(new_n1238_), .A1(new_n1237_), .B0(new_n351_), .Y(new_n1239_));
  AOI22X1  g0976(.A0(new_n1120_), .A1(new_n276_), .B0(new_n1016_), .B1(new_n287_), .Y(new_n1240_));
  AOI22X1  g0977(.A0(new_n1032_), .A1(new_n298_), .B0(new_n1021_), .B1(new_n308_), .Y(new_n1241_));
  AOI21X1  g0978(.A0(new_n1241_), .A1(new_n1240_), .B0(new_n391_), .Y(new_n1242_));
  AOI22X1  g0979(.A0(new_n1027_), .A1(new_n276_), .B0(new_n970_), .B1(new_n287_), .Y(new_n1243_));
  AOI22X1  g0980(.A0(new_n986_), .A1(new_n298_), .B0(new_n975_), .B1(new_n308_), .Y(new_n1244_));
  AOI21X1  g0981(.A0(new_n1244_), .A1(new_n1243_), .B0(new_n431_), .Y(new_n1245_));
  OR4X1    g0982(.A(new_n1245_), .B(new_n1242_), .C(new_n1239_), .D(new_n1236_), .Y(new_n1246_));
  AOI22X1  g0983(.A0(new_n1091_), .A1(new_n308_), .B0(new_n1086_), .B1(new_n287_), .Y(new_n1247_));
  AOI22X1  g0984(.A0(new_n1102_), .A1(new_n298_), .B0(new_n1074_), .B1(new_n276_), .Y(new_n1248_));
  AOI21X1  g0985(.A0(new_n1248_), .A1(new_n1247_), .B0(new_n431_), .Y(new_n1249_));
  AOI22X1  g0986(.A0(new_n1063_), .A1(new_n287_), .B0(new_n1050_), .B1(new_n276_), .Y(new_n1250_));
  AOI22X1  g0987(.A0(new_n1079_), .A1(new_n298_), .B0(new_n1068_), .B1(new_n308_), .Y(new_n1251_));
  AOI21X1  g0988(.A0(new_n1251_), .A1(new_n1250_), .B0(new_n391_), .Y(new_n1252_));
  AOI22X1  g0989(.A0(new_n1132_), .A1(new_n287_), .B0(new_n1097_), .B1(new_n276_), .Y(new_n1253_));
  AOI22X1  g0990(.A0(new_n1148_), .A1(new_n298_), .B0(new_n1137_), .B1(new_n308_), .Y(new_n1254_));
  AOI21X1  g0991(.A0(new_n1254_), .A1(new_n1253_), .B0(new_n351_), .Y(new_n1255_));
  AOI22X1  g0992(.A0(new_n1143_), .A1(new_n276_), .B0(new_n1109_), .B1(new_n287_), .Y(new_n1256_));
  AOI22X1  g0993(.A0(new_n1125_), .A1(new_n298_), .B0(new_n1114_), .B1(new_n308_), .Y(new_n1257_));
  AOI21X1  g0994(.A0(new_n1257_), .A1(new_n1256_), .B0(new_n310_), .Y(new_n1258_));
  OR4X1    g0995(.A(new_n1258_), .B(new_n1255_), .C(new_n1252_), .D(new_n1249_), .Y(new_n1259_));
  MX2X1    g0996(.A(new_n1259_), .B(new_n1246_), .S0(new_n264_), .Y(\result[7] ));
  AOI22X1  g0997(.A0(new_n348_), .A1(new_n276_), .B0(new_n339_), .B1(new_n287_), .Y(new_n1261_));
  AOI22X1  g0998(.A0(new_n308_), .A1(new_n275_), .B0(new_n298_), .B1(new_n285_), .Y(new_n1262_));
  AOI21X1  g0999(.A0(new_n1262_), .A1(new_n1261_), .B0(new_n310_), .Y(new_n1263_));
  AOI22X1  g1000(.A0(new_n429_), .A1(new_n276_), .B0(new_n420_), .B1(new_n287_), .Y(new_n1264_));
  AOI22X1  g1001(.A0(new_n329_), .A1(new_n298_), .B0(new_n320_), .B1(new_n308_), .Y(new_n1265_));
  AOI21X1  g1002(.A0(new_n1265_), .A1(new_n1264_), .B0(new_n351_), .Y(new_n1266_));
  AOI22X1  g1003(.A0(new_n470_), .A1(new_n276_), .B0(new_n461_), .B1(new_n287_), .Y(new_n1267_));
  AOI22X1  g1004(.A0(new_n370_), .A1(new_n298_), .B0(new_n361_), .B1(new_n308_), .Y(new_n1268_));
  AOI21X1  g1005(.A0(new_n1268_), .A1(new_n1267_), .B0(new_n391_), .Y(new_n1269_));
  AOI22X1  g1006(.A0(new_n389_), .A1(new_n276_), .B0(new_n380_), .B1(new_n287_), .Y(new_n1270_));
  AOI22X1  g1007(.A0(new_n410_), .A1(new_n298_), .B0(new_n401_), .B1(new_n308_), .Y(new_n1271_));
  AOI21X1  g1008(.A0(new_n1271_), .A1(new_n1270_), .B0(new_n431_), .Y(new_n1272_));
  OR4X1    g1009(.A(new_n1272_), .B(new_n1269_), .C(new_n1266_), .D(new_n1263_), .Y(new_n1273_));
  AOI22X1  g1010(.A0(new_n548_), .A1(new_n276_), .B0(new_n539_), .B1(new_n287_), .Y(new_n1274_));
  AOI22X1  g1011(.A0(new_n568_), .A1(new_n298_), .B0(new_n559_), .B1(new_n308_), .Y(new_n1275_));
  AOI21X1  g1012(.A0(new_n1275_), .A1(new_n1274_), .B0(new_n431_), .Y(new_n1276_));
  AOI22X1  g1013(.A0(new_n307_), .A1(new_n276_), .B0(new_n297_), .B1(new_n287_), .Y(new_n1277_));
  AOI22X1  g1014(.A0(new_n529_), .A1(new_n298_), .B0(new_n520_), .B1(new_n308_), .Y(new_n1278_));
  AOI21X1  g1015(.A0(new_n1278_), .A1(new_n1277_), .B0(new_n391_), .Y(new_n1279_));
  AOI22X1  g1016(.A0(new_n587_), .A1(new_n276_), .B0(new_n578_), .B1(new_n287_), .Y(new_n1280_));
  AOI22X1  g1017(.A0(new_n490_), .A1(new_n298_), .B0(new_n481_), .B1(new_n308_), .Y(new_n1281_));
  AOI21X1  g1018(.A0(new_n1281_), .A1(new_n1280_), .B0(new_n351_), .Y(new_n1282_));
  AOI22X1  g1019(.A0(new_n509_), .A1(new_n276_), .B0(new_n500_), .B1(new_n287_), .Y(new_n1283_));
  AOI22X1  g1020(.A0(new_n451_), .A1(new_n298_), .B0(new_n442_), .B1(new_n308_), .Y(new_n1284_));
  AOI21X1  g1021(.A0(new_n1284_), .A1(new_n1283_), .B0(new_n310_), .Y(new_n1285_));
  OR4X1    g1022(.A(new_n1285_), .B(new_n1282_), .C(new_n1279_), .D(new_n1276_), .Y(new_n1286_));
  MX2X1    g1023(.A(new_n1286_), .B(new_n1273_), .S0(new_n264_), .Y(\result[8] ));
  AOI22X1  g1024(.A0(new_n635_), .A1(new_n276_), .B0(new_n630_), .B1(new_n287_), .Y(new_n1288_));
  AOI22X1  g1025(.A0(new_n601_), .A1(new_n298_), .B0(new_n596_), .B1(new_n308_), .Y(new_n1289_));
  AOI21X1  g1026(.A0(new_n1289_), .A1(new_n1288_), .B0(new_n310_), .Y(new_n1290_));
  AOI22X1  g1027(.A0(new_n681_), .A1(new_n276_), .B0(new_n676_), .B1(new_n287_), .Y(new_n1291_));
  AOI22X1  g1028(.A0(new_n624_), .A1(new_n298_), .B0(new_n619_), .B1(new_n308_), .Y(new_n1292_));
  AOI21X1  g1029(.A0(new_n1292_), .A1(new_n1291_), .B0(new_n351_), .Y(new_n1293_));
  AOI22X1  g1030(.A0(new_n728_), .A1(new_n276_), .B0(new_n723_), .B1(new_n287_), .Y(new_n1294_));
  AOI22X1  g1031(.A0(new_n647_), .A1(new_n298_), .B0(new_n642_), .B1(new_n308_), .Y(new_n1295_));
  AOI21X1  g1032(.A0(new_n1295_), .A1(new_n1294_), .B0(new_n391_), .Y(new_n1296_));
  AOI22X1  g1033(.A0(new_n658_), .A1(new_n276_), .B0(new_n653_), .B1(new_n287_), .Y(new_n1297_));
  AOI22X1  g1034(.A0(new_n670_), .A1(new_n298_), .B0(new_n665_), .B1(new_n308_), .Y(new_n1298_));
  AOI21X1  g1035(.A0(new_n1298_), .A1(new_n1297_), .B0(new_n431_), .Y(new_n1299_));
  OR4X1    g1036(.A(new_n1299_), .B(new_n1296_), .C(new_n1293_), .D(new_n1290_), .Y(new_n1300_));
  AOI22X1  g1037(.A0(new_n705_), .A1(new_n276_), .B0(new_n700_), .B1(new_n287_), .Y(new_n1301_));
  AOI22X1  g1038(.A0(new_n740_), .A1(new_n298_), .B0(new_n735_), .B1(new_n308_), .Y(new_n1302_));
  AOI21X1  g1039(.A0(new_n1302_), .A1(new_n1301_), .B0(new_n431_), .Y(new_n1303_));
  AOI22X1  g1040(.A0(new_n612_), .A1(new_n276_), .B0(new_n607_), .B1(new_n287_), .Y(new_n1304_));
  AOI22X1  g1041(.A0(new_n694_), .A1(new_n298_), .B0(new_n689_), .B1(new_n308_), .Y(new_n1305_));
  AOI21X1  g1042(.A0(new_n1305_), .A1(new_n1304_), .B0(new_n391_), .Y(new_n1306_));
  AOI22X1  g1043(.A0(new_n751_), .A1(new_n276_), .B0(new_n746_), .B1(new_n287_), .Y(new_n1307_));
  AOI22X1  g1044(.A0(new_n763_), .A1(new_n298_), .B0(new_n758_), .B1(new_n308_), .Y(new_n1308_));
  AOI21X1  g1045(.A0(new_n1308_), .A1(new_n1307_), .B0(new_n351_), .Y(new_n1309_));
  AOI22X1  g1046(.A0(new_n774_), .A1(new_n276_), .B0(new_n769_), .B1(new_n287_), .Y(new_n1310_));
  AOI22X1  g1047(.A0(new_n717_), .A1(new_n298_), .B0(new_n712_), .B1(new_n308_), .Y(new_n1311_));
  AOI21X1  g1048(.A0(new_n1311_), .A1(new_n1310_), .B0(new_n310_), .Y(new_n1312_));
  OR4X1    g1049(.A(new_n1312_), .B(new_n1309_), .C(new_n1306_), .D(new_n1303_), .Y(new_n1313_));
  MX2X1    g1050(.A(new_n1313_), .B(new_n1300_), .S0(new_n264_), .Y(\result[9] ));
  AOI22X1  g1051(.A0(new_n822_), .A1(new_n276_), .B0(new_n817_), .B1(new_n287_), .Y(new_n1315_));
  AOI22X1  g1052(.A0(new_n788_), .A1(new_n298_), .B0(new_n783_), .B1(new_n308_), .Y(new_n1316_));
  AOI21X1  g1053(.A0(new_n1316_), .A1(new_n1315_), .B0(new_n310_), .Y(new_n1317_));
  AOI22X1  g1054(.A0(new_n868_), .A1(new_n276_), .B0(new_n863_), .B1(new_n287_), .Y(new_n1318_));
  AOI22X1  g1055(.A0(new_n811_), .A1(new_n298_), .B0(new_n806_), .B1(new_n308_), .Y(new_n1319_));
  AOI21X1  g1056(.A0(new_n1319_), .A1(new_n1318_), .B0(new_n351_), .Y(new_n1320_));
  AOI22X1  g1057(.A0(new_n915_), .A1(new_n276_), .B0(new_n910_), .B1(new_n287_), .Y(new_n1321_));
  AOI22X1  g1058(.A0(new_n834_), .A1(new_n298_), .B0(new_n829_), .B1(new_n308_), .Y(new_n1322_));
  AOI21X1  g1059(.A0(new_n1322_), .A1(new_n1321_), .B0(new_n391_), .Y(new_n1323_));
  AOI22X1  g1060(.A0(new_n845_), .A1(new_n276_), .B0(new_n840_), .B1(new_n287_), .Y(new_n1324_));
  AOI22X1  g1061(.A0(new_n857_), .A1(new_n298_), .B0(new_n852_), .B1(new_n308_), .Y(new_n1325_));
  AOI21X1  g1062(.A0(new_n1325_), .A1(new_n1324_), .B0(new_n431_), .Y(new_n1326_));
  OR4X1    g1063(.A(new_n1326_), .B(new_n1323_), .C(new_n1320_), .D(new_n1317_), .Y(new_n1327_));
  AOI22X1  g1064(.A0(new_n892_), .A1(new_n276_), .B0(new_n887_), .B1(new_n287_), .Y(new_n1328_));
  AOI22X1  g1065(.A0(new_n927_), .A1(new_n298_), .B0(new_n922_), .B1(new_n308_), .Y(new_n1329_));
  AOI21X1  g1066(.A0(new_n1329_), .A1(new_n1328_), .B0(new_n431_), .Y(new_n1330_));
  AOI22X1  g1067(.A0(new_n799_), .A1(new_n276_), .B0(new_n794_), .B1(new_n287_), .Y(new_n1331_));
  AOI22X1  g1068(.A0(new_n881_), .A1(new_n298_), .B0(new_n876_), .B1(new_n308_), .Y(new_n1332_));
  AOI21X1  g1069(.A0(new_n1332_), .A1(new_n1331_), .B0(new_n391_), .Y(new_n1333_));
  AOI22X1  g1070(.A0(new_n938_), .A1(new_n276_), .B0(new_n933_), .B1(new_n287_), .Y(new_n1334_));
  AOI22X1  g1071(.A0(new_n950_), .A1(new_n298_), .B0(new_n945_), .B1(new_n308_), .Y(new_n1335_));
  AOI21X1  g1072(.A0(new_n1335_), .A1(new_n1334_), .B0(new_n351_), .Y(new_n1336_));
  AOI22X1  g1073(.A0(new_n961_), .A1(new_n276_), .B0(new_n956_), .B1(new_n287_), .Y(new_n1337_));
  AOI22X1  g1074(.A0(new_n904_), .A1(new_n298_), .B0(new_n899_), .B1(new_n308_), .Y(new_n1338_));
  AOI21X1  g1075(.A0(new_n1338_), .A1(new_n1337_), .B0(new_n310_), .Y(new_n1339_));
  OR4X1    g1076(.A(new_n1339_), .B(new_n1336_), .C(new_n1333_), .D(new_n1330_), .Y(new_n1340_));
  MX2X1    g1077(.A(new_n1340_), .B(new_n1327_), .S0(new_n264_), .Y(\result[10] ));
  AOI22X1  g1078(.A0(new_n1009_), .A1(new_n276_), .B0(new_n1004_), .B1(new_n287_), .Y(new_n1342_));
  AOI22X1  g1079(.A0(new_n1044_), .A1(new_n298_), .B0(new_n1039_), .B1(new_n308_), .Y(new_n1343_));
  AOI21X1  g1080(.A0(new_n1343_), .A1(new_n1342_), .B0(new_n310_), .Y(new_n1344_));
  AOI22X1  g1081(.A0(new_n986_), .A1(new_n276_), .B0(new_n981_), .B1(new_n287_), .Y(new_n1345_));
  AOI22X1  g1082(.A0(new_n998_), .A1(new_n298_), .B0(new_n993_), .B1(new_n308_), .Y(new_n1346_));
  AOI21X1  g1083(.A0(new_n1346_), .A1(new_n1345_), .B0(new_n351_), .Y(new_n1347_));
  AOI22X1  g1084(.A0(new_n1125_), .A1(new_n276_), .B0(new_n1120_), .B1(new_n287_), .Y(new_n1348_));
  AOI22X1  g1085(.A0(new_n1021_), .A1(new_n298_), .B0(new_n1016_), .B1(new_n308_), .Y(new_n1349_));
  AOI21X1  g1086(.A0(new_n1349_), .A1(new_n1348_), .B0(new_n391_), .Y(new_n1350_));
  AOI22X1  g1087(.A0(new_n1032_), .A1(new_n276_), .B0(new_n1027_), .B1(new_n287_), .Y(new_n1351_));
  AOI22X1  g1088(.A0(new_n975_), .A1(new_n298_), .B0(new_n970_), .B1(new_n308_), .Y(new_n1352_));
  AOI21X1  g1089(.A0(new_n1352_), .A1(new_n1351_), .B0(new_n431_), .Y(new_n1353_));
  OR4X1    g1090(.A(new_n1353_), .B(new_n1350_), .C(new_n1347_), .D(new_n1344_), .Y(new_n1354_));
  AOI22X1  g1091(.A0(new_n1086_), .A1(new_n308_), .B0(new_n1079_), .B1(new_n276_), .Y(new_n1355_));
  AOI22X1  g1092(.A0(new_n1091_), .A1(new_n298_), .B0(new_n1074_), .B1(new_n287_), .Y(new_n1356_));
  AOI21X1  g1093(.A0(new_n1356_), .A1(new_n1355_), .B0(new_n431_), .Y(new_n1357_));
  AOI22X1  g1094(.A0(new_n1055_), .A1(new_n276_), .B0(new_n1050_), .B1(new_n287_), .Y(new_n1358_));
  AOI22X1  g1095(.A0(new_n1068_), .A1(new_n298_), .B0(new_n1063_), .B1(new_n308_), .Y(new_n1359_));
  AOI21X1  g1096(.A0(new_n1359_), .A1(new_n1358_), .B0(new_n391_), .Y(new_n1360_));
  AOI22X1  g1097(.A0(new_n1102_), .A1(new_n276_), .B0(new_n1097_), .B1(new_n287_), .Y(new_n1361_));
  AOI22X1  g1098(.A0(new_n1137_), .A1(new_n298_), .B0(new_n1132_), .B1(new_n308_), .Y(new_n1362_));
  AOI21X1  g1099(.A0(new_n1362_), .A1(new_n1361_), .B0(new_n351_), .Y(new_n1363_));
  AOI22X1  g1100(.A0(new_n1148_), .A1(new_n276_), .B0(new_n1143_), .B1(new_n287_), .Y(new_n1364_));
  AOI22X1  g1101(.A0(new_n1114_), .A1(new_n298_), .B0(new_n1109_), .B1(new_n308_), .Y(new_n1365_));
  AOI21X1  g1102(.A0(new_n1365_), .A1(new_n1364_), .B0(new_n310_), .Y(new_n1366_));
  OR4X1    g1103(.A(new_n1366_), .B(new_n1363_), .C(new_n1360_), .D(new_n1357_), .Y(new_n1367_));
  MX2X1    g1104(.A(new_n1367_), .B(new_n1354_), .S0(new_n264_), .Y(\result[11] ));
  AOI22X1  g1105(.A0(new_n348_), .A1(new_n287_), .B0(new_n329_), .B1(new_n276_), .Y(new_n1369_));
  AOI22X1  g1106(.A0(new_n339_), .A1(new_n308_), .B0(new_n298_), .B1(new_n275_), .Y(new_n1370_));
  AOI21X1  g1107(.A0(new_n1370_), .A1(new_n1369_), .B0(new_n310_), .Y(new_n1371_));
  AOI22X1  g1108(.A0(new_n429_), .A1(new_n287_), .B0(new_n410_), .B1(new_n276_), .Y(new_n1372_));
  AOI22X1  g1109(.A0(new_n420_), .A1(new_n308_), .B0(new_n320_), .B1(new_n298_), .Y(new_n1373_));
  AOI21X1  g1110(.A0(new_n1373_), .A1(new_n1372_), .B0(new_n351_), .Y(new_n1374_));
  AOI22X1  g1111(.A0(new_n470_), .A1(new_n287_), .B0(new_n451_), .B1(new_n276_), .Y(new_n1375_));
  AOI22X1  g1112(.A0(new_n461_), .A1(new_n308_), .B0(new_n361_), .B1(new_n298_), .Y(new_n1376_));
  AOI21X1  g1113(.A0(new_n1376_), .A1(new_n1375_), .B0(new_n391_), .Y(new_n1377_));
  AOI22X1  g1114(.A0(new_n389_), .A1(new_n287_), .B0(new_n370_), .B1(new_n276_), .Y(new_n1378_));
  AOI22X1  g1115(.A0(new_n401_), .A1(new_n298_), .B0(new_n380_), .B1(new_n308_), .Y(new_n1379_));
  AOI21X1  g1116(.A0(new_n1379_), .A1(new_n1378_), .B0(new_n431_), .Y(new_n1380_));
  OR4X1    g1117(.A(new_n1380_), .B(new_n1377_), .C(new_n1374_), .D(new_n1371_), .Y(new_n1381_));
  AOI22X1  g1118(.A0(new_n548_), .A1(new_n287_), .B0(new_n529_), .B1(new_n276_), .Y(new_n1382_));
  AOI22X1  g1119(.A0(new_n559_), .A1(new_n298_), .B0(new_n539_), .B1(new_n308_), .Y(new_n1383_));
  AOI21X1  g1120(.A0(new_n1383_), .A1(new_n1382_), .B0(new_n431_), .Y(new_n1384_));
  AOI22X1  g1121(.A0(new_n307_), .A1(new_n287_), .B0(new_n285_), .B1(new_n276_), .Y(new_n1385_));
  AOI22X1  g1122(.A0(new_n520_), .A1(new_n298_), .B0(new_n308_), .B1(new_n297_), .Y(new_n1386_));
  AOI21X1  g1123(.A0(new_n1386_), .A1(new_n1385_), .B0(new_n391_), .Y(new_n1387_));
  AOI22X1  g1124(.A0(new_n587_), .A1(new_n287_), .B0(new_n568_), .B1(new_n276_), .Y(new_n1388_));
  AOI22X1  g1125(.A0(new_n578_), .A1(new_n308_), .B0(new_n481_), .B1(new_n298_), .Y(new_n1389_));
  AOI21X1  g1126(.A0(new_n1389_), .A1(new_n1388_), .B0(new_n351_), .Y(new_n1390_));
  AOI22X1  g1127(.A0(new_n509_), .A1(new_n287_), .B0(new_n490_), .B1(new_n276_), .Y(new_n1391_));
  AOI22X1  g1128(.A0(new_n500_), .A1(new_n308_), .B0(new_n442_), .B1(new_n298_), .Y(new_n1392_));
  AOI21X1  g1129(.A0(new_n1392_), .A1(new_n1391_), .B0(new_n310_), .Y(new_n1393_));
  OR4X1    g1130(.A(new_n1393_), .B(new_n1390_), .C(new_n1387_), .D(new_n1384_), .Y(new_n1394_));
  MX2X1    g1131(.A(new_n1394_), .B(new_n1381_), .S0(new_n264_), .Y(\result[12] ));
  AOI22X1  g1132(.A0(new_n635_), .A1(new_n287_), .B0(new_n624_), .B1(new_n276_), .Y(new_n1396_));
  AOI22X1  g1133(.A0(new_n630_), .A1(new_n308_), .B0(new_n596_), .B1(new_n298_), .Y(new_n1397_));
  AOI21X1  g1134(.A0(new_n1397_), .A1(new_n1396_), .B0(new_n310_), .Y(new_n1398_));
  AOI22X1  g1135(.A0(new_n681_), .A1(new_n287_), .B0(new_n670_), .B1(new_n276_), .Y(new_n1399_));
  AOI22X1  g1136(.A0(new_n676_), .A1(new_n308_), .B0(new_n619_), .B1(new_n298_), .Y(new_n1400_));
  AOI21X1  g1137(.A0(new_n1400_), .A1(new_n1399_), .B0(new_n351_), .Y(new_n1401_));
  AOI22X1  g1138(.A0(new_n728_), .A1(new_n287_), .B0(new_n717_), .B1(new_n276_), .Y(new_n1402_));
  AOI22X1  g1139(.A0(new_n723_), .A1(new_n308_), .B0(new_n642_), .B1(new_n298_), .Y(new_n1403_));
  AOI21X1  g1140(.A0(new_n1403_), .A1(new_n1402_), .B0(new_n391_), .Y(new_n1404_));
  AOI22X1  g1141(.A0(new_n658_), .A1(new_n287_), .B0(new_n647_), .B1(new_n276_), .Y(new_n1405_));
  AOI22X1  g1142(.A0(new_n665_), .A1(new_n298_), .B0(new_n653_), .B1(new_n308_), .Y(new_n1406_));
  AOI21X1  g1143(.A0(new_n1406_), .A1(new_n1405_), .B0(new_n431_), .Y(new_n1407_));
  OR4X1    g1144(.A(new_n1407_), .B(new_n1404_), .C(new_n1401_), .D(new_n1398_), .Y(new_n1408_));
  AOI22X1  g1145(.A0(new_n705_), .A1(new_n287_), .B0(new_n694_), .B1(new_n276_), .Y(new_n1409_));
  AOI22X1  g1146(.A0(new_n735_), .A1(new_n298_), .B0(new_n700_), .B1(new_n308_), .Y(new_n1410_));
  AOI21X1  g1147(.A0(new_n1410_), .A1(new_n1409_), .B0(new_n431_), .Y(new_n1411_));
  AOI22X1  g1148(.A0(new_n612_), .A1(new_n287_), .B0(new_n601_), .B1(new_n276_), .Y(new_n1412_));
  AOI22X1  g1149(.A0(new_n689_), .A1(new_n298_), .B0(new_n607_), .B1(new_n308_), .Y(new_n1413_));
  AOI21X1  g1150(.A0(new_n1413_), .A1(new_n1412_), .B0(new_n391_), .Y(new_n1414_));
  AOI22X1  g1151(.A0(new_n751_), .A1(new_n287_), .B0(new_n740_), .B1(new_n276_), .Y(new_n1415_));
  AOI22X1  g1152(.A0(new_n758_), .A1(new_n298_), .B0(new_n746_), .B1(new_n308_), .Y(new_n1416_));
  AOI21X1  g1153(.A0(new_n1416_), .A1(new_n1415_), .B0(new_n351_), .Y(new_n1417_));
  AOI22X1  g1154(.A0(new_n774_), .A1(new_n287_), .B0(new_n763_), .B1(new_n276_), .Y(new_n1418_));
  AOI22X1  g1155(.A0(new_n769_), .A1(new_n308_), .B0(new_n712_), .B1(new_n298_), .Y(new_n1419_));
  AOI21X1  g1156(.A0(new_n1419_), .A1(new_n1418_), .B0(new_n310_), .Y(new_n1420_));
  OR4X1    g1157(.A(new_n1420_), .B(new_n1417_), .C(new_n1414_), .D(new_n1411_), .Y(new_n1421_));
  MX2X1    g1158(.A(new_n1421_), .B(new_n1408_), .S0(new_n264_), .Y(\result[13] ));
  AOI22X1  g1159(.A0(new_n822_), .A1(new_n287_), .B0(new_n811_), .B1(new_n276_), .Y(new_n1423_));
  AOI22X1  g1160(.A0(new_n817_), .A1(new_n308_), .B0(new_n783_), .B1(new_n298_), .Y(new_n1424_));
  AOI21X1  g1161(.A0(new_n1424_), .A1(new_n1423_), .B0(new_n310_), .Y(new_n1425_));
  AOI22X1  g1162(.A0(new_n868_), .A1(new_n287_), .B0(new_n857_), .B1(new_n276_), .Y(new_n1426_));
  AOI22X1  g1163(.A0(new_n863_), .A1(new_n308_), .B0(new_n806_), .B1(new_n298_), .Y(new_n1427_));
  AOI21X1  g1164(.A0(new_n1427_), .A1(new_n1426_), .B0(new_n351_), .Y(new_n1428_));
  AOI22X1  g1165(.A0(new_n915_), .A1(new_n287_), .B0(new_n904_), .B1(new_n276_), .Y(new_n1429_));
  AOI22X1  g1166(.A0(new_n910_), .A1(new_n308_), .B0(new_n829_), .B1(new_n298_), .Y(new_n1430_));
  AOI21X1  g1167(.A0(new_n1430_), .A1(new_n1429_), .B0(new_n391_), .Y(new_n1431_));
  AOI22X1  g1168(.A0(new_n845_), .A1(new_n287_), .B0(new_n834_), .B1(new_n276_), .Y(new_n1432_));
  AOI22X1  g1169(.A0(new_n852_), .A1(new_n298_), .B0(new_n840_), .B1(new_n308_), .Y(new_n1433_));
  AOI21X1  g1170(.A0(new_n1433_), .A1(new_n1432_), .B0(new_n431_), .Y(new_n1434_));
  OR4X1    g1171(.A(new_n1434_), .B(new_n1431_), .C(new_n1428_), .D(new_n1425_), .Y(new_n1435_));
  AOI22X1  g1172(.A0(new_n892_), .A1(new_n287_), .B0(new_n881_), .B1(new_n276_), .Y(new_n1436_));
  AOI22X1  g1173(.A0(new_n922_), .A1(new_n298_), .B0(new_n887_), .B1(new_n308_), .Y(new_n1437_));
  AOI21X1  g1174(.A0(new_n1437_), .A1(new_n1436_), .B0(new_n431_), .Y(new_n1438_));
  AOI22X1  g1175(.A0(new_n799_), .A1(new_n287_), .B0(new_n788_), .B1(new_n276_), .Y(new_n1439_));
  AOI22X1  g1176(.A0(new_n876_), .A1(new_n298_), .B0(new_n794_), .B1(new_n308_), .Y(new_n1440_));
  AOI21X1  g1177(.A0(new_n1440_), .A1(new_n1439_), .B0(new_n391_), .Y(new_n1441_));
  AOI22X1  g1178(.A0(new_n938_), .A1(new_n287_), .B0(new_n927_), .B1(new_n276_), .Y(new_n1442_));
  AOI22X1  g1179(.A0(new_n945_), .A1(new_n298_), .B0(new_n933_), .B1(new_n308_), .Y(new_n1443_));
  AOI21X1  g1180(.A0(new_n1443_), .A1(new_n1442_), .B0(new_n351_), .Y(new_n1444_));
  AOI22X1  g1181(.A0(new_n961_), .A1(new_n287_), .B0(new_n950_), .B1(new_n276_), .Y(new_n1445_));
  AOI22X1  g1182(.A0(new_n956_), .A1(new_n308_), .B0(new_n899_), .B1(new_n298_), .Y(new_n1446_));
  AOI21X1  g1183(.A0(new_n1446_), .A1(new_n1445_), .B0(new_n310_), .Y(new_n1447_));
  OR4X1    g1184(.A(new_n1447_), .B(new_n1444_), .C(new_n1441_), .D(new_n1438_), .Y(new_n1448_));
  MX2X1    g1185(.A(new_n1448_), .B(new_n1435_), .S0(new_n264_), .Y(\result[14] ));
  AOI22X1  g1186(.A0(new_n1009_), .A1(new_n287_), .B0(new_n998_), .B1(new_n276_), .Y(new_n1450_));
  AOI22X1  g1187(.A0(new_n1039_), .A1(new_n298_), .B0(new_n1004_), .B1(new_n308_), .Y(new_n1451_));
  AOI21X1  g1188(.A0(new_n1451_), .A1(new_n1450_), .B0(new_n310_), .Y(new_n1452_));
  AOI22X1  g1189(.A0(new_n986_), .A1(new_n287_), .B0(new_n975_), .B1(new_n276_), .Y(new_n1453_));
  AOI22X1  g1190(.A0(new_n993_), .A1(new_n298_), .B0(new_n981_), .B1(new_n308_), .Y(new_n1454_));
  AOI21X1  g1191(.A0(new_n1454_), .A1(new_n1453_), .B0(new_n351_), .Y(new_n1455_));
  AOI22X1  g1192(.A0(new_n1125_), .A1(new_n287_), .B0(new_n1114_), .B1(new_n276_), .Y(new_n1456_));
  AOI22X1  g1193(.A0(new_n1120_), .A1(new_n308_), .B0(new_n1016_), .B1(new_n298_), .Y(new_n1457_));
  AOI21X1  g1194(.A0(new_n1457_), .A1(new_n1456_), .B0(new_n391_), .Y(new_n1458_));
  AOI22X1  g1195(.A0(new_n1032_), .A1(new_n287_), .B0(new_n1021_), .B1(new_n276_), .Y(new_n1459_));
  AOI22X1  g1196(.A0(new_n1027_), .A1(new_n308_), .B0(new_n970_), .B1(new_n298_), .Y(new_n1460_));
  AOI21X1  g1197(.A0(new_n1460_), .A1(new_n1459_), .B0(new_n431_), .Y(new_n1461_));
  OR4X1    g1198(.A(new_n1461_), .B(new_n1458_), .C(new_n1455_), .D(new_n1452_), .Y(new_n1462_));
  AOI22X1  g1199(.A0(new_n1079_), .A1(new_n287_), .B0(new_n1068_), .B1(new_n276_), .Y(new_n1463_));
  AOI22X1  g1200(.A0(new_n1086_), .A1(new_n298_), .B0(new_n1074_), .B1(new_n308_), .Y(new_n1464_));
  AOI21X1  g1201(.A0(new_n1464_), .A1(new_n1463_), .B0(new_n431_), .Y(new_n1465_));
  AOI22X1  g1202(.A0(new_n1055_), .A1(new_n287_), .B0(new_n1044_), .B1(new_n276_), .Y(new_n1466_));
  AOI22X1  g1203(.A0(new_n1063_), .A1(new_n298_), .B0(new_n1050_), .B1(new_n308_), .Y(new_n1467_));
  AOI21X1  g1204(.A0(new_n1467_), .A1(new_n1466_), .B0(new_n391_), .Y(new_n1468_));
  AOI22X1  g1205(.A0(new_n1102_), .A1(new_n287_), .B0(new_n1091_), .B1(new_n276_), .Y(new_n1469_));
  AOI22X1  g1206(.A0(new_n1132_), .A1(new_n298_), .B0(new_n1097_), .B1(new_n308_), .Y(new_n1470_));
  AOI21X1  g1207(.A0(new_n1470_), .A1(new_n1469_), .B0(new_n351_), .Y(new_n1471_));
  AOI22X1  g1208(.A0(new_n1148_), .A1(new_n287_), .B0(new_n1137_), .B1(new_n276_), .Y(new_n1472_));
  AOI22X1  g1209(.A0(new_n1143_), .A1(new_n308_), .B0(new_n1109_), .B1(new_n298_), .Y(new_n1473_));
  AOI21X1  g1210(.A0(new_n1473_), .A1(new_n1472_), .B0(new_n310_), .Y(new_n1474_));
  OR4X1    g1211(.A(new_n1474_), .B(new_n1471_), .C(new_n1468_), .D(new_n1465_), .Y(new_n1475_));
  MX2X1    g1212(.A(new_n1475_), .B(new_n1462_), .S0(new_n264_), .Y(\result[15] ));
  AOI21X1  g1213(.A0(new_n349_), .A1(new_n330_), .B0(new_n310_), .Y(new_n1477_));
  AOI21X1  g1214(.A0(new_n430_), .A1(new_n411_), .B0(new_n351_), .Y(new_n1478_));
  AOI21X1  g1215(.A0(new_n471_), .A1(new_n452_), .B0(new_n391_), .Y(new_n1479_));
  AOI21X1  g1216(.A0(new_n390_), .A1(new_n371_), .B0(new_n431_), .Y(new_n1480_));
  OR4X1    g1217(.A(new_n1480_), .B(new_n1479_), .C(new_n1478_), .D(new_n1477_), .Y(new_n1481_));
  AOI21X1  g1218(.A0(new_n309_), .A1(new_n288_), .B0(new_n391_), .Y(new_n1482_));
  AOI21X1  g1219(.A0(new_n510_), .A1(new_n491_), .B0(new_n310_), .Y(new_n1483_));
  AOI21X1  g1220(.A0(new_n549_), .A1(new_n530_), .B0(new_n431_), .Y(new_n1484_));
  AOI21X1  g1221(.A0(new_n588_), .A1(new_n569_), .B0(new_n351_), .Y(new_n1485_));
  OR4X1    g1222(.A(new_n1485_), .B(new_n1484_), .C(new_n1483_), .D(new_n1482_), .Y(new_n1486_));
  MX2X1    g1223(.A(new_n1486_), .B(new_n1481_), .S0(new_n264_), .Y(\result[16] ));
  AOI21X1  g1224(.A0(new_n636_), .A1(new_n625_), .B0(new_n310_), .Y(new_n1488_));
  AOI21X1  g1225(.A0(new_n682_), .A1(new_n671_), .B0(new_n351_), .Y(new_n1489_));
  AOI21X1  g1226(.A0(new_n729_), .A1(new_n718_), .B0(new_n391_), .Y(new_n1490_));
  AOI21X1  g1227(.A0(new_n659_), .A1(new_n648_), .B0(new_n431_), .Y(new_n1491_));
  OR4X1    g1228(.A(new_n1491_), .B(new_n1490_), .C(new_n1489_), .D(new_n1488_), .Y(new_n1492_));
  AOI21X1  g1229(.A0(new_n706_), .A1(new_n695_), .B0(new_n431_), .Y(new_n1493_));
  AOI21X1  g1230(.A0(new_n613_), .A1(new_n602_), .B0(new_n391_), .Y(new_n1494_));
  AOI21X1  g1231(.A0(new_n752_), .A1(new_n741_), .B0(new_n351_), .Y(new_n1495_));
  AOI21X1  g1232(.A0(new_n775_), .A1(new_n764_), .B0(new_n310_), .Y(new_n1496_));
  OR4X1    g1233(.A(new_n1496_), .B(new_n1495_), .C(new_n1494_), .D(new_n1493_), .Y(new_n1497_));
  MX2X1    g1234(.A(new_n1497_), .B(new_n1492_), .S0(new_n264_), .Y(\result[17] ));
  AOI21X1  g1235(.A0(new_n823_), .A1(new_n812_), .B0(new_n310_), .Y(new_n1499_));
  AOI21X1  g1236(.A0(new_n869_), .A1(new_n858_), .B0(new_n351_), .Y(new_n1500_));
  AOI21X1  g1237(.A0(new_n916_), .A1(new_n905_), .B0(new_n391_), .Y(new_n1501_));
  AOI21X1  g1238(.A0(new_n846_), .A1(new_n835_), .B0(new_n431_), .Y(new_n1502_));
  OR4X1    g1239(.A(new_n1502_), .B(new_n1501_), .C(new_n1500_), .D(new_n1499_), .Y(new_n1503_));
  AOI21X1  g1240(.A0(new_n893_), .A1(new_n882_), .B0(new_n431_), .Y(new_n1504_));
  AOI21X1  g1241(.A0(new_n800_), .A1(new_n789_), .B0(new_n391_), .Y(new_n1505_));
  AOI21X1  g1242(.A0(new_n939_), .A1(new_n928_), .B0(new_n351_), .Y(new_n1506_));
  AOI21X1  g1243(.A0(new_n962_), .A1(new_n951_), .B0(new_n310_), .Y(new_n1507_));
  OR4X1    g1244(.A(new_n1507_), .B(new_n1506_), .C(new_n1505_), .D(new_n1504_), .Y(new_n1508_));
  MX2X1    g1245(.A(new_n1508_), .B(new_n1503_), .S0(new_n264_), .Y(\result[18] ));
  AOI21X1  g1246(.A0(new_n987_), .A1(new_n976_), .B0(new_n351_), .Y(new_n1510_));
  AOI21X1  g1247(.A0(new_n1010_), .A1(new_n999_), .B0(new_n310_), .Y(new_n1511_));
  AOI21X1  g1248(.A0(new_n1033_), .A1(new_n1022_), .B0(new_n431_), .Y(new_n1512_));
  AOI21X1  g1249(.A0(new_n1126_), .A1(new_n1115_), .B0(new_n391_), .Y(new_n1513_));
  OR4X1    g1250(.A(new_n1513_), .B(new_n1512_), .C(new_n1511_), .D(new_n1510_), .Y(new_n1514_));
  AOI21X1  g1251(.A0(new_n1080_), .A1(new_n1069_), .B0(new_n431_), .Y(new_n1515_));
  AOI21X1  g1252(.A0(new_n1056_), .A1(new_n1045_), .B0(new_n391_), .Y(new_n1516_));
  AOI21X1  g1253(.A0(new_n1149_), .A1(new_n1138_), .B0(new_n310_), .Y(new_n1517_));
  AOI21X1  g1254(.A0(new_n1103_), .A1(new_n1092_), .B0(new_n351_), .Y(new_n1518_));
  OR4X1    g1255(.A(new_n1518_), .B(new_n1517_), .C(new_n1516_), .D(new_n1515_), .Y(new_n1519_));
  MX2X1    g1256(.A(new_n1519_), .B(new_n1514_), .S0(new_n264_), .Y(\result[19] ));
  AOI21X1  g1257(.A0(new_n1157_), .A1(new_n1156_), .B0(new_n310_), .Y(new_n1521_));
  AOI21X1  g1258(.A0(new_n1163_), .A1(new_n1162_), .B0(new_n351_), .Y(new_n1522_));
  AOI21X1  g1259(.A0(new_n1176_), .A1(new_n1175_), .B0(new_n391_), .Y(new_n1523_));
  AOI21X1  g1260(.A0(new_n1160_), .A1(new_n1159_), .B0(new_n431_), .Y(new_n1524_));
  OR4X1    g1261(.A(new_n1524_), .B(new_n1523_), .C(new_n1522_), .D(new_n1521_), .Y(new_n1525_));
  AOI21X1  g1262(.A0(new_n1154_), .A1(new_n1153_), .B0(new_n391_), .Y(new_n1526_));
  AOI21X1  g1263(.A0(new_n1167_), .A1(new_n1166_), .B0(new_n351_), .Y(new_n1527_));
  AOI21X1  g1264(.A0(new_n1173_), .A1(new_n1172_), .B0(new_n310_), .Y(new_n1528_));
  AOI21X1  g1265(.A0(new_n1170_), .A1(new_n1169_), .B0(new_n431_), .Y(new_n1529_));
  OR4X1    g1266(.A(new_n1529_), .B(new_n1528_), .C(new_n1527_), .D(new_n1526_), .Y(new_n1530_));
  MX2X1    g1267(.A(new_n1530_), .B(new_n1525_), .S0(new_n264_), .Y(\result[20] ));
  AOI21X1  g1268(.A0(new_n1184_), .A1(new_n1183_), .B0(new_n310_), .Y(new_n1532_));
  AOI21X1  g1269(.A0(new_n1190_), .A1(new_n1189_), .B0(new_n351_), .Y(new_n1533_));
  AOI21X1  g1270(.A0(new_n1203_), .A1(new_n1202_), .B0(new_n391_), .Y(new_n1534_));
  AOI21X1  g1271(.A0(new_n1187_), .A1(new_n1186_), .B0(new_n431_), .Y(new_n1535_));
  OR4X1    g1272(.A(new_n1535_), .B(new_n1534_), .C(new_n1533_), .D(new_n1532_), .Y(new_n1536_));
  AOI21X1  g1273(.A0(new_n1181_), .A1(new_n1180_), .B0(new_n391_), .Y(new_n1537_));
  AOI21X1  g1274(.A0(new_n1194_), .A1(new_n1193_), .B0(new_n351_), .Y(new_n1538_));
  AOI21X1  g1275(.A0(new_n1200_), .A1(new_n1199_), .B0(new_n310_), .Y(new_n1539_));
  AOI21X1  g1276(.A0(new_n1197_), .A1(new_n1196_), .B0(new_n431_), .Y(new_n1540_));
  OR4X1    g1277(.A(new_n1540_), .B(new_n1539_), .C(new_n1538_), .D(new_n1537_), .Y(new_n1541_));
  MX2X1    g1278(.A(new_n1541_), .B(new_n1536_), .S0(new_n264_), .Y(\result[21] ));
  AOI21X1  g1279(.A0(new_n1211_), .A1(new_n1210_), .B0(new_n310_), .Y(new_n1543_));
  AOI21X1  g1280(.A0(new_n1217_), .A1(new_n1216_), .B0(new_n351_), .Y(new_n1544_));
  AOI21X1  g1281(.A0(new_n1230_), .A1(new_n1229_), .B0(new_n391_), .Y(new_n1545_));
  AOI21X1  g1282(.A0(new_n1214_), .A1(new_n1213_), .B0(new_n431_), .Y(new_n1546_));
  OR4X1    g1283(.A(new_n1546_), .B(new_n1545_), .C(new_n1544_), .D(new_n1543_), .Y(new_n1547_));
  AOI21X1  g1284(.A0(new_n1208_), .A1(new_n1207_), .B0(new_n391_), .Y(new_n1548_));
  AOI21X1  g1285(.A0(new_n1221_), .A1(new_n1220_), .B0(new_n351_), .Y(new_n1549_));
  AOI21X1  g1286(.A0(new_n1227_), .A1(new_n1226_), .B0(new_n310_), .Y(new_n1550_));
  AOI21X1  g1287(.A0(new_n1224_), .A1(new_n1223_), .B0(new_n431_), .Y(new_n1551_));
  OR4X1    g1288(.A(new_n1551_), .B(new_n1550_), .C(new_n1549_), .D(new_n1548_), .Y(new_n1552_));
  MX2X1    g1289(.A(new_n1552_), .B(new_n1547_), .S0(new_n264_), .Y(\result[22] ));
  AOI21X1  g1290(.A0(new_n1238_), .A1(new_n1237_), .B0(new_n310_), .Y(new_n1554_));
  AOI21X1  g1291(.A0(new_n1257_), .A1(new_n1256_), .B0(new_n391_), .Y(new_n1555_));
  AOI21X1  g1292(.A0(new_n1241_), .A1(new_n1240_), .B0(new_n431_), .Y(new_n1556_));
  AOI21X1  g1293(.A0(new_n1244_), .A1(new_n1243_), .B0(new_n351_), .Y(new_n1557_));
  OR4X1    g1294(.A(new_n1557_), .B(new_n1556_), .C(new_n1555_), .D(new_n1554_), .Y(new_n1558_));
  AOI21X1  g1295(.A0(new_n1248_), .A1(new_n1247_), .B0(new_n351_), .Y(new_n1559_));
  AOI21X1  g1296(.A0(new_n1251_), .A1(new_n1250_), .B0(new_n431_), .Y(new_n1560_));
  AOI21X1  g1297(.A0(new_n1254_), .A1(new_n1253_), .B0(new_n310_), .Y(new_n1561_));
  AOI21X1  g1298(.A0(new_n1235_), .A1(new_n1234_), .B0(new_n391_), .Y(new_n1562_));
  OR4X1    g1299(.A(new_n1562_), .B(new_n1561_), .C(new_n1560_), .D(new_n1559_), .Y(new_n1563_));
  MX2X1    g1300(.A(new_n1563_), .B(new_n1558_), .S0(new_n264_), .Y(\result[23] ));
  AOI21X1  g1301(.A0(new_n1265_), .A1(new_n1264_), .B0(new_n310_), .Y(new_n1565_));
  AOI21X1  g1302(.A0(new_n1284_), .A1(new_n1283_), .B0(new_n391_), .Y(new_n1566_));
  AOI21X1  g1303(.A0(new_n1268_), .A1(new_n1267_), .B0(new_n431_), .Y(new_n1567_));
  AOI21X1  g1304(.A0(new_n1271_), .A1(new_n1270_), .B0(new_n351_), .Y(new_n1568_));
  OR4X1    g1305(.A(new_n1568_), .B(new_n1567_), .C(new_n1566_), .D(new_n1565_), .Y(new_n1569_));
  AOI21X1  g1306(.A0(new_n1275_), .A1(new_n1274_), .B0(new_n351_), .Y(new_n1570_));
  AOI21X1  g1307(.A0(new_n1278_), .A1(new_n1277_), .B0(new_n431_), .Y(new_n1571_));
  AOI21X1  g1308(.A0(new_n1281_), .A1(new_n1280_), .B0(new_n310_), .Y(new_n1572_));
  AOI21X1  g1309(.A0(new_n1262_), .A1(new_n1261_), .B0(new_n391_), .Y(new_n1573_));
  OR4X1    g1310(.A(new_n1573_), .B(new_n1572_), .C(new_n1571_), .D(new_n1570_), .Y(new_n1574_));
  MX2X1    g1311(.A(new_n1574_), .B(new_n1569_), .S0(new_n264_), .Y(\result[24] ));
  AOI21X1  g1312(.A0(new_n1292_), .A1(new_n1291_), .B0(new_n310_), .Y(new_n1576_));
  AOI21X1  g1313(.A0(new_n1311_), .A1(new_n1310_), .B0(new_n391_), .Y(new_n1577_));
  AOI21X1  g1314(.A0(new_n1295_), .A1(new_n1294_), .B0(new_n431_), .Y(new_n1578_));
  AOI21X1  g1315(.A0(new_n1298_), .A1(new_n1297_), .B0(new_n351_), .Y(new_n1579_));
  OR4X1    g1316(.A(new_n1579_), .B(new_n1578_), .C(new_n1577_), .D(new_n1576_), .Y(new_n1580_));
  AOI21X1  g1317(.A0(new_n1302_), .A1(new_n1301_), .B0(new_n351_), .Y(new_n1581_));
  AOI21X1  g1318(.A0(new_n1305_), .A1(new_n1304_), .B0(new_n431_), .Y(new_n1582_));
  AOI21X1  g1319(.A0(new_n1308_), .A1(new_n1307_), .B0(new_n310_), .Y(new_n1583_));
  AOI21X1  g1320(.A0(new_n1289_), .A1(new_n1288_), .B0(new_n391_), .Y(new_n1584_));
  OR4X1    g1321(.A(new_n1584_), .B(new_n1583_), .C(new_n1582_), .D(new_n1581_), .Y(new_n1585_));
  MX2X1    g1322(.A(new_n1585_), .B(new_n1580_), .S0(new_n264_), .Y(\result[25] ));
  AOI21X1  g1323(.A0(new_n1319_), .A1(new_n1318_), .B0(new_n310_), .Y(new_n1587_));
  AOI21X1  g1324(.A0(new_n1325_), .A1(new_n1324_), .B0(new_n351_), .Y(new_n1588_));
  AOI21X1  g1325(.A0(new_n1338_), .A1(new_n1337_), .B0(new_n391_), .Y(new_n1589_));
  AOI21X1  g1326(.A0(new_n1322_), .A1(new_n1321_), .B0(new_n431_), .Y(new_n1590_));
  OR4X1    g1327(.A(new_n1590_), .B(new_n1589_), .C(new_n1588_), .D(new_n1587_), .Y(new_n1591_));
  AOI21X1  g1328(.A0(new_n1329_), .A1(new_n1328_), .B0(new_n351_), .Y(new_n1592_));
  AOI21X1  g1329(.A0(new_n1332_), .A1(new_n1331_), .B0(new_n431_), .Y(new_n1593_));
  AOI21X1  g1330(.A0(new_n1335_), .A1(new_n1334_), .B0(new_n310_), .Y(new_n1594_));
  AOI21X1  g1331(.A0(new_n1316_), .A1(new_n1315_), .B0(new_n391_), .Y(new_n1595_));
  OR4X1    g1332(.A(new_n1595_), .B(new_n1594_), .C(new_n1593_), .D(new_n1592_), .Y(new_n1596_));
  MX2X1    g1333(.A(new_n1596_), .B(new_n1591_), .S0(new_n264_), .Y(\result[26] ));
  AOI21X1  g1334(.A0(new_n1346_), .A1(new_n1345_), .B0(new_n310_), .Y(new_n1598_));
  AOI21X1  g1335(.A0(new_n1352_), .A1(new_n1351_), .B0(new_n351_), .Y(new_n1599_));
  AOI21X1  g1336(.A0(new_n1365_), .A1(new_n1364_), .B0(new_n391_), .Y(new_n1600_));
  AOI21X1  g1337(.A0(new_n1349_), .A1(new_n1348_), .B0(new_n431_), .Y(new_n1601_));
  OR4X1    g1338(.A(new_n1601_), .B(new_n1600_), .C(new_n1599_), .D(new_n1598_), .Y(new_n1602_));
  AOI21X1  g1339(.A0(new_n1356_), .A1(new_n1355_), .B0(new_n351_), .Y(new_n1603_));
  AOI21X1  g1340(.A0(new_n1359_), .A1(new_n1358_), .B0(new_n431_), .Y(new_n1604_));
  AOI21X1  g1341(.A0(new_n1362_), .A1(new_n1361_), .B0(new_n310_), .Y(new_n1605_));
  AOI21X1  g1342(.A0(new_n1343_), .A1(new_n1342_), .B0(new_n391_), .Y(new_n1606_));
  OR4X1    g1343(.A(new_n1606_), .B(new_n1605_), .C(new_n1604_), .D(new_n1603_), .Y(new_n1607_));
  MX2X1    g1344(.A(new_n1607_), .B(new_n1602_), .S0(new_n264_), .Y(\result[27] ));
  AOI21X1  g1345(.A0(new_n1373_), .A1(new_n1372_), .B0(new_n310_), .Y(new_n1609_));
  AOI21X1  g1346(.A0(new_n1379_), .A1(new_n1378_), .B0(new_n351_), .Y(new_n1610_));
  AOI21X1  g1347(.A0(new_n1392_), .A1(new_n1391_), .B0(new_n391_), .Y(new_n1611_));
  AOI21X1  g1348(.A0(new_n1376_), .A1(new_n1375_), .B0(new_n431_), .Y(new_n1612_));
  OR4X1    g1349(.A(new_n1612_), .B(new_n1611_), .C(new_n1610_), .D(new_n1609_), .Y(new_n1613_));
  AOI21X1  g1350(.A0(new_n1383_), .A1(new_n1382_), .B0(new_n351_), .Y(new_n1614_));
  AOI21X1  g1351(.A0(new_n1386_), .A1(new_n1385_), .B0(new_n431_), .Y(new_n1615_));
  AOI21X1  g1352(.A0(new_n1389_), .A1(new_n1388_), .B0(new_n310_), .Y(new_n1616_));
  AOI21X1  g1353(.A0(new_n1370_), .A1(new_n1369_), .B0(new_n391_), .Y(new_n1617_));
  OR4X1    g1354(.A(new_n1617_), .B(new_n1616_), .C(new_n1615_), .D(new_n1614_), .Y(new_n1618_));
  MX2X1    g1355(.A(new_n1618_), .B(new_n1613_), .S0(new_n264_), .Y(\result[28] ));
  AOI21X1  g1356(.A0(new_n1400_), .A1(new_n1399_), .B0(new_n310_), .Y(new_n1620_));
  AOI21X1  g1357(.A0(new_n1406_), .A1(new_n1405_), .B0(new_n351_), .Y(new_n1621_));
  AOI21X1  g1358(.A0(new_n1419_), .A1(new_n1418_), .B0(new_n391_), .Y(new_n1622_));
  AOI21X1  g1359(.A0(new_n1403_), .A1(new_n1402_), .B0(new_n431_), .Y(new_n1623_));
  OR4X1    g1360(.A(new_n1623_), .B(new_n1622_), .C(new_n1621_), .D(new_n1620_), .Y(new_n1624_));
  AOI21X1  g1361(.A0(new_n1410_), .A1(new_n1409_), .B0(new_n351_), .Y(new_n1625_));
  AOI21X1  g1362(.A0(new_n1413_), .A1(new_n1412_), .B0(new_n431_), .Y(new_n1626_));
  AOI21X1  g1363(.A0(new_n1416_), .A1(new_n1415_), .B0(new_n310_), .Y(new_n1627_));
  AOI21X1  g1364(.A0(new_n1397_), .A1(new_n1396_), .B0(new_n391_), .Y(new_n1628_));
  OR4X1    g1365(.A(new_n1628_), .B(new_n1627_), .C(new_n1626_), .D(new_n1625_), .Y(new_n1629_));
  MX2X1    g1366(.A(new_n1629_), .B(new_n1624_), .S0(new_n264_), .Y(\result[29] ));
  AOI21X1  g1367(.A0(new_n1427_), .A1(new_n1426_), .B0(new_n310_), .Y(new_n1631_));
  AOI21X1  g1368(.A0(new_n1433_), .A1(new_n1432_), .B0(new_n351_), .Y(new_n1632_));
  AOI21X1  g1369(.A0(new_n1446_), .A1(new_n1445_), .B0(new_n391_), .Y(new_n1633_));
  AOI21X1  g1370(.A0(new_n1430_), .A1(new_n1429_), .B0(new_n431_), .Y(new_n1634_));
  OR4X1    g1371(.A(new_n1634_), .B(new_n1633_), .C(new_n1632_), .D(new_n1631_), .Y(new_n1635_));
  AOI21X1  g1372(.A0(new_n1437_), .A1(new_n1436_), .B0(new_n351_), .Y(new_n1636_));
  AOI21X1  g1373(.A0(new_n1440_), .A1(new_n1439_), .B0(new_n431_), .Y(new_n1637_));
  AOI21X1  g1374(.A0(new_n1443_), .A1(new_n1442_), .B0(new_n310_), .Y(new_n1638_));
  AOI21X1  g1375(.A0(new_n1424_), .A1(new_n1423_), .B0(new_n391_), .Y(new_n1639_));
  OR4X1    g1376(.A(new_n1639_), .B(new_n1638_), .C(new_n1637_), .D(new_n1636_), .Y(new_n1640_));
  MX2X1    g1377(.A(new_n1640_), .B(new_n1635_), .S0(new_n264_), .Y(\result[30] ));
  AOI21X1  g1378(.A0(new_n1454_), .A1(new_n1453_), .B0(new_n310_), .Y(new_n1642_));
  AOI21X1  g1379(.A0(new_n1460_), .A1(new_n1459_), .B0(new_n351_), .Y(new_n1643_));
  AOI21X1  g1380(.A0(new_n1473_), .A1(new_n1472_), .B0(new_n391_), .Y(new_n1644_));
  AOI21X1  g1381(.A0(new_n1457_), .A1(new_n1456_), .B0(new_n431_), .Y(new_n1645_));
  OR4X1    g1382(.A(new_n1645_), .B(new_n1644_), .C(new_n1643_), .D(new_n1642_), .Y(new_n1646_));
  AOI21X1  g1383(.A0(new_n1464_), .A1(new_n1463_), .B0(new_n351_), .Y(new_n1647_));
  AOI21X1  g1384(.A0(new_n1467_), .A1(new_n1466_), .B0(new_n431_), .Y(new_n1648_));
  AOI21X1  g1385(.A0(new_n1470_), .A1(new_n1469_), .B0(new_n310_), .Y(new_n1649_));
  AOI21X1  g1386(.A0(new_n1451_), .A1(new_n1450_), .B0(new_n391_), .Y(new_n1650_));
  OR4X1    g1387(.A(new_n1650_), .B(new_n1649_), .C(new_n1648_), .D(new_n1647_), .Y(new_n1651_));
  MX2X1    g1388(.A(new_n1651_), .B(new_n1646_), .S0(new_n264_), .Y(\result[31] ));
  AOI21X1  g1389(.A0(new_n430_), .A1(new_n411_), .B0(new_n310_), .Y(new_n1653_));
  AOI21X1  g1390(.A0(new_n390_), .A1(new_n371_), .B0(new_n351_), .Y(new_n1654_));
  AOI21X1  g1391(.A0(new_n510_), .A1(new_n491_), .B0(new_n391_), .Y(new_n1655_));
  AOI21X1  g1392(.A0(new_n471_), .A1(new_n452_), .B0(new_n431_), .Y(new_n1656_));
  OR4X1    g1393(.A(new_n1656_), .B(new_n1655_), .C(new_n1654_), .D(new_n1653_), .Y(new_n1657_));
  AOI21X1  g1394(.A0(new_n309_), .A1(new_n288_), .B0(new_n431_), .Y(new_n1658_));
  AOI21X1  g1395(.A0(new_n349_), .A1(new_n330_), .B0(new_n391_), .Y(new_n1659_));
  AOI21X1  g1396(.A0(new_n549_), .A1(new_n530_), .B0(new_n351_), .Y(new_n1660_));
  AOI21X1  g1397(.A0(new_n588_), .A1(new_n569_), .B0(new_n310_), .Y(new_n1661_));
  OR4X1    g1398(.A(new_n1661_), .B(new_n1660_), .C(new_n1659_), .D(new_n1658_), .Y(new_n1662_));
  MX2X1    g1399(.A(new_n1662_), .B(new_n1657_), .S0(new_n264_), .Y(\result[32] ));
  AOI21X1  g1400(.A0(new_n682_), .A1(new_n671_), .B0(new_n310_), .Y(new_n1664_));
  AOI21X1  g1401(.A0(new_n659_), .A1(new_n648_), .B0(new_n351_), .Y(new_n1665_));
  AOI21X1  g1402(.A0(new_n775_), .A1(new_n764_), .B0(new_n391_), .Y(new_n1666_));
  AOI21X1  g1403(.A0(new_n729_), .A1(new_n718_), .B0(new_n431_), .Y(new_n1667_));
  OR4X1    g1404(.A(new_n1667_), .B(new_n1666_), .C(new_n1665_), .D(new_n1664_), .Y(new_n1668_));
  AOI21X1  g1405(.A0(new_n706_), .A1(new_n695_), .B0(new_n351_), .Y(new_n1669_));
  AOI21X1  g1406(.A0(new_n613_), .A1(new_n602_), .B0(new_n431_), .Y(new_n1670_));
  AOI21X1  g1407(.A0(new_n752_), .A1(new_n741_), .B0(new_n310_), .Y(new_n1671_));
  AOI21X1  g1408(.A0(new_n636_), .A1(new_n625_), .B0(new_n391_), .Y(new_n1672_));
  OR4X1    g1409(.A(new_n1672_), .B(new_n1671_), .C(new_n1670_), .D(new_n1669_), .Y(new_n1673_));
  MX2X1    g1410(.A(new_n1673_), .B(new_n1668_), .S0(new_n264_), .Y(\result[33] ));
  AOI21X1  g1411(.A0(new_n869_), .A1(new_n858_), .B0(new_n310_), .Y(new_n1675_));
  AOI21X1  g1412(.A0(new_n846_), .A1(new_n835_), .B0(new_n351_), .Y(new_n1676_));
  AOI21X1  g1413(.A0(new_n962_), .A1(new_n951_), .B0(new_n391_), .Y(new_n1677_));
  AOI21X1  g1414(.A0(new_n916_), .A1(new_n905_), .B0(new_n431_), .Y(new_n1678_));
  OR4X1    g1415(.A(new_n1678_), .B(new_n1677_), .C(new_n1676_), .D(new_n1675_), .Y(new_n1679_));
  AOI21X1  g1416(.A0(new_n893_), .A1(new_n882_), .B0(new_n351_), .Y(new_n1680_));
  AOI21X1  g1417(.A0(new_n800_), .A1(new_n789_), .B0(new_n431_), .Y(new_n1681_));
  AOI21X1  g1418(.A0(new_n939_), .A1(new_n928_), .B0(new_n310_), .Y(new_n1682_));
  AOI21X1  g1419(.A0(new_n823_), .A1(new_n812_), .B0(new_n391_), .Y(new_n1683_));
  OR4X1    g1420(.A(new_n1683_), .B(new_n1682_), .C(new_n1681_), .D(new_n1680_), .Y(new_n1684_));
  MX2X1    g1421(.A(new_n1684_), .B(new_n1679_), .S0(new_n264_), .Y(\result[34] ));
  AOI21X1  g1422(.A0(new_n987_), .A1(new_n976_), .B0(new_n310_), .Y(new_n1686_));
  AOI21X1  g1423(.A0(new_n1149_), .A1(new_n1138_), .B0(new_n391_), .Y(new_n1687_));
  AOI21X1  g1424(.A0(new_n1033_), .A1(new_n1022_), .B0(new_n351_), .Y(new_n1688_));
  AOI21X1  g1425(.A0(new_n1126_), .A1(new_n1115_), .B0(new_n431_), .Y(new_n1689_));
  OR4X1    g1426(.A(new_n1689_), .B(new_n1688_), .C(new_n1687_), .D(new_n1686_), .Y(new_n1690_));
  AOI21X1  g1427(.A0(new_n1080_), .A1(new_n1069_), .B0(new_n351_), .Y(new_n1691_));
  AOI21X1  g1428(.A0(new_n1010_), .A1(new_n999_), .B0(new_n391_), .Y(new_n1692_));
  AOI21X1  g1429(.A0(new_n1103_), .A1(new_n1092_), .B0(new_n310_), .Y(new_n1693_));
  AOI21X1  g1430(.A0(new_n1056_), .A1(new_n1045_), .B0(new_n431_), .Y(new_n1694_));
  OR4X1    g1431(.A(new_n1694_), .B(new_n1693_), .C(new_n1692_), .D(new_n1691_), .Y(new_n1695_));
  MX2X1    g1432(.A(new_n1695_), .B(new_n1690_), .S0(new_n264_), .Y(\result[35] ));
  AOI21X1  g1433(.A0(new_n1163_), .A1(new_n1162_), .B0(new_n310_), .Y(new_n1697_));
  AOI21X1  g1434(.A0(new_n1160_), .A1(new_n1159_), .B0(new_n351_), .Y(new_n1698_));
  AOI21X1  g1435(.A0(new_n1173_), .A1(new_n1172_), .B0(new_n391_), .Y(new_n1699_));
  AOI21X1  g1436(.A0(new_n1176_), .A1(new_n1175_), .B0(new_n431_), .Y(new_n1700_));
  OR4X1    g1437(.A(new_n1700_), .B(new_n1699_), .C(new_n1698_), .D(new_n1697_), .Y(new_n1701_));
  AOI21X1  g1438(.A0(new_n1154_), .A1(new_n1153_), .B0(new_n431_), .Y(new_n1702_));
  AOI21X1  g1439(.A0(new_n1157_), .A1(new_n1156_), .B0(new_n391_), .Y(new_n1703_));
  AOI21X1  g1440(.A0(new_n1170_), .A1(new_n1169_), .B0(new_n351_), .Y(new_n1704_));
  AOI21X1  g1441(.A0(new_n1167_), .A1(new_n1166_), .B0(new_n310_), .Y(new_n1705_));
  OR4X1    g1442(.A(new_n1705_), .B(new_n1704_), .C(new_n1703_), .D(new_n1702_), .Y(new_n1706_));
  MX2X1    g1443(.A(new_n1706_), .B(new_n1701_), .S0(new_n264_), .Y(\result[36] ));
  AOI21X1  g1444(.A0(new_n1190_), .A1(new_n1189_), .B0(new_n310_), .Y(new_n1708_));
  AOI21X1  g1445(.A0(new_n1187_), .A1(new_n1186_), .B0(new_n351_), .Y(new_n1709_));
  AOI21X1  g1446(.A0(new_n1200_), .A1(new_n1199_), .B0(new_n391_), .Y(new_n1710_));
  AOI21X1  g1447(.A0(new_n1203_), .A1(new_n1202_), .B0(new_n431_), .Y(new_n1711_));
  OR4X1    g1448(.A(new_n1711_), .B(new_n1710_), .C(new_n1709_), .D(new_n1708_), .Y(new_n1712_));
  AOI21X1  g1449(.A0(new_n1181_), .A1(new_n1180_), .B0(new_n431_), .Y(new_n1713_));
  AOI21X1  g1450(.A0(new_n1184_), .A1(new_n1183_), .B0(new_n391_), .Y(new_n1714_));
  AOI21X1  g1451(.A0(new_n1197_), .A1(new_n1196_), .B0(new_n351_), .Y(new_n1715_));
  AOI21X1  g1452(.A0(new_n1194_), .A1(new_n1193_), .B0(new_n310_), .Y(new_n1716_));
  OR4X1    g1453(.A(new_n1716_), .B(new_n1715_), .C(new_n1714_), .D(new_n1713_), .Y(new_n1717_));
  MX2X1    g1454(.A(new_n1717_), .B(new_n1712_), .S0(new_n264_), .Y(\result[37] ));
  AOI21X1  g1455(.A0(new_n1217_), .A1(new_n1216_), .B0(new_n310_), .Y(new_n1719_));
  AOI21X1  g1456(.A0(new_n1214_), .A1(new_n1213_), .B0(new_n351_), .Y(new_n1720_));
  AOI21X1  g1457(.A0(new_n1227_), .A1(new_n1226_), .B0(new_n391_), .Y(new_n1721_));
  AOI21X1  g1458(.A0(new_n1230_), .A1(new_n1229_), .B0(new_n431_), .Y(new_n1722_));
  OR4X1    g1459(.A(new_n1722_), .B(new_n1721_), .C(new_n1720_), .D(new_n1719_), .Y(new_n1723_));
  AOI21X1  g1460(.A0(new_n1208_), .A1(new_n1207_), .B0(new_n431_), .Y(new_n1724_));
  AOI21X1  g1461(.A0(new_n1211_), .A1(new_n1210_), .B0(new_n391_), .Y(new_n1725_));
  AOI21X1  g1462(.A0(new_n1224_), .A1(new_n1223_), .B0(new_n351_), .Y(new_n1726_));
  AOI21X1  g1463(.A0(new_n1221_), .A1(new_n1220_), .B0(new_n310_), .Y(new_n1727_));
  OR4X1    g1464(.A(new_n1727_), .B(new_n1726_), .C(new_n1725_), .D(new_n1724_), .Y(new_n1728_));
  MX2X1    g1465(.A(new_n1728_), .B(new_n1723_), .S0(new_n264_), .Y(\result[38] ));
  AOI21X1  g1466(.A0(new_n1257_), .A1(new_n1256_), .B0(new_n431_), .Y(new_n1730_));
  AOI21X1  g1467(.A0(new_n1254_), .A1(new_n1253_), .B0(new_n391_), .Y(new_n1731_));
  AOI21X1  g1468(.A0(new_n1241_), .A1(new_n1240_), .B0(new_n351_), .Y(new_n1732_));
  AOI21X1  g1469(.A0(new_n1244_), .A1(new_n1243_), .B0(new_n310_), .Y(new_n1733_));
  OR4X1    g1470(.A(new_n1733_), .B(new_n1732_), .C(new_n1731_), .D(new_n1730_), .Y(new_n1734_));
  AOI21X1  g1471(.A0(new_n1248_), .A1(new_n1247_), .B0(new_n310_), .Y(new_n1735_));
  AOI21X1  g1472(.A0(new_n1251_), .A1(new_n1250_), .B0(new_n351_), .Y(new_n1736_));
  AOI21X1  g1473(.A0(new_n1238_), .A1(new_n1237_), .B0(new_n391_), .Y(new_n1737_));
  AOI21X1  g1474(.A0(new_n1235_), .A1(new_n1234_), .B0(new_n431_), .Y(new_n1738_));
  OR4X1    g1475(.A(new_n1738_), .B(new_n1737_), .C(new_n1736_), .D(new_n1735_), .Y(new_n1739_));
  MX2X1    g1476(.A(new_n1739_), .B(new_n1734_), .S0(new_n264_), .Y(\result[39] ));
  AOI21X1  g1477(.A0(new_n1284_), .A1(new_n1283_), .B0(new_n431_), .Y(new_n1741_));
  AOI21X1  g1478(.A0(new_n1281_), .A1(new_n1280_), .B0(new_n391_), .Y(new_n1742_));
  AOI21X1  g1479(.A0(new_n1268_), .A1(new_n1267_), .B0(new_n351_), .Y(new_n1743_));
  AOI21X1  g1480(.A0(new_n1271_), .A1(new_n1270_), .B0(new_n310_), .Y(new_n1744_));
  OR4X1    g1481(.A(new_n1744_), .B(new_n1743_), .C(new_n1742_), .D(new_n1741_), .Y(new_n1745_));
  AOI21X1  g1482(.A0(new_n1275_), .A1(new_n1274_), .B0(new_n310_), .Y(new_n1746_));
  AOI21X1  g1483(.A0(new_n1278_), .A1(new_n1277_), .B0(new_n351_), .Y(new_n1747_));
  AOI21X1  g1484(.A0(new_n1265_), .A1(new_n1264_), .B0(new_n391_), .Y(new_n1748_));
  AOI21X1  g1485(.A0(new_n1262_), .A1(new_n1261_), .B0(new_n431_), .Y(new_n1749_));
  OR4X1    g1486(.A(new_n1749_), .B(new_n1748_), .C(new_n1747_), .D(new_n1746_), .Y(new_n1750_));
  MX2X1    g1487(.A(new_n1750_), .B(new_n1745_), .S0(new_n264_), .Y(\result[40] ));
  AOI21X1  g1488(.A0(new_n1311_), .A1(new_n1310_), .B0(new_n431_), .Y(new_n1752_));
  AOI21X1  g1489(.A0(new_n1308_), .A1(new_n1307_), .B0(new_n391_), .Y(new_n1753_));
  AOI21X1  g1490(.A0(new_n1295_), .A1(new_n1294_), .B0(new_n351_), .Y(new_n1754_));
  AOI21X1  g1491(.A0(new_n1298_), .A1(new_n1297_), .B0(new_n310_), .Y(new_n1755_));
  OR4X1    g1492(.A(new_n1755_), .B(new_n1754_), .C(new_n1753_), .D(new_n1752_), .Y(new_n1756_));
  AOI21X1  g1493(.A0(new_n1302_), .A1(new_n1301_), .B0(new_n310_), .Y(new_n1757_));
  AOI21X1  g1494(.A0(new_n1305_), .A1(new_n1304_), .B0(new_n351_), .Y(new_n1758_));
  AOI21X1  g1495(.A0(new_n1292_), .A1(new_n1291_), .B0(new_n391_), .Y(new_n1759_));
  AOI21X1  g1496(.A0(new_n1289_), .A1(new_n1288_), .B0(new_n431_), .Y(new_n1760_));
  OR4X1    g1497(.A(new_n1760_), .B(new_n1759_), .C(new_n1758_), .D(new_n1757_), .Y(new_n1761_));
  MX2X1    g1498(.A(new_n1761_), .B(new_n1756_), .S0(new_n264_), .Y(\result[41] ));
  AOI21X1  g1499(.A0(new_n1325_), .A1(new_n1324_), .B0(new_n310_), .Y(new_n1763_));
  AOI21X1  g1500(.A0(new_n1322_), .A1(new_n1321_), .B0(new_n351_), .Y(new_n1764_));
  AOI21X1  g1501(.A0(new_n1335_), .A1(new_n1334_), .B0(new_n391_), .Y(new_n1765_));
  AOI21X1  g1502(.A0(new_n1338_), .A1(new_n1337_), .B0(new_n431_), .Y(new_n1766_));
  OR4X1    g1503(.A(new_n1766_), .B(new_n1765_), .C(new_n1764_), .D(new_n1763_), .Y(new_n1767_));
  AOI21X1  g1504(.A0(new_n1329_), .A1(new_n1328_), .B0(new_n310_), .Y(new_n1768_));
  AOI21X1  g1505(.A0(new_n1332_), .A1(new_n1331_), .B0(new_n351_), .Y(new_n1769_));
  AOI21X1  g1506(.A0(new_n1319_), .A1(new_n1318_), .B0(new_n391_), .Y(new_n1770_));
  AOI21X1  g1507(.A0(new_n1316_), .A1(new_n1315_), .B0(new_n431_), .Y(new_n1771_));
  OR4X1    g1508(.A(new_n1771_), .B(new_n1770_), .C(new_n1769_), .D(new_n1768_), .Y(new_n1772_));
  MX2X1    g1509(.A(new_n1772_), .B(new_n1767_), .S0(new_n264_), .Y(\result[42] ));
  AOI21X1  g1510(.A0(new_n1352_), .A1(new_n1351_), .B0(new_n310_), .Y(new_n1774_));
  AOI21X1  g1511(.A0(new_n1349_), .A1(new_n1348_), .B0(new_n351_), .Y(new_n1775_));
  AOI21X1  g1512(.A0(new_n1362_), .A1(new_n1361_), .B0(new_n391_), .Y(new_n1776_));
  AOI21X1  g1513(.A0(new_n1365_), .A1(new_n1364_), .B0(new_n431_), .Y(new_n1777_));
  OR4X1    g1514(.A(new_n1777_), .B(new_n1776_), .C(new_n1775_), .D(new_n1774_), .Y(new_n1778_));
  AOI21X1  g1515(.A0(new_n1356_), .A1(new_n1355_), .B0(new_n310_), .Y(new_n1779_));
  AOI21X1  g1516(.A0(new_n1359_), .A1(new_n1358_), .B0(new_n351_), .Y(new_n1780_));
  AOI21X1  g1517(.A0(new_n1346_), .A1(new_n1345_), .B0(new_n391_), .Y(new_n1781_));
  AOI21X1  g1518(.A0(new_n1343_), .A1(new_n1342_), .B0(new_n431_), .Y(new_n1782_));
  OR4X1    g1519(.A(new_n1782_), .B(new_n1781_), .C(new_n1780_), .D(new_n1779_), .Y(new_n1783_));
  MX2X1    g1520(.A(new_n1783_), .B(new_n1778_), .S0(new_n264_), .Y(\result[43] ));
  AOI21X1  g1521(.A0(new_n1379_), .A1(new_n1378_), .B0(new_n310_), .Y(new_n1785_));
  AOI21X1  g1522(.A0(new_n1376_), .A1(new_n1375_), .B0(new_n351_), .Y(new_n1786_));
  AOI21X1  g1523(.A0(new_n1389_), .A1(new_n1388_), .B0(new_n391_), .Y(new_n1787_));
  AOI21X1  g1524(.A0(new_n1392_), .A1(new_n1391_), .B0(new_n431_), .Y(new_n1788_));
  OR4X1    g1525(.A(new_n1788_), .B(new_n1787_), .C(new_n1786_), .D(new_n1785_), .Y(new_n1789_));
  AOI21X1  g1526(.A0(new_n1383_), .A1(new_n1382_), .B0(new_n310_), .Y(new_n1790_));
  AOI21X1  g1527(.A0(new_n1386_), .A1(new_n1385_), .B0(new_n351_), .Y(new_n1791_));
  AOI21X1  g1528(.A0(new_n1373_), .A1(new_n1372_), .B0(new_n391_), .Y(new_n1792_));
  AOI21X1  g1529(.A0(new_n1370_), .A1(new_n1369_), .B0(new_n431_), .Y(new_n1793_));
  OR4X1    g1530(.A(new_n1793_), .B(new_n1792_), .C(new_n1791_), .D(new_n1790_), .Y(new_n1794_));
  MX2X1    g1531(.A(new_n1794_), .B(new_n1789_), .S0(new_n264_), .Y(\result[44] ));
  AOI21X1  g1532(.A0(new_n1406_), .A1(new_n1405_), .B0(new_n310_), .Y(new_n1796_));
  AOI21X1  g1533(.A0(new_n1403_), .A1(new_n1402_), .B0(new_n351_), .Y(new_n1797_));
  AOI21X1  g1534(.A0(new_n1416_), .A1(new_n1415_), .B0(new_n391_), .Y(new_n1798_));
  AOI21X1  g1535(.A0(new_n1419_), .A1(new_n1418_), .B0(new_n431_), .Y(new_n1799_));
  OR4X1    g1536(.A(new_n1799_), .B(new_n1798_), .C(new_n1797_), .D(new_n1796_), .Y(new_n1800_));
  AOI21X1  g1537(.A0(new_n1410_), .A1(new_n1409_), .B0(new_n310_), .Y(new_n1801_));
  AOI21X1  g1538(.A0(new_n1413_), .A1(new_n1412_), .B0(new_n351_), .Y(new_n1802_));
  AOI21X1  g1539(.A0(new_n1400_), .A1(new_n1399_), .B0(new_n391_), .Y(new_n1803_));
  AOI21X1  g1540(.A0(new_n1397_), .A1(new_n1396_), .B0(new_n431_), .Y(new_n1804_));
  OR4X1    g1541(.A(new_n1804_), .B(new_n1803_), .C(new_n1802_), .D(new_n1801_), .Y(new_n1805_));
  MX2X1    g1542(.A(new_n1805_), .B(new_n1800_), .S0(new_n264_), .Y(\result[45] ));
  AOI21X1  g1543(.A0(new_n1433_), .A1(new_n1432_), .B0(new_n310_), .Y(new_n1807_));
  AOI21X1  g1544(.A0(new_n1430_), .A1(new_n1429_), .B0(new_n351_), .Y(new_n1808_));
  AOI21X1  g1545(.A0(new_n1443_), .A1(new_n1442_), .B0(new_n391_), .Y(new_n1809_));
  AOI21X1  g1546(.A0(new_n1446_), .A1(new_n1445_), .B0(new_n431_), .Y(new_n1810_));
  OR4X1    g1547(.A(new_n1810_), .B(new_n1809_), .C(new_n1808_), .D(new_n1807_), .Y(new_n1811_));
  AOI21X1  g1548(.A0(new_n1437_), .A1(new_n1436_), .B0(new_n310_), .Y(new_n1812_));
  AOI21X1  g1549(.A0(new_n1440_), .A1(new_n1439_), .B0(new_n351_), .Y(new_n1813_));
  AOI21X1  g1550(.A0(new_n1427_), .A1(new_n1426_), .B0(new_n391_), .Y(new_n1814_));
  AOI21X1  g1551(.A0(new_n1424_), .A1(new_n1423_), .B0(new_n431_), .Y(new_n1815_));
  OR4X1    g1552(.A(new_n1815_), .B(new_n1814_), .C(new_n1813_), .D(new_n1812_), .Y(new_n1816_));
  MX2X1    g1553(.A(new_n1816_), .B(new_n1811_), .S0(new_n264_), .Y(\result[46] ));
  AOI21X1  g1554(.A0(new_n1460_), .A1(new_n1459_), .B0(new_n310_), .Y(new_n1818_));
  AOI21X1  g1555(.A0(new_n1457_), .A1(new_n1456_), .B0(new_n351_), .Y(new_n1819_));
  AOI21X1  g1556(.A0(new_n1470_), .A1(new_n1469_), .B0(new_n391_), .Y(new_n1820_));
  AOI21X1  g1557(.A0(new_n1473_), .A1(new_n1472_), .B0(new_n431_), .Y(new_n1821_));
  OR4X1    g1558(.A(new_n1821_), .B(new_n1820_), .C(new_n1819_), .D(new_n1818_), .Y(new_n1822_));
  AOI21X1  g1559(.A0(new_n1464_), .A1(new_n1463_), .B0(new_n310_), .Y(new_n1823_));
  AOI21X1  g1560(.A0(new_n1467_), .A1(new_n1466_), .B0(new_n351_), .Y(new_n1824_));
  AOI21X1  g1561(.A0(new_n1454_), .A1(new_n1453_), .B0(new_n391_), .Y(new_n1825_));
  AOI21X1  g1562(.A0(new_n1451_), .A1(new_n1450_), .B0(new_n431_), .Y(new_n1826_));
  OR4X1    g1563(.A(new_n1826_), .B(new_n1825_), .C(new_n1824_), .D(new_n1823_), .Y(new_n1827_));
  MX2X1    g1564(.A(new_n1827_), .B(new_n1822_), .S0(new_n264_), .Y(\result[47] ));
  AOI21X1  g1565(.A0(new_n390_), .A1(new_n371_), .B0(new_n310_), .Y(new_n1829_));
  AOI21X1  g1566(.A0(new_n471_), .A1(new_n452_), .B0(new_n351_), .Y(new_n1830_));
  AOI21X1  g1567(.A0(new_n588_), .A1(new_n569_), .B0(new_n391_), .Y(new_n1831_));
  AOI21X1  g1568(.A0(new_n510_), .A1(new_n491_), .B0(new_n431_), .Y(new_n1832_));
  OR4X1    g1569(.A(new_n1832_), .B(new_n1831_), .C(new_n1830_), .D(new_n1829_), .Y(new_n1833_));
  AOI21X1  g1570(.A0(new_n309_), .A1(new_n288_), .B0(new_n351_), .Y(new_n1834_));
  AOI21X1  g1571(.A0(new_n349_), .A1(new_n330_), .B0(new_n431_), .Y(new_n1835_));
  AOI21X1  g1572(.A0(new_n549_), .A1(new_n530_), .B0(new_n310_), .Y(new_n1836_));
  AOI21X1  g1573(.A0(new_n430_), .A1(new_n411_), .B0(new_n391_), .Y(new_n1837_));
  OR4X1    g1574(.A(new_n1837_), .B(new_n1836_), .C(new_n1835_), .D(new_n1834_), .Y(new_n1838_));
  MX2X1    g1575(.A(new_n1838_), .B(new_n1833_), .S0(new_n264_), .Y(\result[48] ));
  AOI21X1  g1576(.A0(new_n659_), .A1(new_n648_), .B0(new_n310_), .Y(new_n1840_));
  AOI21X1  g1577(.A0(new_n729_), .A1(new_n718_), .B0(new_n351_), .Y(new_n1841_));
  AOI21X1  g1578(.A0(new_n752_), .A1(new_n741_), .B0(new_n391_), .Y(new_n1842_));
  AOI21X1  g1579(.A0(new_n775_), .A1(new_n764_), .B0(new_n431_), .Y(new_n1843_));
  OR4X1    g1580(.A(new_n1843_), .B(new_n1842_), .C(new_n1841_), .D(new_n1840_), .Y(new_n1844_));
  AOI21X1  g1581(.A0(new_n706_), .A1(new_n695_), .B0(new_n310_), .Y(new_n1845_));
  AOI21X1  g1582(.A0(new_n613_), .A1(new_n602_), .B0(new_n351_), .Y(new_n1846_));
  AOI21X1  g1583(.A0(new_n682_), .A1(new_n671_), .B0(new_n391_), .Y(new_n1847_));
  AOI21X1  g1584(.A0(new_n636_), .A1(new_n625_), .B0(new_n431_), .Y(new_n1848_));
  OR4X1    g1585(.A(new_n1848_), .B(new_n1847_), .C(new_n1846_), .D(new_n1845_), .Y(new_n1849_));
  MX2X1    g1586(.A(new_n1849_), .B(new_n1844_), .S0(new_n264_), .Y(\result[49] ));
  AOI21X1  g1587(.A0(new_n846_), .A1(new_n835_), .B0(new_n310_), .Y(new_n1851_));
  AOI21X1  g1588(.A0(new_n916_), .A1(new_n905_), .B0(new_n351_), .Y(new_n1852_));
  AOI21X1  g1589(.A0(new_n939_), .A1(new_n928_), .B0(new_n391_), .Y(new_n1853_));
  AOI21X1  g1590(.A0(new_n962_), .A1(new_n951_), .B0(new_n431_), .Y(new_n1854_));
  OR4X1    g1591(.A(new_n1854_), .B(new_n1853_), .C(new_n1852_), .D(new_n1851_), .Y(new_n1855_));
  AOI21X1  g1592(.A0(new_n893_), .A1(new_n882_), .B0(new_n310_), .Y(new_n1856_));
  AOI21X1  g1593(.A0(new_n800_), .A1(new_n789_), .B0(new_n351_), .Y(new_n1857_));
  AOI21X1  g1594(.A0(new_n869_), .A1(new_n858_), .B0(new_n391_), .Y(new_n1858_));
  AOI21X1  g1595(.A0(new_n823_), .A1(new_n812_), .B0(new_n431_), .Y(new_n1859_));
  OR4X1    g1596(.A(new_n1859_), .B(new_n1858_), .C(new_n1857_), .D(new_n1856_), .Y(new_n1860_));
  MX2X1    g1597(.A(new_n1860_), .B(new_n1855_), .S0(new_n264_), .Y(\result[50] ));
  AOI21X1  g1598(.A0(new_n1103_), .A1(new_n1092_), .B0(new_n391_), .Y(new_n1862_));
  AOI21X1  g1599(.A0(new_n1149_), .A1(new_n1138_), .B0(new_n431_), .Y(new_n1863_));
  AOI21X1  g1600(.A0(new_n1033_), .A1(new_n1022_), .B0(new_n310_), .Y(new_n1864_));
  AOI21X1  g1601(.A0(new_n1126_), .A1(new_n1115_), .B0(new_n351_), .Y(new_n1865_));
  OR4X1    g1602(.A(new_n1865_), .B(new_n1864_), .C(new_n1863_), .D(new_n1862_), .Y(new_n1866_));
  AOI21X1  g1603(.A0(new_n1080_), .A1(new_n1069_), .B0(new_n310_), .Y(new_n1867_));
  AOI21X1  g1604(.A0(new_n987_), .A1(new_n976_), .B0(new_n391_), .Y(new_n1868_));
  AOI21X1  g1605(.A0(new_n1056_), .A1(new_n1045_), .B0(new_n351_), .Y(new_n1869_));
  AOI21X1  g1606(.A0(new_n1010_), .A1(new_n999_), .B0(new_n431_), .Y(new_n1870_));
  OR4X1    g1607(.A(new_n1870_), .B(new_n1869_), .C(new_n1868_), .D(new_n1867_), .Y(new_n1871_));
  MX2X1    g1608(.A(new_n1871_), .B(new_n1866_), .S0(new_n264_), .Y(\result[51] ));
  AOI21X1  g1609(.A0(new_n1167_), .A1(new_n1166_), .B0(new_n391_), .Y(new_n1873_));
  AOI21X1  g1610(.A0(new_n1160_), .A1(new_n1159_), .B0(new_n310_), .Y(new_n1874_));
  AOI21X1  g1611(.A0(new_n1173_), .A1(new_n1172_), .B0(new_n431_), .Y(new_n1875_));
  AOI21X1  g1612(.A0(new_n1176_), .A1(new_n1175_), .B0(new_n351_), .Y(new_n1876_));
  OR4X1    g1613(.A(new_n1876_), .B(new_n1875_), .C(new_n1874_), .D(new_n1873_), .Y(new_n1877_));
  AOI21X1  g1614(.A0(new_n1154_), .A1(new_n1153_), .B0(new_n351_), .Y(new_n1878_));
  AOI21X1  g1615(.A0(new_n1157_), .A1(new_n1156_), .B0(new_n431_), .Y(new_n1879_));
  AOI21X1  g1616(.A0(new_n1163_), .A1(new_n1162_), .B0(new_n391_), .Y(new_n1880_));
  AOI21X1  g1617(.A0(new_n1170_), .A1(new_n1169_), .B0(new_n310_), .Y(new_n1881_));
  OR4X1    g1618(.A(new_n1881_), .B(new_n1880_), .C(new_n1879_), .D(new_n1878_), .Y(new_n1882_));
  MX2X1    g1619(.A(new_n1882_), .B(new_n1877_), .S0(new_n264_), .Y(\result[52] ));
  AOI21X1  g1620(.A0(new_n1194_), .A1(new_n1193_), .B0(new_n391_), .Y(new_n1884_));
  AOI21X1  g1621(.A0(new_n1187_), .A1(new_n1186_), .B0(new_n310_), .Y(new_n1885_));
  AOI21X1  g1622(.A0(new_n1200_), .A1(new_n1199_), .B0(new_n431_), .Y(new_n1886_));
  AOI21X1  g1623(.A0(new_n1203_), .A1(new_n1202_), .B0(new_n351_), .Y(new_n1887_));
  OR4X1    g1624(.A(new_n1887_), .B(new_n1886_), .C(new_n1885_), .D(new_n1884_), .Y(new_n1888_));
  AOI21X1  g1625(.A0(new_n1181_), .A1(new_n1180_), .B0(new_n351_), .Y(new_n1889_));
  AOI21X1  g1626(.A0(new_n1184_), .A1(new_n1183_), .B0(new_n431_), .Y(new_n1890_));
  AOI21X1  g1627(.A0(new_n1190_), .A1(new_n1189_), .B0(new_n391_), .Y(new_n1891_));
  AOI21X1  g1628(.A0(new_n1197_), .A1(new_n1196_), .B0(new_n310_), .Y(new_n1892_));
  OR4X1    g1629(.A(new_n1892_), .B(new_n1891_), .C(new_n1890_), .D(new_n1889_), .Y(new_n1893_));
  MX2X1    g1630(.A(new_n1893_), .B(new_n1888_), .S0(new_n264_), .Y(\result[53] ));
  AOI21X1  g1631(.A0(new_n1221_), .A1(new_n1220_), .B0(new_n391_), .Y(new_n1895_));
  AOI21X1  g1632(.A0(new_n1214_), .A1(new_n1213_), .B0(new_n310_), .Y(new_n1896_));
  AOI21X1  g1633(.A0(new_n1227_), .A1(new_n1226_), .B0(new_n431_), .Y(new_n1897_));
  AOI21X1  g1634(.A0(new_n1230_), .A1(new_n1229_), .B0(new_n351_), .Y(new_n1898_));
  OR4X1    g1635(.A(new_n1898_), .B(new_n1897_), .C(new_n1896_), .D(new_n1895_), .Y(new_n1899_));
  AOI21X1  g1636(.A0(new_n1208_), .A1(new_n1207_), .B0(new_n351_), .Y(new_n1900_));
  AOI21X1  g1637(.A0(new_n1211_), .A1(new_n1210_), .B0(new_n431_), .Y(new_n1901_));
  AOI21X1  g1638(.A0(new_n1217_), .A1(new_n1216_), .B0(new_n391_), .Y(new_n1902_));
  AOI21X1  g1639(.A0(new_n1224_), .A1(new_n1223_), .B0(new_n310_), .Y(new_n1903_));
  OR4X1    g1640(.A(new_n1903_), .B(new_n1902_), .C(new_n1901_), .D(new_n1900_), .Y(new_n1904_));
  MX2X1    g1641(.A(new_n1904_), .B(new_n1899_), .S0(new_n264_), .Y(\result[54] ));
  AOI21X1  g1642(.A0(new_n1248_), .A1(new_n1247_), .B0(new_n391_), .Y(new_n1906_));
  AOI21X1  g1643(.A0(new_n1257_), .A1(new_n1256_), .B0(new_n351_), .Y(new_n1907_));
  AOI21X1  g1644(.A0(new_n1241_), .A1(new_n1240_), .B0(new_n310_), .Y(new_n1908_));
  AOI21X1  g1645(.A0(new_n1254_), .A1(new_n1253_), .B0(new_n431_), .Y(new_n1909_));
  OR4X1    g1646(.A(new_n1909_), .B(new_n1908_), .C(new_n1907_), .D(new_n1906_), .Y(new_n1910_));
  AOI21X1  g1647(.A0(new_n1251_), .A1(new_n1250_), .B0(new_n310_), .Y(new_n1911_));
  AOI21X1  g1648(.A0(new_n1235_), .A1(new_n1234_), .B0(new_n351_), .Y(new_n1912_));
  AOI21X1  g1649(.A0(new_n1244_), .A1(new_n1243_), .B0(new_n391_), .Y(new_n1913_));
  AOI21X1  g1650(.A0(new_n1238_), .A1(new_n1237_), .B0(new_n431_), .Y(new_n1914_));
  OR4X1    g1651(.A(new_n1914_), .B(new_n1913_), .C(new_n1912_), .D(new_n1911_), .Y(new_n1915_));
  MX2X1    g1652(.A(new_n1915_), .B(new_n1910_), .S0(new_n264_), .Y(\result[55] ));
  AOI21X1  g1653(.A0(new_n1275_), .A1(new_n1274_), .B0(new_n391_), .Y(new_n1917_));
  AOI21X1  g1654(.A0(new_n1284_), .A1(new_n1283_), .B0(new_n351_), .Y(new_n1918_));
  AOI21X1  g1655(.A0(new_n1268_), .A1(new_n1267_), .B0(new_n310_), .Y(new_n1919_));
  AOI21X1  g1656(.A0(new_n1281_), .A1(new_n1280_), .B0(new_n431_), .Y(new_n1920_));
  OR4X1    g1657(.A(new_n1920_), .B(new_n1919_), .C(new_n1918_), .D(new_n1917_), .Y(new_n1921_));
  AOI21X1  g1658(.A0(new_n1278_), .A1(new_n1277_), .B0(new_n310_), .Y(new_n1922_));
  AOI21X1  g1659(.A0(new_n1262_), .A1(new_n1261_), .B0(new_n351_), .Y(new_n1923_));
  AOI21X1  g1660(.A0(new_n1271_), .A1(new_n1270_), .B0(new_n391_), .Y(new_n1924_));
  AOI21X1  g1661(.A0(new_n1265_), .A1(new_n1264_), .B0(new_n431_), .Y(new_n1925_));
  OR4X1    g1662(.A(new_n1925_), .B(new_n1924_), .C(new_n1923_), .D(new_n1922_), .Y(new_n1926_));
  MX2X1    g1663(.A(new_n1926_), .B(new_n1921_), .S0(new_n264_), .Y(\result[56] ));
  AOI21X1  g1664(.A0(new_n1302_), .A1(new_n1301_), .B0(new_n391_), .Y(new_n1928_));
  AOI21X1  g1665(.A0(new_n1311_), .A1(new_n1310_), .B0(new_n351_), .Y(new_n1929_));
  AOI21X1  g1666(.A0(new_n1295_), .A1(new_n1294_), .B0(new_n310_), .Y(new_n1930_));
  AOI21X1  g1667(.A0(new_n1308_), .A1(new_n1307_), .B0(new_n431_), .Y(new_n1931_));
  OR4X1    g1668(.A(new_n1931_), .B(new_n1930_), .C(new_n1929_), .D(new_n1928_), .Y(new_n1932_));
  AOI21X1  g1669(.A0(new_n1305_), .A1(new_n1304_), .B0(new_n310_), .Y(new_n1933_));
  AOI21X1  g1670(.A0(new_n1289_), .A1(new_n1288_), .B0(new_n351_), .Y(new_n1934_));
  AOI21X1  g1671(.A0(new_n1298_), .A1(new_n1297_), .B0(new_n391_), .Y(new_n1935_));
  AOI21X1  g1672(.A0(new_n1292_), .A1(new_n1291_), .B0(new_n431_), .Y(new_n1936_));
  OR4X1    g1673(.A(new_n1936_), .B(new_n1935_), .C(new_n1934_), .D(new_n1933_), .Y(new_n1937_));
  MX2X1    g1674(.A(new_n1937_), .B(new_n1932_), .S0(new_n264_), .Y(\result[57] ));
  AOI21X1  g1675(.A0(new_n1329_), .A1(new_n1328_), .B0(new_n391_), .Y(new_n1939_));
  AOI21X1  g1676(.A0(new_n1322_), .A1(new_n1321_), .B0(new_n310_), .Y(new_n1940_));
  AOI21X1  g1677(.A0(new_n1335_), .A1(new_n1334_), .B0(new_n431_), .Y(new_n1941_));
  AOI21X1  g1678(.A0(new_n1338_), .A1(new_n1337_), .B0(new_n351_), .Y(new_n1942_));
  OR4X1    g1679(.A(new_n1942_), .B(new_n1941_), .C(new_n1940_), .D(new_n1939_), .Y(new_n1943_));
  AOI21X1  g1680(.A0(new_n1332_), .A1(new_n1331_), .B0(new_n310_), .Y(new_n1944_));
  AOI21X1  g1681(.A0(new_n1316_), .A1(new_n1315_), .B0(new_n351_), .Y(new_n1945_));
  AOI21X1  g1682(.A0(new_n1325_), .A1(new_n1324_), .B0(new_n391_), .Y(new_n1946_));
  AOI21X1  g1683(.A0(new_n1319_), .A1(new_n1318_), .B0(new_n431_), .Y(new_n1947_));
  OR4X1    g1684(.A(new_n1947_), .B(new_n1946_), .C(new_n1945_), .D(new_n1944_), .Y(new_n1948_));
  MX2X1    g1685(.A(new_n1948_), .B(new_n1943_), .S0(new_n264_), .Y(\result[58] ));
  AOI21X1  g1686(.A0(new_n1356_), .A1(new_n1355_), .B0(new_n391_), .Y(new_n1950_));
  AOI21X1  g1687(.A0(new_n1349_), .A1(new_n1348_), .B0(new_n310_), .Y(new_n1951_));
  AOI21X1  g1688(.A0(new_n1362_), .A1(new_n1361_), .B0(new_n431_), .Y(new_n1952_));
  AOI21X1  g1689(.A0(new_n1365_), .A1(new_n1364_), .B0(new_n351_), .Y(new_n1953_));
  OR4X1    g1690(.A(new_n1953_), .B(new_n1952_), .C(new_n1951_), .D(new_n1950_), .Y(new_n1954_));
  AOI21X1  g1691(.A0(new_n1359_), .A1(new_n1358_), .B0(new_n310_), .Y(new_n1955_));
  AOI21X1  g1692(.A0(new_n1343_), .A1(new_n1342_), .B0(new_n351_), .Y(new_n1956_));
  AOI21X1  g1693(.A0(new_n1352_), .A1(new_n1351_), .B0(new_n391_), .Y(new_n1957_));
  AOI21X1  g1694(.A0(new_n1346_), .A1(new_n1345_), .B0(new_n431_), .Y(new_n1958_));
  OR4X1    g1695(.A(new_n1958_), .B(new_n1957_), .C(new_n1956_), .D(new_n1955_), .Y(new_n1959_));
  MX2X1    g1696(.A(new_n1959_), .B(new_n1954_), .S0(new_n264_), .Y(\result[59] ));
  AOI21X1  g1697(.A0(new_n1383_), .A1(new_n1382_), .B0(new_n391_), .Y(new_n1961_));
  AOI21X1  g1698(.A0(new_n1376_), .A1(new_n1375_), .B0(new_n310_), .Y(new_n1962_));
  AOI21X1  g1699(.A0(new_n1389_), .A1(new_n1388_), .B0(new_n431_), .Y(new_n1963_));
  AOI21X1  g1700(.A0(new_n1392_), .A1(new_n1391_), .B0(new_n351_), .Y(new_n1964_));
  OR4X1    g1701(.A(new_n1964_), .B(new_n1963_), .C(new_n1962_), .D(new_n1961_), .Y(new_n1965_));
  AOI21X1  g1702(.A0(new_n1386_), .A1(new_n1385_), .B0(new_n310_), .Y(new_n1966_));
  AOI21X1  g1703(.A0(new_n1370_), .A1(new_n1369_), .B0(new_n351_), .Y(new_n1967_));
  AOI21X1  g1704(.A0(new_n1379_), .A1(new_n1378_), .B0(new_n391_), .Y(new_n1968_));
  AOI21X1  g1705(.A0(new_n1373_), .A1(new_n1372_), .B0(new_n431_), .Y(new_n1969_));
  OR4X1    g1706(.A(new_n1969_), .B(new_n1968_), .C(new_n1967_), .D(new_n1966_), .Y(new_n1970_));
  MX2X1    g1707(.A(new_n1970_), .B(new_n1965_), .S0(new_n264_), .Y(\result[60] ));
  AOI21X1  g1708(.A0(new_n1410_), .A1(new_n1409_), .B0(new_n391_), .Y(new_n1972_));
  AOI21X1  g1709(.A0(new_n1403_), .A1(new_n1402_), .B0(new_n310_), .Y(new_n1973_));
  AOI21X1  g1710(.A0(new_n1416_), .A1(new_n1415_), .B0(new_n431_), .Y(new_n1974_));
  AOI21X1  g1711(.A0(new_n1419_), .A1(new_n1418_), .B0(new_n351_), .Y(new_n1975_));
  OR4X1    g1712(.A(new_n1975_), .B(new_n1974_), .C(new_n1973_), .D(new_n1972_), .Y(new_n1976_));
  AOI21X1  g1713(.A0(new_n1413_), .A1(new_n1412_), .B0(new_n310_), .Y(new_n1977_));
  AOI21X1  g1714(.A0(new_n1397_), .A1(new_n1396_), .B0(new_n351_), .Y(new_n1978_));
  AOI21X1  g1715(.A0(new_n1406_), .A1(new_n1405_), .B0(new_n391_), .Y(new_n1979_));
  AOI21X1  g1716(.A0(new_n1400_), .A1(new_n1399_), .B0(new_n431_), .Y(new_n1980_));
  OR4X1    g1717(.A(new_n1980_), .B(new_n1979_), .C(new_n1978_), .D(new_n1977_), .Y(new_n1981_));
  MX2X1    g1718(.A(new_n1981_), .B(new_n1976_), .S0(new_n264_), .Y(\result[61] ));
  AOI21X1  g1719(.A0(new_n1437_), .A1(new_n1436_), .B0(new_n391_), .Y(new_n1983_));
  AOI21X1  g1720(.A0(new_n1430_), .A1(new_n1429_), .B0(new_n310_), .Y(new_n1984_));
  AOI21X1  g1721(.A0(new_n1443_), .A1(new_n1442_), .B0(new_n431_), .Y(new_n1985_));
  AOI21X1  g1722(.A0(new_n1446_), .A1(new_n1445_), .B0(new_n351_), .Y(new_n1986_));
  OR4X1    g1723(.A(new_n1986_), .B(new_n1985_), .C(new_n1984_), .D(new_n1983_), .Y(new_n1987_));
  AOI21X1  g1724(.A0(new_n1440_), .A1(new_n1439_), .B0(new_n310_), .Y(new_n1988_));
  AOI21X1  g1725(.A0(new_n1424_), .A1(new_n1423_), .B0(new_n351_), .Y(new_n1989_));
  AOI21X1  g1726(.A0(new_n1433_), .A1(new_n1432_), .B0(new_n391_), .Y(new_n1990_));
  AOI21X1  g1727(.A0(new_n1427_), .A1(new_n1426_), .B0(new_n431_), .Y(new_n1991_));
  OR4X1    g1728(.A(new_n1991_), .B(new_n1990_), .C(new_n1989_), .D(new_n1988_), .Y(new_n1992_));
  MX2X1    g1729(.A(new_n1992_), .B(new_n1987_), .S0(new_n264_), .Y(\result[62] ));
  AOI21X1  g1730(.A0(new_n1464_), .A1(new_n1463_), .B0(new_n391_), .Y(new_n1994_));
  AOI21X1  g1731(.A0(new_n1457_), .A1(new_n1456_), .B0(new_n310_), .Y(new_n1995_));
  AOI21X1  g1732(.A0(new_n1470_), .A1(new_n1469_), .B0(new_n431_), .Y(new_n1996_));
  AOI21X1  g1733(.A0(new_n1473_), .A1(new_n1472_), .B0(new_n351_), .Y(new_n1997_));
  OR4X1    g1734(.A(new_n1997_), .B(new_n1996_), .C(new_n1995_), .D(new_n1994_), .Y(new_n1998_));
  AOI21X1  g1735(.A0(new_n1467_), .A1(new_n1466_), .B0(new_n310_), .Y(new_n1999_));
  AOI21X1  g1736(.A0(new_n1451_), .A1(new_n1450_), .B0(new_n351_), .Y(new_n2000_));
  AOI21X1  g1737(.A0(new_n1460_), .A1(new_n1459_), .B0(new_n391_), .Y(new_n2001_));
  AOI21X1  g1738(.A0(new_n1454_), .A1(new_n1453_), .B0(new_n431_), .Y(new_n2002_));
  OR4X1    g1739(.A(new_n2002_), .B(new_n2001_), .C(new_n2000_), .D(new_n1999_), .Y(new_n2003_));
  MX2X1    g1740(.A(new_n2003_), .B(new_n1998_), .S0(new_n264_), .Y(\result[63] ));
  MX2X1    g1741(.A(new_n590_), .B(new_n433_), .S0(\shift[6] ), .Y(\result[64] ));
  MX2X1    g1742(.A(new_n777_), .B(new_n684_), .S0(\shift[6] ), .Y(\result[65] ));
  MX2X1    g1743(.A(new_n964_), .B(new_n871_), .S0(\shift[6] ), .Y(\result[66] ));
  MX2X1    g1744(.A(new_n1151_), .B(new_n1058_), .S0(\shift[6] ), .Y(\result[67] ));
  MX2X1    g1745(.A(new_n1178_), .B(new_n1165_), .S0(\shift[6] ), .Y(\result[68] ));
  MX2X1    g1746(.A(new_n1205_), .B(new_n1192_), .S0(\shift[6] ), .Y(\result[69] ));
  MX2X1    g1747(.A(new_n1232_), .B(new_n1219_), .S0(\shift[6] ), .Y(\result[70] ));
  MX2X1    g1748(.A(new_n1259_), .B(new_n1246_), .S0(\shift[6] ), .Y(\result[71] ));
  MX2X1    g1749(.A(new_n1286_), .B(new_n1273_), .S0(\shift[6] ), .Y(\result[72] ));
  MX2X1    g1750(.A(new_n1313_), .B(new_n1300_), .S0(\shift[6] ), .Y(\result[73] ));
  MX2X1    g1751(.A(new_n1340_), .B(new_n1327_), .S0(\shift[6] ), .Y(\result[74] ));
  MX2X1    g1752(.A(new_n1367_), .B(new_n1354_), .S0(\shift[6] ), .Y(\result[75] ));
  MX2X1    g1753(.A(new_n1394_), .B(new_n1381_), .S0(\shift[6] ), .Y(\result[76] ));
  MX2X1    g1754(.A(new_n1421_), .B(new_n1408_), .S0(\shift[6] ), .Y(\result[77] ));
  MX2X1    g1755(.A(new_n1448_), .B(new_n1435_), .S0(\shift[6] ), .Y(\result[78] ));
  MX2X1    g1756(.A(new_n1475_), .B(new_n1462_), .S0(\shift[6] ), .Y(\result[79] ));
  MX2X1    g1757(.A(new_n1486_), .B(new_n1481_), .S0(\shift[6] ), .Y(\result[80] ));
  MX2X1    g1758(.A(new_n1497_), .B(new_n1492_), .S0(\shift[6] ), .Y(\result[81] ));
  MX2X1    g1759(.A(new_n1508_), .B(new_n1503_), .S0(\shift[6] ), .Y(\result[82] ));
  MX2X1    g1760(.A(new_n1519_), .B(new_n1514_), .S0(\shift[6] ), .Y(\result[83] ));
  MX2X1    g1761(.A(new_n1530_), .B(new_n1525_), .S0(\shift[6] ), .Y(\result[84] ));
  MX2X1    g1762(.A(new_n1541_), .B(new_n1536_), .S0(\shift[6] ), .Y(\result[85] ));
  MX2X1    g1763(.A(new_n1552_), .B(new_n1547_), .S0(\shift[6] ), .Y(\result[86] ));
  MX2X1    g1764(.A(new_n1563_), .B(new_n1558_), .S0(\shift[6] ), .Y(\result[87] ));
  MX2X1    g1765(.A(new_n1574_), .B(new_n1569_), .S0(\shift[6] ), .Y(\result[88] ));
  MX2X1    g1766(.A(new_n1585_), .B(new_n1580_), .S0(\shift[6] ), .Y(\result[89] ));
  MX2X1    g1767(.A(new_n1596_), .B(new_n1591_), .S0(\shift[6] ), .Y(\result[90] ));
  MX2X1    g1768(.A(new_n1607_), .B(new_n1602_), .S0(\shift[6] ), .Y(\result[91] ));
  MX2X1    g1769(.A(new_n1618_), .B(new_n1613_), .S0(\shift[6] ), .Y(\result[92] ));
  MX2X1    g1770(.A(new_n1629_), .B(new_n1624_), .S0(\shift[6] ), .Y(\result[93] ));
  MX2X1    g1771(.A(new_n1640_), .B(new_n1635_), .S0(\shift[6] ), .Y(\result[94] ));
  MX2X1    g1772(.A(new_n1651_), .B(new_n1646_), .S0(\shift[6] ), .Y(\result[95] ));
  MX2X1    g1773(.A(new_n1662_), .B(new_n1657_), .S0(\shift[6] ), .Y(\result[96] ));
  MX2X1    g1774(.A(new_n1673_), .B(new_n1668_), .S0(\shift[6] ), .Y(\result[97] ));
  MX2X1    g1775(.A(new_n1684_), .B(new_n1679_), .S0(\shift[6] ), .Y(\result[98] ));
  MX2X1    g1776(.A(new_n1695_), .B(new_n1690_), .S0(\shift[6] ), .Y(\result[99] ));
  MX2X1    g1777(.A(new_n1706_), .B(new_n1701_), .S0(\shift[6] ), .Y(\result[100] ));
  MX2X1    g1778(.A(new_n1717_), .B(new_n1712_), .S0(\shift[6] ), .Y(\result[101] ));
  MX2X1    g1779(.A(new_n1728_), .B(new_n1723_), .S0(\shift[6] ), .Y(\result[102] ));
  MX2X1    g1780(.A(new_n1739_), .B(new_n1734_), .S0(\shift[6] ), .Y(\result[103] ));
  MX2X1    g1781(.A(new_n1750_), .B(new_n1745_), .S0(\shift[6] ), .Y(\result[104] ));
  MX2X1    g1782(.A(new_n1761_), .B(new_n1756_), .S0(\shift[6] ), .Y(\result[105] ));
  MX2X1    g1783(.A(new_n1772_), .B(new_n1767_), .S0(\shift[6] ), .Y(\result[106] ));
  MX2X1    g1784(.A(new_n1783_), .B(new_n1778_), .S0(\shift[6] ), .Y(\result[107] ));
  MX2X1    g1785(.A(new_n1794_), .B(new_n1789_), .S0(\shift[6] ), .Y(\result[108] ));
  MX2X1    g1786(.A(new_n1805_), .B(new_n1800_), .S0(\shift[6] ), .Y(\result[109] ));
  MX2X1    g1787(.A(new_n1816_), .B(new_n1811_), .S0(\shift[6] ), .Y(\result[110] ));
  MX2X1    g1788(.A(new_n1827_), .B(new_n1822_), .S0(\shift[6] ), .Y(\result[111] ));
  MX2X1    g1789(.A(new_n1838_), .B(new_n1833_), .S0(\shift[6] ), .Y(\result[112] ));
  MX2X1    g1790(.A(new_n1849_), .B(new_n1844_), .S0(\shift[6] ), .Y(\result[113] ));
  MX2X1    g1791(.A(new_n1860_), .B(new_n1855_), .S0(\shift[6] ), .Y(\result[114] ));
  MX2X1    g1792(.A(new_n1871_), .B(new_n1866_), .S0(\shift[6] ), .Y(\result[115] ));
  MX2X1    g1793(.A(new_n1882_), .B(new_n1877_), .S0(\shift[6] ), .Y(\result[116] ));
  MX2X1    g1794(.A(new_n1893_), .B(new_n1888_), .S0(\shift[6] ), .Y(\result[117] ));
  MX2X1    g1795(.A(new_n1904_), .B(new_n1899_), .S0(\shift[6] ), .Y(\result[118] ));
  MX2X1    g1796(.A(new_n1915_), .B(new_n1910_), .S0(\shift[6] ), .Y(\result[119] ));
  MX2X1    g1797(.A(new_n1926_), .B(new_n1921_), .S0(\shift[6] ), .Y(\result[120] ));
  MX2X1    g1798(.A(new_n1937_), .B(new_n1932_), .S0(\shift[6] ), .Y(\result[121] ));
  MX2X1    g1799(.A(new_n1948_), .B(new_n1943_), .S0(\shift[6] ), .Y(\result[122] ));
  MX2X1    g1800(.A(new_n1959_), .B(new_n1954_), .S0(\shift[6] ), .Y(\result[123] ));
  MX2X1    g1801(.A(new_n1970_), .B(new_n1965_), .S0(\shift[6] ), .Y(\result[124] ));
  MX2X1    g1802(.A(new_n1981_), .B(new_n1976_), .S0(\shift[6] ), .Y(\result[125] ));
  MX2X1    g1803(.A(new_n1992_), .B(new_n1987_), .S0(\shift[6] ), .Y(\result[126] ));
  MX2X1    g1804(.A(new_n2003_), .B(new_n1998_), .S0(\shift[6] ), .Y(\result[127] ));
endmodule


