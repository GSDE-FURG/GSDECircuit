//Converted to Combinational (Partial output: n1879) , Module name: s35932_n1879 , Timestamp: 2018-12-03T15:51:08.913058 
module s35932_n1879 ( RESET, TM1, TM0, WX1810, WX2034, WX2162, WX3327, WX3455, WX1970, WX2098, WX3263, WX3391, WX2164, WX2166, WX2168, WX2170, WX2172, WX2130, WX2174, WX2132, WX2176, WX2134, WX2178, WX2136, WX2180, WX2138, WX2182, WX2140, WX2184, WX2142, WX2186, WX2144, WX2188, WX2146, WX2190, WX2148, WX2192, WX2150, WX2152, WX2154, WX2156, WX2158, WX2160, n1879 );
input RESET, TM1, TM0, WX1810, WX2034, WX2162, WX3327, WX3455, WX1970, WX2098, WX3263, WX3391, WX2164, WX2166, WX2168, WX2170, WX2172, WX2130, WX2174, WX2132, WX2176, WX2134, WX2178, WX2136, WX2180, WX2138, WX2182, WX2140, WX2184, WX2142, WX2186, WX2144, WX2188, WX2146, WX2190, WX2148, WX2192, WX2150, WX2152, WX2154, WX2156, WX2158, WX2160;
output n1879;
wire n5827, n6610, n6609_1, n6607, n5539, n6026_1, n6608, n6605, n6600, n6023, n6025, n6602, n6604_1, CRC_OUT_8_15, n6022, n6024, n6601, n6603, n6920, CRC_OUT_8_14, n6918, CRC_OUT_8_13, n6916, CRC_OUT_8_12, n6914_1, CRC_OUT_8_11, n6912, CRC_OUT_8_10, n6911, n6909_1, CRC_OUT_8_31, CRC_OUT_8_9, n6953, n6907, CRC_OUT_8_30, CRC_OUT_8_8, n6951, n6905, CRC_OUT_8_29, CRC_OUT_8_7, n6949_1, n6903, CRC_OUT_8_28, CRC_OUT_8_6, n6947, n6901, CRC_OUT_8_27, CRC_OUT_8_5, n6945, n6899_1, CRC_OUT_8_26, CRC_OUT_8_4, n6943, n6897, CRC_OUT_8_25, CRC_OUT_8_3, n6896, n6941, n6894_1, CRC_OUT_8_24, CRC_OUT_8_2, n6939_1, n6892, CRC_OUT_8_23, CRC_OUT_8_1, n6937, n6890, CRC_OUT_8_22, CRC_OUT_8_0, n6935, n6888, CRC_OUT_8_21, n6933, CRC_OUT_8_20, n6931, CRC_OUT_8_19, n6929_1, CRC_OUT_8_18, n6927, CRC_OUT_8_17, n6925, CRC_OUT_8_16, n6923, n6922;
NOR2X1   g1023(.A(n6610), .B(n5827), .Y(n1879));
INVX1    g0288(.A(RESET), .Y(n5827));
MX2X1    g1022(.A(n6607), .B(n6609_1), .S0(TM1), .Y(n6610));
MX2X1    g1021(.A(n6608), .B(n6026_1), .S0(n5539), .Y(n6609_1));
MX2X1    g1019(.A(n6600), .B(n6605), .S0(n5539), .Y(n6607));
INVX1    g0000(.A(TM0), .Y(n5539));
XOR2X1   g0471(.A(n6025), .B(n6023), .Y(n6026_1));
INVX1    g1020(.A(WX1810), .Y(n6608));
XOR2X1   g1018(.A(n6604_1), .B(n6602), .Y(n6605));
INVX1    g1013(.A(CRC_OUT_8_15), .Y(n6600));
XOR2X1   g0468(.A(n6022), .B(WX2034), .Y(n6023));
XOR2X1   g0470(.A(WX2162), .B(n6024), .Y(n6025));
XOR2X1   g1015(.A(n6601), .B(WX3327), .Y(n6602));
XOR2X1   g1017(.A(WX3455), .B(n6603), .Y(n6604_1));
NOR2X1   g1318(.A(n6920), .B(n5827), .Y(CRC_OUT_8_15));
XOR2X1   g0467(.A(WX1970), .B(TM0), .Y(n6022));
INVX1    g0469(.A(WX2098), .Y(n6024));
XOR2X1   g1014(.A(WX3263), .B(TM0), .Y(n6601));
INVX1    g1016(.A(WX3391), .Y(n6603));
XOR2X1   g1317(.A(CRC_OUT_8_14), .B(WX2162), .Y(n6920));
NOR2X1   g1316(.A(n6918), .B(n5827), .Y(CRC_OUT_8_14));
XOR2X1   g1315(.A(CRC_OUT_8_13), .B(WX2164), .Y(n6918));
NOR2X1   g1314(.A(n6916), .B(n5827), .Y(CRC_OUT_8_13));
XOR2X1   g1313(.A(CRC_OUT_8_12), .B(WX2166), .Y(n6916));
NOR2X1   g1312(.A(n6914_1), .B(n5827), .Y(CRC_OUT_8_12));
XOR2X1   g1311(.A(CRC_OUT_8_11), .B(WX2168), .Y(n6914_1));
NOR2X1   g1310(.A(n6912), .B(n5827), .Y(CRC_OUT_8_11));
XOR2X1   g1309(.A(n6911), .B(CRC_OUT_8_10), .Y(n6912));
NOR2X1   g1307(.A(n6909_1), .B(n5827), .Y(CRC_OUT_8_10));
XOR2X1   g1308(.A(CRC_OUT_8_31), .B(WX2170), .Y(n6911));
XOR2X1   g1306(.A(CRC_OUT_8_9), .B(WX2172), .Y(n6909_1));
NOR2X1   g1351(.A(n6953), .B(n5827), .Y(CRC_OUT_8_31));
NOR2X1   g1305(.A(n6907), .B(n5827), .Y(CRC_OUT_8_9));
XOR2X1   g1350(.A(CRC_OUT_8_30), .B(WX2130), .Y(n6953));
XOR2X1   g1304(.A(CRC_OUT_8_8), .B(WX2174), .Y(n6907));
NOR2X1   g1349(.A(n6951), .B(n5827), .Y(CRC_OUT_8_30));
NOR2X1   g1303(.A(n6905), .B(n5827), .Y(CRC_OUT_8_8));
XOR2X1   g1348(.A(CRC_OUT_8_29), .B(WX2132), .Y(n6951));
XOR2X1   g1302(.A(CRC_OUT_8_7), .B(WX2176), .Y(n6905));
NOR2X1   g1347(.A(n6949_1), .B(n5827), .Y(CRC_OUT_8_29));
NOR2X1   g1301(.A(n6903), .B(n5827), .Y(CRC_OUT_8_7));
XOR2X1   g1346(.A(CRC_OUT_8_28), .B(WX2134), .Y(n6949_1));
XOR2X1   g1300(.A(CRC_OUT_8_6), .B(WX2178), .Y(n6903));
NOR2X1   g1345(.A(n6947), .B(n5827), .Y(CRC_OUT_8_28));
NOR2X1   g1299(.A(n6901), .B(n5827), .Y(CRC_OUT_8_6));
XOR2X1   g1344(.A(CRC_OUT_8_27), .B(WX2136), .Y(n6947));
XOR2X1   g1298(.A(CRC_OUT_8_5), .B(WX2180), .Y(n6901));
NOR2X1   g1343(.A(n6945), .B(n5827), .Y(CRC_OUT_8_27));
NOR2X1   g1297(.A(n6899_1), .B(n5827), .Y(CRC_OUT_8_5));
XOR2X1   g1342(.A(CRC_OUT_8_26), .B(WX2138), .Y(n6945));
XOR2X1   g1296(.A(CRC_OUT_8_4), .B(WX2182), .Y(n6899_1));
NOR2X1   g1341(.A(n6943), .B(n5827), .Y(CRC_OUT_8_26));
NOR2X1   g1295(.A(n6897), .B(n5827), .Y(CRC_OUT_8_4));
XOR2X1   g1340(.A(CRC_OUT_8_25), .B(WX2140), .Y(n6943));
XOR2X1   g1294(.A(n6896), .B(CRC_OUT_8_3), .Y(n6897));
NOR2X1   g1339(.A(n6941), .B(n5827), .Y(CRC_OUT_8_25));
NOR2X1   g1292(.A(n6894_1), .B(n5827), .Y(CRC_OUT_8_3));
XOR2X1   g1293(.A(CRC_OUT_8_31), .B(WX2184), .Y(n6896));
XOR2X1   g1338(.A(CRC_OUT_8_24), .B(WX2142), .Y(n6941));
XOR2X1   g1291(.A(CRC_OUT_8_2), .B(WX2186), .Y(n6894_1));
NOR2X1   g1337(.A(n6939_1), .B(n5827), .Y(CRC_OUT_8_24));
NOR2X1   g1290(.A(n6892), .B(n5827), .Y(CRC_OUT_8_2));
XOR2X1   g1336(.A(CRC_OUT_8_23), .B(WX2144), .Y(n6939_1));
XOR2X1   g1289(.A(CRC_OUT_8_1), .B(WX2188), .Y(n6892));
NOR2X1   g1335(.A(n6937), .B(n5827), .Y(CRC_OUT_8_23));
NOR2X1   g1288(.A(n6890), .B(n5827), .Y(CRC_OUT_8_1));
XOR2X1   g1334(.A(CRC_OUT_8_22), .B(WX2146), .Y(n6937));
XOR2X1   g1287(.A(CRC_OUT_8_0), .B(WX2190), .Y(n6890));
NOR2X1   g1333(.A(n6935), .B(n5827), .Y(CRC_OUT_8_22));
NOR2X1   g1286(.A(n6888), .B(n5827), .Y(CRC_OUT_8_0));
XOR2X1   g1332(.A(CRC_OUT_8_21), .B(WX2148), .Y(n6935));
XOR2X1   g1285(.A(CRC_OUT_8_31), .B(WX2192), .Y(n6888));
NOR2X1   g1331(.A(n6933), .B(n5827), .Y(CRC_OUT_8_21));
XOR2X1   g1330(.A(CRC_OUT_8_20), .B(WX2150), .Y(n6933));
NOR2X1   g1329(.A(n6931), .B(n5827), .Y(CRC_OUT_8_20));
XOR2X1   g1328(.A(CRC_OUT_8_19), .B(WX2152), .Y(n6931));
NOR2X1   g1327(.A(n6929_1), .B(n5827), .Y(CRC_OUT_8_19));
XOR2X1   g1326(.A(CRC_OUT_8_18), .B(WX2154), .Y(n6929_1));
NOR2X1   g1325(.A(n6927), .B(n5827), .Y(CRC_OUT_8_18));
XOR2X1   g1324(.A(CRC_OUT_8_17), .B(WX2156), .Y(n6927));
NOR2X1   g1323(.A(n6925), .B(n5827), .Y(CRC_OUT_8_17));
XOR2X1   g1322(.A(CRC_OUT_8_16), .B(WX2158), .Y(n6925));
NOR2X1   g1321(.A(n6923), .B(n5827), .Y(CRC_OUT_8_16));
XOR2X1   g1320(.A(n6922), .B(CRC_OUT_8_15), .Y(n6923));
XOR2X1   g1319(.A(CRC_OUT_8_31), .B(WX2160), .Y(n6922));

endmodule
