//Converted to Combinational (Partial output: n2809) , Module name: s38584_n2809 , Timestamp: 2018-12-03T15:51:16.598848 
module s38584_n2809 ( g6049, g35, g5990, g93, g4358, g4349, g4311, g113, g4681, g4801, g4793, g4785, g134, g99, g37, g4776, g4653, g4669, g4659, g4754, g4709, g4322, g4332, g72, g73, n2809 );
input g6049, g35, g5990, g93, g4358, g4349, g4311, g113, g4681, g4801, g4793, g4785, g134, g99, g37, g4776, g4653, g4669, g4659, g4754, g4709, g4322, g4332, g72, g73;
output n2809;
wire n7703, n4620, n7702, n7699, n7700, n7701, n6747_1, n7697, n7698, n6466, n6951, n6944, n6746, n5174, n4957, n5506, n6744, n4721, n6745, n4952, n4955, n4809, n4720, n4723, n4814, n4815, n4951, n4954_1, n4950, n4953;
OAI21X1  g3059(.A0(n7702), .A1(n4620), .B0(n7703), .Y(n2809));
NAND2X1  g3058(.A(g6049), .B(n4620), .Y(n7703));
INVX1    g0000(.A(g35), .Y(n4620));
OAI21X1  g3057(.A0(n7701), .A1(n7700), .B0(n7699), .Y(n7702));
OR4X1    g3054(.A(n6466), .B(n7698), .C(n7697), .D(n6747_1), .Y(n7699));
NOR3X1   g3055(.A(n6747_1), .B(n6951), .C(g5990), .Y(n7700));
AOI21X1  g3056(.A0(n6746), .A1(g6049), .B0(n6944), .Y(n7701));
INVX1    g2106(.A(n6746), .Y(n6747_1));
INVX1    g3052(.A(g93), .Y(n7697));
NAND3X1  g3053(.A(n4957), .B(g4358), .C(n5174), .Y(n7698));
INVX1    g1826(.A(n5506), .Y(n6466));
INVX1    g2308(.A(g6049), .Y(n6951));
INVX1    g2301(.A(g5990), .Y(n6944));
AOI21X1  g2105(.A0(n6745), .A1(n4721), .B0(n6744), .Y(n6746));
INVX1    g0541(.A(g4349), .Y(n5174));
NOR3X1   g0337(.A(n4955), .B(n4952), .C(g4311), .Y(n4957));
NOR2X1   g0866(.A(n4809), .B(g113), .Y(n5506));
INVX1    g2103(.A(g4681), .Y(n6744));
NOR3X1   g0101(.A(g4793), .B(g4801), .C(n4720), .Y(n4721));
NOR4X1   g2104(.A(g4785), .B(n4815), .C(n4814), .D(n4723), .Y(n6745));
INVX1    g0332(.A(n4951), .Y(n4952));
INVX1    g0335(.A(n4954_1), .Y(n4955));
AOI21X1  g0189(.A0(g37), .A1(g99), .B0(g134), .Y(n4809));
INVX1    g0100(.A(g4776), .Y(n4720));
NAND3X1  g0103(.A(g4659), .B(g4669), .C(g4653), .Y(n4723));
INVX1    g0194(.A(g4754), .Y(n4814));
INVX1    g0195(.A(g4709), .Y(n4815));
XOR2X1   g0331(.A(g4322), .B(n4950), .Y(n4951));
XOR2X1   g0334(.A(g4332), .B(n4953), .Y(n4954_1));
INVX1    g0330(.A(g72), .Y(n4950));
INVX1    g0333(.A(g73), .Y(n4953));

endmodule
