// Benchmark "top" written by ABC on Mon Sep 21 03:40:48 2020

module top ( 
    \in0[0] , \in0[1] , \in0[2] , \in0[3] , \in0[4] , \in0[5] , \in0[6] ,
    \in0[7] , \in0[8] , \in0[9] , \in0[10] , \in0[11] , \in0[12] ,
    \in0[13] , \in0[14] , \in0[15] , \in0[16] , \in0[17] , \in0[18] ,
    \in0[19] , \in0[20] , \in0[21] , \in0[22] , \in0[23] , \in0[24] ,
    \in0[25] , \in0[26] , \in0[27] , \in0[28] , \in0[29] , \in0[30] ,
    \in0[31] , \in0[32] , \in0[33] , \in0[34] , \in0[35] , \in0[36] ,
    \in0[37] , \in0[38] , \in0[39] , \in0[40] , \in0[41] , \in0[42] ,
    \in0[43] , \in0[44] , \in0[45] , \in0[46] , \in0[47] , \in0[48] ,
    \in0[49] , \in0[50] , \in0[51] , \in0[52] , \in0[53] , \in0[54] ,
    \in0[55] , \in0[56] , \in0[57] , \in0[58] , \in0[59] , \in0[60] ,
    \in0[61] , \in0[62] , \in0[63] , \in0[64] , \in0[65] , \in0[66] ,
    \in0[67] , \in0[68] , \in0[69] , \in0[70] , \in0[71] , \in0[72] ,
    \in0[73] , \in0[74] , \in0[75] , \in0[76] , \in0[77] , \in0[78] ,
    \in0[79] , \in0[80] , \in0[81] , \in0[82] , \in0[83] , \in0[84] ,
    \in0[85] , \in0[86] , \in0[87] , \in0[88] , \in0[89] , \in0[90] ,
    \in0[91] , \in0[92] , \in0[93] , \in0[94] , \in0[95] , \in0[96] ,
    \in0[97] , \in0[98] , \in0[99] , \in0[100] , \in0[101] , \in0[102] ,
    \in0[103] , \in0[104] , \in0[105] , \in0[106] , \in0[107] , \in0[108] ,
    \in0[109] , \in0[110] , \in0[111] , \in0[112] , \in0[113] , \in0[114] ,
    \in0[115] , \in0[116] , \in0[117] , \in0[118] , \in0[119] , \in0[120] ,
    \in0[121] , \in0[122] , \in0[123] , \in0[124] , \in0[125] , \in0[126] ,
    \in0[127] , \in1[0] , \in1[1] , \in1[2] , \in1[3] , \in1[4] , \in1[5] ,
    \in1[6] , \in1[7] , \in1[8] , \in1[9] , \in1[10] , \in1[11] ,
    \in1[12] , \in1[13] , \in1[14] , \in1[15] , \in1[16] , \in1[17] ,
    \in1[18] , \in1[19] , \in1[20] , \in1[21] , \in1[22] , \in1[23] ,
    \in1[24] , \in1[25] , \in1[26] , \in1[27] , \in1[28] , \in1[29] ,
    \in1[30] , \in1[31] , \in1[32] , \in1[33] , \in1[34] , \in1[35] ,
    \in1[36] , \in1[37] , \in1[38] , \in1[39] , \in1[40] , \in1[41] ,
    \in1[42] , \in1[43] , \in1[44] , \in1[45] , \in1[46] , \in1[47] ,
    \in1[48] , \in1[49] , \in1[50] , \in1[51] , \in1[52] , \in1[53] ,
    \in1[54] , \in1[55] , \in1[56] , \in1[57] , \in1[58] , \in1[59] ,
    \in1[60] , \in1[61] , \in1[62] , \in1[63] , \in1[64] , \in1[65] ,
    \in1[66] , \in1[67] , \in1[68] , \in1[69] , \in1[70] , \in1[71] ,
    \in1[72] , \in1[73] , \in1[74] , \in1[75] , \in1[76] , \in1[77] ,
    \in1[78] , \in1[79] , \in1[80] , \in1[81] , \in1[82] , \in1[83] ,
    \in1[84] , \in1[85] , \in1[86] , \in1[87] , \in1[88] , \in1[89] ,
    \in1[90] , \in1[91] , \in1[92] , \in1[93] , \in1[94] , \in1[95] ,
    \in1[96] , \in1[97] , \in1[98] , \in1[99] , \in1[100] , \in1[101] ,
    \in1[102] , \in1[103] , \in1[104] , \in1[105] , \in1[106] , \in1[107] ,
    \in1[108] , \in1[109] , \in1[110] , \in1[111] , \in1[112] , \in1[113] ,
    \in1[114] , \in1[115] , \in1[116] , \in1[117] , \in1[118] , \in1[119] ,
    \in1[120] , \in1[121] , \in1[122] , \in1[123] , \in1[124] , \in1[125] ,
    \in1[126] , \in1[127] , \in2[0] , \in2[1] , \in2[2] , \in2[3] ,
    \in2[4] , \in2[5] , \in2[6] , \in2[7] , \in2[8] , \in2[9] , \in2[10] ,
    \in2[11] , \in2[12] , \in2[13] , \in2[14] , \in2[15] , \in2[16] ,
    \in2[17] , \in2[18] , \in2[19] , \in2[20] , \in2[21] , \in2[22] ,
    \in2[23] , \in2[24] , \in2[25] , \in2[26] , \in2[27] , \in2[28] ,
    \in2[29] , \in2[30] , \in2[31] , \in2[32] , \in2[33] , \in2[34] ,
    \in2[35] , \in2[36] , \in2[37] , \in2[38] , \in2[39] , \in2[40] ,
    \in2[41] , \in2[42] , \in2[43] , \in2[44] , \in2[45] , \in2[46] ,
    \in2[47] , \in2[48] , \in2[49] , \in2[50] , \in2[51] , \in2[52] ,
    \in2[53] , \in2[54] , \in2[55] , \in2[56] , \in2[57] , \in2[58] ,
    \in2[59] , \in2[60] , \in2[61] , \in2[62] , \in2[63] , \in2[64] ,
    \in2[65] , \in2[66] , \in2[67] , \in2[68] , \in2[69] , \in2[70] ,
    \in2[71] , \in2[72] , \in2[73] , \in2[74] , \in2[75] , \in2[76] ,
    \in2[77] , \in2[78] , \in2[79] , \in2[80] , \in2[81] , \in2[82] ,
    \in2[83] , \in2[84] , \in2[85] , \in2[86] , \in2[87] , \in2[88] ,
    \in2[89] , \in2[90] , \in2[91] , \in2[92] , \in2[93] , \in2[94] ,
    \in2[95] , \in2[96] , \in2[97] , \in2[98] , \in2[99] , \in2[100] ,
    \in2[101] , \in2[102] , \in2[103] , \in2[104] , \in2[105] , \in2[106] ,
    \in2[107] , \in2[108] , \in2[109] , \in2[110] , \in2[111] , \in2[112] ,
    \in2[113] , \in2[114] , \in2[115] , \in2[116] , \in2[117] , \in2[118] ,
    \in2[119] , \in2[120] , \in2[121] , \in2[122] , \in2[123] , \in2[124] ,
    \in2[125] , \in2[126] , \in2[127] , \in3[0] , \in3[1] , \in3[2] ,
    \in3[3] , \in3[4] , \in3[5] , \in3[6] , \in3[7] , \in3[8] , \in3[9] ,
    \in3[10] , \in3[11] , \in3[12] , \in3[13] , \in3[14] , \in3[15] ,
    \in3[16] , \in3[17] , \in3[18] , \in3[19] , \in3[20] , \in3[21] ,
    \in3[22] , \in3[23] , \in3[24] , \in3[25] , \in3[26] , \in3[27] ,
    \in3[28] , \in3[29] , \in3[30] , \in3[31] , \in3[32] , \in3[33] ,
    \in3[34] , \in3[35] , \in3[36] , \in3[37] , \in3[38] , \in3[39] ,
    \in3[40] , \in3[41] , \in3[42] , \in3[43] , \in3[44] , \in3[45] ,
    \in3[46] , \in3[47] , \in3[48] , \in3[49] , \in3[50] , \in3[51] ,
    \in3[52] , \in3[53] , \in3[54] , \in3[55] , \in3[56] , \in3[57] ,
    \in3[58] , \in3[59] , \in3[60] , \in3[61] , \in3[62] , \in3[63] ,
    \in3[64] , \in3[65] , \in3[66] , \in3[67] , \in3[68] , \in3[69] ,
    \in3[70] , \in3[71] , \in3[72] , \in3[73] , \in3[74] , \in3[75] ,
    \in3[76] , \in3[77] , \in3[78] , \in3[79] , \in3[80] , \in3[81] ,
    \in3[82] , \in3[83] , \in3[84] , \in3[85] , \in3[86] , \in3[87] ,
    \in3[88] , \in3[89] , \in3[90] , \in3[91] , \in3[92] , \in3[93] ,
    \in3[94] , \in3[95] , \in3[96] , \in3[97] , \in3[98] , \in3[99] ,
    \in3[100] , \in3[101] , \in3[102] , \in3[103] , \in3[104] , \in3[105] ,
    \in3[106] , \in3[107] , \in3[108] , \in3[109] , \in3[110] , \in3[111] ,
    \in3[112] , \in3[113] , \in3[114] , \in3[115] , \in3[116] , \in3[117] ,
    \in3[118] , \in3[119] , \in3[120] , \in3[121] , \in3[122] , \in3[123] ,
    \in3[124] , \in3[125] , \in3[126] , \in3[127] ,
    \result[0] , \result[1] , \result[2] , \result[3] , \result[4] ,
    \result[5] , \result[6] , \result[7] , \result[8] , \result[9] ,
    \result[10] , \result[11] , \result[12] , \result[13] , \result[14] ,
    \result[15] , \result[16] , \result[17] , \result[18] , \result[19] ,
    \result[20] , \result[21] , \result[22] , \result[23] , \result[24] ,
    \result[25] , \result[26] , \result[27] , \result[28] , \result[29] ,
    \result[30] , \result[31] , \result[32] , \result[33] , \result[34] ,
    \result[35] , \result[36] , \result[37] , \result[38] , \result[39] ,
    \result[40] , \result[41] , \result[42] , \result[43] , \result[44] ,
    \result[45] , \result[46] , \result[47] , \result[48] , \result[49] ,
    \result[50] , \result[51] , \result[52] , \result[53] , \result[54] ,
    \result[55] , \result[56] , \result[57] , \result[58] , \result[59] ,
    \result[60] , \result[61] , \result[62] , \result[63] , \result[64] ,
    \result[65] , \result[66] , \result[67] , \result[68] , \result[69] ,
    \result[70] , \result[71] , \result[72] , \result[73] , \result[74] ,
    \result[75] , \result[76] , \result[77] , \result[78] , \result[79] ,
    \result[80] , \result[81] , \result[82] , \result[83] , \result[84] ,
    \result[85] , \result[86] , \result[87] , \result[88] , \result[89] ,
    \result[90] , \result[91] , \result[92] , \result[93] , \result[94] ,
    \result[95] , \result[96] , \result[97] , \result[98] , \result[99] ,
    \result[100] , \result[101] , \result[102] , \result[103] ,
    \result[104] , \result[105] , \result[106] , \result[107] ,
    \result[108] , \result[109] , \result[110] , \result[111] ,
    \result[112] , \result[113] , \result[114] , \result[115] ,
    \result[116] , \result[117] , \result[118] , \result[119] ,
    \result[120] , \result[121] , \result[122] , \result[123] ,
    \result[124] , \result[125] , \result[126] , \result[127] ,
    \address[0] , \address[1]   );
  input  \in0[0] , \in0[1] , \in0[2] , \in0[3] , \in0[4] , \in0[5] ,
    \in0[6] , \in0[7] , \in0[8] , \in0[9] , \in0[10] , \in0[11] ,
    \in0[12] , \in0[13] , \in0[14] , \in0[15] , \in0[16] , \in0[17] ,
    \in0[18] , \in0[19] , \in0[20] , \in0[21] , \in0[22] , \in0[23] ,
    \in0[24] , \in0[25] , \in0[26] , \in0[27] , \in0[28] , \in0[29] ,
    \in0[30] , \in0[31] , \in0[32] , \in0[33] , \in0[34] , \in0[35] ,
    \in0[36] , \in0[37] , \in0[38] , \in0[39] , \in0[40] , \in0[41] ,
    \in0[42] , \in0[43] , \in0[44] , \in0[45] , \in0[46] , \in0[47] ,
    \in0[48] , \in0[49] , \in0[50] , \in0[51] , \in0[52] , \in0[53] ,
    \in0[54] , \in0[55] , \in0[56] , \in0[57] , \in0[58] , \in0[59] ,
    \in0[60] , \in0[61] , \in0[62] , \in0[63] , \in0[64] , \in0[65] ,
    \in0[66] , \in0[67] , \in0[68] , \in0[69] , \in0[70] , \in0[71] ,
    \in0[72] , \in0[73] , \in0[74] , \in0[75] , \in0[76] , \in0[77] ,
    \in0[78] , \in0[79] , \in0[80] , \in0[81] , \in0[82] , \in0[83] ,
    \in0[84] , \in0[85] , \in0[86] , \in0[87] , \in0[88] , \in0[89] ,
    \in0[90] , \in0[91] , \in0[92] , \in0[93] , \in0[94] , \in0[95] ,
    \in0[96] , \in0[97] , \in0[98] , \in0[99] , \in0[100] , \in0[101] ,
    \in0[102] , \in0[103] , \in0[104] , \in0[105] , \in0[106] , \in0[107] ,
    \in0[108] , \in0[109] , \in0[110] , \in0[111] , \in0[112] , \in0[113] ,
    \in0[114] , \in0[115] , \in0[116] , \in0[117] , \in0[118] , \in0[119] ,
    \in0[120] , \in0[121] , \in0[122] , \in0[123] , \in0[124] , \in0[125] ,
    \in0[126] , \in0[127] , \in1[0] , \in1[1] , \in1[2] , \in1[3] ,
    \in1[4] , \in1[5] , \in1[6] , \in1[7] , \in1[8] , \in1[9] , \in1[10] ,
    \in1[11] , \in1[12] , \in1[13] , \in1[14] , \in1[15] , \in1[16] ,
    \in1[17] , \in1[18] , \in1[19] , \in1[20] , \in1[21] , \in1[22] ,
    \in1[23] , \in1[24] , \in1[25] , \in1[26] , \in1[27] , \in1[28] ,
    \in1[29] , \in1[30] , \in1[31] , \in1[32] , \in1[33] , \in1[34] ,
    \in1[35] , \in1[36] , \in1[37] , \in1[38] , \in1[39] , \in1[40] ,
    \in1[41] , \in1[42] , \in1[43] , \in1[44] , \in1[45] , \in1[46] ,
    \in1[47] , \in1[48] , \in1[49] , \in1[50] , \in1[51] , \in1[52] ,
    \in1[53] , \in1[54] , \in1[55] , \in1[56] , \in1[57] , \in1[58] ,
    \in1[59] , \in1[60] , \in1[61] , \in1[62] , \in1[63] , \in1[64] ,
    \in1[65] , \in1[66] , \in1[67] , \in1[68] , \in1[69] , \in1[70] ,
    \in1[71] , \in1[72] , \in1[73] , \in1[74] , \in1[75] , \in1[76] ,
    \in1[77] , \in1[78] , \in1[79] , \in1[80] , \in1[81] , \in1[82] ,
    \in1[83] , \in1[84] , \in1[85] , \in1[86] , \in1[87] , \in1[88] ,
    \in1[89] , \in1[90] , \in1[91] , \in1[92] , \in1[93] , \in1[94] ,
    \in1[95] , \in1[96] , \in1[97] , \in1[98] , \in1[99] , \in1[100] ,
    \in1[101] , \in1[102] , \in1[103] , \in1[104] , \in1[105] , \in1[106] ,
    \in1[107] , \in1[108] , \in1[109] , \in1[110] , \in1[111] , \in1[112] ,
    \in1[113] , \in1[114] , \in1[115] , \in1[116] , \in1[117] , \in1[118] ,
    \in1[119] , \in1[120] , \in1[121] , \in1[122] , \in1[123] , \in1[124] ,
    \in1[125] , \in1[126] , \in1[127] , \in2[0] , \in2[1] , \in2[2] ,
    \in2[3] , \in2[4] , \in2[5] , \in2[6] , \in2[7] , \in2[8] , \in2[9] ,
    \in2[10] , \in2[11] , \in2[12] , \in2[13] , \in2[14] , \in2[15] ,
    \in2[16] , \in2[17] , \in2[18] , \in2[19] , \in2[20] , \in2[21] ,
    \in2[22] , \in2[23] , \in2[24] , \in2[25] , \in2[26] , \in2[27] ,
    \in2[28] , \in2[29] , \in2[30] , \in2[31] , \in2[32] , \in2[33] ,
    \in2[34] , \in2[35] , \in2[36] , \in2[37] , \in2[38] , \in2[39] ,
    \in2[40] , \in2[41] , \in2[42] , \in2[43] , \in2[44] , \in2[45] ,
    \in2[46] , \in2[47] , \in2[48] , \in2[49] , \in2[50] , \in2[51] ,
    \in2[52] , \in2[53] , \in2[54] , \in2[55] , \in2[56] , \in2[57] ,
    \in2[58] , \in2[59] , \in2[60] , \in2[61] , \in2[62] , \in2[63] ,
    \in2[64] , \in2[65] , \in2[66] , \in2[67] , \in2[68] , \in2[69] ,
    \in2[70] , \in2[71] , \in2[72] , \in2[73] , \in2[74] , \in2[75] ,
    \in2[76] , \in2[77] , \in2[78] , \in2[79] , \in2[80] , \in2[81] ,
    \in2[82] , \in2[83] , \in2[84] , \in2[85] , \in2[86] , \in2[87] ,
    \in2[88] , \in2[89] , \in2[90] , \in2[91] , \in2[92] , \in2[93] ,
    \in2[94] , \in2[95] , \in2[96] , \in2[97] , \in2[98] , \in2[99] ,
    \in2[100] , \in2[101] , \in2[102] , \in2[103] , \in2[104] , \in2[105] ,
    \in2[106] , \in2[107] , \in2[108] , \in2[109] , \in2[110] , \in2[111] ,
    \in2[112] , \in2[113] , \in2[114] , \in2[115] , \in2[116] , \in2[117] ,
    \in2[118] , \in2[119] , \in2[120] , \in2[121] , \in2[122] , \in2[123] ,
    \in2[124] , \in2[125] , \in2[126] , \in2[127] , \in3[0] , \in3[1] ,
    \in3[2] , \in3[3] , \in3[4] , \in3[5] , \in3[6] , \in3[7] , \in3[8] ,
    \in3[9] , \in3[10] , \in3[11] , \in3[12] , \in3[13] , \in3[14] ,
    \in3[15] , \in3[16] , \in3[17] , \in3[18] , \in3[19] , \in3[20] ,
    \in3[21] , \in3[22] , \in3[23] , \in3[24] , \in3[25] , \in3[26] ,
    \in3[27] , \in3[28] , \in3[29] , \in3[30] , \in3[31] , \in3[32] ,
    \in3[33] , \in3[34] , \in3[35] , \in3[36] , \in3[37] , \in3[38] ,
    \in3[39] , \in3[40] , \in3[41] , \in3[42] , \in3[43] , \in3[44] ,
    \in3[45] , \in3[46] , \in3[47] , \in3[48] , \in3[49] , \in3[50] ,
    \in3[51] , \in3[52] , \in3[53] , \in3[54] , \in3[55] , \in3[56] ,
    \in3[57] , \in3[58] , \in3[59] , \in3[60] , \in3[61] , \in3[62] ,
    \in3[63] , \in3[64] , \in3[65] , \in3[66] , \in3[67] , \in3[68] ,
    \in3[69] , \in3[70] , \in3[71] , \in3[72] , \in3[73] , \in3[74] ,
    \in3[75] , \in3[76] , \in3[77] , \in3[78] , \in3[79] , \in3[80] ,
    \in3[81] , \in3[82] , \in3[83] , \in3[84] , \in3[85] , \in3[86] ,
    \in3[87] , \in3[88] , \in3[89] , \in3[90] , \in3[91] , \in3[92] ,
    \in3[93] , \in3[94] , \in3[95] , \in3[96] , \in3[97] , \in3[98] ,
    \in3[99] , \in3[100] , \in3[101] , \in3[102] , \in3[103] , \in3[104] ,
    \in3[105] , \in3[106] , \in3[107] , \in3[108] , \in3[109] , \in3[110] ,
    \in3[111] , \in3[112] , \in3[113] , \in3[114] , \in3[115] , \in3[116] ,
    \in3[117] , \in3[118] , \in3[119] , \in3[120] , \in3[121] , \in3[122] ,
    \in3[123] , \in3[124] , \in3[125] , \in3[126] , \in3[127] ;
  output \result[0] , \result[1] , \result[2] , \result[3] , \result[4] ,
    \result[5] , \result[6] , \result[7] , \result[8] , \result[9] ,
    \result[10] , \result[11] , \result[12] , \result[13] , \result[14] ,
    \result[15] , \result[16] , \result[17] , \result[18] , \result[19] ,
    \result[20] , \result[21] , \result[22] , \result[23] , \result[24] ,
    \result[25] , \result[26] , \result[27] , \result[28] , \result[29] ,
    \result[30] , \result[31] , \result[32] , \result[33] , \result[34] ,
    \result[35] , \result[36] , \result[37] , \result[38] , \result[39] ,
    \result[40] , \result[41] , \result[42] , \result[43] , \result[44] ,
    \result[45] , \result[46] , \result[47] , \result[48] , \result[49] ,
    \result[50] , \result[51] , \result[52] , \result[53] , \result[54] ,
    \result[55] , \result[56] , \result[57] , \result[58] , \result[59] ,
    \result[60] , \result[61] , \result[62] , \result[63] , \result[64] ,
    \result[65] , \result[66] , \result[67] , \result[68] , \result[69] ,
    \result[70] , \result[71] , \result[72] , \result[73] , \result[74] ,
    \result[75] , \result[76] , \result[77] , \result[78] , \result[79] ,
    \result[80] , \result[81] , \result[82] , \result[83] , \result[84] ,
    \result[85] , \result[86] , \result[87] , \result[88] , \result[89] ,
    \result[90] , \result[91] , \result[92] , \result[93] , \result[94] ,
    \result[95] , \result[96] , \result[97] , \result[98] , \result[99] ,
    \result[100] , \result[101] , \result[102] , \result[103] ,
    \result[104] , \result[105] , \result[106] , \result[107] ,
    \result[108] , \result[109] , \result[110] , \result[111] ,
    \result[112] , \result[113] , \result[114] , \result[115] ,
    \result[116] , \result[117] , \result[118] , \result[119] ,
    \result[120] , \result[121] , \result[122] , \result[123] ,
    \result[124] , \result[125] , \result[126] , \result[127] ,
    \address[0] , \address[1] ;
  wire new_n643_, new_n644_, new_n645_, new_n646_, new_n647_, new_n648_,
    new_n649_, new_n650_, new_n651_, new_n652_, new_n653_, new_n654_,
    new_n655_, new_n656_, new_n657_, new_n658_, new_n659_, new_n660_,
    new_n661_, new_n662_, new_n663_, new_n664_, new_n665_, new_n666_,
    new_n667_, new_n668_, new_n669_, new_n670_, new_n671_, new_n672_,
    new_n673_, new_n674_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n687_, new_n688_, new_n689_, new_n690_,
    new_n691_, new_n692_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n817_, new_n818_, new_n819_, new_n820_, new_n821_, new_n822_,
    new_n823_, new_n824_, new_n825_, new_n826_, new_n827_, new_n828_,
    new_n829_, new_n830_, new_n831_, new_n832_, new_n833_, new_n834_,
    new_n835_, new_n836_, new_n837_, new_n838_, new_n839_, new_n840_,
    new_n841_, new_n842_, new_n843_, new_n844_, new_n845_, new_n846_,
    new_n847_, new_n848_, new_n849_, new_n850_, new_n851_, new_n852_,
    new_n853_, new_n854_, new_n855_, new_n856_, new_n857_, new_n858_,
    new_n859_, new_n860_, new_n861_, new_n862_, new_n863_, new_n864_,
    new_n865_, new_n866_, new_n867_, new_n868_, new_n869_, new_n870_,
    new_n871_, new_n872_, new_n873_, new_n874_, new_n875_, new_n876_,
    new_n877_, new_n878_, new_n879_, new_n880_, new_n881_, new_n882_,
    new_n883_, new_n884_, new_n885_, new_n886_, new_n887_, new_n888_,
    new_n889_, new_n890_, new_n891_, new_n892_, new_n893_, new_n894_,
    new_n895_, new_n896_, new_n897_, new_n898_, new_n899_, new_n900_,
    new_n901_, new_n902_, new_n903_, new_n904_, new_n905_, new_n906_,
    new_n907_, new_n908_, new_n909_, new_n910_, new_n911_, new_n912_,
    new_n913_, new_n914_, new_n915_, new_n916_, new_n917_, new_n918_,
    new_n919_, new_n920_, new_n921_, new_n922_, new_n923_, new_n924_,
    new_n925_, new_n926_, new_n927_, new_n928_, new_n929_, new_n930_,
    new_n931_, new_n932_, new_n933_, new_n934_, new_n935_, new_n936_,
    new_n937_, new_n938_, new_n939_, new_n940_, new_n941_, new_n942_,
    new_n943_, new_n944_, new_n945_, new_n946_, new_n947_, new_n948_,
    new_n949_, new_n950_, new_n951_, new_n952_, new_n953_, new_n954_,
    new_n955_, new_n956_, new_n957_, new_n958_, new_n959_, new_n960_,
    new_n961_, new_n962_, new_n963_, new_n964_, new_n965_, new_n966_,
    new_n967_, new_n968_, new_n969_, new_n970_, new_n971_, new_n972_,
    new_n973_, new_n974_, new_n975_, new_n976_, new_n977_, new_n978_,
    new_n979_, new_n980_, new_n981_, new_n982_, new_n983_, new_n984_,
    new_n985_, new_n986_, new_n987_, new_n988_, new_n989_, new_n990_,
    new_n991_, new_n992_, new_n993_, new_n994_, new_n995_, new_n996_,
    new_n997_, new_n998_, new_n999_, new_n1000_, new_n1001_, new_n1002_,
    new_n1003_, new_n1004_, new_n1005_, new_n1006_, new_n1007_, new_n1008_,
    new_n1009_, new_n1010_, new_n1011_, new_n1012_, new_n1013_, new_n1014_,
    new_n1015_, new_n1016_, new_n1017_, new_n1018_, new_n1019_, new_n1020_,
    new_n1021_, new_n1022_, new_n1023_, new_n1024_, new_n1025_, new_n1026_,
    new_n1027_, new_n1028_, new_n1029_, new_n1030_, new_n1031_, new_n1032_,
    new_n1033_, new_n1034_, new_n1035_, new_n1036_, new_n1037_, new_n1038_,
    new_n1039_, new_n1040_, new_n1041_, new_n1042_, new_n1043_, new_n1044_,
    new_n1045_, new_n1046_, new_n1047_, new_n1048_, new_n1049_, new_n1050_,
    new_n1051_, new_n1052_, new_n1053_, new_n1054_, new_n1055_, new_n1056_,
    new_n1057_, new_n1058_, new_n1059_, new_n1060_, new_n1061_, new_n1062_,
    new_n1063_, new_n1064_, new_n1065_, new_n1066_, new_n1067_, new_n1068_,
    new_n1069_, new_n1070_, new_n1071_, new_n1072_, new_n1073_, new_n1074_,
    new_n1075_, new_n1076_, new_n1077_, new_n1078_, new_n1079_, new_n1080_,
    new_n1081_, new_n1082_, new_n1083_, new_n1084_, new_n1085_, new_n1086_,
    new_n1087_, new_n1088_, new_n1089_, new_n1090_, new_n1091_, new_n1092_,
    new_n1093_, new_n1094_, new_n1095_, new_n1096_, new_n1097_, new_n1098_,
    new_n1099_, new_n1100_, new_n1101_, new_n1102_, new_n1103_, new_n1104_,
    new_n1105_, new_n1106_, new_n1107_, new_n1108_, new_n1109_, new_n1110_,
    new_n1111_, new_n1112_, new_n1113_, new_n1114_, new_n1115_, new_n1116_,
    new_n1117_, new_n1118_, new_n1119_, new_n1120_, new_n1121_, new_n1122_,
    new_n1123_, new_n1124_, new_n1125_, new_n1126_, new_n1127_, new_n1128_,
    new_n1129_, new_n1130_, new_n1131_, new_n1132_, new_n1133_, new_n1134_,
    new_n1135_, new_n1136_, new_n1137_, new_n1138_, new_n1139_, new_n1140_,
    new_n1141_, new_n1142_, new_n1143_, new_n1144_, new_n1145_, new_n1146_,
    new_n1147_, new_n1148_, new_n1149_, new_n1150_, new_n1151_, new_n1152_,
    new_n1153_, new_n1154_, new_n1155_, new_n1156_, new_n1157_, new_n1158_,
    new_n1159_, new_n1160_, new_n1161_, new_n1162_, new_n1163_, new_n1164_,
    new_n1165_, new_n1166_, new_n1167_, new_n1168_, new_n1169_, new_n1170_,
    new_n1171_, new_n1172_, new_n1173_, new_n1174_, new_n1175_, new_n1176_,
    new_n1177_, new_n1178_, new_n1179_, new_n1180_, new_n1181_, new_n1182_,
    new_n1183_, new_n1184_, new_n1185_, new_n1186_, new_n1187_, new_n1188_,
    new_n1189_, new_n1190_, new_n1191_, new_n1192_, new_n1193_, new_n1194_,
    new_n1195_, new_n1196_, new_n1197_, new_n1198_, new_n1199_, new_n1200_,
    new_n1201_, new_n1202_, new_n1203_, new_n1204_, new_n1205_, new_n1206_,
    new_n1207_, new_n1208_, new_n1209_, new_n1210_, new_n1211_, new_n1212_,
    new_n1213_, new_n1214_, new_n1215_, new_n1216_, new_n1217_, new_n1218_,
    new_n1219_, new_n1220_, new_n1221_, new_n1222_, new_n1223_, new_n1224_,
    new_n1225_, new_n1226_, new_n1227_, new_n1228_, new_n1229_, new_n1230_,
    new_n1231_, new_n1232_, new_n1233_, new_n1234_, new_n1235_, new_n1236_,
    new_n1237_, new_n1238_, new_n1239_, new_n1240_, new_n1241_, new_n1242_,
    new_n1243_, new_n1244_, new_n1245_, new_n1246_, new_n1247_, new_n1248_,
    new_n1249_, new_n1250_, new_n1251_, new_n1252_, new_n1253_, new_n1254_,
    new_n1255_, new_n1256_, new_n1257_, new_n1258_, new_n1259_, new_n1260_,
    new_n1261_, new_n1262_, new_n1263_, new_n1264_, new_n1265_, new_n1266_,
    new_n1267_, new_n1268_, new_n1269_, new_n1270_, new_n1271_, new_n1272_,
    new_n1273_, new_n1274_, new_n1275_, new_n1276_, new_n1277_, new_n1278_,
    new_n1279_, new_n1280_, new_n1281_, new_n1282_, new_n1283_, new_n1284_,
    new_n1285_, new_n1286_, new_n1287_, new_n1288_, new_n1289_, new_n1290_,
    new_n1291_, new_n1292_, new_n1293_, new_n1294_, new_n1295_, new_n1296_,
    new_n1297_, new_n1298_, new_n1299_, new_n1300_, new_n1301_, new_n1302_,
    new_n1303_, new_n1304_, new_n1305_, new_n1306_, new_n1307_, new_n1308_,
    new_n1309_, new_n1310_, new_n1311_, new_n1312_, new_n1313_, new_n1314_,
    new_n1315_, new_n1316_, new_n1317_, new_n1318_, new_n1319_, new_n1320_,
    new_n1321_, new_n1322_, new_n1323_, new_n1324_, new_n1325_, new_n1326_,
    new_n1327_, new_n1328_, new_n1329_, new_n1330_, new_n1331_, new_n1332_,
    new_n1333_, new_n1334_, new_n1335_, new_n1336_, new_n1337_, new_n1338_,
    new_n1339_, new_n1340_, new_n1341_, new_n1342_, new_n1343_, new_n1344_,
    new_n1345_, new_n1346_, new_n1347_, new_n1348_, new_n1349_, new_n1350_,
    new_n1351_, new_n1352_, new_n1353_, new_n1354_, new_n1355_, new_n1356_,
    new_n1357_, new_n1358_, new_n1359_, new_n1360_, new_n1361_, new_n1362_,
    new_n1363_, new_n1364_, new_n1365_, new_n1366_, new_n1367_, new_n1368_,
    new_n1369_, new_n1370_, new_n1371_, new_n1372_, new_n1373_, new_n1374_,
    new_n1375_, new_n1376_, new_n1377_, new_n1378_, new_n1379_, new_n1380_,
    new_n1381_, new_n1382_, new_n1383_, new_n1384_, new_n1385_, new_n1386_,
    new_n1387_, new_n1388_, new_n1389_, new_n1390_, new_n1391_, new_n1392_,
    new_n1393_, new_n1394_, new_n1395_, new_n1396_, new_n1397_, new_n1398_,
    new_n1399_, new_n1400_, new_n1401_, new_n1402_, new_n1403_, new_n1404_,
    new_n1405_, new_n1406_, new_n1407_, new_n1408_, new_n1409_, new_n1410_,
    new_n1411_, new_n1412_, new_n1413_, new_n1414_, new_n1415_, new_n1416_,
    new_n1417_, new_n1418_, new_n1419_, new_n1420_, new_n1421_, new_n1422_,
    new_n1423_, new_n1424_, new_n1425_, new_n1426_, new_n1427_, new_n1428_,
    new_n1429_, new_n1430_, new_n1431_, new_n1432_, new_n1433_, new_n1434_,
    new_n1435_, new_n1436_, new_n1437_, new_n1438_, new_n1439_, new_n1440_,
    new_n1441_, new_n1442_, new_n1443_, new_n1444_, new_n1445_, new_n1446_,
    new_n1447_, new_n1448_, new_n1449_, new_n1450_, new_n1451_, new_n1452_,
    new_n1453_, new_n1454_, new_n1455_, new_n1456_, new_n1457_, new_n1458_,
    new_n1459_, new_n1460_, new_n1461_, new_n1462_, new_n1463_, new_n1464_,
    new_n1465_, new_n1466_, new_n1467_, new_n1468_, new_n1469_, new_n1470_,
    new_n1471_, new_n1472_, new_n1473_, new_n1474_, new_n1475_, new_n1476_,
    new_n1477_, new_n1478_, new_n1479_, new_n1480_, new_n1481_, new_n1482_,
    new_n1483_, new_n1484_, new_n1485_, new_n1486_, new_n1487_, new_n1488_,
    new_n1489_, new_n1490_, new_n1491_, new_n1492_, new_n1493_, new_n1494_,
    new_n1495_, new_n1496_, new_n1497_, new_n1498_, new_n1499_, new_n1500_,
    new_n1501_, new_n1502_, new_n1503_, new_n1504_, new_n1505_, new_n1506_,
    new_n1507_, new_n1508_, new_n1509_, new_n1510_, new_n1511_, new_n1512_,
    new_n1513_, new_n1514_, new_n1515_, new_n1516_, new_n1517_, new_n1518_,
    new_n1519_, new_n1520_, new_n1521_, new_n1522_, new_n1523_, new_n1524_,
    new_n1525_, new_n1526_, new_n1527_, new_n1528_, new_n1529_, new_n1530_,
    new_n1531_, new_n1532_, new_n1533_, new_n1534_, new_n1535_, new_n1536_,
    new_n1537_, new_n1538_, new_n1539_, new_n1540_, new_n1541_, new_n1542_,
    new_n1543_, new_n1544_, new_n1545_, new_n1546_, new_n1547_, new_n1548_,
    new_n1549_, new_n1550_, new_n1551_, new_n1552_, new_n1553_, new_n1554_,
    new_n1555_, new_n1556_, new_n1557_, new_n1558_, new_n1559_, new_n1560_,
    new_n1561_, new_n1562_, new_n1563_, new_n1564_, new_n1565_, new_n1566_,
    new_n1567_, new_n1568_, new_n1569_, new_n1570_, new_n1571_, new_n1572_,
    new_n1573_, new_n1574_, new_n1575_, new_n1576_, new_n1577_, new_n1578_,
    new_n1579_, new_n1580_, new_n1581_, new_n1582_, new_n1583_, new_n1584_,
    new_n1585_, new_n1586_, new_n1587_, new_n1588_, new_n1589_, new_n1590_,
    new_n1591_, new_n1592_, new_n1593_, new_n1594_, new_n1595_, new_n1596_,
    new_n1597_, new_n1598_, new_n1599_, new_n1600_, new_n1601_, new_n1602_,
    new_n1603_, new_n1604_, new_n1605_, new_n1606_, new_n1607_, new_n1608_,
    new_n1609_, new_n1610_, new_n1611_, new_n1612_, new_n1613_, new_n1614_,
    new_n1615_, new_n1616_, new_n1617_, new_n1618_, new_n1619_, new_n1620_,
    new_n1621_, new_n1622_, new_n1623_, new_n1624_, new_n1625_, new_n1626_,
    new_n1627_, new_n1628_, new_n1629_, new_n1630_, new_n1631_, new_n1632_,
    new_n1633_, new_n1634_, new_n1635_, new_n1636_, new_n1637_, new_n1638_,
    new_n1639_, new_n1640_, new_n1641_, new_n1642_, new_n1643_, new_n1644_,
    new_n1645_, new_n1646_, new_n1647_, new_n1648_, new_n1649_, new_n1650_,
    new_n1651_, new_n1652_, new_n1653_, new_n1654_, new_n1655_, new_n1656_,
    new_n1657_, new_n1658_, new_n1659_, new_n1660_, new_n1661_, new_n1662_,
    new_n1663_, new_n1664_, new_n1665_, new_n1666_, new_n1667_, new_n1668_,
    new_n1669_, new_n1670_, new_n1671_, new_n1672_, new_n1673_, new_n1674_,
    new_n1675_, new_n1676_, new_n1677_, new_n1678_, new_n1679_, new_n1680_,
    new_n1681_, new_n1682_, new_n1683_, new_n1684_, new_n1685_, new_n1686_,
    new_n1687_, new_n1688_, new_n1689_, new_n1690_, new_n1691_, new_n1692_,
    new_n1693_, new_n1694_, new_n1695_, new_n1696_, new_n1697_, new_n1698_,
    new_n1699_, new_n1700_, new_n1701_, new_n1702_, new_n1703_, new_n1704_,
    new_n1705_, new_n1706_, new_n1707_, new_n1708_, new_n1709_, new_n1710_,
    new_n1711_, new_n1712_, new_n1713_, new_n1714_, new_n1715_, new_n1716_,
    new_n1717_, new_n1718_, new_n1719_, new_n1720_, new_n1721_, new_n1722_,
    new_n1723_, new_n1724_, new_n1725_, new_n1726_, new_n1727_, new_n1728_,
    new_n1729_, new_n1730_, new_n1731_, new_n1732_, new_n1733_, new_n1734_,
    new_n1735_, new_n1736_, new_n1737_, new_n1738_, new_n1739_, new_n1740_,
    new_n1741_, new_n1742_, new_n1743_, new_n1744_, new_n1745_, new_n1746_,
    new_n1747_, new_n1748_, new_n1749_, new_n1750_, new_n1751_, new_n1752_,
    new_n1753_, new_n1754_, new_n1755_, new_n1756_, new_n1757_, new_n1758_,
    new_n1759_, new_n1760_, new_n1761_, new_n1762_, new_n1763_, new_n1764_,
    new_n1765_, new_n1766_, new_n1767_, new_n1768_, new_n1769_, new_n1770_,
    new_n1771_, new_n1772_, new_n1773_, new_n1774_, new_n1775_, new_n1776_,
    new_n1777_, new_n1778_, new_n1779_, new_n1780_, new_n1781_, new_n1782_,
    new_n1783_, new_n1784_, new_n1785_, new_n1786_, new_n1787_, new_n1788_,
    new_n1789_, new_n1790_, new_n1791_, new_n1792_, new_n1793_, new_n1794_,
    new_n1795_, new_n1796_, new_n1797_, new_n1798_, new_n1799_, new_n1800_,
    new_n1801_, new_n1802_, new_n1803_, new_n1804_, new_n1805_, new_n1806_,
    new_n1807_, new_n1808_, new_n1809_, new_n1810_, new_n1811_, new_n1812_,
    new_n1813_, new_n1814_, new_n1815_, new_n1816_, new_n1817_, new_n1818_,
    new_n1819_, new_n1820_, new_n1821_, new_n1822_, new_n1823_, new_n1824_,
    new_n1825_, new_n1826_, new_n1827_, new_n1828_, new_n1829_, new_n1830_,
    new_n1831_, new_n1832_, new_n1833_, new_n1834_, new_n1835_, new_n1836_,
    new_n1837_, new_n1838_, new_n1839_, new_n1840_, new_n1841_, new_n1842_,
    new_n1843_, new_n1844_, new_n1845_, new_n1846_, new_n1847_, new_n1848_,
    new_n1849_, new_n1850_, new_n1851_, new_n1852_, new_n1853_, new_n1854_,
    new_n1855_, new_n1856_, new_n1857_, new_n1858_, new_n1859_, new_n1860_,
    new_n1861_, new_n1862_, new_n1863_, new_n1864_, new_n1865_, new_n1866_,
    new_n1867_, new_n1868_, new_n1869_, new_n1870_, new_n1871_, new_n1872_,
    new_n1873_, new_n1874_, new_n1875_, new_n1876_, new_n1877_, new_n1878_,
    new_n1879_, new_n1880_, new_n1881_, new_n1882_, new_n1883_, new_n1884_,
    new_n1885_, new_n1886_, new_n1887_, new_n1888_, new_n1889_, new_n1890_,
    new_n1891_, new_n1892_, new_n1893_, new_n1894_, new_n1895_, new_n1896_,
    new_n1897_, new_n1898_, new_n1899_, new_n1900_, new_n1901_, new_n1902_,
    new_n1903_, new_n1904_, new_n1905_, new_n1906_, new_n1907_, new_n1908_,
    new_n1909_, new_n1910_, new_n1911_, new_n1912_, new_n1913_, new_n1914_,
    new_n1915_, new_n1916_, new_n1917_, new_n1918_, new_n1919_, new_n1920_,
    new_n1921_, new_n1922_, new_n1923_, new_n1924_, new_n1925_, new_n1926_,
    new_n1927_, new_n1928_, new_n1929_, new_n1930_, new_n1931_, new_n1932_,
    new_n1933_, new_n1934_, new_n1935_, new_n1936_, new_n1937_, new_n1938_,
    new_n1939_, new_n1940_, new_n1941_, new_n1942_, new_n1943_, new_n1944_,
    new_n1945_, new_n1946_, new_n1947_, new_n1948_, new_n1949_, new_n1950_,
    new_n1951_, new_n1952_, new_n1953_, new_n1954_, new_n1955_, new_n1956_,
    new_n1957_, new_n1958_, new_n1959_, new_n1960_, new_n1961_, new_n1962_,
    new_n1963_, new_n1964_, new_n1965_, new_n1966_, new_n1967_, new_n1968_,
    new_n1969_, new_n1970_, new_n1971_, new_n1972_, new_n1973_, new_n1974_,
    new_n1975_, new_n1976_, new_n1977_, new_n1978_, new_n1979_, new_n1980_,
    new_n1981_, new_n1982_, new_n1983_, new_n1984_, new_n1985_, new_n1986_,
    new_n1987_, new_n1988_, new_n1989_, new_n1990_, new_n1991_, new_n1992_,
    new_n1993_, new_n1994_, new_n1995_, new_n1996_, new_n1997_, new_n1998_,
    new_n1999_, new_n2000_, new_n2001_, new_n2002_, new_n2003_, new_n2004_,
    new_n2005_, new_n2006_, new_n2007_, new_n2008_, new_n2009_, new_n2010_,
    new_n2011_, new_n2012_, new_n2013_, new_n2014_, new_n2015_, new_n2016_,
    new_n2017_, new_n2018_, new_n2019_, new_n2020_, new_n2021_, new_n2022_,
    new_n2023_, new_n2024_, new_n2025_, new_n2026_, new_n2027_, new_n2028_,
    new_n2029_, new_n2030_, new_n2031_, new_n2032_, new_n2033_, new_n2034_,
    new_n2035_, new_n2036_, new_n2037_, new_n2038_, new_n2039_, new_n2040_,
    new_n2041_, new_n2042_, new_n2043_, new_n2044_, new_n2045_, new_n2046_,
    new_n2047_, new_n2048_, new_n2049_, new_n2050_, new_n2051_, new_n2052_,
    new_n2053_, new_n2054_, new_n2055_, new_n2056_, new_n2057_, new_n2058_,
    new_n2059_, new_n2060_, new_n2061_, new_n2062_, new_n2063_, new_n2064_,
    new_n2065_, new_n2066_, new_n2067_, new_n2068_, new_n2069_, new_n2070_,
    new_n2071_, new_n2072_, new_n2073_, new_n2074_, new_n2075_, new_n2076_,
    new_n2077_, new_n2078_, new_n2079_, new_n2080_, new_n2081_, new_n2082_,
    new_n2083_, new_n2084_, new_n2085_, new_n2086_, new_n2087_, new_n2088_,
    new_n2089_, new_n2090_, new_n2091_, new_n2092_, new_n2093_, new_n2094_,
    new_n2095_, new_n2096_, new_n2097_, new_n2098_, new_n2099_, new_n2100_,
    new_n2101_, new_n2102_, new_n2103_, new_n2104_, new_n2105_, new_n2106_,
    new_n2107_, new_n2108_, new_n2109_, new_n2110_, new_n2111_, new_n2112_,
    new_n2113_, new_n2114_, new_n2115_, new_n2116_, new_n2117_, new_n2118_,
    new_n2119_, new_n2120_, new_n2121_, new_n2122_, new_n2123_, new_n2124_,
    new_n2125_, new_n2126_, new_n2127_, new_n2128_, new_n2129_, new_n2130_,
    new_n2131_, new_n2132_, new_n2133_, new_n2134_, new_n2135_, new_n2136_,
    new_n2137_, new_n2138_, new_n2139_, new_n2140_, new_n2141_, new_n2142_,
    new_n2143_, new_n2144_, new_n2145_, new_n2146_, new_n2147_, new_n2148_,
    new_n2149_, new_n2150_, new_n2151_, new_n2152_, new_n2153_, new_n2154_,
    new_n2155_, new_n2156_, new_n2157_, new_n2158_, new_n2159_, new_n2160_,
    new_n2161_, new_n2162_, new_n2163_, new_n2164_, new_n2165_, new_n2166_,
    new_n2167_, new_n2168_, new_n2169_, new_n2170_, new_n2171_, new_n2172_,
    new_n2173_, new_n2174_, new_n2175_, new_n2176_, new_n2177_, new_n2178_,
    new_n2179_, new_n2180_, new_n2181_, new_n2182_, new_n2183_, new_n2184_,
    new_n2185_, new_n2186_, new_n2187_, new_n2188_, new_n2189_, new_n2190_,
    new_n2191_, new_n2192_, new_n2193_, new_n2194_, new_n2195_, new_n2196_,
    new_n2197_, new_n2198_, new_n2199_, new_n2200_, new_n2201_, new_n2202_,
    new_n2203_, new_n2204_, new_n2205_, new_n2206_, new_n2207_, new_n2208_,
    new_n2209_, new_n2210_, new_n2211_, new_n2212_, new_n2213_, new_n2214_,
    new_n2215_, new_n2216_, new_n2217_, new_n2218_, new_n2219_, new_n2220_,
    new_n2221_, new_n2222_, new_n2223_, new_n2224_, new_n2225_, new_n2226_,
    new_n2227_, new_n2228_, new_n2229_, new_n2230_, new_n2231_, new_n2232_,
    new_n2233_, new_n2234_, new_n2235_, new_n2236_, new_n2237_, new_n2238_,
    new_n2239_, new_n2240_, new_n2241_, new_n2242_, new_n2243_, new_n2244_,
    new_n2245_, new_n2246_, new_n2247_, new_n2248_, new_n2249_, new_n2250_,
    new_n2251_, new_n2252_, new_n2253_, new_n2254_, new_n2255_, new_n2256_,
    new_n2257_, new_n2258_, new_n2259_, new_n2260_, new_n2261_, new_n2262_,
    new_n2263_, new_n2264_, new_n2265_, new_n2266_, new_n2267_, new_n2268_,
    new_n2269_, new_n2270_, new_n2271_, new_n2272_, new_n2273_, new_n2274_,
    new_n2275_, new_n2276_, new_n2277_, new_n2278_, new_n2279_, new_n2280_,
    new_n2281_, new_n2282_, new_n2283_, new_n2284_, new_n2285_, new_n2286_,
    new_n2287_, new_n2288_, new_n2289_, new_n2290_, new_n2291_, new_n2292_,
    new_n2293_, new_n2294_, new_n2295_, new_n2296_, new_n2297_, new_n2298_,
    new_n2299_, new_n2300_, new_n2301_, new_n2302_, new_n2303_, new_n2304_,
    new_n2305_, new_n2306_, new_n2307_, new_n2308_, new_n2309_, new_n2310_,
    new_n2311_, new_n2312_, new_n2313_, new_n2314_, new_n2315_, new_n2316_,
    new_n2317_, new_n2318_, new_n2319_, new_n2320_, new_n2321_, new_n2322_,
    new_n2323_, new_n2324_, new_n2325_, new_n2326_, new_n2327_, new_n2328_,
    new_n2329_, new_n2330_, new_n2331_, new_n2332_, new_n2333_, new_n2334_,
    new_n2335_, new_n2336_, new_n2337_, new_n2338_, new_n2339_, new_n2340_,
    new_n2341_, new_n2342_, new_n2343_, new_n2344_, new_n2345_, new_n2346_,
    new_n2347_, new_n2348_, new_n2349_, new_n2350_, new_n2351_, new_n2352_,
    new_n2353_, new_n2354_, new_n2355_, new_n2356_, new_n2357_, new_n2358_,
    new_n2359_, new_n2360_, new_n2361_, new_n2362_, new_n2363_, new_n2364_,
    new_n2365_, new_n2366_, new_n2367_, new_n2368_, new_n2369_, new_n2370_,
    new_n2371_, new_n2372_, new_n2373_, new_n2374_, new_n2375_, new_n2376_,
    new_n2377_, new_n2378_, new_n2379_, new_n2380_, new_n2381_, new_n2382_,
    new_n2383_, new_n2384_, new_n2385_, new_n2386_, new_n2387_, new_n2388_,
    new_n2389_, new_n2390_, new_n2391_, new_n2392_, new_n2393_, new_n2394_,
    new_n2395_, new_n2396_, new_n2397_, new_n2398_, new_n2399_, new_n2400_,
    new_n2401_, new_n2402_, new_n2403_, new_n2404_, new_n2405_, new_n2406_,
    new_n2407_, new_n2408_, new_n2409_, new_n2410_, new_n2411_, new_n2412_,
    new_n2413_, new_n2414_, new_n2415_, new_n2416_, new_n2417_, new_n2418_,
    new_n2419_, new_n2420_, new_n2421_, new_n2422_, new_n2423_, new_n2424_,
    new_n2425_, new_n2426_, new_n2427_, new_n2428_, new_n2429_, new_n2430_,
    new_n2431_, new_n2432_, new_n2433_, new_n2434_, new_n2435_, new_n2436_,
    new_n2437_, new_n2438_, new_n2439_, new_n2440_, new_n2441_, new_n2442_,
    new_n2443_, new_n2444_, new_n2445_, new_n2446_, new_n2447_, new_n2448_,
    new_n2449_, new_n2450_, new_n2451_, new_n2452_, new_n2453_, new_n2454_,
    new_n2455_, new_n2456_, new_n2457_, new_n2458_, new_n2459_, new_n2460_,
    new_n2461_, new_n2462_, new_n2463_, new_n2464_, new_n2465_, new_n2466_,
    new_n2467_, new_n2468_, new_n2469_, new_n2470_, new_n2471_, new_n2472_,
    new_n2473_, new_n2474_, new_n2475_, new_n2476_, new_n2477_, new_n2478_,
    new_n2479_, new_n2480_, new_n2481_, new_n2482_, new_n2483_, new_n2484_,
    new_n2485_, new_n2486_, new_n2487_, new_n2488_, new_n2489_, new_n2490_,
    new_n2491_, new_n2492_, new_n2493_, new_n2494_, new_n2495_, new_n2496_,
    new_n2497_, new_n2498_, new_n2499_, new_n2500_, new_n2501_, new_n2502_,
    new_n2503_, new_n2504_, new_n2505_, new_n2506_, new_n2507_, new_n2508_,
    new_n2509_, new_n2510_, new_n2511_, new_n2512_, new_n2513_, new_n2514_,
    new_n2515_, new_n2516_, new_n2517_, new_n2518_, new_n2519_, new_n2520_,
    new_n2521_, new_n2522_, new_n2523_, new_n2524_, new_n2525_, new_n2526_,
    new_n2527_, new_n2528_, new_n2529_, new_n2530_, new_n2531_, new_n2532_,
    new_n2533_, new_n2534_, new_n2535_, new_n2536_, new_n2537_, new_n2538_,
    new_n2539_, new_n2540_, new_n2541_, new_n2542_, new_n2543_, new_n2544_,
    new_n2545_, new_n2546_, new_n2547_, new_n2548_, new_n2549_, new_n2550_,
    new_n2551_, new_n2552_, new_n2553_, new_n2554_, new_n2555_, new_n2556_,
    new_n2557_, new_n2558_, new_n2559_, new_n2560_, new_n2561_, new_n2562_,
    new_n2563_, new_n2564_, new_n2565_, new_n2566_, new_n2567_, new_n2568_,
    new_n2569_, new_n2570_, new_n2571_, new_n2572_, new_n2573_, new_n2574_,
    new_n2575_, new_n2576_, new_n2577_, new_n2578_, new_n2579_, new_n2580_,
    new_n2581_, new_n2582_, new_n2583_, new_n2584_, new_n2585_, new_n2586_,
    new_n2587_, new_n2588_, new_n2589_, new_n2590_, new_n2591_, new_n2592_,
    new_n2593_, new_n2594_, new_n2595_, new_n2596_, new_n2597_, new_n2598_,
    new_n2599_, new_n2600_, new_n2601_, new_n2602_, new_n2603_, new_n2604_,
    new_n2605_, new_n2606_, new_n2607_, new_n2608_, new_n2609_, new_n2610_,
    new_n2611_, new_n2612_, new_n2613_, new_n2614_, new_n2615_, new_n2616_,
    new_n2617_, new_n2618_, new_n2619_, new_n2620_, new_n2621_, new_n2622_,
    new_n2623_, new_n2624_, new_n2625_, new_n2626_, new_n2627_, new_n2628_,
    new_n2629_, new_n2630_, new_n2631_, new_n2632_, new_n2633_, new_n2634_,
    new_n2635_, new_n2636_, new_n2637_, new_n2638_, new_n2639_, new_n2640_,
    new_n2641_, new_n2642_, new_n2643_, new_n2644_, new_n2645_, new_n2646_,
    new_n2647_, new_n2648_, new_n2649_, new_n2650_, new_n2651_, new_n2652_,
    new_n2653_, new_n2654_, new_n2655_, new_n2656_, new_n2657_, new_n2658_,
    new_n2659_, new_n2660_, new_n2661_, new_n2662_, new_n2663_, new_n2664_,
    new_n2665_, new_n2666_, new_n2667_, new_n2668_, new_n2669_, new_n2670_,
    new_n2671_, new_n2672_, new_n2673_, new_n2674_, new_n2675_, new_n2676_,
    new_n2677_, new_n2678_, new_n2679_, new_n2680_, new_n2681_, new_n2682_,
    new_n2683_, new_n2684_, new_n2685_, new_n2686_, new_n2687_, new_n2688_,
    new_n2689_, new_n2690_, new_n2691_, new_n2692_, new_n2693_, new_n2694_,
    new_n2695_, new_n2696_, new_n2697_, new_n2698_, new_n2699_, new_n2700_,
    new_n2701_, new_n2702_, new_n2703_, new_n2704_, new_n2705_, new_n2706_,
    new_n2707_, new_n2708_, new_n2709_, new_n2710_, new_n2711_, new_n2712_,
    new_n2713_, new_n2714_, new_n2715_, new_n2716_, new_n2717_, new_n2718_,
    new_n2719_, new_n2720_, new_n2721_, new_n2722_, new_n2723_, new_n2724_,
    new_n2725_, new_n2726_, new_n2727_, new_n2728_, new_n2729_, new_n2730_,
    new_n2731_, new_n2732_, new_n2733_, new_n2734_, new_n2735_, new_n2736_,
    new_n2737_, new_n2738_, new_n2739_, new_n2740_, new_n2741_, new_n2742_,
    new_n2743_, new_n2744_, new_n2745_, new_n2746_, new_n2747_, new_n2748_,
    new_n2749_, new_n2750_, new_n2751_, new_n2752_, new_n2753_, new_n2754_,
    new_n2755_, new_n2756_, new_n2757_, new_n2758_, new_n2759_, new_n2760_,
    new_n2761_, new_n2762_, new_n2763_, new_n2764_, new_n2765_, new_n2769_,
    new_n2773_, new_n2777_, new_n2780_, new_n2783_, new_n2786_, new_n2788_,
    new_n2791_, new_n2794_, new_n2797_, new_n2801_, new_n2804_, new_n2807_,
    new_n2810_, new_n2812_, new_n2814_, new_n2816_, new_n2819_, new_n2821_,
    new_n2824_, new_n2830_, new_n2832_, new_n2835_, new_n2837_, new_n2839_,
    new_n2841_, new_n2844_, new_n2846_, new_n2854_, new_n2856_, new_n2859_,
    new_n2862_, new_n2867_, new_n2870_, new_n2873_, new_n2878_, new_n2881_,
    new_n2884_, new_n2889_, new_n2892_, new_n2895_, new_n2900_, new_n2903_,
    new_n2906_, new_n2911_, new_n2914_, new_n2917_, new_n2922_, new_n2925_,
    new_n2928_, new_n2933_, new_n2936_, new_n2939_, new_n2945_, new_n2947_,
    new_n2949_, new_n2950_, new_n2952_;
  INVX1    g0000(.A(\in3[0] ), .Y(new_n643_));
  INVX1    g0001(.A(\in2[31] ), .Y(new_n644_));
  AND2X1   g0002(.A(\in3[31] ), .B(new_n644_), .Y(new_n645_));
  INVX1    g0003(.A(\in2[30] ), .Y(new_n646_));
  AND2X1   g0004(.A(\in3[30] ), .B(new_n646_), .Y(new_n647_));
  INVX1    g0005(.A(new_n647_), .Y(new_n648_));
  INVX1    g0006(.A(\in2[29] ), .Y(new_n649_));
  AND2X1   g0007(.A(\in3[29] ), .B(new_n649_), .Y(new_n650_));
  INVX1    g0008(.A(\in2[28] ), .Y(new_n651_));
  AND2X1   g0009(.A(\in3[28] ), .B(new_n651_), .Y(new_n652_));
  INVX1    g0010(.A(new_n652_), .Y(new_n653_));
  INVX1    g0011(.A(\in2[27] ), .Y(new_n654_));
  AND2X1   g0012(.A(\in3[27] ), .B(new_n654_), .Y(new_n655_));
  INVX1    g0013(.A(\in2[26] ), .Y(new_n656_));
  AND2X1   g0014(.A(\in3[26] ), .B(new_n656_), .Y(new_n657_));
  INVX1    g0015(.A(new_n657_), .Y(new_n658_));
  INVX1    g0016(.A(\in2[24] ), .Y(new_n659_));
  INVX1    g0017(.A(\in2[23] ), .Y(new_n660_));
  AND2X1   g0018(.A(\in3[23] ), .B(new_n660_), .Y(new_n661_));
  INVX1    g0019(.A(new_n661_), .Y(new_n662_));
  INVX1    g0020(.A(\in2[22] ), .Y(new_n663_));
  AND2X1   g0021(.A(\in3[22] ), .B(new_n663_), .Y(new_n664_));
  INVX1    g0022(.A(\in2[21] ), .Y(new_n665_));
  AND2X1   g0023(.A(\in3[21] ), .B(new_n665_), .Y(new_n666_));
  INVX1    g0024(.A(new_n666_), .Y(new_n667_));
  INVX1    g0025(.A(\in2[20] ), .Y(new_n668_));
  AND2X1   g0026(.A(\in3[20] ), .B(new_n668_), .Y(new_n669_));
  INVX1    g0027(.A(\in2[19] ), .Y(new_n670_));
  AND2X1   g0028(.A(\in3[19] ), .B(new_n670_), .Y(new_n671_));
  INVX1    g0029(.A(new_n671_), .Y(new_n672_));
  INVX1    g0030(.A(\in2[18] ), .Y(new_n673_));
  AND2X1   g0031(.A(\in3[18] ), .B(new_n673_), .Y(new_n674_));
  INVX1    g0032(.A(\in3[17] ), .Y(new_n675_));
  INVX1    g0033(.A(\in2[17] ), .Y(new_n676_));
  INVX1    g0034(.A(\in3[16] ), .Y(new_n677_));
  INVX1    g0035(.A(\in2[15] ), .Y(new_n678_));
  AND2X1   g0036(.A(\in3[15] ), .B(new_n678_), .Y(new_n679_));
  INVX1    g0037(.A(\in2[14] ), .Y(new_n680_));
  AND2X1   g0038(.A(\in3[14] ), .B(new_n680_), .Y(new_n681_));
  INVX1    g0039(.A(new_n681_), .Y(new_n682_));
  INVX1    g0040(.A(\in2[13] ), .Y(new_n683_));
  AND2X1   g0041(.A(\in3[13] ), .B(new_n683_), .Y(new_n684_));
  INVX1    g0042(.A(\in2[12] ), .Y(new_n685_));
  AND2X1   g0043(.A(\in3[12] ), .B(new_n685_), .Y(new_n686_));
  INVX1    g0044(.A(new_n686_), .Y(new_n687_));
  INVX1    g0045(.A(\in2[11] ), .Y(new_n688_));
  AND2X1   g0046(.A(\in3[11] ), .B(new_n688_), .Y(new_n689_));
  INVX1    g0047(.A(\in2[10] ), .Y(new_n690_));
  AND2X1   g0048(.A(\in3[10] ), .B(new_n690_), .Y(new_n691_));
  INVX1    g0049(.A(new_n691_), .Y(new_n692_));
  INVX1    g0050(.A(\in2[8] ), .Y(new_n693_));
  INVX1    g0051(.A(\in2[7] ), .Y(new_n694_));
  AND2X1   g0052(.A(\in3[7] ), .B(new_n694_), .Y(new_n695_));
  INVX1    g0053(.A(new_n695_), .Y(new_n696_));
  INVX1    g0054(.A(\in2[6] ), .Y(new_n697_));
  AND2X1   g0055(.A(\in3[6] ), .B(new_n697_), .Y(new_n698_));
  INVX1    g0056(.A(\in3[5] ), .Y(new_n699_));
  INVX1    g0057(.A(\in2[5] ), .Y(new_n700_));
  INVX1    g0058(.A(\in3[4] ), .Y(new_n701_));
  INVX1    g0059(.A(\in2[3] ), .Y(new_n702_));
  AND2X1   g0060(.A(\in3[3] ), .B(new_n702_), .Y(new_n703_));
  INVX1    g0061(.A(\in3[2] ), .Y(new_n704_));
  INVX1    g0062(.A(\in2[1] ), .Y(new_n705_));
  INVX1    g0063(.A(\in2[0] ), .Y(new_n706_));
  OR2X1    g0064(.A(\in3[0] ), .B(new_n706_), .Y(new_n707_));
  OAI21X1  g0065(.A0(new_n707_), .A1(new_n705_), .B0(\in3[1] ), .Y(new_n708_));
  INVX1    g0066(.A(\in2[2] ), .Y(new_n709_));
  AOI22X1  g0067(.A0(new_n707_), .A1(new_n705_), .B0(\in3[2] ), .B1(new_n709_), .Y(new_n710_));
  AOI22X1  g0068(.A0(new_n710_), .A1(new_n708_), .B0(new_n704_), .B1(\in2[2] ), .Y(new_n711_));
  INVX1    g0069(.A(\in3[3] ), .Y(new_n712_));
  AND2X1   g0070(.A(new_n712_), .B(\in2[3] ), .Y(new_n713_));
  INVX1    g0071(.A(new_n713_), .Y(new_n714_));
  OAI21X1  g0072(.A0(new_n711_), .A1(new_n703_), .B0(new_n714_), .Y(new_n715_));
  OAI21X1  g0073(.A0(new_n715_), .A1(\in2[4] ), .B0(new_n701_), .Y(new_n716_));
  INVX1    g0074(.A(\in2[4] ), .Y(new_n717_));
  INVX1    g0075(.A(new_n703_), .Y(new_n718_));
  INVX1    g0076(.A(\in3[1] ), .Y(new_n719_));
  AND2X1   g0077(.A(new_n643_), .B(\in2[0] ), .Y(new_n720_));
  AOI21X1  g0078(.A0(new_n720_), .A1(\in2[1] ), .B0(new_n719_), .Y(new_n721_));
  OAI22X1  g0079(.A0(new_n720_), .A1(\in2[1] ), .B0(new_n704_), .B1(\in2[2] ), .Y(new_n722_));
  OAI22X1  g0080(.A0(new_n722_), .A1(new_n721_), .B0(\in3[2] ), .B1(new_n709_), .Y(new_n723_));
  AOI21X1  g0081(.A0(new_n723_), .A1(new_n718_), .B0(new_n713_), .Y(new_n724_));
  OR2X1    g0082(.A(new_n724_), .B(new_n717_), .Y(new_n725_));
  NAND3X1  g0083(.A(new_n725_), .B(new_n716_), .C(new_n700_), .Y(new_n726_));
  AOI21X1  g0084(.A0(new_n725_), .A1(new_n716_), .B0(new_n700_), .Y(new_n727_));
  AOI21X1  g0085(.A0(new_n726_), .A1(new_n699_), .B0(new_n727_), .Y(new_n728_));
  INVX1    g0086(.A(\in3[6] ), .Y(new_n729_));
  AND2X1   g0087(.A(new_n729_), .B(\in2[6] ), .Y(new_n730_));
  INVX1    g0088(.A(new_n730_), .Y(new_n731_));
  OAI21X1  g0089(.A0(new_n728_), .A1(new_n698_), .B0(new_n731_), .Y(new_n732_));
  INVX1    g0090(.A(\in3[7] ), .Y(new_n733_));
  AND2X1   g0091(.A(new_n733_), .B(\in2[7] ), .Y(new_n734_));
  AOI21X1  g0092(.A0(new_n732_), .A1(new_n696_), .B0(new_n734_), .Y(new_n735_));
  AOI21X1  g0093(.A0(new_n735_), .A1(new_n693_), .B0(\in3[8] ), .Y(new_n736_));
  INVX1    g0094(.A(new_n698_), .Y(new_n737_));
  AOI21X1  g0095(.A0(new_n724_), .A1(new_n717_), .B0(\in3[4] ), .Y(new_n738_));
  AND2X1   g0096(.A(new_n715_), .B(\in2[4] ), .Y(new_n739_));
  NOR3X1   g0097(.A(new_n739_), .B(new_n738_), .C(\in2[5] ), .Y(new_n740_));
  OAI21X1  g0098(.A0(new_n739_), .A1(new_n738_), .B0(\in2[5] ), .Y(new_n741_));
  OAI21X1  g0099(.A0(new_n740_), .A1(\in3[5] ), .B0(new_n741_), .Y(new_n742_));
  AOI21X1  g0100(.A0(new_n742_), .A1(new_n737_), .B0(new_n730_), .Y(new_n743_));
  INVX1    g0101(.A(new_n734_), .Y(new_n744_));
  OAI21X1  g0102(.A0(new_n743_), .A1(new_n695_), .B0(new_n744_), .Y(new_n745_));
  AND2X1   g0103(.A(new_n745_), .B(\in2[8] ), .Y(new_n746_));
  NOR3X1   g0104(.A(new_n746_), .B(new_n736_), .C(\in2[9] ), .Y(new_n747_));
  OAI21X1  g0105(.A0(new_n746_), .A1(new_n736_), .B0(\in2[9] ), .Y(new_n748_));
  OAI21X1  g0106(.A0(new_n747_), .A1(\in3[9] ), .B0(new_n748_), .Y(new_n749_));
  INVX1    g0107(.A(\in3[10] ), .Y(new_n750_));
  AND2X1   g0108(.A(new_n750_), .B(\in2[10] ), .Y(new_n751_));
  AOI21X1  g0109(.A0(new_n749_), .A1(new_n692_), .B0(new_n751_), .Y(new_n752_));
  INVX1    g0110(.A(\in3[11] ), .Y(new_n753_));
  AND2X1   g0111(.A(new_n753_), .B(\in2[11] ), .Y(new_n754_));
  INVX1    g0112(.A(new_n754_), .Y(new_n755_));
  OAI21X1  g0113(.A0(new_n752_), .A1(new_n689_), .B0(new_n755_), .Y(new_n756_));
  INVX1    g0114(.A(\in3[12] ), .Y(new_n757_));
  AND2X1   g0115(.A(new_n757_), .B(\in2[12] ), .Y(new_n758_));
  AOI21X1  g0116(.A0(new_n756_), .A1(new_n687_), .B0(new_n758_), .Y(new_n759_));
  INVX1    g0117(.A(\in3[13] ), .Y(new_n760_));
  AND2X1   g0118(.A(new_n760_), .B(\in2[13] ), .Y(new_n761_));
  INVX1    g0119(.A(new_n761_), .Y(new_n762_));
  OAI21X1  g0120(.A0(new_n759_), .A1(new_n684_), .B0(new_n762_), .Y(new_n763_));
  INVX1    g0121(.A(\in3[14] ), .Y(new_n764_));
  AND2X1   g0122(.A(new_n764_), .B(\in2[14] ), .Y(new_n765_));
  AOI21X1  g0123(.A0(new_n763_), .A1(new_n682_), .B0(new_n765_), .Y(new_n766_));
  INVX1    g0124(.A(\in3[15] ), .Y(new_n767_));
  AND2X1   g0125(.A(new_n767_), .B(\in2[15] ), .Y(new_n768_));
  INVX1    g0126(.A(new_n768_), .Y(new_n769_));
  OAI21X1  g0127(.A0(new_n766_), .A1(new_n679_), .B0(new_n769_), .Y(new_n770_));
  OAI21X1  g0128(.A0(new_n770_), .A1(\in2[16] ), .B0(new_n677_), .Y(new_n771_));
  INVX1    g0129(.A(\in2[16] ), .Y(new_n772_));
  INVX1    g0130(.A(new_n679_), .Y(new_n773_));
  INVX1    g0131(.A(new_n684_), .Y(new_n774_));
  INVX1    g0132(.A(new_n689_), .Y(new_n775_));
  INVX1    g0133(.A(\in3[9] ), .Y(new_n776_));
  INVX1    g0134(.A(\in2[9] ), .Y(new_n777_));
  INVX1    g0135(.A(\in3[8] ), .Y(new_n778_));
  OAI21X1  g0136(.A0(new_n745_), .A1(\in2[8] ), .B0(new_n778_), .Y(new_n779_));
  OR2X1    g0137(.A(new_n735_), .B(new_n693_), .Y(new_n780_));
  NAND3X1  g0138(.A(new_n780_), .B(new_n779_), .C(new_n777_), .Y(new_n781_));
  AOI21X1  g0139(.A0(new_n780_), .A1(new_n779_), .B0(new_n777_), .Y(new_n782_));
  AOI21X1  g0140(.A0(new_n781_), .A1(new_n776_), .B0(new_n782_), .Y(new_n783_));
  INVX1    g0141(.A(new_n751_), .Y(new_n784_));
  OAI21X1  g0142(.A0(new_n783_), .A1(new_n691_), .B0(new_n784_), .Y(new_n785_));
  AOI21X1  g0143(.A0(new_n785_), .A1(new_n775_), .B0(new_n754_), .Y(new_n786_));
  INVX1    g0144(.A(new_n758_), .Y(new_n787_));
  OAI21X1  g0145(.A0(new_n786_), .A1(new_n686_), .B0(new_n787_), .Y(new_n788_));
  AOI21X1  g0146(.A0(new_n788_), .A1(new_n774_), .B0(new_n761_), .Y(new_n789_));
  INVX1    g0147(.A(new_n765_), .Y(new_n790_));
  OAI21X1  g0148(.A0(new_n789_), .A1(new_n681_), .B0(new_n790_), .Y(new_n791_));
  AOI21X1  g0149(.A0(new_n791_), .A1(new_n773_), .B0(new_n768_), .Y(new_n792_));
  OR2X1    g0150(.A(new_n792_), .B(new_n772_), .Y(new_n793_));
  NAND3X1  g0151(.A(new_n793_), .B(new_n771_), .C(new_n676_), .Y(new_n794_));
  AOI21X1  g0152(.A0(new_n793_), .A1(new_n771_), .B0(new_n676_), .Y(new_n795_));
  AOI21X1  g0153(.A0(new_n794_), .A1(new_n675_), .B0(new_n795_), .Y(new_n796_));
  INVX1    g0154(.A(\in3[18] ), .Y(new_n797_));
  AND2X1   g0155(.A(new_n797_), .B(\in2[18] ), .Y(new_n798_));
  INVX1    g0156(.A(new_n798_), .Y(new_n799_));
  OAI21X1  g0157(.A0(new_n796_), .A1(new_n674_), .B0(new_n799_), .Y(new_n800_));
  INVX1    g0158(.A(\in3[19] ), .Y(new_n801_));
  AND2X1   g0159(.A(new_n801_), .B(\in2[19] ), .Y(new_n802_));
  AOI21X1  g0160(.A0(new_n800_), .A1(new_n672_), .B0(new_n802_), .Y(new_n803_));
  INVX1    g0161(.A(\in3[20] ), .Y(new_n804_));
  AND2X1   g0162(.A(new_n804_), .B(\in2[20] ), .Y(new_n805_));
  INVX1    g0163(.A(new_n805_), .Y(new_n806_));
  OAI21X1  g0164(.A0(new_n803_), .A1(new_n669_), .B0(new_n806_), .Y(new_n807_));
  INVX1    g0165(.A(\in3[21] ), .Y(new_n808_));
  AND2X1   g0166(.A(new_n808_), .B(\in2[21] ), .Y(new_n809_));
  AOI21X1  g0167(.A0(new_n807_), .A1(new_n667_), .B0(new_n809_), .Y(new_n810_));
  INVX1    g0168(.A(\in3[22] ), .Y(new_n811_));
  AND2X1   g0169(.A(new_n811_), .B(\in2[22] ), .Y(new_n812_));
  INVX1    g0170(.A(new_n812_), .Y(new_n813_));
  OAI21X1  g0171(.A0(new_n810_), .A1(new_n664_), .B0(new_n813_), .Y(new_n814_));
  INVX1    g0172(.A(\in3[23] ), .Y(new_n815_));
  AND2X1   g0173(.A(new_n815_), .B(\in2[23] ), .Y(new_n816_));
  AOI21X1  g0174(.A0(new_n814_), .A1(new_n662_), .B0(new_n816_), .Y(new_n817_));
  AOI21X1  g0175(.A0(new_n817_), .A1(new_n659_), .B0(\in3[24] ), .Y(new_n818_));
  INVX1    g0176(.A(new_n664_), .Y(new_n819_));
  INVX1    g0177(.A(new_n669_), .Y(new_n820_));
  INVX1    g0178(.A(new_n674_), .Y(new_n821_));
  AOI21X1  g0179(.A0(new_n792_), .A1(new_n772_), .B0(\in3[16] ), .Y(new_n822_));
  AND2X1   g0180(.A(new_n770_), .B(\in2[16] ), .Y(new_n823_));
  NOR3X1   g0181(.A(new_n823_), .B(new_n822_), .C(\in2[17] ), .Y(new_n824_));
  OAI21X1  g0182(.A0(new_n823_), .A1(new_n822_), .B0(\in2[17] ), .Y(new_n825_));
  OAI21X1  g0183(.A0(new_n824_), .A1(\in3[17] ), .B0(new_n825_), .Y(new_n826_));
  AOI21X1  g0184(.A0(new_n826_), .A1(new_n821_), .B0(new_n798_), .Y(new_n827_));
  INVX1    g0185(.A(new_n802_), .Y(new_n828_));
  OAI21X1  g0186(.A0(new_n827_), .A1(new_n671_), .B0(new_n828_), .Y(new_n829_));
  AOI21X1  g0187(.A0(new_n829_), .A1(new_n820_), .B0(new_n805_), .Y(new_n830_));
  INVX1    g0188(.A(new_n809_), .Y(new_n831_));
  OAI21X1  g0189(.A0(new_n830_), .A1(new_n666_), .B0(new_n831_), .Y(new_n832_));
  AOI21X1  g0190(.A0(new_n832_), .A1(new_n819_), .B0(new_n812_), .Y(new_n833_));
  INVX1    g0191(.A(new_n816_), .Y(new_n834_));
  OAI21X1  g0192(.A0(new_n833_), .A1(new_n661_), .B0(new_n834_), .Y(new_n835_));
  AND2X1   g0193(.A(new_n835_), .B(\in2[24] ), .Y(new_n836_));
  NOR3X1   g0194(.A(new_n836_), .B(new_n818_), .C(\in2[25] ), .Y(new_n837_));
  OAI21X1  g0195(.A0(new_n836_), .A1(new_n818_), .B0(\in2[25] ), .Y(new_n838_));
  OAI21X1  g0196(.A0(new_n837_), .A1(\in3[25] ), .B0(new_n838_), .Y(new_n839_));
  INVX1    g0197(.A(\in3[26] ), .Y(new_n840_));
  AND2X1   g0198(.A(new_n840_), .B(\in2[26] ), .Y(new_n841_));
  AOI21X1  g0199(.A0(new_n839_), .A1(new_n658_), .B0(new_n841_), .Y(new_n842_));
  INVX1    g0200(.A(\in3[27] ), .Y(new_n843_));
  AND2X1   g0201(.A(new_n843_), .B(\in2[27] ), .Y(new_n844_));
  INVX1    g0202(.A(new_n844_), .Y(new_n845_));
  OAI21X1  g0203(.A0(new_n842_), .A1(new_n655_), .B0(new_n845_), .Y(new_n846_));
  INVX1    g0204(.A(\in3[28] ), .Y(new_n847_));
  AND2X1   g0205(.A(new_n847_), .B(\in2[28] ), .Y(new_n848_));
  AOI21X1  g0206(.A0(new_n846_), .A1(new_n653_), .B0(new_n848_), .Y(new_n849_));
  INVX1    g0207(.A(\in3[29] ), .Y(new_n850_));
  AND2X1   g0208(.A(new_n850_), .B(\in2[29] ), .Y(new_n851_));
  INVX1    g0209(.A(new_n851_), .Y(new_n852_));
  OAI21X1  g0210(.A0(new_n849_), .A1(new_n650_), .B0(new_n852_), .Y(new_n853_));
  INVX1    g0211(.A(\in3[30] ), .Y(new_n854_));
  AND2X1   g0212(.A(new_n854_), .B(\in2[30] ), .Y(new_n855_));
  AOI21X1  g0213(.A0(new_n853_), .A1(new_n648_), .B0(new_n855_), .Y(new_n856_));
  INVX1    g0214(.A(\in3[31] ), .Y(new_n857_));
  AND2X1   g0215(.A(new_n857_), .B(\in2[31] ), .Y(new_n858_));
  INVX1    g0216(.A(new_n858_), .Y(new_n859_));
  OAI21X1  g0217(.A0(new_n856_), .A1(new_n645_), .B0(new_n859_), .Y(new_n860_));
  INVX1    g0218(.A(\in2[38] ), .Y(new_n861_));
  INVX1    g0219(.A(\in2[39] ), .Y(new_n862_));
  AOI22X1  g0220(.A0(\in3[39] ), .A1(new_n862_), .B0(\in3[38] ), .B1(new_n861_), .Y(new_n863_));
  INVX1    g0221(.A(new_n863_), .Y(new_n864_));
  INVX1    g0222(.A(\in3[36] ), .Y(new_n865_));
  INVX1    g0223(.A(\in3[37] ), .Y(new_n866_));
  OAI22X1  g0224(.A0(new_n866_), .A1(\in2[37] ), .B0(new_n865_), .B1(\in2[36] ), .Y(new_n867_));
  INVX1    g0225(.A(\in2[34] ), .Y(new_n868_));
  INVX1    g0226(.A(\in2[35] ), .Y(new_n869_));
  AOI22X1  g0227(.A0(\in3[35] ), .A1(new_n869_), .B0(\in3[34] ), .B1(new_n868_), .Y(new_n870_));
  INVX1    g0228(.A(new_n870_), .Y(new_n871_));
  INVX1    g0229(.A(\in3[32] ), .Y(new_n872_));
  INVX1    g0230(.A(\in3[33] ), .Y(new_n873_));
  OAI22X1  g0231(.A0(new_n873_), .A1(\in2[33] ), .B0(new_n872_), .B1(\in2[32] ), .Y(new_n874_));
  NOR4X1   g0232(.A(new_n874_), .B(new_n871_), .C(new_n867_), .D(new_n864_), .Y(new_n875_));
  NOR2X1   g0233(.A(new_n867_), .B(new_n864_), .Y(new_n876_));
  AND2X1   g0234(.A(new_n872_), .B(\in2[32] ), .Y(new_n877_));
  OAI21X1  g0235(.A0(new_n873_), .A1(\in2[33] ), .B0(new_n877_), .Y(new_n878_));
  INVX1    g0236(.A(\in3[34] ), .Y(new_n879_));
  AOI22X1  g0237(.A0(new_n879_), .A1(\in2[34] ), .B0(new_n873_), .B1(\in2[33] ), .Y(new_n880_));
  AND2X1   g0238(.A(new_n880_), .B(new_n878_), .Y(new_n881_));
  OAI22X1  g0239(.A0(new_n881_), .A1(new_n871_), .B0(\in3[35] ), .B1(new_n869_), .Y(new_n882_));
  INVX1    g0240(.A(\in2[36] ), .Y(new_n883_));
  INVX1    g0241(.A(\in2[37] ), .Y(new_n884_));
  AND2X1   g0242(.A(\in3[37] ), .B(new_n884_), .Y(new_n885_));
  NOR3X1   g0243(.A(new_n885_), .B(\in3[36] ), .C(new_n883_), .Y(new_n886_));
  AOI21X1  g0244(.A0(new_n866_), .A1(\in2[37] ), .B0(new_n886_), .Y(new_n887_));
  INVX1    g0245(.A(\in3[39] ), .Y(new_n888_));
  AND2X1   g0246(.A(\in3[39] ), .B(new_n862_), .Y(new_n889_));
  NOR3X1   g0247(.A(new_n889_), .B(\in3[38] ), .C(new_n861_), .Y(new_n890_));
  AOI21X1  g0248(.A0(new_n888_), .A1(\in2[39] ), .B0(new_n890_), .Y(new_n891_));
  OAI21X1  g0249(.A0(new_n887_), .A1(new_n864_), .B0(new_n891_), .Y(new_n892_));
  AOI21X1  g0250(.A0(new_n882_), .A1(new_n876_), .B0(new_n892_), .Y(new_n893_));
  INVX1    g0251(.A(new_n893_), .Y(new_n894_));
  AOI21X1  g0252(.A0(new_n875_), .A1(new_n860_), .B0(new_n894_), .Y(new_n895_));
  INVX1    g0253(.A(\in2[46] ), .Y(new_n896_));
  INVX1    g0254(.A(\in2[47] ), .Y(new_n897_));
  AOI22X1  g0255(.A0(\in3[47] ), .A1(new_n897_), .B0(\in3[46] ), .B1(new_n896_), .Y(new_n898_));
  INVX1    g0256(.A(new_n898_), .Y(new_n899_));
  INVX1    g0257(.A(\in3[44] ), .Y(new_n900_));
  INVX1    g0258(.A(\in3[45] ), .Y(new_n901_));
  OAI22X1  g0259(.A0(new_n901_), .A1(\in2[45] ), .B0(new_n900_), .B1(\in2[44] ), .Y(new_n902_));
  INVX1    g0260(.A(\in2[42] ), .Y(new_n903_));
  INVX1    g0261(.A(\in2[43] ), .Y(new_n904_));
  AOI22X1  g0262(.A0(\in3[43] ), .A1(new_n904_), .B0(\in3[42] ), .B1(new_n903_), .Y(new_n905_));
  INVX1    g0263(.A(new_n905_), .Y(new_n906_));
  INVX1    g0264(.A(\in3[40] ), .Y(new_n907_));
  INVX1    g0265(.A(\in3[41] ), .Y(new_n908_));
  OAI22X1  g0266(.A0(new_n908_), .A1(\in2[41] ), .B0(new_n907_), .B1(\in2[40] ), .Y(new_n909_));
  NOR4X1   g0267(.A(new_n909_), .B(new_n906_), .C(new_n902_), .D(new_n899_), .Y(new_n910_));
  INVX1    g0268(.A(new_n910_), .Y(new_n911_));
  NOR2X1   g0269(.A(new_n902_), .B(new_n899_), .Y(new_n912_));
  AND2X1   g0270(.A(new_n907_), .B(\in2[40] ), .Y(new_n913_));
  OAI21X1  g0271(.A0(new_n908_), .A1(\in2[41] ), .B0(new_n913_), .Y(new_n914_));
  INVX1    g0272(.A(\in3[42] ), .Y(new_n915_));
  AOI22X1  g0273(.A0(new_n915_), .A1(\in2[42] ), .B0(new_n908_), .B1(\in2[41] ), .Y(new_n916_));
  AND2X1   g0274(.A(new_n916_), .B(new_n914_), .Y(new_n917_));
  OAI22X1  g0275(.A0(new_n917_), .A1(new_n906_), .B0(\in3[43] ), .B1(new_n904_), .Y(new_n918_));
  INVX1    g0276(.A(\in2[44] ), .Y(new_n919_));
  INVX1    g0277(.A(\in2[45] ), .Y(new_n920_));
  AND2X1   g0278(.A(\in3[45] ), .B(new_n920_), .Y(new_n921_));
  NOR3X1   g0279(.A(new_n921_), .B(\in3[44] ), .C(new_n919_), .Y(new_n922_));
  AOI21X1  g0280(.A0(new_n901_), .A1(\in2[45] ), .B0(new_n922_), .Y(new_n923_));
  INVX1    g0281(.A(\in3[47] ), .Y(new_n924_));
  AND2X1   g0282(.A(\in3[47] ), .B(new_n897_), .Y(new_n925_));
  NOR3X1   g0283(.A(new_n925_), .B(\in3[46] ), .C(new_n896_), .Y(new_n926_));
  AOI21X1  g0284(.A0(new_n924_), .A1(\in2[47] ), .B0(new_n926_), .Y(new_n927_));
  OAI21X1  g0285(.A0(new_n923_), .A1(new_n899_), .B0(new_n927_), .Y(new_n928_));
  AOI21X1  g0286(.A0(new_n918_), .A1(new_n912_), .B0(new_n928_), .Y(new_n929_));
  OAI21X1  g0287(.A0(new_n911_), .A1(new_n895_), .B0(new_n929_), .Y(new_n930_));
  INVX1    g0288(.A(\in2[54] ), .Y(new_n931_));
  INVX1    g0289(.A(\in2[55] ), .Y(new_n932_));
  AOI22X1  g0290(.A0(\in3[55] ), .A1(new_n932_), .B0(\in3[54] ), .B1(new_n931_), .Y(new_n933_));
  INVX1    g0291(.A(new_n933_), .Y(new_n934_));
  INVX1    g0292(.A(\in3[52] ), .Y(new_n935_));
  INVX1    g0293(.A(\in3[53] ), .Y(new_n936_));
  OAI22X1  g0294(.A0(new_n936_), .A1(\in2[53] ), .B0(new_n935_), .B1(\in2[52] ), .Y(new_n937_));
  INVX1    g0295(.A(\in2[50] ), .Y(new_n938_));
  INVX1    g0296(.A(\in2[51] ), .Y(new_n939_));
  AOI22X1  g0297(.A0(\in3[51] ), .A1(new_n939_), .B0(\in3[50] ), .B1(new_n938_), .Y(new_n940_));
  INVX1    g0298(.A(new_n940_), .Y(new_n941_));
  INVX1    g0299(.A(\in3[48] ), .Y(new_n942_));
  INVX1    g0300(.A(\in3[49] ), .Y(new_n943_));
  OAI22X1  g0301(.A0(new_n943_), .A1(\in2[49] ), .B0(new_n942_), .B1(\in2[48] ), .Y(new_n944_));
  NOR4X1   g0302(.A(new_n944_), .B(new_n941_), .C(new_n937_), .D(new_n934_), .Y(new_n945_));
  NOR2X1   g0303(.A(new_n937_), .B(new_n934_), .Y(new_n946_));
  AND2X1   g0304(.A(new_n942_), .B(\in2[48] ), .Y(new_n947_));
  OAI21X1  g0305(.A0(new_n943_), .A1(\in2[49] ), .B0(new_n947_), .Y(new_n948_));
  INVX1    g0306(.A(\in3[50] ), .Y(new_n949_));
  AOI22X1  g0307(.A0(new_n949_), .A1(\in2[50] ), .B0(new_n943_), .B1(\in2[49] ), .Y(new_n950_));
  AND2X1   g0308(.A(new_n950_), .B(new_n948_), .Y(new_n951_));
  OAI22X1  g0309(.A0(new_n951_), .A1(new_n941_), .B0(\in3[51] ), .B1(new_n939_), .Y(new_n952_));
  AND2X1   g0310(.A(new_n935_), .B(\in2[52] ), .Y(new_n953_));
  OAI21X1  g0311(.A0(new_n936_), .A1(\in2[53] ), .B0(new_n953_), .Y(new_n954_));
  INVX1    g0312(.A(\in3[54] ), .Y(new_n955_));
  AOI22X1  g0313(.A0(new_n955_), .A1(\in2[54] ), .B0(new_n936_), .B1(\in2[53] ), .Y(new_n956_));
  AND2X1   g0314(.A(new_n956_), .B(new_n954_), .Y(new_n957_));
  OAI22X1  g0315(.A0(new_n957_), .A1(new_n934_), .B0(\in3[55] ), .B1(new_n932_), .Y(new_n958_));
  AOI21X1  g0316(.A0(new_n952_), .A1(new_n946_), .B0(new_n958_), .Y(new_n959_));
  INVX1    g0317(.A(new_n959_), .Y(new_n960_));
  AOI21X1  g0318(.A0(new_n945_), .A1(new_n930_), .B0(new_n960_), .Y(new_n961_));
  INVX1    g0319(.A(\in2[62] ), .Y(new_n962_));
  INVX1    g0320(.A(\in2[63] ), .Y(new_n963_));
  AOI22X1  g0321(.A0(\in3[63] ), .A1(new_n963_), .B0(\in3[62] ), .B1(new_n962_), .Y(new_n964_));
  INVX1    g0322(.A(new_n964_), .Y(new_n965_));
  INVX1    g0323(.A(\in3[60] ), .Y(new_n966_));
  INVX1    g0324(.A(\in3[61] ), .Y(new_n967_));
  OAI22X1  g0325(.A0(new_n967_), .A1(\in2[61] ), .B0(new_n966_), .B1(\in2[60] ), .Y(new_n968_));
  INVX1    g0326(.A(\in2[58] ), .Y(new_n969_));
  INVX1    g0327(.A(\in2[59] ), .Y(new_n970_));
  AOI22X1  g0328(.A0(\in3[59] ), .A1(new_n970_), .B0(\in3[58] ), .B1(new_n969_), .Y(new_n971_));
  INVX1    g0329(.A(new_n971_), .Y(new_n972_));
  INVX1    g0330(.A(\in3[56] ), .Y(new_n973_));
  INVX1    g0331(.A(\in3[57] ), .Y(new_n974_));
  OAI22X1  g0332(.A0(new_n974_), .A1(\in2[57] ), .B0(new_n973_), .B1(\in2[56] ), .Y(new_n975_));
  NOR4X1   g0333(.A(new_n975_), .B(new_n972_), .C(new_n968_), .D(new_n965_), .Y(new_n976_));
  INVX1    g0334(.A(new_n976_), .Y(new_n977_));
  NOR2X1   g0335(.A(new_n968_), .B(new_n965_), .Y(new_n978_));
  AND2X1   g0336(.A(new_n973_), .B(\in2[56] ), .Y(new_n979_));
  OAI21X1  g0337(.A0(new_n974_), .A1(\in2[57] ), .B0(new_n979_), .Y(new_n980_));
  INVX1    g0338(.A(\in3[58] ), .Y(new_n981_));
  AOI22X1  g0339(.A0(new_n981_), .A1(\in2[58] ), .B0(new_n974_), .B1(\in2[57] ), .Y(new_n982_));
  AND2X1   g0340(.A(new_n982_), .B(new_n980_), .Y(new_n983_));
  OAI22X1  g0341(.A0(new_n983_), .A1(new_n972_), .B0(\in3[59] ), .B1(new_n970_), .Y(new_n984_));
  INVX1    g0342(.A(\in2[60] ), .Y(new_n985_));
  INVX1    g0343(.A(\in2[61] ), .Y(new_n986_));
  AND2X1   g0344(.A(\in3[61] ), .B(new_n986_), .Y(new_n987_));
  NOR3X1   g0345(.A(new_n987_), .B(\in3[60] ), .C(new_n985_), .Y(new_n988_));
  AOI21X1  g0346(.A0(new_n967_), .A1(\in2[61] ), .B0(new_n988_), .Y(new_n989_));
  INVX1    g0347(.A(\in3[63] ), .Y(new_n990_));
  AND2X1   g0348(.A(\in3[63] ), .B(new_n963_), .Y(new_n991_));
  NOR3X1   g0349(.A(new_n991_), .B(\in3[62] ), .C(new_n962_), .Y(new_n992_));
  AOI21X1  g0350(.A0(new_n990_), .A1(\in2[63] ), .B0(new_n992_), .Y(new_n993_));
  OAI21X1  g0351(.A0(new_n989_), .A1(new_n965_), .B0(new_n993_), .Y(new_n994_));
  AOI21X1  g0352(.A0(new_n984_), .A1(new_n978_), .B0(new_n994_), .Y(new_n995_));
  OAI21X1  g0353(.A0(new_n977_), .A1(new_n961_), .B0(new_n995_), .Y(new_n996_));
  INVX1    g0354(.A(\in2[66] ), .Y(new_n997_));
  INVX1    g0355(.A(\in2[67] ), .Y(new_n998_));
  AOI22X1  g0356(.A0(\in3[67] ), .A1(new_n998_), .B0(\in3[66] ), .B1(new_n997_), .Y(new_n999_));
  INVX1    g0357(.A(\in2[64] ), .Y(new_n1000_));
  INVX1    g0358(.A(\in2[65] ), .Y(new_n1001_));
  AOI22X1  g0359(.A0(\in3[65] ), .A1(new_n1001_), .B0(\in3[64] ), .B1(new_n1000_), .Y(new_n1002_));
  AND2X1   g0360(.A(new_n1002_), .B(new_n999_), .Y(new_n1003_));
  OR2X1    g0361(.A(\in3[67] ), .B(new_n998_), .Y(new_n1004_));
  AND2X1   g0362(.A(\in3[65] ), .B(new_n1001_), .Y(new_n1005_));
  NOR3X1   g0363(.A(new_n1005_), .B(\in3[64] ), .C(new_n1000_), .Y(new_n1006_));
  INVX1    g0364(.A(\in3[65] ), .Y(new_n1007_));
  INVX1    g0365(.A(\in3[66] ), .Y(new_n1008_));
  AOI22X1  g0366(.A0(new_n1008_), .A1(\in2[66] ), .B0(new_n1007_), .B1(\in2[65] ), .Y(new_n1009_));
  INVX1    g0367(.A(new_n1009_), .Y(new_n1010_));
  OAI21X1  g0368(.A0(new_n1010_), .A1(new_n1006_), .B0(new_n999_), .Y(new_n1011_));
  AND2X1   g0369(.A(new_n1011_), .B(new_n1004_), .Y(new_n1012_));
  INVX1    g0370(.A(new_n1012_), .Y(new_n1013_));
  AOI21X1  g0371(.A0(new_n1003_), .A1(new_n996_), .B0(new_n1013_), .Y(new_n1014_));
  INVX1    g0372(.A(\in2[70] ), .Y(new_n1015_));
  INVX1    g0373(.A(\in2[71] ), .Y(new_n1016_));
  AOI22X1  g0374(.A0(\in3[71] ), .A1(new_n1016_), .B0(\in3[70] ), .B1(new_n1015_), .Y(new_n1017_));
  INVX1    g0375(.A(\in2[68] ), .Y(new_n1018_));
  INVX1    g0376(.A(\in2[69] ), .Y(new_n1019_));
  AOI22X1  g0377(.A0(\in3[69] ), .A1(new_n1019_), .B0(\in3[68] ), .B1(new_n1018_), .Y(new_n1020_));
  AND2X1   g0378(.A(new_n1020_), .B(new_n1017_), .Y(new_n1021_));
  INVX1    g0379(.A(new_n1021_), .Y(new_n1022_));
  AND2X1   g0380(.A(\in3[69] ), .B(new_n1019_), .Y(new_n1023_));
  NOR3X1   g0381(.A(new_n1023_), .B(\in3[68] ), .C(new_n1018_), .Y(new_n1024_));
  INVX1    g0382(.A(\in3[69] ), .Y(new_n1025_));
  AND2X1   g0383(.A(new_n1025_), .B(\in2[69] ), .Y(new_n1026_));
  OAI21X1  g0384(.A0(new_n1026_), .A1(new_n1024_), .B0(new_n1017_), .Y(new_n1027_));
  INVX1    g0385(.A(\in3[71] ), .Y(new_n1028_));
  AND2X1   g0386(.A(\in3[71] ), .B(new_n1016_), .Y(new_n1029_));
  NOR3X1   g0387(.A(new_n1029_), .B(\in3[70] ), .C(new_n1015_), .Y(new_n1030_));
  AOI21X1  g0388(.A0(new_n1028_), .A1(\in2[71] ), .B0(new_n1030_), .Y(new_n1031_));
  AND2X1   g0389(.A(new_n1031_), .B(new_n1027_), .Y(new_n1032_));
  OAI21X1  g0390(.A0(new_n1022_), .A1(new_n1014_), .B0(new_n1032_), .Y(new_n1033_));
  INVX1    g0391(.A(\in2[74] ), .Y(new_n1034_));
  INVX1    g0392(.A(\in2[75] ), .Y(new_n1035_));
  AOI22X1  g0393(.A0(\in3[75] ), .A1(new_n1035_), .B0(\in3[74] ), .B1(new_n1034_), .Y(new_n1036_));
  INVX1    g0394(.A(\in2[72] ), .Y(new_n1037_));
  INVX1    g0395(.A(\in2[73] ), .Y(new_n1038_));
  AOI22X1  g0396(.A0(\in3[73] ), .A1(new_n1038_), .B0(\in3[72] ), .B1(new_n1037_), .Y(new_n1039_));
  AND2X1   g0397(.A(new_n1039_), .B(new_n1036_), .Y(new_n1040_));
  OR2X1    g0398(.A(\in3[75] ), .B(new_n1035_), .Y(new_n1041_));
  AND2X1   g0399(.A(\in3[73] ), .B(new_n1038_), .Y(new_n1042_));
  NOR3X1   g0400(.A(new_n1042_), .B(\in3[72] ), .C(new_n1037_), .Y(new_n1043_));
  INVX1    g0401(.A(\in3[73] ), .Y(new_n1044_));
  INVX1    g0402(.A(\in3[74] ), .Y(new_n1045_));
  AOI22X1  g0403(.A0(new_n1045_), .A1(\in2[74] ), .B0(new_n1044_), .B1(\in2[73] ), .Y(new_n1046_));
  INVX1    g0404(.A(new_n1046_), .Y(new_n1047_));
  OAI21X1  g0405(.A0(new_n1047_), .A1(new_n1043_), .B0(new_n1036_), .Y(new_n1048_));
  AND2X1   g0406(.A(new_n1048_), .B(new_n1041_), .Y(new_n1049_));
  INVX1    g0407(.A(new_n1049_), .Y(new_n1050_));
  AOI21X1  g0408(.A0(new_n1040_), .A1(new_n1033_), .B0(new_n1050_), .Y(new_n1051_));
  INVX1    g0409(.A(\in2[78] ), .Y(new_n1052_));
  INVX1    g0410(.A(\in2[79] ), .Y(new_n1053_));
  AOI22X1  g0411(.A0(\in3[79] ), .A1(new_n1053_), .B0(\in3[78] ), .B1(new_n1052_), .Y(new_n1054_));
  INVX1    g0412(.A(\in2[76] ), .Y(new_n1055_));
  INVX1    g0413(.A(\in2[77] ), .Y(new_n1056_));
  AOI22X1  g0414(.A0(\in3[77] ), .A1(new_n1056_), .B0(\in3[76] ), .B1(new_n1055_), .Y(new_n1057_));
  AND2X1   g0415(.A(new_n1057_), .B(new_n1054_), .Y(new_n1058_));
  INVX1    g0416(.A(new_n1058_), .Y(new_n1059_));
  AND2X1   g0417(.A(\in3[77] ), .B(new_n1056_), .Y(new_n1060_));
  NOR3X1   g0418(.A(new_n1060_), .B(\in3[76] ), .C(new_n1055_), .Y(new_n1061_));
  INVX1    g0419(.A(\in3[77] ), .Y(new_n1062_));
  AND2X1   g0420(.A(new_n1062_), .B(\in2[77] ), .Y(new_n1063_));
  OAI21X1  g0421(.A0(new_n1063_), .A1(new_n1061_), .B0(new_n1054_), .Y(new_n1064_));
  INVX1    g0422(.A(\in3[79] ), .Y(new_n1065_));
  AND2X1   g0423(.A(\in3[79] ), .B(new_n1053_), .Y(new_n1066_));
  NOR3X1   g0424(.A(new_n1066_), .B(\in3[78] ), .C(new_n1052_), .Y(new_n1067_));
  AOI21X1  g0425(.A0(new_n1065_), .A1(\in2[79] ), .B0(new_n1067_), .Y(new_n1068_));
  AND2X1   g0426(.A(new_n1068_), .B(new_n1064_), .Y(new_n1069_));
  OAI21X1  g0427(.A0(new_n1059_), .A1(new_n1051_), .B0(new_n1069_), .Y(new_n1070_));
  INVX1    g0428(.A(\in2[82] ), .Y(new_n1071_));
  INVX1    g0429(.A(\in2[83] ), .Y(new_n1072_));
  AOI22X1  g0430(.A0(\in3[83] ), .A1(new_n1072_), .B0(\in3[82] ), .B1(new_n1071_), .Y(new_n1073_));
  INVX1    g0431(.A(\in2[80] ), .Y(new_n1074_));
  INVX1    g0432(.A(\in2[81] ), .Y(new_n1075_));
  AOI22X1  g0433(.A0(\in3[81] ), .A1(new_n1075_), .B0(\in3[80] ), .B1(new_n1074_), .Y(new_n1076_));
  AND2X1   g0434(.A(new_n1076_), .B(new_n1073_), .Y(new_n1077_));
  OR2X1    g0435(.A(\in3[83] ), .B(new_n1072_), .Y(new_n1078_));
  AND2X1   g0436(.A(\in3[81] ), .B(new_n1075_), .Y(new_n1079_));
  NOR3X1   g0437(.A(new_n1079_), .B(\in3[80] ), .C(new_n1074_), .Y(new_n1080_));
  INVX1    g0438(.A(\in3[81] ), .Y(new_n1081_));
  INVX1    g0439(.A(\in3[82] ), .Y(new_n1082_));
  AOI22X1  g0440(.A0(new_n1082_), .A1(\in2[82] ), .B0(new_n1081_), .B1(\in2[81] ), .Y(new_n1083_));
  INVX1    g0441(.A(new_n1083_), .Y(new_n1084_));
  OAI21X1  g0442(.A0(new_n1084_), .A1(new_n1080_), .B0(new_n1073_), .Y(new_n1085_));
  AND2X1   g0443(.A(new_n1085_), .B(new_n1078_), .Y(new_n1086_));
  INVX1    g0444(.A(new_n1086_), .Y(new_n1087_));
  AOI21X1  g0445(.A0(new_n1077_), .A1(new_n1070_), .B0(new_n1087_), .Y(new_n1088_));
  INVX1    g0446(.A(\in2[86] ), .Y(new_n1089_));
  INVX1    g0447(.A(\in2[87] ), .Y(new_n1090_));
  AOI22X1  g0448(.A0(\in3[87] ), .A1(new_n1090_), .B0(\in3[86] ), .B1(new_n1089_), .Y(new_n1091_));
  INVX1    g0449(.A(\in2[84] ), .Y(new_n1092_));
  INVX1    g0450(.A(\in2[85] ), .Y(new_n1093_));
  AOI22X1  g0451(.A0(\in3[85] ), .A1(new_n1093_), .B0(\in3[84] ), .B1(new_n1092_), .Y(new_n1094_));
  AND2X1   g0452(.A(new_n1094_), .B(new_n1091_), .Y(new_n1095_));
  INVX1    g0453(.A(new_n1095_), .Y(new_n1096_));
  AND2X1   g0454(.A(\in3[85] ), .B(new_n1093_), .Y(new_n1097_));
  NOR3X1   g0455(.A(new_n1097_), .B(\in3[84] ), .C(new_n1092_), .Y(new_n1098_));
  INVX1    g0456(.A(\in3[85] ), .Y(new_n1099_));
  AND2X1   g0457(.A(new_n1099_), .B(\in2[85] ), .Y(new_n1100_));
  OAI21X1  g0458(.A0(new_n1100_), .A1(new_n1098_), .B0(new_n1091_), .Y(new_n1101_));
  INVX1    g0459(.A(\in3[87] ), .Y(new_n1102_));
  AND2X1   g0460(.A(\in3[87] ), .B(new_n1090_), .Y(new_n1103_));
  NOR3X1   g0461(.A(new_n1103_), .B(\in3[86] ), .C(new_n1089_), .Y(new_n1104_));
  AOI21X1  g0462(.A0(new_n1102_), .A1(\in2[87] ), .B0(new_n1104_), .Y(new_n1105_));
  AND2X1   g0463(.A(new_n1105_), .B(new_n1101_), .Y(new_n1106_));
  OAI21X1  g0464(.A0(new_n1096_), .A1(new_n1088_), .B0(new_n1106_), .Y(new_n1107_));
  INVX1    g0465(.A(\in2[90] ), .Y(new_n1108_));
  INVX1    g0466(.A(\in2[91] ), .Y(new_n1109_));
  AOI22X1  g0467(.A0(\in3[91] ), .A1(new_n1109_), .B0(\in3[90] ), .B1(new_n1108_), .Y(new_n1110_));
  INVX1    g0468(.A(\in2[88] ), .Y(new_n1111_));
  INVX1    g0469(.A(\in2[89] ), .Y(new_n1112_));
  AOI22X1  g0470(.A0(\in3[89] ), .A1(new_n1112_), .B0(\in3[88] ), .B1(new_n1111_), .Y(new_n1113_));
  AND2X1   g0471(.A(new_n1113_), .B(new_n1110_), .Y(new_n1114_));
  OR2X1    g0472(.A(\in3[91] ), .B(new_n1109_), .Y(new_n1115_));
  AND2X1   g0473(.A(\in3[89] ), .B(new_n1112_), .Y(new_n1116_));
  NOR3X1   g0474(.A(new_n1116_), .B(\in3[88] ), .C(new_n1111_), .Y(new_n1117_));
  INVX1    g0475(.A(\in3[89] ), .Y(new_n1118_));
  INVX1    g0476(.A(\in3[90] ), .Y(new_n1119_));
  AOI22X1  g0477(.A0(new_n1119_), .A1(\in2[90] ), .B0(new_n1118_), .B1(\in2[89] ), .Y(new_n1120_));
  INVX1    g0478(.A(new_n1120_), .Y(new_n1121_));
  OAI21X1  g0479(.A0(new_n1121_), .A1(new_n1117_), .B0(new_n1110_), .Y(new_n1122_));
  AND2X1   g0480(.A(new_n1122_), .B(new_n1115_), .Y(new_n1123_));
  INVX1    g0481(.A(new_n1123_), .Y(new_n1124_));
  AOI21X1  g0482(.A0(new_n1114_), .A1(new_n1107_), .B0(new_n1124_), .Y(new_n1125_));
  INVX1    g0483(.A(\in2[94] ), .Y(new_n1126_));
  INVX1    g0484(.A(\in2[95] ), .Y(new_n1127_));
  AOI22X1  g0485(.A0(\in3[95] ), .A1(new_n1127_), .B0(\in3[94] ), .B1(new_n1126_), .Y(new_n1128_));
  INVX1    g0486(.A(\in2[92] ), .Y(new_n1129_));
  INVX1    g0487(.A(\in2[93] ), .Y(new_n1130_));
  AOI22X1  g0488(.A0(\in3[93] ), .A1(new_n1130_), .B0(\in3[92] ), .B1(new_n1129_), .Y(new_n1131_));
  AND2X1   g0489(.A(new_n1131_), .B(new_n1128_), .Y(new_n1132_));
  INVX1    g0490(.A(new_n1132_), .Y(new_n1133_));
  AND2X1   g0491(.A(\in3[93] ), .B(new_n1130_), .Y(new_n1134_));
  NOR3X1   g0492(.A(new_n1134_), .B(\in3[92] ), .C(new_n1129_), .Y(new_n1135_));
  INVX1    g0493(.A(\in3[93] ), .Y(new_n1136_));
  AND2X1   g0494(.A(new_n1136_), .B(\in2[93] ), .Y(new_n1137_));
  OAI21X1  g0495(.A0(new_n1137_), .A1(new_n1135_), .B0(new_n1128_), .Y(new_n1138_));
  INVX1    g0496(.A(\in3[95] ), .Y(new_n1139_));
  AND2X1   g0497(.A(\in3[95] ), .B(new_n1127_), .Y(new_n1140_));
  NOR3X1   g0498(.A(new_n1140_), .B(\in3[94] ), .C(new_n1126_), .Y(new_n1141_));
  AOI21X1  g0499(.A0(new_n1139_), .A1(\in2[95] ), .B0(new_n1141_), .Y(new_n1142_));
  AND2X1   g0500(.A(new_n1142_), .B(new_n1138_), .Y(new_n1143_));
  OAI21X1  g0501(.A0(new_n1133_), .A1(new_n1125_), .B0(new_n1143_), .Y(new_n1144_));
  INVX1    g0502(.A(\in2[98] ), .Y(new_n1145_));
  INVX1    g0503(.A(\in2[99] ), .Y(new_n1146_));
  AOI22X1  g0504(.A0(\in3[99] ), .A1(new_n1146_), .B0(\in3[98] ), .B1(new_n1145_), .Y(new_n1147_));
  INVX1    g0505(.A(\in2[96] ), .Y(new_n1148_));
  INVX1    g0506(.A(\in2[97] ), .Y(new_n1149_));
  AOI22X1  g0507(.A0(\in3[97] ), .A1(new_n1149_), .B0(\in3[96] ), .B1(new_n1148_), .Y(new_n1150_));
  AND2X1   g0508(.A(new_n1150_), .B(new_n1147_), .Y(new_n1151_));
  OR2X1    g0509(.A(\in3[99] ), .B(new_n1146_), .Y(new_n1152_));
  AND2X1   g0510(.A(\in3[97] ), .B(new_n1149_), .Y(new_n1153_));
  NOR3X1   g0511(.A(new_n1153_), .B(\in3[96] ), .C(new_n1148_), .Y(new_n1154_));
  INVX1    g0512(.A(\in3[97] ), .Y(new_n1155_));
  INVX1    g0513(.A(\in3[98] ), .Y(new_n1156_));
  AOI22X1  g0514(.A0(new_n1156_), .A1(\in2[98] ), .B0(new_n1155_), .B1(\in2[97] ), .Y(new_n1157_));
  INVX1    g0515(.A(new_n1157_), .Y(new_n1158_));
  OAI21X1  g0516(.A0(new_n1158_), .A1(new_n1154_), .B0(new_n1147_), .Y(new_n1159_));
  AND2X1   g0517(.A(new_n1159_), .B(new_n1152_), .Y(new_n1160_));
  INVX1    g0518(.A(new_n1160_), .Y(new_n1161_));
  AOI21X1  g0519(.A0(new_n1151_), .A1(new_n1144_), .B0(new_n1161_), .Y(new_n1162_));
  INVX1    g0520(.A(\in2[102] ), .Y(new_n1163_));
  INVX1    g0521(.A(\in2[103] ), .Y(new_n1164_));
  AOI22X1  g0522(.A0(\in3[103] ), .A1(new_n1164_), .B0(\in3[102] ), .B1(new_n1163_), .Y(new_n1165_));
  INVX1    g0523(.A(\in2[100] ), .Y(new_n1166_));
  INVX1    g0524(.A(\in2[101] ), .Y(new_n1167_));
  AOI22X1  g0525(.A0(\in3[101] ), .A1(new_n1167_), .B0(\in3[100] ), .B1(new_n1166_), .Y(new_n1168_));
  AND2X1   g0526(.A(new_n1168_), .B(new_n1165_), .Y(new_n1169_));
  INVX1    g0527(.A(new_n1169_), .Y(new_n1170_));
  AND2X1   g0528(.A(\in3[101] ), .B(new_n1167_), .Y(new_n1171_));
  NOR3X1   g0529(.A(new_n1171_), .B(\in3[100] ), .C(new_n1166_), .Y(new_n1172_));
  INVX1    g0530(.A(\in3[101] ), .Y(new_n1173_));
  AND2X1   g0531(.A(new_n1173_), .B(\in2[101] ), .Y(new_n1174_));
  OAI21X1  g0532(.A0(new_n1174_), .A1(new_n1172_), .B0(new_n1165_), .Y(new_n1175_));
  INVX1    g0533(.A(\in3[103] ), .Y(new_n1176_));
  AND2X1   g0534(.A(\in3[103] ), .B(new_n1164_), .Y(new_n1177_));
  NOR3X1   g0535(.A(new_n1177_), .B(\in3[102] ), .C(new_n1163_), .Y(new_n1178_));
  AOI21X1  g0536(.A0(new_n1176_), .A1(\in2[103] ), .B0(new_n1178_), .Y(new_n1179_));
  AND2X1   g0537(.A(new_n1179_), .B(new_n1175_), .Y(new_n1180_));
  OAI21X1  g0538(.A0(new_n1170_), .A1(new_n1162_), .B0(new_n1180_), .Y(new_n1181_));
  INVX1    g0539(.A(\in2[106] ), .Y(new_n1182_));
  INVX1    g0540(.A(\in2[107] ), .Y(new_n1183_));
  AOI22X1  g0541(.A0(\in3[107] ), .A1(new_n1183_), .B0(\in3[106] ), .B1(new_n1182_), .Y(new_n1184_));
  INVX1    g0542(.A(\in2[104] ), .Y(new_n1185_));
  INVX1    g0543(.A(\in2[105] ), .Y(new_n1186_));
  AOI22X1  g0544(.A0(\in3[105] ), .A1(new_n1186_), .B0(\in3[104] ), .B1(new_n1185_), .Y(new_n1187_));
  AND2X1   g0545(.A(new_n1187_), .B(new_n1184_), .Y(new_n1188_));
  OR2X1    g0546(.A(\in3[107] ), .B(new_n1183_), .Y(new_n1189_));
  AND2X1   g0547(.A(\in3[105] ), .B(new_n1186_), .Y(new_n1190_));
  NOR3X1   g0548(.A(new_n1190_), .B(\in3[104] ), .C(new_n1185_), .Y(new_n1191_));
  INVX1    g0549(.A(\in3[105] ), .Y(new_n1192_));
  INVX1    g0550(.A(\in3[106] ), .Y(new_n1193_));
  AOI22X1  g0551(.A0(new_n1193_), .A1(\in2[106] ), .B0(new_n1192_), .B1(\in2[105] ), .Y(new_n1194_));
  INVX1    g0552(.A(new_n1194_), .Y(new_n1195_));
  OAI21X1  g0553(.A0(new_n1195_), .A1(new_n1191_), .B0(new_n1184_), .Y(new_n1196_));
  AND2X1   g0554(.A(new_n1196_), .B(new_n1189_), .Y(new_n1197_));
  INVX1    g0555(.A(new_n1197_), .Y(new_n1198_));
  AOI21X1  g0556(.A0(new_n1188_), .A1(new_n1181_), .B0(new_n1198_), .Y(new_n1199_));
  INVX1    g0557(.A(\in2[110] ), .Y(new_n1200_));
  INVX1    g0558(.A(\in2[111] ), .Y(new_n1201_));
  AOI22X1  g0559(.A0(\in3[111] ), .A1(new_n1201_), .B0(\in3[110] ), .B1(new_n1200_), .Y(new_n1202_));
  INVX1    g0560(.A(\in2[108] ), .Y(new_n1203_));
  INVX1    g0561(.A(\in2[109] ), .Y(new_n1204_));
  AOI22X1  g0562(.A0(\in3[109] ), .A1(new_n1204_), .B0(\in3[108] ), .B1(new_n1203_), .Y(new_n1205_));
  AND2X1   g0563(.A(new_n1205_), .B(new_n1202_), .Y(new_n1206_));
  INVX1    g0564(.A(new_n1206_), .Y(new_n1207_));
  AND2X1   g0565(.A(\in3[109] ), .B(new_n1204_), .Y(new_n1208_));
  NOR3X1   g0566(.A(new_n1208_), .B(\in3[108] ), .C(new_n1203_), .Y(new_n1209_));
  INVX1    g0567(.A(\in3[109] ), .Y(new_n1210_));
  AND2X1   g0568(.A(new_n1210_), .B(\in2[109] ), .Y(new_n1211_));
  OAI21X1  g0569(.A0(new_n1211_), .A1(new_n1209_), .B0(new_n1202_), .Y(new_n1212_));
  INVX1    g0570(.A(\in3[111] ), .Y(new_n1213_));
  AND2X1   g0571(.A(\in3[111] ), .B(new_n1201_), .Y(new_n1214_));
  NOR3X1   g0572(.A(new_n1214_), .B(\in3[110] ), .C(new_n1200_), .Y(new_n1215_));
  AOI21X1  g0573(.A0(new_n1213_), .A1(\in2[111] ), .B0(new_n1215_), .Y(new_n1216_));
  AND2X1   g0574(.A(new_n1216_), .B(new_n1212_), .Y(new_n1217_));
  OAI21X1  g0575(.A0(new_n1207_), .A1(new_n1199_), .B0(new_n1217_), .Y(new_n1218_));
  INVX1    g0576(.A(\in2[114] ), .Y(new_n1219_));
  INVX1    g0577(.A(\in2[115] ), .Y(new_n1220_));
  AOI22X1  g0578(.A0(\in3[115] ), .A1(new_n1220_), .B0(\in3[114] ), .B1(new_n1219_), .Y(new_n1221_));
  INVX1    g0579(.A(\in2[112] ), .Y(new_n1222_));
  INVX1    g0580(.A(\in2[113] ), .Y(new_n1223_));
  AOI22X1  g0581(.A0(\in3[113] ), .A1(new_n1223_), .B0(\in3[112] ), .B1(new_n1222_), .Y(new_n1224_));
  AND2X1   g0582(.A(new_n1224_), .B(new_n1221_), .Y(new_n1225_));
  OR2X1    g0583(.A(\in3[115] ), .B(new_n1220_), .Y(new_n1226_));
  AND2X1   g0584(.A(\in3[113] ), .B(new_n1223_), .Y(new_n1227_));
  NOR3X1   g0585(.A(new_n1227_), .B(\in3[112] ), .C(new_n1222_), .Y(new_n1228_));
  INVX1    g0586(.A(\in3[113] ), .Y(new_n1229_));
  INVX1    g0587(.A(\in3[114] ), .Y(new_n1230_));
  AOI22X1  g0588(.A0(new_n1230_), .A1(\in2[114] ), .B0(new_n1229_), .B1(\in2[113] ), .Y(new_n1231_));
  INVX1    g0589(.A(new_n1231_), .Y(new_n1232_));
  OAI21X1  g0590(.A0(new_n1232_), .A1(new_n1228_), .B0(new_n1221_), .Y(new_n1233_));
  AND2X1   g0591(.A(new_n1233_), .B(new_n1226_), .Y(new_n1234_));
  INVX1    g0592(.A(new_n1234_), .Y(new_n1235_));
  AOI21X1  g0593(.A0(new_n1225_), .A1(new_n1218_), .B0(new_n1235_), .Y(new_n1236_));
  INVX1    g0594(.A(\in2[118] ), .Y(new_n1237_));
  INVX1    g0595(.A(\in2[119] ), .Y(new_n1238_));
  AOI22X1  g0596(.A0(\in3[119] ), .A1(new_n1238_), .B0(\in3[118] ), .B1(new_n1237_), .Y(new_n1239_));
  INVX1    g0597(.A(\in2[116] ), .Y(new_n1240_));
  INVX1    g0598(.A(\in2[117] ), .Y(new_n1241_));
  AOI22X1  g0599(.A0(\in3[117] ), .A1(new_n1241_), .B0(\in3[116] ), .B1(new_n1240_), .Y(new_n1242_));
  AND2X1   g0600(.A(new_n1242_), .B(new_n1239_), .Y(new_n1243_));
  INVX1    g0601(.A(new_n1243_), .Y(new_n1244_));
  AND2X1   g0602(.A(\in3[117] ), .B(new_n1241_), .Y(new_n1245_));
  NOR3X1   g0603(.A(new_n1245_), .B(\in3[116] ), .C(new_n1240_), .Y(new_n1246_));
  INVX1    g0604(.A(\in3[117] ), .Y(new_n1247_));
  AND2X1   g0605(.A(new_n1247_), .B(\in2[117] ), .Y(new_n1248_));
  OAI21X1  g0606(.A0(new_n1248_), .A1(new_n1246_), .B0(new_n1239_), .Y(new_n1249_));
  INVX1    g0607(.A(\in3[119] ), .Y(new_n1250_));
  AND2X1   g0608(.A(\in3[119] ), .B(new_n1238_), .Y(new_n1251_));
  NOR3X1   g0609(.A(new_n1251_), .B(\in3[118] ), .C(new_n1237_), .Y(new_n1252_));
  AOI21X1  g0610(.A0(new_n1250_), .A1(\in2[119] ), .B0(new_n1252_), .Y(new_n1253_));
  AND2X1   g0611(.A(new_n1253_), .B(new_n1249_), .Y(new_n1254_));
  OAI21X1  g0612(.A0(new_n1244_), .A1(new_n1236_), .B0(new_n1254_), .Y(new_n1255_));
  INVX1    g0613(.A(\in2[122] ), .Y(new_n1256_));
  INVX1    g0614(.A(\in2[123] ), .Y(new_n1257_));
  AOI22X1  g0615(.A0(\in3[123] ), .A1(new_n1257_), .B0(\in3[122] ), .B1(new_n1256_), .Y(new_n1258_));
  INVX1    g0616(.A(\in2[120] ), .Y(new_n1259_));
  INVX1    g0617(.A(\in2[121] ), .Y(new_n1260_));
  AOI22X1  g0618(.A0(\in3[121] ), .A1(new_n1260_), .B0(\in3[120] ), .B1(new_n1259_), .Y(new_n1261_));
  AND2X1   g0619(.A(new_n1261_), .B(new_n1258_), .Y(new_n1262_));
  OR2X1    g0620(.A(\in3[123] ), .B(new_n1257_), .Y(new_n1263_));
  AND2X1   g0621(.A(\in3[121] ), .B(new_n1260_), .Y(new_n1264_));
  NOR3X1   g0622(.A(new_n1264_), .B(\in3[120] ), .C(new_n1259_), .Y(new_n1265_));
  INVX1    g0623(.A(\in3[121] ), .Y(new_n1266_));
  INVX1    g0624(.A(\in3[122] ), .Y(new_n1267_));
  AOI22X1  g0625(.A0(new_n1267_), .A1(\in2[122] ), .B0(new_n1266_), .B1(\in2[121] ), .Y(new_n1268_));
  INVX1    g0626(.A(new_n1268_), .Y(new_n1269_));
  OAI21X1  g0627(.A0(new_n1269_), .A1(new_n1265_), .B0(new_n1258_), .Y(new_n1270_));
  AND2X1   g0628(.A(new_n1270_), .B(new_n1263_), .Y(new_n1271_));
  INVX1    g0629(.A(new_n1271_), .Y(new_n1272_));
  AOI21X1  g0630(.A0(new_n1262_), .A1(new_n1255_), .B0(new_n1272_), .Y(new_n1273_));
  INVX1    g0631(.A(\in3[127] ), .Y(new_n1274_));
  AND2X1   g0632(.A(new_n1274_), .B(\in2[127] ), .Y(new_n1275_));
  INVX1    g0633(.A(\in2[125] ), .Y(new_n1276_));
  INVX1    g0634(.A(\in2[126] ), .Y(new_n1277_));
  AOI22X1  g0635(.A0(\in3[126] ), .A1(new_n1277_), .B0(\in3[125] ), .B1(new_n1276_), .Y(new_n1278_));
  INVX1    g0636(.A(\in2[124] ), .Y(new_n1279_));
  AOI22X1  g0637(.A0(new_n1274_), .A1(\in2[127] ), .B0(\in3[124] ), .B1(new_n1279_), .Y(new_n1280_));
  AND2X1   g0638(.A(new_n1280_), .B(new_n1278_), .Y(new_n1281_));
  INVX1    g0639(.A(new_n1281_), .Y(new_n1282_));
  INVX1    g0640(.A(\in3[126] ), .Y(new_n1283_));
  INVX1    g0641(.A(\in3[124] ), .Y(new_n1284_));
  INVX1    g0642(.A(\in3[125] ), .Y(new_n1285_));
  AOI22X1  g0643(.A0(new_n1285_), .A1(\in2[125] ), .B0(new_n1284_), .B1(\in2[124] ), .Y(new_n1286_));
  INVX1    g0644(.A(new_n1286_), .Y(new_n1287_));
  AOI22X1  g0645(.A0(new_n1287_), .A1(new_n1278_), .B0(new_n1283_), .B1(\in2[126] ), .Y(new_n1288_));
  OAI22X1  g0646(.A0(new_n1288_), .A1(new_n1275_), .B0(new_n1282_), .B1(new_n1273_), .Y(new_n1289_));
  INVX1    g0647(.A(\in2[127] ), .Y(new_n1290_));
  AND2X1   g0648(.A(\in3[127] ), .B(new_n1290_), .Y(new_n1291_));
  NOR3X1   g0649(.A(new_n1291_), .B(new_n1289_), .C(new_n643_), .Y(new_n1292_));
  INVX1    g0650(.A(new_n645_), .Y(new_n1293_));
  INVX1    g0651(.A(new_n650_), .Y(new_n1294_));
  INVX1    g0652(.A(new_n655_), .Y(new_n1295_));
  INVX1    g0653(.A(\in3[25] ), .Y(new_n1296_));
  INVX1    g0654(.A(\in2[25] ), .Y(new_n1297_));
  INVX1    g0655(.A(\in3[24] ), .Y(new_n1298_));
  OAI21X1  g0656(.A0(new_n835_), .A1(\in2[24] ), .B0(new_n1298_), .Y(new_n1299_));
  OR2X1    g0657(.A(new_n817_), .B(new_n659_), .Y(new_n1300_));
  NAND3X1  g0658(.A(new_n1300_), .B(new_n1299_), .C(new_n1297_), .Y(new_n1301_));
  AOI21X1  g0659(.A0(new_n1300_), .A1(new_n1299_), .B0(new_n1297_), .Y(new_n1302_));
  AOI21X1  g0660(.A0(new_n1301_), .A1(new_n1296_), .B0(new_n1302_), .Y(new_n1303_));
  INVX1    g0661(.A(new_n841_), .Y(new_n1304_));
  OAI21X1  g0662(.A0(new_n1303_), .A1(new_n657_), .B0(new_n1304_), .Y(new_n1305_));
  AOI21X1  g0663(.A0(new_n1305_), .A1(new_n1295_), .B0(new_n844_), .Y(new_n1306_));
  INVX1    g0664(.A(new_n848_), .Y(new_n1307_));
  OAI21X1  g0665(.A0(new_n1306_), .A1(new_n652_), .B0(new_n1307_), .Y(new_n1308_));
  AOI21X1  g0666(.A0(new_n1308_), .A1(new_n1294_), .B0(new_n851_), .Y(new_n1309_));
  INVX1    g0667(.A(new_n855_), .Y(new_n1310_));
  OAI21X1  g0668(.A0(new_n1309_), .A1(new_n647_), .B0(new_n1310_), .Y(new_n1311_));
  AOI21X1  g0669(.A0(new_n1311_), .A1(new_n1293_), .B0(new_n858_), .Y(new_n1312_));
  INVX1    g0670(.A(new_n875_), .Y(new_n1313_));
  OAI21X1  g0671(.A0(new_n1313_), .A1(new_n1312_), .B0(new_n893_), .Y(new_n1314_));
  INVX1    g0672(.A(new_n929_), .Y(new_n1315_));
  AOI21X1  g0673(.A0(new_n910_), .A1(new_n1314_), .B0(new_n1315_), .Y(new_n1316_));
  INVX1    g0674(.A(new_n945_), .Y(new_n1317_));
  OAI21X1  g0675(.A0(new_n1317_), .A1(new_n1316_), .B0(new_n959_), .Y(new_n1318_));
  INVX1    g0676(.A(new_n995_), .Y(new_n1319_));
  AOI21X1  g0677(.A0(new_n976_), .A1(new_n1318_), .B0(new_n1319_), .Y(new_n1320_));
  INVX1    g0678(.A(new_n1003_), .Y(new_n1321_));
  OAI21X1  g0679(.A0(new_n1321_), .A1(new_n1320_), .B0(new_n1012_), .Y(new_n1322_));
  INVX1    g0680(.A(new_n1032_), .Y(new_n1323_));
  AOI21X1  g0681(.A0(new_n1021_), .A1(new_n1322_), .B0(new_n1323_), .Y(new_n1324_));
  INVX1    g0682(.A(new_n1040_), .Y(new_n1325_));
  OAI21X1  g0683(.A0(new_n1325_), .A1(new_n1324_), .B0(new_n1049_), .Y(new_n1326_));
  INVX1    g0684(.A(new_n1069_), .Y(new_n1327_));
  AOI21X1  g0685(.A0(new_n1058_), .A1(new_n1326_), .B0(new_n1327_), .Y(new_n1328_));
  INVX1    g0686(.A(new_n1077_), .Y(new_n1329_));
  OAI21X1  g0687(.A0(new_n1329_), .A1(new_n1328_), .B0(new_n1086_), .Y(new_n1330_));
  INVX1    g0688(.A(new_n1106_), .Y(new_n1331_));
  AOI21X1  g0689(.A0(new_n1095_), .A1(new_n1330_), .B0(new_n1331_), .Y(new_n1332_));
  INVX1    g0690(.A(new_n1114_), .Y(new_n1333_));
  OAI21X1  g0691(.A0(new_n1333_), .A1(new_n1332_), .B0(new_n1123_), .Y(new_n1334_));
  INVX1    g0692(.A(new_n1143_), .Y(new_n1335_));
  AOI21X1  g0693(.A0(new_n1132_), .A1(new_n1334_), .B0(new_n1335_), .Y(new_n1336_));
  INVX1    g0694(.A(new_n1151_), .Y(new_n1337_));
  OAI21X1  g0695(.A0(new_n1337_), .A1(new_n1336_), .B0(new_n1160_), .Y(new_n1338_));
  INVX1    g0696(.A(new_n1180_), .Y(new_n1339_));
  AOI21X1  g0697(.A0(new_n1169_), .A1(new_n1338_), .B0(new_n1339_), .Y(new_n1340_));
  INVX1    g0698(.A(new_n1188_), .Y(new_n1341_));
  OAI21X1  g0699(.A0(new_n1341_), .A1(new_n1340_), .B0(new_n1197_), .Y(new_n1342_));
  INVX1    g0700(.A(new_n1217_), .Y(new_n1343_));
  AOI21X1  g0701(.A0(new_n1206_), .A1(new_n1342_), .B0(new_n1343_), .Y(new_n1344_));
  INVX1    g0702(.A(new_n1225_), .Y(new_n1345_));
  OAI21X1  g0703(.A0(new_n1345_), .A1(new_n1344_), .B0(new_n1234_), .Y(new_n1346_));
  INVX1    g0704(.A(new_n1254_), .Y(new_n1347_));
  AOI21X1  g0705(.A0(new_n1243_), .A1(new_n1346_), .B0(new_n1347_), .Y(new_n1348_));
  INVX1    g0706(.A(new_n1262_), .Y(new_n1349_));
  OAI21X1  g0707(.A0(new_n1349_), .A1(new_n1348_), .B0(new_n1271_), .Y(new_n1350_));
  NOR2X1   g0708(.A(new_n1288_), .B(new_n1275_), .Y(new_n1351_));
  AOI21X1  g0709(.A0(new_n1281_), .A1(new_n1350_), .B0(new_n1351_), .Y(new_n1352_));
  INVX1    g0710(.A(new_n1291_), .Y(new_n1353_));
  AOI21X1  g0711(.A0(new_n1353_), .A1(new_n1352_), .B0(new_n706_), .Y(new_n1354_));
  OR2X1    g0712(.A(new_n1354_), .B(new_n1292_), .Y(new_n1355_));
  INVX1    g0713(.A(\in1[127] ), .Y(new_n1356_));
  INVX1    g0714(.A(\in0[31] ), .Y(new_n1357_));
  AND2X1   g0715(.A(\in1[31] ), .B(new_n1357_), .Y(new_n1358_));
  INVX1    g0716(.A(new_n1358_), .Y(new_n1359_));
  INVX1    g0717(.A(\in0[30] ), .Y(new_n1360_));
  AND2X1   g0718(.A(\in1[30] ), .B(new_n1360_), .Y(new_n1361_));
  INVX1    g0719(.A(\in0[29] ), .Y(new_n1362_));
  AND2X1   g0720(.A(\in1[29] ), .B(new_n1362_), .Y(new_n1363_));
  INVX1    g0721(.A(new_n1363_), .Y(new_n1364_));
  INVX1    g0722(.A(\in0[28] ), .Y(new_n1365_));
  AND2X1   g0723(.A(\in1[28] ), .B(new_n1365_), .Y(new_n1366_));
  INVX1    g0724(.A(\in0[27] ), .Y(new_n1367_));
  AND2X1   g0725(.A(\in1[27] ), .B(new_n1367_), .Y(new_n1368_));
  INVX1    g0726(.A(new_n1368_), .Y(new_n1369_));
  INVX1    g0727(.A(\in0[26] ), .Y(new_n1370_));
  AND2X1   g0728(.A(\in1[26] ), .B(new_n1370_), .Y(new_n1371_));
  INVX1    g0729(.A(\in1[25] ), .Y(new_n1372_));
  INVX1    g0730(.A(\in0[25] ), .Y(new_n1373_));
  INVX1    g0731(.A(\in1[24] ), .Y(new_n1374_));
  INVX1    g0732(.A(\in0[23] ), .Y(new_n1375_));
  AND2X1   g0733(.A(\in1[23] ), .B(new_n1375_), .Y(new_n1376_));
  INVX1    g0734(.A(\in0[22] ), .Y(new_n1377_));
  AND2X1   g0735(.A(\in1[22] ), .B(new_n1377_), .Y(new_n1378_));
  INVX1    g0736(.A(new_n1378_), .Y(new_n1379_));
  INVX1    g0737(.A(\in0[21] ), .Y(new_n1380_));
  AND2X1   g0738(.A(\in1[21] ), .B(new_n1380_), .Y(new_n1381_));
  INVX1    g0739(.A(\in0[20] ), .Y(new_n1382_));
  AND2X1   g0740(.A(\in1[20] ), .B(new_n1382_), .Y(new_n1383_));
  INVX1    g0741(.A(new_n1383_), .Y(new_n1384_));
  INVX1    g0742(.A(\in0[19] ), .Y(new_n1385_));
  AND2X1   g0743(.A(\in1[19] ), .B(new_n1385_), .Y(new_n1386_));
  INVX1    g0744(.A(\in0[18] ), .Y(new_n1387_));
  AND2X1   g0745(.A(\in1[18] ), .B(new_n1387_), .Y(new_n1388_));
  INVX1    g0746(.A(new_n1388_), .Y(new_n1389_));
  INVX1    g0747(.A(\in0[16] ), .Y(new_n1390_));
  INVX1    g0748(.A(\in0[15] ), .Y(new_n1391_));
  AND2X1   g0749(.A(\in1[15] ), .B(new_n1391_), .Y(new_n1392_));
  INVX1    g0750(.A(new_n1392_), .Y(new_n1393_));
  INVX1    g0751(.A(\in0[14] ), .Y(new_n1394_));
  AND2X1   g0752(.A(\in1[14] ), .B(new_n1394_), .Y(new_n1395_));
  INVX1    g0753(.A(\in0[13] ), .Y(new_n1396_));
  AND2X1   g0754(.A(\in1[13] ), .B(new_n1396_), .Y(new_n1397_));
  INVX1    g0755(.A(new_n1397_), .Y(new_n1398_));
  INVX1    g0756(.A(\in0[12] ), .Y(new_n1399_));
  AND2X1   g0757(.A(\in1[12] ), .B(new_n1399_), .Y(new_n1400_));
  INVX1    g0758(.A(\in0[11] ), .Y(new_n1401_));
  AND2X1   g0759(.A(\in1[11] ), .B(new_n1401_), .Y(new_n1402_));
  INVX1    g0760(.A(new_n1402_), .Y(new_n1403_));
  INVX1    g0761(.A(\in0[10] ), .Y(new_n1404_));
  AND2X1   g0762(.A(\in1[10] ), .B(new_n1404_), .Y(new_n1405_));
  INVX1    g0763(.A(\in1[9] ), .Y(new_n1406_));
  INVX1    g0764(.A(\in0[9] ), .Y(new_n1407_));
  INVX1    g0765(.A(\in1[8] ), .Y(new_n1408_));
  INVX1    g0766(.A(\in0[7] ), .Y(new_n1409_));
  AND2X1   g0767(.A(\in1[7] ), .B(new_n1409_), .Y(new_n1410_));
  INVX1    g0768(.A(\in0[6] ), .Y(new_n1411_));
  AND2X1   g0769(.A(\in1[6] ), .B(new_n1411_), .Y(new_n1412_));
  INVX1    g0770(.A(new_n1412_), .Y(new_n1413_));
  INVX1    g0771(.A(\in0[4] ), .Y(new_n1414_));
  INVX1    g0772(.A(\in1[3] ), .Y(new_n1415_));
  OR2X1    g0773(.A(new_n1415_), .B(\in0[3] ), .Y(new_n1416_));
  INVX1    g0774(.A(\in0[2] ), .Y(new_n1417_));
  INVX1    g0775(.A(\in1[0] ), .Y(new_n1418_));
  INVX1    g0776(.A(\in1[1] ), .Y(new_n1419_));
  AOI22X1  g0777(.A0(new_n1419_), .A1(\in0[1] ), .B0(new_n1418_), .B1(\in0[0] ), .Y(new_n1420_));
  INVX1    g0778(.A(\in1[2] ), .Y(new_n1421_));
  OAI22X1  g0779(.A0(new_n1421_), .A1(\in0[2] ), .B0(new_n1419_), .B1(\in0[1] ), .Y(new_n1422_));
  OAI22X1  g0780(.A0(new_n1422_), .A1(new_n1420_), .B0(\in1[2] ), .B1(new_n1417_), .Y(new_n1423_));
  AND2X1   g0781(.A(new_n1415_), .B(\in0[3] ), .Y(new_n1424_));
  AOI21X1  g0782(.A0(new_n1423_), .A1(new_n1416_), .B0(new_n1424_), .Y(new_n1425_));
  AOI21X1  g0783(.A0(new_n1425_), .A1(new_n1414_), .B0(\in1[4] ), .Y(new_n1426_));
  INVX1    g0784(.A(\in0[3] ), .Y(new_n1427_));
  AND2X1   g0785(.A(\in1[3] ), .B(new_n1427_), .Y(new_n1428_));
  INVX1    g0786(.A(\in0[0] ), .Y(new_n1429_));
  INVX1    g0787(.A(\in0[1] ), .Y(new_n1430_));
  OAI22X1  g0788(.A0(\in1[1] ), .A1(new_n1430_), .B0(\in1[0] ), .B1(new_n1429_), .Y(new_n1431_));
  AOI22X1  g0789(.A0(\in1[2] ), .A1(new_n1417_), .B0(\in1[1] ), .B1(new_n1430_), .Y(new_n1432_));
  AOI22X1  g0790(.A0(new_n1432_), .A1(new_n1431_), .B0(new_n1421_), .B1(\in0[2] ), .Y(new_n1433_));
  OR2X1    g0791(.A(\in1[3] ), .B(new_n1427_), .Y(new_n1434_));
  OAI21X1  g0792(.A0(new_n1433_), .A1(new_n1428_), .B0(new_n1434_), .Y(new_n1435_));
  AND2X1   g0793(.A(new_n1435_), .B(\in0[4] ), .Y(new_n1436_));
  NOR3X1   g0794(.A(new_n1436_), .B(new_n1426_), .C(\in0[5] ), .Y(new_n1437_));
  OAI21X1  g0795(.A0(new_n1436_), .A1(new_n1426_), .B0(\in0[5] ), .Y(new_n1438_));
  OAI21X1  g0796(.A0(new_n1437_), .A1(\in1[5] ), .B0(new_n1438_), .Y(new_n1439_));
  INVX1    g0797(.A(\in1[6] ), .Y(new_n1440_));
  AND2X1   g0798(.A(new_n1440_), .B(\in0[6] ), .Y(new_n1441_));
  AOI21X1  g0799(.A0(new_n1439_), .A1(new_n1413_), .B0(new_n1441_), .Y(new_n1442_));
  INVX1    g0800(.A(\in1[7] ), .Y(new_n1443_));
  AND2X1   g0801(.A(new_n1443_), .B(\in0[7] ), .Y(new_n1444_));
  INVX1    g0802(.A(new_n1444_), .Y(new_n1445_));
  OAI21X1  g0803(.A0(new_n1442_), .A1(new_n1410_), .B0(new_n1445_), .Y(new_n1446_));
  OAI21X1  g0804(.A0(new_n1446_), .A1(\in0[8] ), .B0(new_n1408_), .Y(new_n1447_));
  INVX1    g0805(.A(\in0[8] ), .Y(new_n1448_));
  INVX1    g0806(.A(new_n1410_), .Y(new_n1449_));
  INVX1    g0807(.A(\in1[5] ), .Y(new_n1450_));
  INVX1    g0808(.A(\in0[5] ), .Y(new_n1451_));
  INVX1    g0809(.A(\in1[4] ), .Y(new_n1452_));
  OAI21X1  g0810(.A0(new_n1435_), .A1(\in0[4] ), .B0(new_n1452_), .Y(new_n1453_));
  OR2X1    g0811(.A(new_n1425_), .B(new_n1414_), .Y(new_n1454_));
  NAND3X1  g0812(.A(new_n1454_), .B(new_n1453_), .C(new_n1451_), .Y(new_n1455_));
  AOI21X1  g0813(.A0(new_n1454_), .A1(new_n1453_), .B0(new_n1451_), .Y(new_n1456_));
  AOI21X1  g0814(.A0(new_n1455_), .A1(new_n1450_), .B0(new_n1456_), .Y(new_n1457_));
  INVX1    g0815(.A(new_n1441_), .Y(new_n1458_));
  OAI21X1  g0816(.A0(new_n1457_), .A1(new_n1412_), .B0(new_n1458_), .Y(new_n1459_));
  AOI21X1  g0817(.A0(new_n1459_), .A1(new_n1449_), .B0(new_n1444_), .Y(new_n1460_));
  OR2X1    g0818(.A(new_n1460_), .B(new_n1448_), .Y(new_n1461_));
  NAND3X1  g0819(.A(new_n1461_), .B(new_n1447_), .C(new_n1407_), .Y(new_n1462_));
  AOI21X1  g0820(.A0(new_n1461_), .A1(new_n1447_), .B0(new_n1407_), .Y(new_n1463_));
  AOI21X1  g0821(.A0(new_n1462_), .A1(new_n1406_), .B0(new_n1463_), .Y(new_n1464_));
  INVX1    g0822(.A(\in1[10] ), .Y(new_n1465_));
  AND2X1   g0823(.A(new_n1465_), .B(\in0[10] ), .Y(new_n1466_));
  INVX1    g0824(.A(new_n1466_), .Y(new_n1467_));
  OAI21X1  g0825(.A0(new_n1464_), .A1(new_n1405_), .B0(new_n1467_), .Y(new_n1468_));
  INVX1    g0826(.A(\in1[11] ), .Y(new_n1469_));
  AND2X1   g0827(.A(new_n1469_), .B(\in0[11] ), .Y(new_n1470_));
  AOI21X1  g0828(.A0(new_n1468_), .A1(new_n1403_), .B0(new_n1470_), .Y(new_n1471_));
  INVX1    g0829(.A(\in1[12] ), .Y(new_n1472_));
  AND2X1   g0830(.A(new_n1472_), .B(\in0[12] ), .Y(new_n1473_));
  INVX1    g0831(.A(new_n1473_), .Y(new_n1474_));
  OAI21X1  g0832(.A0(new_n1471_), .A1(new_n1400_), .B0(new_n1474_), .Y(new_n1475_));
  INVX1    g0833(.A(\in1[13] ), .Y(new_n1476_));
  AND2X1   g0834(.A(new_n1476_), .B(\in0[13] ), .Y(new_n1477_));
  AOI21X1  g0835(.A0(new_n1475_), .A1(new_n1398_), .B0(new_n1477_), .Y(new_n1478_));
  INVX1    g0836(.A(\in1[14] ), .Y(new_n1479_));
  AND2X1   g0837(.A(new_n1479_), .B(\in0[14] ), .Y(new_n1480_));
  INVX1    g0838(.A(new_n1480_), .Y(new_n1481_));
  OAI21X1  g0839(.A0(new_n1478_), .A1(new_n1395_), .B0(new_n1481_), .Y(new_n1482_));
  INVX1    g0840(.A(\in1[15] ), .Y(new_n1483_));
  AND2X1   g0841(.A(new_n1483_), .B(\in0[15] ), .Y(new_n1484_));
  AOI21X1  g0842(.A0(new_n1482_), .A1(new_n1393_), .B0(new_n1484_), .Y(new_n1485_));
  AOI21X1  g0843(.A0(new_n1485_), .A1(new_n1390_), .B0(\in1[16] ), .Y(new_n1486_));
  NOR2X1   g0844(.A(new_n1485_), .B(new_n1390_), .Y(new_n1487_));
  NOR3X1   g0845(.A(new_n1487_), .B(new_n1486_), .C(\in0[17] ), .Y(new_n1488_));
  OAI21X1  g0846(.A0(new_n1487_), .A1(new_n1486_), .B0(\in0[17] ), .Y(new_n1489_));
  OAI21X1  g0847(.A0(new_n1488_), .A1(\in1[17] ), .B0(new_n1489_), .Y(new_n1490_));
  INVX1    g0848(.A(\in1[18] ), .Y(new_n1491_));
  AND2X1   g0849(.A(new_n1491_), .B(\in0[18] ), .Y(new_n1492_));
  AOI21X1  g0850(.A0(new_n1490_), .A1(new_n1389_), .B0(new_n1492_), .Y(new_n1493_));
  INVX1    g0851(.A(\in1[19] ), .Y(new_n1494_));
  AND2X1   g0852(.A(new_n1494_), .B(\in0[19] ), .Y(new_n1495_));
  INVX1    g0853(.A(new_n1495_), .Y(new_n1496_));
  OAI21X1  g0854(.A0(new_n1493_), .A1(new_n1386_), .B0(new_n1496_), .Y(new_n1497_));
  INVX1    g0855(.A(\in1[20] ), .Y(new_n1498_));
  AND2X1   g0856(.A(new_n1498_), .B(\in0[20] ), .Y(new_n1499_));
  AOI21X1  g0857(.A0(new_n1497_), .A1(new_n1384_), .B0(new_n1499_), .Y(new_n1500_));
  INVX1    g0858(.A(\in1[21] ), .Y(new_n1501_));
  AND2X1   g0859(.A(new_n1501_), .B(\in0[21] ), .Y(new_n1502_));
  INVX1    g0860(.A(new_n1502_), .Y(new_n1503_));
  OAI21X1  g0861(.A0(new_n1500_), .A1(new_n1381_), .B0(new_n1503_), .Y(new_n1504_));
  INVX1    g0862(.A(\in1[22] ), .Y(new_n1505_));
  AND2X1   g0863(.A(new_n1505_), .B(\in0[22] ), .Y(new_n1506_));
  AOI21X1  g0864(.A0(new_n1504_), .A1(new_n1379_), .B0(new_n1506_), .Y(new_n1507_));
  INVX1    g0865(.A(\in1[23] ), .Y(new_n1508_));
  AND2X1   g0866(.A(new_n1508_), .B(\in0[23] ), .Y(new_n1509_));
  INVX1    g0867(.A(new_n1509_), .Y(new_n1510_));
  OAI21X1  g0868(.A0(new_n1507_), .A1(new_n1376_), .B0(new_n1510_), .Y(new_n1511_));
  OAI21X1  g0869(.A0(new_n1511_), .A1(\in0[24] ), .B0(new_n1374_), .Y(new_n1512_));
  NAND2X1  g0870(.A(new_n1511_), .B(\in0[24] ), .Y(new_n1513_));
  NAND3X1  g0871(.A(new_n1513_), .B(new_n1512_), .C(new_n1373_), .Y(new_n1514_));
  AOI21X1  g0872(.A0(new_n1513_), .A1(new_n1512_), .B0(new_n1373_), .Y(new_n1515_));
  AOI21X1  g0873(.A0(new_n1514_), .A1(new_n1372_), .B0(new_n1515_), .Y(new_n1516_));
  INVX1    g0874(.A(\in1[26] ), .Y(new_n1517_));
  AND2X1   g0875(.A(new_n1517_), .B(\in0[26] ), .Y(new_n1518_));
  INVX1    g0876(.A(new_n1518_), .Y(new_n1519_));
  OAI21X1  g0877(.A0(new_n1516_), .A1(new_n1371_), .B0(new_n1519_), .Y(new_n1520_));
  INVX1    g0878(.A(\in1[27] ), .Y(new_n1521_));
  AND2X1   g0879(.A(new_n1521_), .B(\in0[27] ), .Y(new_n1522_));
  AOI21X1  g0880(.A0(new_n1520_), .A1(new_n1369_), .B0(new_n1522_), .Y(new_n1523_));
  INVX1    g0881(.A(\in1[28] ), .Y(new_n1524_));
  AND2X1   g0882(.A(new_n1524_), .B(\in0[28] ), .Y(new_n1525_));
  INVX1    g0883(.A(new_n1525_), .Y(new_n1526_));
  OAI21X1  g0884(.A0(new_n1523_), .A1(new_n1366_), .B0(new_n1526_), .Y(new_n1527_));
  INVX1    g0885(.A(\in1[29] ), .Y(new_n1528_));
  AND2X1   g0886(.A(new_n1528_), .B(\in0[29] ), .Y(new_n1529_));
  AOI21X1  g0887(.A0(new_n1527_), .A1(new_n1364_), .B0(new_n1529_), .Y(new_n1530_));
  INVX1    g0888(.A(\in1[30] ), .Y(new_n1531_));
  AND2X1   g0889(.A(new_n1531_), .B(\in0[30] ), .Y(new_n1532_));
  INVX1    g0890(.A(new_n1532_), .Y(new_n1533_));
  OAI21X1  g0891(.A0(new_n1530_), .A1(new_n1361_), .B0(new_n1533_), .Y(new_n1534_));
  INVX1    g0892(.A(\in1[31] ), .Y(new_n1535_));
  AND2X1   g0893(.A(new_n1535_), .B(\in0[31] ), .Y(new_n1536_));
  AOI21X1  g0894(.A0(new_n1534_), .A1(new_n1359_), .B0(new_n1536_), .Y(new_n1537_));
  INVX1    g0895(.A(\in0[38] ), .Y(new_n1538_));
  INVX1    g0896(.A(\in0[39] ), .Y(new_n1539_));
  AOI22X1  g0897(.A0(\in1[39] ), .A1(new_n1539_), .B0(\in1[38] ), .B1(new_n1538_), .Y(new_n1540_));
  INVX1    g0898(.A(new_n1540_), .Y(new_n1541_));
  INVX1    g0899(.A(\in1[36] ), .Y(new_n1542_));
  INVX1    g0900(.A(\in1[37] ), .Y(new_n1543_));
  OAI22X1  g0901(.A0(new_n1543_), .A1(\in0[37] ), .B0(new_n1542_), .B1(\in0[36] ), .Y(new_n1544_));
  INVX1    g0902(.A(\in0[34] ), .Y(new_n1545_));
  INVX1    g0903(.A(\in0[35] ), .Y(new_n1546_));
  AOI22X1  g0904(.A0(\in1[35] ), .A1(new_n1546_), .B0(\in1[34] ), .B1(new_n1545_), .Y(new_n1547_));
  INVX1    g0905(.A(new_n1547_), .Y(new_n1548_));
  INVX1    g0906(.A(\in1[32] ), .Y(new_n1549_));
  INVX1    g0907(.A(\in1[33] ), .Y(new_n1550_));
  OAI22X1  g0908(.A0(new_n1550_), .A1(\in0[33] ), .B0(new_n1549_), .B1(\in0[32] ), .Y(new_n1551_));
  NOR4X1   g0909(.A(new_n1551_), .B(new_n1548_), .C(new_n1544_), .D(new_n1541_), .Y(new_n1552_));
  INVX1    g0910(.A(new_n1552_), .Y(new_n1553_));
  NOR2X1   g0911(.A(new_n1544_), .B(new_n1541_), .Y(new_n1554_));
  INVX1    g0912(.A(\in0[32] ), .Y(new_n1555_));
  INVX1    g0913(.A(\in0[33] ), .Y(new_n1556_));
  AND2X1   g0914(.A(\in1[33] ), .B(new_n1556_), .Y(new_n1557_));
  NOR3X1   g0915(.A(new_n1557_), .B(\in1[32] ), .C(new_n1555_), .Y(new_n1558_));
  OAI22X1  g0916(.A0(\in1[34] ), .A1(new_n1545_), .B0(\in1[33] ), .B1(new_n1556_), .Y(new_n1559_));
  OAI21X1  g0917(.A0(new_n1559_), .A1(new_n1558_), .B0(new_n1547_), .Y(new_n1560_));
  OAI21X1  g0918(.A0(\in1[35] ), .A1(new_n1546_), .B0(new_n1560_), .Y(new_n1561_));
  AND2X1   g0919(.A(new_n1561_), .B(new_n1554_), .Y(new_n1562_));
  INVX1    g0920(.A(\in0[36] ), .Y(new_n1563_));
  NOR2X1   g0921(.A(new_n1543_), .B(\in0[37] ), .Y(new_n1564_));
  NOR3X1   g0922(.A(new_n1564_), .B(\in1[36] ), .C(new_n1563_), .Y(new_n1565_));
  AOI21X1  g0923(.A0(new_n1543_), .A1(\in0[37] ), .B0(new_n1565_), .Y(new_n1566_));
  NOR2X1   g0924(.A(new_n1566_), .B(new_n1541_), .Y(new_n1567_));
  AND2X1   g0925(.A(\in1[39] ), .B(new_n1539_), .Y(new_n1568_));
  OR2X1    g0926(.A(\in1[39] ), .B(new_n1539_), .Y(new_n1569_));
  OR2X1    g0927(.A(\in1[38] ), .B(new_n1538_), .Y(new_n1570_));
  OAI21X1  g0928(.A0(new_n1570_), .A1(new_n1568_), .B0(new_n1569_), .Y(new_n1571_));
  NOR3X1   g0929(.A(new_n1571_), .B(new_n1567_), .C(new_n1562_), .Y(new_n1572_));
  OAI21X1  g0930(.A0(new_n1553_), .A1(new_n1537_), .B0(new_n1572_), .Y(new_n1573_));
  INVX1    g0931(.A(\in0[46] ), .Y(new_n1574_));
  INVX1    g0932(.A(\in0[47] ), .Y(new_n1575_));
  AOI22X1  g0933(.A0(\in1[47] ), .A1(new_n1575_), .B0(\in1[46] ), .B1(new_n1574_), .Y(new_n1576_));
  INVX1    g0934(.A(new_n1576_), .Y(new_n1577_));
  INVX1    g0935(.A(\in1[44] ), .Y(new_n1578_));
  INVX1    g0936(.A(\in1[45] ), .Y(new_n1579_));
  OAI22X1  g0937(.A0(new_n1579_), .A1(\in0[45] ), .B0(new_n1578_), .B1(\in0[44] ), .Y(new_n1580_));
  INVX1    g0938(.A(\in0[42] ), .Y(new_n1581_));
  INVX1    g0939(.A(\in0[43] ), .Y(new_n1582_));
  AOI22X1  g0940(.A0(\in1[43] ), .A1(new_n1582_), .B0(\in1[42] ), .B1(new_n1581_), .Y(new_n1583_));
  INVX1    g0941(.A(new_n1583_), .Y(new_n1584_));
  INVX1    g0942(.A(\in1[40] ), .Y(new_n1585_));
  INVX1    g0943(.A(\in1[41] ), .Y(new_n1586_));
  OAI22X1  g0944(.A0(new_n1586_), .A1(\in0[41] ), .B0(new_n1585_), .B1(\in0[40] ), .Y(new_n1587_));
  NOR4X1   g0945(.A(new_n1587_), .B(new_n1584_), .C(new_n1580_), .D(new_n1577_), .Y(new_n1588_));
  NOR2X1   g0946(.A(new_n1580_), .B(new_n1577_), .Y(new_n1589_));
  AND2X1   g0947(.A(new_n1585_), .B(\in0[40] ), .Y(new_n1590_));
  OAI21X1  g0948(.A0(new_n1586_), .A1(\in0[41] ), .B0(new_n1590_), .Y(new_n1591_));
  INVX1    g0949(.A(\in1[42] ), .Y(new_n1592_));
  AOI22X1  g0950(.A0(new_n1592_), .A1(\in0[42] ), .B0(new_n1586_), .B1(\in0[41] ), .Y(new_n1593_));
  AND2X1   g0951(.A(new_n1593_), .B(new_n1591_), .Y(new_n1594_));
  OAI22X1  g0952(.A0(new_n1594_), .A1(new_n1584_), .B0(\in1[43] ), .B1(new_n1582_), .Y(new_n1595_));
  AND2X1   g0953(.A(new_n1595_), .B(new_n1589_), .Y(new_n1596_));
  NOR2X1   g0954(.A(new_n1579_), .B(\in0[45] ), .Y(new_n1597_));
  NAND2X1  g0955(.A(new_n1578_), .B(\in0[44] ), .Y(new_n1598_));
  NOR2X1   g0956(.A(new_n1598_), .B(new_n1597_), .Y(new_n1599_));
  AOI21X1  g0957(.A0(new_n1579_), .A1(\in0[45] ), .B0(new_n1599_), .Y(new_n1600_));
  NOR2X1   g0958(.A(new_n1600_), .B(new_n1577_), .Y(new_n1601_));
  AND2X1   g0959(.A(\in1[47] ), .B(new_n1575_), .Y(new_n1602_));
  OR2X1    g0960(.A(\in1[47] ), .B(new_n1575_), .Y(new_n1603_));
  OR2X1    g0961(.A(\in1[46] ), .B(new_n1574_), .Y(new_n1604_));
  OAI21X1  g0962(.A0(new_n1604_), .A1(new_n1602_), .B0(new_n1603_), .Y(new_n1605_));
  NOR3X1   g0963(.A(new_n1605_), .B(new_n1601_), .C(new_n1596_), .Y(new_n1606_));
  INVX1    g0964(.A(new_n1606_), .Y(new_n1607_));
  AOI21X1  g0965(.A0(new_n1588_), .A1(new_n1573_), .B0(new_n1607_), .Y(new_n1608_));
  INVX1    g0966(.A(\in0[54] ), .Y(new_n1609_));
  INVX1    g0967(.A(\in0[55] ), .Y(new_n1610_));
  AOI22X1  g0968(.A0(\in1[55] ), .A1(new_n1610_), .B0(\in1[54] ), .B1(new_n1609_), .Y(new_n1611_));
  INVX1    g0969(.A(new_n1611_), .Y(new_n1612_));
  INVX1    g0970(.A(\in1[52] ), .Y(new_n1613_));
  INVX1    g0971(.A(\in1[53] ), .Y(new_n1614_));
  OAI22X1  g0972(.A0(new_n1614_), .A1(\in0[53] ), .B0(new_n1613_), .B1(\in0[52] ), .Y(new_n1615_));
  INVX1    g0973(.A(\in0[50] ), .Y(new_n1616_));
  INVX1    g0974(.A(\in0[51] ), .Y(new_n1617_));
  AOI22X1  g0975(.A0(\in1[51] ), .A1(new_n1617_), .B0(\in1[50] ), .B1(new_n1616_), .Y(new_n1618_));
  INVX1    g0976(.A(new_n1618_), .Y(new_n1619_));
  INVX1    g0977(.A(\in1[48] ), .Y(new_n1620_));
  INVX1    g0978(.A(\in1[49] ), .Y(new_n1621_));
  OAI22X1  g0979(.A0(new_n1621_), .A1(\in0[49] ), .B0(new_n1620_), .B1(\in0[48] ), .Y(new_n1622_));
  NOR4X1   g0980(.A(new_n1622_), .B(new_n1619_), .C(new_n1615_), .D(new_n1612_), .Y(new_n1623_));
  INVX1    g0981(.A(new_n1623_), .Y(new_n1624_));
  NOR2X1   g0982(.A(new_n1615_), .B(new_n1612_), .Y(new_n1625_));
  INVX1    g0983(.A(\in0[48] ), .Y(new_n1626_));
  INVX1    g0984(.A(\in0[49] ), .Y(new_n1627_));
  AND2X1   g0985(.A(\in1[49] ), .B(new_n1627_), .Y(new_n1628_));
  NOR3X1   g0986(.A(new_n1628_), .B(\in1[48] ), .C(new_n1626_), .Y(new_n1629_));
  OAI22X1  g0987(.A0(\in1[50] ), .A1(new_n1616_), .B0(\in1[49] ), .B1(new_n1627_), .Y(new_n1630_));
  OAI21X1  g0988(.A0(new_n1630_), .A1(new_n1629_), .B0(new_n1618_), .Y(new_n1631_));
  OAI21X1  g0989(.A0(\in1[51] ), .A1(new_n1617_), .B0(new_n1631_), .Y(new_n1632_));
  AND2X1   g0990(.A(new_n1613_), .B(\in0[52] ), .Y(new_n1633_));
  OAI21X1  g0991(.A0(new_n1614_), .A1(\in0[53] ), .B0(new_n1633_), .Y(new_n1634_));
  INVX1    g0992(.A(\in1[54] ), .Y(new_n1635_));
  AOI22X1  g0993(.A0(new_n1635_), .A1(\in0[54] ), .B0(new_n1614_), .B1(\in0[53] ), .Y(new_n1636_));
  AND2X1   g0994(.A(new_n1636_), .B(new_n1634_), .Y(new_n1637_));
  OAI22X1  g0995(.A0(new_n1637_), .A1(new_n1612_), .B0(\in1[55] ), .B1(new_n1610_), .Y(new_n1638_));
  AOI21X1  g0996(.A0(new_n1632_), .A1(new_n1625_), .B0(new_n1638_), .Y(new_n1639_));
  OAI21X1  g0997(.A0(new_n1624_), .A1(new_n1608_), .B0(new_n1639_), .Y(new_n1640_));
  INVX1    g0998(.A(\in0[62] ), .Y(new_n1641_));
  INVX1    g0999(.A(\in0[63] ), .Y(new_n1642_));
  AOI22X1  g1000(.A0(\in1[63] ), .A1(new_n1642_), .B0(\in1[62] ), .B1(new_n1641_), .Y(new_n1643_));
  INVX1    g1001(.A(new_n1643_), .Y(new_n1644_));
  INVX1    g1002(.A(\in1[60] ), .Y(new_n1645_));
  INVX1    g1003(.A(\in1[61] ), .Y(new_n1646_));
  OAI22X1  g1004(.A0(new_n1646_), .A1(\in0[61] ), .B0(new_n1645_), .B1(\in0[60] ), .Y(new_n1647_));
  INVX1    g1005(.A(\in0[58] ), .Y(new_n1648_));
  INVX1    g1006(.A(\in0[59] ), .Y(new_n1649_));
  AOI22X1  g1007(.A0(\in1[59] ), .A1(new_n1649_), .B0(\in1[58] ), .B1(new_n1648_), .Y(new_n1650_));
  INVX1    g1008(.A(new_n1650_), .Y(new_n1651_));
  INVX1    g1009(.A(\in1[56] ), .Y(new_n1652_));
  INVX1    g1010(.A(\in1[57] ), .Y(new_n1653_));
  OAI22X1  g1011(.A0(new_n1653_), .A1(\in0[57] ), .B0(new_n1652_), .B1(\in0[56] ), .Y(new_n1654_));
  NOR4X1   g1012(.A(new_n1654_), .B(new_n1651_), .C(new_n1647_), .D(new_n1644_), .Y(new_n1655_));
  NOR2X1   g1013(.A(new_n1647_), .B(new_n1644_), .Y(new_n1656_));
  AND2X1   g1014(.A(new_n1652_), .B(\in0[56] ), .Y(new_n1657_));
  OAI21X1  g1015(.A0(new_n1653_), .A1(\in0[57] ), .B0(new_n1657_), .Y(new_n1658_));
  INVX1    g1016(.A(\in1[58] ), .Y(new_n1659_));
  AOI22X1  g1017(.A0(new_n1659_), .A1(\in0[58] ), .B0(new_n1653_), .B1(\in0[57] ), .Y(new_n1660_));
  AND2X1   g1018(.A(new_n1660_), .B(new_n1658_), .Y(new_n1661_));
  OAI22X1  g1019(.A0(new_n1661_), .A1(new_n1651_), .B0(\in1[59] ), .B1(new_n1649_), .Y(new_n1662_));
  AND2X1   g1020(.A(new_n1662_), .B(new_n1656_), .Y(new_n1663_));
  NOR2X1   g1021(.A(new_n1646_), .B(\in0[61] ), .Y(new_n1664_));
  NAND2X1  g1022(.A(new_n1645_), .B(\in0[60] ), .Y(new_n1665_));
  NOR2X1   g1023(.A(new_n1665_), .B(new_n1664_), .Y(new_n1666_));
  AOI21X1  g1024(.A0(new_n1646_), .A1(\in0[61] ), .B0(new_n1666_), .Y(new_n1667_));
  NOR2X1   g1025(.A(new_n1667_), .B(new_n1644_), .Y(new_n1668_));
  AND2X1   g1026(.A(\in1[63] ), .B(new_n1642_), .Y(new_n1669_));
  OR2X1    g1027(.A(\in1[63] ), .B(new_n1642_), .Y(new_n1670_));
  OR2X1    g1028(.A(\in1[62] ), .B(new_n1641_), .Y(new_n1671_));
  OAI21X1  g1029(.A0(new_n1671_), .A1(new_n1669_), .B0(new_n1670_), .Y(new_n1672_));
  NOR3X1   g1030(.A(new_n1672_), .B(new_n1668_), .C(new_n1663_), .Y(new_n1673_));
  INVX1    g1031(.A(new_n1673_), .Y(new_n1674_));
  AOI21X1  g1032(.A0(new_n1655_), .A1(new_n1640_), .B0(new_n1674_), .Y(new_n1675_));
  INVX1    g1033(.A(\in0[66] ), .Y(new_n1676_));
  INVX1    g1034(.A(\in0[67] ), .Y(new_n1677_));
  AOI22X1  g1035(.A0(\in1[67] ), .A1(new_n1677_), .B0(\in1[66] ), .B1(new_n1676_), .Y(new_n1678_));
  INVX1    g1036(.A(\in0[64] ), .Y(new_n1679_));
  INVX1    g1037(.A(\in0[65] ), .Y(new_n1680_));
  AOI22X1  g1038(.A0(\in1[65] ), .A1(new_n1680_), .B0(\in1[64] ), .B1(new_n1679_), .Y(new_n1681_));
  AND2X1   g1039(.A(new_n1681_), .B(new_n1678_), .Y(new_n1682_));
  INVX1    g1040(.A(new_n1682_), .Y(new_n1683_));
  OR2X1    g1041(.A(\in1[67] ), .B(new_n1677_), .Y(new_n1684_));
  AND2X1   g1042(.A(\in1[65] ), .B(new_n1680_), .Y(new_n1685_));
  NOR3X1   g1043(.A(new_n1685_), .B(\in1[64] ), .C(new_n1679_), .Y(new_n1686_));
  INVX1    g1044(.A(\in1[65] ), .Y(new_n1687_));
  INVX1    g1045(.A(\in1[66] ), .Y(new_n1688_));
  AOI22X1  g1046(.A0(new_n1688_), .A1(\in0[66] ), .B0(new_n1687_), .B1(\in0[65] ), .Y(new_n1689_));
  INVX1    g1047(.A(new_n1689_), .Y(new_n1690_));
  OAI21X1  g1048(.A0(new_n1690_), .A1(new_n1686_), .B0(new_n1678_), .Y(new_n1691_));
  AND2X1   g1049(.A(new_n1691_), .B(new_n1684_), .Y(new_n1692_));
  OAI21X1  g1050(.A0(new_n1683_), .A1(new_n1675_), .B0(new_n1692_), .Y(new_n1693_));
  INVX1    g1051(.A(\in0[70] ), .Y(new_n1694_));
  INVX1    g1052(.A(\in0[71] ), .Y(new_n1695_));
  AOI22X1  g1053(.A0(\in1[71] ), .A1(new_n1695_), .B0(\in1[70] ), .B1(new_n1694_), .Y(new_n1696_));
  INVX1    g1054(.A(\in0[68] ), .Y(new_n1697_));
  INVX1    g1055(.A(\in0[69] ), .Y(new_n1698_));
  AOI22X1  g1056(.A0(\in1[69] ), .A1(new_n1698_), .B0(\in1[68] ), .B1(new_n1697_), .Y(new_n1699_));
  AND2X1   g1057(.A(new_n1699_), .B(new_n1696_), .Y(new_n1700_));
  AND2X1   g1058(.A(\in1[69] ), .B(new_n1698_), .Y(new_n1701_));
  OR2X1    g1059(.A(\in1[68] ), .B(new_n1697_), .Y(new_n1702_));
  OR2X1    g1060(.A(\in1[69] ), .B(new_n1698_), .Y(new_n1703_));
  OAI21X1  g1061(.A0(new_n1702_), .A1(new_n1701_), .B0(new_n1703_), .Y(new_n1704_));
  AND2X1   g1062(.A(\in1[71] ), .B(new_n1695_), .Y(new_n1705_));
  OR2X1    g1063(.A(\in1[71] ), .B(new_n1695_), .Y(new_n1706_));
  OR2X1    g1064(.A(\in1[70] ), .B(new_n1694_), .Y(new_n1707_));
  OAI21X1  g1065(.A0(new_n1707_), .A1(new_n1705_), .B0(new_n1706_), .Y(new_n1708_));
  AOI21X1  g1066(.A0(new_n1704_), .A1(new_n1696_), .B0(new_n1708_), .Y(new_n1709_));
  INVX1    g1067(.A(new_n1709_), .Y(new_n1710_));
  AOI21X1  g1068(.A0(new_n1700_), .A1(new_n1693_), .B0(new_n1710_), .Y(new_n1711_));
  INVX1    g1069(.A(\in0[74] ), .Y(new_n1712_));
  INVX1    g1070(.A(\in0[75] ), .Y(new_n1713_));
  AOI22X1  g1071(.A0(\in1[75] ), .A1(new_n1713_), .B0(\in1[74] ), .B1(new_n1712_), .Y(new_n1714_));
  INVX1    g1072(.A(\in0[72] ), .Y(new_n1715_));
  INVX1    g1073(.A(\in0[73] ), .Y(new_n1716_));
  AOI22X1  g1074(.A0(\in1[73] ), .A1(new_n1716_), .B0(\in1[72] ), .B1(new_n1715_), .Y(new_n1717_));
  AND2X1   g1075(.A(new_n1717_), .B(new_n1714_), .Y(new_n1718_));
  INVX1    g1076(.A(new_n1718_), .Y(new_n1719_));
  OR2X1    g1077(.A(\in1[75] ), .B(new_n1713_), .Y(new_n1720_));
  AND2X1   g1078(.A(\in1[73] ), .B(new_n1716_), .Y(new_n1721_));
  NOR3X1   g1079(.A(new_n1721_), .B(\in1[72] ), .C(new_n1715_), .Y(new_n1722_));
  INVX1    g1080(.A(\in1[73] ), .Y(new_n1723_));
  INVX1    g1081(.A(\in1[74] ), .Y(new_n1724_));
  AOI22X1  g1082(.A0(new_n1724_), .A1(\in0[74] ), .B0(new_n1723_), .B1(\in0[73] ), .Y(new_n1725_));
  INVX1    g1083(.A(new_n1725_), .Y(new_n1726_));
  OAI21X1  g1084(.A0(new_n1726_), .A1(new_n1722_), .B0(new_n1714_), .Y(new_n1727_));
  AND2X1   g1085(.A(new_n1727_), .B(new_n1720_), .Y(new_n1728_));
  OAI21X1  g1086(.A0(new_n1719_), .A1(new_n1711_), .B0(new_n1728_), .Y(new_n1729_));
  INVX1    g1087(.A(\in0[78] ), .Y(new_n1730_));
  INVX1    g1088(.A(\in0[79] ), .Y(new_n1731_));
  AOI22X1  g1089(.A0(\in1[79] ), .A1(new_n1731_), .B0(\in1[78] ), .B1(new_n1730_), .Y(new_n1732_));
  INVX1    g1090(.A(\in0[76] ), .Y(new_n1733_));
  INVX1    g1091(.A(\in0[77] ), .Y(new_n1734_));
  AOI22X1  g1092(.A0(\in1[77] ), .A1(new_n1734_), .B0(\in1[76] ), .B1(new_n1733_), .Y(new_n1735_));
  AND2X1   g1093(.A(new_n1735_), .B(new_n1732_), .Y(new_n1736_));
  AND2X1   g1094(.A(\in1[77] ), .B(new_n1734_), .Y(new_n1737_));
  OR2X1    g1095(.A(\in1[76] ), .B(new_n1733_), .Y(new_n1738_));
  OR2X1    g1096(.A(\in1[77] ), .B(new_n1734_), .Y(new_n1739_));
  OAI21X1  g1097(.A0(new_n1738_), .A1(new_n1737_), .B0(new_n1739_), .Y(new_n1740_));
  AND2X1   g1098(.A(\in1[79] ), .B(new_n1731_), .Y(new_n1741_));
  OR2X1    g1099(.A(\in1[79] ), .B(new_n1731_), .Y(new_n1742_));
  OR2X1    g1100(.A(\in1[78] ), .B(new_n1730_), .Y(new_n1743_));
  OAI21X1  g1101(.A0(new_n1743_), .A1(new_n1741_), .B0(new_n1742_), .Y(new_n1744_));
  AOI21X1  g1102(.A0(new_n1740_), .A1(new_n1732_), .B0(new_n1744_), .Y(new_n1745_));
  INVX1    g1103(.A(new_n1745_), .Y(new_n1746_));
  AOI21X1  g1104(.A0(new_n1736_), .A1(new_n1729_), .B0(new_n1746_), .Y(new_n1747_));
  INVX1    g1105(.A(\in0[82] ), .Y(new_n1748_));
  INVX1    g1106(.A(\in0[83] ), .Y(new_n1749_));
  AOI22X1  g1107(.A0(\in1[83] ), .A1(new_n1749_), .B0(\in1[82] ), .B1(new_n1748_), .Y(new_n1750_));
  INVX1    g1108(.A(\in0[80] ), .Y(new_n1751_));
  INVX1    g1109(.A(\in0[81] ), .Y(new_n1752_));
  AOI22X1  g1110(.A0(\in1[81] ), .A1(new_n1752_), .B0(\in1[80] ), .B1(new_n1751_), .Y(new_n1753_));
  AND2X1   g1111(.A(new_n1753_), .B(new_n1750_), .Y(new_n1754_));
  INVX1    g1112(.A(new_n1754_), .Y(new_n1755_));
  OR2X1    g1113(.A(\in1[83] ), .B(new_n1749_), .Y(new_n1756_));
  AND2X1   g1114(.A(\in1[81] ), .B(new_n1752_), .Y(new_n1757_));
  NOR3X1   g1115(.A(new_n1757_), .B(\in1[80] ), .C(new_n1751_), .Y(new_n1758_));
  INVX1    g1116(.A(\in1[81] ), .Y(new_n1759_));
  INVX1    g1117(.A(\in1[82] ), .Y(new_n1760_));
  AOI22X1  g1118(.A0(new_n1760_), .A1(\in0[82] ), .B0(new_n1759_), .B1(\in0[81] ), .Y(new_n1761_));
  INVX1    g1119(.A(new_n1761_), .Y(new_n1762_));
  OAI21X1  g1120(.A0(new_n1762_), .A1(new_n1758_), .B0(new_n1750_), .Y(new_n1763_));
  AND2X1   g1121(.A(new_n1763_), .B(new_n1756_), .Y(new_n1764_));
  OAI21X1  g1122(.A0(new_n1755_), .A1(new_n1747_), .B0(new_n1764_), .Y(new_n1765_));
  INVX1    g1123(.A(\in0[86] ), .Y(new_n1766_));
  INVX1    g1124(.A(\in0[87] ), .Y(new_n1767_));
  AOI22X1  g1125(.A0(\in1[87] ), .A1(new_n1767_), .B0(\in1[86] ), .B1(new_n1766_), .Y(new_n1768_));
  INVX1    g1126(.A(\in0[84] ), .Y(new_n1769_));
  INVX1    g1127(.A(\in0[85] ), .Y(new_n1770_));
  AOI22X1  g1128(.A0(\in1[85] ), .A1(new_n1770_), .B0(\in1[84] ), .B1(new_n1769_), .Y(new_n1771_));
  AND2X1   g1129(.A(new_n1771_), .B(new_n1768_), .Y(new_n1772_));
  AND2X1   g1130(.A(\in1[85] ), .B(new_n1770_), .Y(new_n1773_));
  OR2X1    g1131(.A(\in1[84] ), .B(new_n1769_), .Y(new_n1774_));
  OR2X1    g1132(.A(\in1[85] ), .B(new_n1770_), .Y(new_n1775_));
  OAI21X1  g1133(.A0(new_n1774_), .A1(new_n1773_), .B0(new_n1775_), .Y(new_n1776_));
  AND2X1   g1134(.A(\in1[87] ), .B(new_n1767_), .Y(new_n1777_));
  OR2X1    g1135(.A(\in1[87] ), .B(new_n1767_), .Y(new_n1778_));
  OR2X1    g1136(.A(\in1[86] ), .B(new_n1766_), .Y(new_n1779_));
  OAI21X1  g1137(.A0(new_n1779_), .A1(new_n1777_), .B0(new_n1778_), .Y(new_n1780_));
  AOI21X1  g1138(.A0(new_n1776_), .A1(new_n1768_), .B0(new_n1780_), .Y(new_n1781_));
  INVX1    g1139(.A(new_n1781_), .Y(new_n1782_));
  AOI21X1  g1140(.A0(new_n1772_), .A1(new_n1765_), .B0(new_n1782_), .Y(new_n1783_));
  INVX1    g1141(.A(\in0[90] ), .Y(new_n1784_));
  INVX1    g1142(.A(\in0[91] ), .Y(new_n1785_));
  AOI22X1  g1143(.A0(\in1[91] ), .A1(new_n1785_), .B0(\in1[90] ), .B1(new_n1784_), .Y(new_n1786_));
  INVX1    g1144(.A(\in0[88] ), .Y(new_n1787_));
  INVX1    g1145(.A(\in0[89] ), .Y(new_n1788_));
  AOI22X1  g1146(.A0(\in1[89] ), .A1(new_n1788_), .B0(\in1[88] ), .B1(new_n1787_), .Y(new_n1789_));
  AND2X1   g1147(.A(new_n1789_), .B(new_n1786_), .Y(new_n1790_));
  INVX1    g1148(.A(new_n1790_), .Y(new_n1791_));
  OR2X1    g1149(.A(\in1[91] ), .B(new_n1785_), .Y(new_n1792_));
  AND2X1   g1150(.A(\in1[89] ), .B(new_n1788_), .Y(new_n1793_));
  NOR3X1   g1151(.A(new_n1793_), .B(\in1[88] ), .C(new_n1787_), .Y(new_n1794_));
  INVX1    g1152(.A(\in1[89] ), .Y(new_n1795_));
  INVX1    g1153(.A(\in1[90] ), .Y(new_n1796_));
  AOI22X1  g1154(.A0(new_n1796_), .A1(\in0[90] ), .B0(new_n1795_), .B1(\in0[89] ), .Y(new_n1797_));
  INVX1    g1155(.A(new_n1797_), .Y(new_n1798_));
  OAI21X1  g1156(.A0(new_n1798_), .A1(new_n1794_), .B0(new_n1786_), .Y(new_n1799_));
  AND2X1   g1157(.A(new_n1799_), .B(new_n1792_), .Y(new_n1800_));
  OAI21X1  g1158(.A0(new_n1791_), .A1(new_n1783_), .B0(new_n1800_), .Y(new_n1801_));
  INVX1    g1159(.A(\in0[94] ), .Y(new_n1802_));
  INVX1    g1160(.A(\in0[95] ), .Y(new_n1803_));
  AOI22X1  g1161(.A0(\in1[95] ), .A1(new_n1803_), .B0(\in1[94] ), .B1(new_n1802_), .Y(new_n1804_));
  INVX1    g1162(.A(\in0[92] ), .Y(new_n1805_));
  INVX1    g1163(.A(\in0[93] ), .Y(new_n1806_));
  AOI22X1  g1164(.A0(\in1[93] ), .A1(new_n1806_), .B0(\in1[92] ), .B1(new_n1805_), .Y(new_n1807_));
  AND2X1   g1165(.A(new_n1807_), .B(new_n1804_), .Y(new_n1808_));
  AND2X1   g1166(.A(\in1[93] ), .B(new_n1806_), .Y(new_n1809_));
  OR2X1    g1167(.A(\in1[92] ), .B(new_n1805_), .Y(new_n1810_));
  OR2X1    g1168(.A(\in1[93] ), .B(new_n1806_), .Y(new_n1811_));
  OAI21X1  g1169(.A0(new_n1810_), .A1(new_n1809_), .B0(new_n1811_), .Y(new_n1812_));
  AND2X1   g1170(.A(\in1[95] ), .B(new_n1803_), .Y(new_n1813_));
  OR2X1    g1171(.A(\in1[95] ), .B(new_n1803_), .Y(new_n1814_));
  OR2X1    g1172(.A(\in1[94] ), .B(new_n1802_), .Y(new_n1815_));
  OAI21X1  g1173(.A0(new_n1815_), .A1(new_n1813_), .B0(new_n1814_), .Y(new_n1816_));
  AOI21X1  g1174(.A0(new_n1812_), .A1(new_n1804_), .B0(new_n1816_), .Y(new_n1817_));
  INVX1    g1175(.A(new_n1817_), .Y(new_n1818_));
  AOI21X1  g1176(.A0(new_n1808_), .A1(new_n1801_), .B0(new_n1818_), .Y(new_n1819_));
  INVX1    g1177(.A(\in0[98] ), .Y(new_n1820_));
  INVX1    g1178(.A(\in0[99] ), .Y(new_n1821_));
  AOI22X1  g1179(.A0(\in1[99] ), .A1(new_n1821_), .B0(\in1[98] ), .B1(new_n1820_), .Y(new_n1822_));
  INVX1    g1180(.A(\in0[96] ), .Y(new_n1823_));
  INVX1    g1181(.A(\in0[97] ), .Y(new_n1824_));
  AOI22X1  g1182(.A0(\in1[97] ), .A1(new_n1824_), .B0(\in1[96] ), .B1(new_n1823_), .Y(new_n1825_));
  AND2X1   g1183(.A(new_n1825_), .B(new_n1822_), .Y(new_n1826_));
  INVX1    g1184(.A(new_n1826_), .Y(new_n1827_));
  OR2X1    g1185(.A(\in1[99] ), .B(new_n1821_), .Y(new_n1828_));
  AND2X1   g1186(.A(\in1[97] ), .B(new_n1824_), .Y(new_n1829_));
  NOR3X1   g1187(.A(new_n1829_), .B(\in1[96] ), .C(new_n1823_), .Y(new_n1830_));
  INVX1    g1188(.A(\in1[97] ), .Y(new_n1831_));
  INVX1    g1189(.A(\in1[98] ), .Y(new_n1832_));
  AOI22X1  g1190(.A0(new_n1832_), .A1(\in0[98] ), .B0(new_n1831_), .B1(\in0[97] ), .Y(new_n1833_));
  INVX1    g1191(.A(new_n1833_), .Y(new_n1834_));
  OAI21X1  g1192(.A0(new_n1834_), .A1(new_n1830_), .B0(new_n1822_), .Y(new_n1835_));
  AND2X1   g1193(.A(new_n1835_), .B(new_n1828_), .Y(new_n1836_));
  OAI21X1  g1194(.A0(new_n1827_), .A1(new_n1819_), .B0(new_n1836_), .Y(new_n1837_));
  INVX1    g1195(.A(\in0[102] ), .Y(new_n1838_));
  INVX1    g1196(.A(\in0[103] ), .Y(new_n1839_));
  AOI22X1  g1197(.A0(\in1[103] ), .A1(new_n1839_), .B0(\in1[102] ), .B1(new_n1838_), .Y(new_n1840_));
  INVX1    g1198(.A(\in0[100] ), .Y(new_n1841_));
  INVX1    g1199(.A(\in0[101] ), .Y(new_n1842_));
  AOI22X1  g1200(.A0(\in1[101] ), .A1(new_n1842_), .B0(\in1[100] ), .B1(new_n1841_), .Y(new_n1843_));
  AND2X1   g1201(.A(new_n1843_), .B(new_n1840_), .Y(new_n1844_));
  AND2X1   g1202(.A(\in1[101] ), .B(new_n1842_), .Y(new_n1845_));
  OR2X1    g1203(.A(\in1[100] ), .B(new_n1841_), .Y(new_n1846_));
  OR2X1    g1204(.A(\in1[101] ), .B(new_n1842_), .Y(new_n1847_));
  OAI21X1  g1205(.A0(new_n1846_), .A1(new_n1845_), .B0(new_n1847_), .Y(new_n1848_));
  AND2X1   g1206(.A(\in1[103] ), .B(new_n1839_), .Y(new_n1849_));
  OR2X1    g1207(.A(\in1[103] ), .B(new_n1839_), .Y(new_n1850_));
  OR2X1    g1208(.A(\in1[102] ), .B(new_n1838_), .Y(new_n1851_));
  OAI21X1  g1209(.A0(new_n1851_), .A1(new_n1849_), .B0(new_n1850_), .Y(new_n1852_));
  AOI21X1  g1210(.A0(new_n1848_), .A1(new_n1840_), .B0(new_n1852_), .Y(new_n1853_));
  INVX1    g1211(.A(new_n1853_), .Y(new_n1854_));
  AOI21X1  g1212(.A0(new_n1844_), .A1(new_n1837_), .B0(new_n1854_), .Y(new_n1855_));
  INVX1    g1213(.A(\in0[106] ), .Y(new_n1856_));
  INVX1    g1214(.A(\in0[107] ), .Y(new_n1857_));
  AOI22X1  g1215(.A0(\in1[107] ), .A1(new_n1857_), .B0(\in1[106] ), .B1(new_n1856_), .Y(new_n1858_));
  INVX1    g1216(.A(\in0[104] ), .Y(new_n1859_));
  INVX1    g1217(.A(\in0[105] ), .Y(new_n1860_));
  AOI22X1  g1218(.A0(\in1[105] ), .A1(new_n1860_), .B0(\in1[104] ), .B1(new_n1859_), .Y(new_n1861_));
  AND2X1   g1219(.A(new_n1861_), .B(new_n1858_), .Y(new_n1862_));
  INVX1    g1220(.A(new_n1862_), .Y(new_n1863_));
  OR2X1    g1221(.A(\in1[107] ), .B(new_n1857_), .Y(new_n1864_));
  AND2X1   g1222(.A(\in1[105] ), .B(new_n1860_), .Y(new_n1865_));
  NOR3X1   g1223(.A(new_n1865_), .B(\in1[104] ), .C(new_n1859_), .Y(new_n1866_));
  INVX1    g1224(.A(\in1[105] ), .Y(new_n1867_));
  INVX1    g1225(.A(\in1[106] ), .Y(new_n1868_));
  AOI22X1  g1226(.A0(new_n1868_), .A1(\in0[106] ), .B0(new_n1867_), .B1(\in0[105] ), .Y(new_n1869_));
  INVX1    g1227(.A(new_n1869_), .Y(new_n1870_));
  OAI21X1  g1228(.A0(new_n1870_), .A1(new_n1866_), .B0(new_n1858_), .Y(new_n1871_));
  AND2X1   g1229(.A(new_n1871_), .B(new_n1864_), .Y(new_n1872_));
  OAI21X1  g1230(.A0(new_n1863_), .A1(new_n1855_), .B0(new_n1872_), .Y(new_n1873_));
  INVX1    g1231(.A(\in0[110] ), .Y(new_n1874_));
  INVX1    g1232(.A(\in0[111] ), .Y(new_n1875_));
  AOI22X1  g1233(.A0(\in1[111] ), .A1(new_n1875_), .B0(\in1[110] ), .B1(new_n1874_), .Y(new_n1876_));
  INVX1    g1234(.A(\in0[108] ), .Y(new_n1877_));
  INVX1    g1235(.A(\in0[109] ), .Y(new_n1878_));
  AOI22X1  g1236(.A0(\in1[109] ), .A1(new_n1878_), .B0(\in1[108] ), .B1(new_n1877_), .Y(new_n1879_));
  AND2X1   g1237(.A(new_n1879_), .B(new_n1876_), .Y(new_n1880_));
  AND2X1   g1238(.A(\in1[109] ), .B(new_n1878_), .Y(new_n1881_));
  OR2X1    g1239(.A(\in1[108] ), .B(new_n1877_), .Y(new_n1882_));
  OR2X1    g1240(.A(\in1[109] ), .B(new_n1878_), .Y(new_n1883_));
  OAI21X1  g1241(.A0(new_n1882_), .A1(new_n1881_), .B0(new_n1883_), .Y(new_n1884_));
  AND2X1   g1242(.A(\in1[111] ), .B(new_n1875_), .Y(new_n1885_));
  OR2X1    g1243(.A(\in1[111] ), .B(new_n1875_), .Y(new_n1886_));
  OR2X1    g1244(.A(\in1[110] ), .B(new_n1874_), .Y(new_n1887_));
  OAI21X1  g1245(.A0(new_n1887_), .A1(new_n1885_), .B0(new_n1886_), .Y(new_n1888_));
  AOI21X1  g1246(.A0(new_n1884_), .A1(new_n1876_), .B0(new_n1888_), .Y(new_n1889_));
  INVX1    g1247(.A(new_n1889_), .Y(new_n1890_));
  AOI21X1  g1248(.A0(new_n1880_), .A1(new_n1873_), .B0(new_n1890_), .Y(new_n1891_));
  INVX1    g1249(.A(\in0[114] ), .Y(new_n1892_));
  INVX1    g1250(.A(\in0[115] ), .Y(new_n1893_));
  AOI22X1  g1251(.A0(\in1[115] ), .A1(new_n1893_), .B0(\in1[114] ), .B1(new_n1892_), .Y(new_n1894_));
  INVX1    g1252(.A(\in0[112] ), .Y(new_n1895_));
  INVX1    g1253(.A(\in0[113] ), .Y(new_n1896_));
  AOI22X1  g1254(.A0(\in1[113] ), .A1(new_n1896_), .B0(\in1[112] ), .B1(new_n1895_), .Y(new_n1897_));
  AND2X1   g1255(.A(new_n1897_), .B(new_n1894_), .Y(new_n1898_));
  INVX1    g1256(.A(new_n1898_), .Y(new_n1899_));
  OR2X1    g1257(.A(\in1[115] ), .B(new_n1893_), .Y(new_n1900_));
  AND2X1   g1258(.A(\in1[113] ), .B(new_n1896_), .Y(new_n1901_));
  NOR3X1   g1259(.A(new_n1901_), .B(\in1[112] ), .C(new_n1895_), .Y(new_n1902_));
  INVX1    g1260(.A(\in1[113] ), .Y(new_n1903_));
  INVX1    g1261(.A(\in1[114] ), .Y(new_n1904_));
  AOI22X1  g1262(.A0(new_n1904_), .A1(\in0[114] ), .B0(new_n1903_), .B1(\in0[113] ), .Y(new_n1905_));
  INVX1    g1263(.A(new_n1905_), .Y(new_n1906_));
  OAI21X1  g1264(.A0(new_n1906_), .A1(new_n1902_), .B0(new_n1894_), .Y(new_n1907_));
  AND2X1   g1265(.A(new_n1907_), .B(new_n1900_), .Y(new_n1908_));
  OAI21X1  g1266(.A0(new_n1899_), .A1(new_n1891_), .B0(new_n1908_), .Y(new_n1909_));
  INVX1    g1267(.A(\in0[118] ), .Y(new_n1910_));
  INVX1    g1268(.A(\in0[119] ), .Y(new_n1911_));
  AOI22X1  g1269(.A0(\in1[119] ), .A1(new_n1911_), .B0(\in1[118] ), .B1(new_n1910_), .Y(new_n1912_));
  INVX1    g1270(.A(\in0[116] ), .Y(new_n1913_));
  INVX1    g1271(.A(\in0[117] ), .Y(new_n1914_));
  AOI22X1  g1272(.A0(\in1[117] ), .A1(new_n1914_), .B0(\in1[116] ), .B1(new_n1913_), .Y(new_n1915_));
  AND2X1   g1273(.A(new_n1915_), .B(new_n1912_), .Y(new_n1916_));
  AND2X1   g1274(.A(\in1[117] ), .B(new_n1914_), .Y(new_n1917_));
  OR2X1    g1275(.A(\in1[116] ), .B(new_n1913_), .Y(new_n1918_));
  OR2X1    g1276(.A(\in1[117] ), .B(new_n1914_), .Y(new_n1919_));
  OAI21X1  g1277(.A0(new_n1918_), .A1(new_n1917_), .B0(new_n1919_), .Y(new_n1920_));
  AND2X1   g1278(.A(\in1[119] ), .B(new_n1911_), .Y(new_n1921_));
  OR2X1    g1279(.A(\in1[119] ), .B(new_n1911_), .Y(new_n1922_));
  OR2X1    g1280(.A(\in1[118] ), .B(new_n1910_), .Y(new_n1923_));
  OAI21X1  g1281(.A0(new_n1923_), .A1(new_n1921_), .B0(new_n1922_), .Y(new_n1924_));
  AOI21X1  g1282(.A0(new_n1920_), .A1(new_n1912_), .B0(new_n1924_), .Y(new_n1925_));
  INVX1    g1283(.A(new_n1925_), .Y(new_n1926_));
  AOI21X1  g1284(.A0(new_n1916_), .A1(new_n1909_), .B0(new_n1926_), .Y(new_n1927_));
  INVX1    g1285(.A(\in0[122] ), .Y(new_n1928_));
  INVX1    g1286(.A(\in0[123] ), .Y(new_n1929_));
  AOI22X1  g1287(.A0(\in1[123] ), .A1(new_n1929_), .B0(\in1[122] ), .B1(new_n1928_), .Y(new_n1930_));
  INVX1    g1288(.A(\in0[120] ), .Y(new_n1931_));
  INVX1    g1289(.A(\in0[121] ), .Y(new_n1932_));
  AOI22X1  g1290(.A0(\in1[121] ), .A1(new_n1932_), .B0(\in1[120] ), .B1(new_n1931_), .Y(new_n1933_));
  AND2X1   g1291(.A(new_n1933_), .B(new_n1930_), .Y(new_n1934_));
  INVX1    g1292(.A(new_n1934_), .Y(new_n1935_));
  OR2X1    g1293(.A(\in1[123] ), .B(new_n1929_), .Y(new_n1936_));
  AND2X1   g1294(.A(\in1[121] ), .B(new_n1932_), .Y(new_n1937_));
  NOR3X1   g1295(.A(new_n1937_), .B(\in1[120] ), .C(new_n1931_), .Y(new_n1938_));
  INVX1    g1296(.A(\in1[121] ), .Y(new_n1939_));
  INVX1    g1297(.A(\in1[122] ), .Y(new_n1940_));
  AOI22X1  g1298(.A0(new_n1940_), .A1(\in0[122] ), .B0(new_n1939_), .B1(\in0[121] ), .Y(new_n1941_));
  INVX1    g1299(.A(new_n1941_), .Y(new_n1942_));
  OAI21X1  g1300(.A0(new_n1942_), .A1(new_n1938_), .B0(new_n1930_), .Y(new_n1943_));
  AND2X1   g1301(.A(new_n1943_), .B(new_n1936_), .Y(new_n1944_));
  OAI21X1  g1302(.A0(new_n1935_), .A1(new_n1927_), .B0(new_n1944_), .Y(new_n1945_));
  INVX1    g1303(.A(\in0[125] ), .Y(new_n1946_));
  INVX1    g1304(.A(\in0[126] ), .Y(new_n1947_));
  AOI22X1  g1305(.A0(\in1[126] ), .A1(new_n1947_), .B0(\in1[125] ), .B1(new_n1946_), .Y(new_n1948_));
  INVX1    g1306(.A(\in0[124] ), .Y(new_n1949_));
  AOI22X1  g1307(.A0(new_n1356_), .A1(\in0[127] ), .B0(\in1[124] ), .B1(new_n1949_), .Y(new_n1950_));
  AND2X1   g1308(.A(new_n1950_), .B(new_n1948_), .Y(new_n1951_));
  INVX1    g1309(.A(\in1[126] ), .Y(new_n1952_));
  INVX1    g1310(.A(\in1[124] ), .Y(new_n1953_));
  INVX1    g1311(.A(\in1[125] ), .Y(new_n1954_));
  AOI22X1  g1312(.A0(new_n1954_), .A1(\in0[125] ), .B0(new_n1953_), .B1(\in0[124] ), .Y(new_n1955_));
  INVX1    g1313(.A(new_n1955_), .Y(new_n1956_));
  AOI22X1  g1314(.A0(new_n1956_), .A1(new_n1948_), .B0(new_n1952_), .B1(\in0[126] ), .Y(new_n1957_));
  AOI21X1  g1315(.A0(new_n1356_), .A1(\in0[127] ), .B0(new_n1957_), .Y(new_n1958_));
  AOI21X1  g1316(.A0(new_n1951_), .A1(new_n1945_), .B0(new_n1958_), .Y(new_n1959_));
  OAI21X1  g1317(.A0(new_n1356_), .A1(\in0[127] ), .B0(new_n1959_), .Y(new_n1960_));
  MX2X1    g1318(.A(\in1[0] ), .B(\in0[0] ), .S0(new_n1960_), .Y(new_n1961_));
  AOI21X1  g1319(.A0(new_n1352_), .A1(new_n1274_), .B0(new_n1290_), .Y(new_n1962_));
  AND2X1   g1320(.A(new_n1951_), .B(new_n1945_), .Y(new_n1963_));
  OAI21X1  g1321(.A0(new_n1963_), .A1(\in1[127] ), .B0(\in0[127] ), .Y(new_n1964_));
  AND2X1   g1322(.A(new_n1964_), .B(new_n1962_), .Y(new_n1965_));
  INVX1    g1323(.A(new_n1965_), .Y(new_n1966_));
  MX2X1    g1324(.A(new_n1535_), .B(new_n1357_), .S0(new_n1960_), .Y(new_n1967_));
  INVX1    g1325(.A(new_n1967_), .Y(new_n1968_));
  OR2X1    g1326(.A(new_n1291_), .B(new_n1289_), .Y(new_n1969_));
  MX2X1    g1327(.A(new_n857_), .B(new_n644_), .S0(new_n1969_), .Y(new_n1970_));
  MX2X1    g1328(.A(new_n1531_), .B(new_n1360_), .S0(new_n1960_), .Y(new_n1971_));
  MX2X1    g1329(.A(new_n854_), .B(new_n646_), .S0(new_n1969_), .Y(new_n1972_));
  INVX1    g1330(.A(new_n1972_), .Y(new_n1973_));
  MX2X1    g1331(.A(new_n1528_), .B(new_n1362_), .S0(new_n1960_), .Y(new_n1974_));
  INVX1    g1332(.A(new_n1974_), .Y(new_n1975_));
  MX2X1    g1333(.A(new_n850_), .B(new_n649_), .S0(new_n1969_), .Y(new_n1976_));
  MX2X1    g1334(.A(new_n1524_), .B(new_n1365_), .S0(new_n1960_), .Y(new_n1977_));
  MX2X1    g1335(.A(new_n847_), .B(new_n651_), .S0(new_n1969_), .Y(new_n1978_));
  INVX1    g1336(.A(new_n1978_), .Y(new_n1979_));
  MX2X1    g1337(.A(new_n1521_), .B(new_n1367_), .S0(new_n1960_), .Y(new_n1980_));
  INVX1    g1338(.A(new_n1980_), .Y(new_n1981_));
  MX2X1    g1339(.A(new_n843_), .B(new_n654_), .S0(new_n1969_), .Y(new_n1982_));
  MX2X1    g1340(.A(new_n1517_), .B(new_n1370_), .S0(new_n1960_), .Y(new_n1983_));
  MX2X1    g1341(.A(new_n840_), .B(new_n656_), .S0(new_n1969_), .Y(new_n1984_));
  INVX1    g1342(.A(new_n1984_), .Y(new_n1985_));
  MX2X1    g1343(.A(new_n1296_), .B(new_n1297_), .S0(new_n1969_), .Y(new_n1986_));
  MX2X1    g1344(.A(new_n1298_), .B(new_n659_), .S0(new_n1969_), .Y(new_n1987_));
  INVX1    g1345(.A(new_n1987_), .Y(new_n1988_));
  MX2X1    g1346(.A(new_n1508_), .B(new_n1375_), .S0(new_n1960_), .Y(new_n1989_));
  MX2X1    g1347(.A(new_n815_), .B(new_n660_), .S0(new_n1969_), .Y(new_n1990_));
  INVX1    g1348(.A(new_n1990_), .Y(new_n1991_));
  MX2X1    g1349(.A(new_n1505_), .B(new_n1377_), .S0(new_n1960_), .Y(new_n1992_));
  INVX1    g1350(.A(new_n1992_), .Y(new_n1993_));
  MX2X1    g1351(.A(new_n811_), .B(new_n663_), .S0(new_n1969_), .Y(new_n1994_));
  MX2X1    g1352(.A(new_n1501_), .B(new_n1380_), .S0(new_n1960_), .Y(new_n1995_));
  MX2X1    g1353(.A(new_n808_), .B(new_n665_), .S0(new_n1969_), .Y(new_n1996_));
  INVX1    g1354(.A(new_n1996_), .Y(new_n1997_));
  MX2X1    g1355(.A(new_n1498_), .B(new_n1382_), .S0(new_n1960_), .Y(new_n1998_));
  INVX1    g1356(.A(new_n1998_), .Y(new_n1999_));
  MX2X1    g1357(.A(new_n804_), .B(new_n668_), .S0(new_n1969_), .Y(new_n2000_));
  MX2X1    g1358(.A(new_n1494_), .B(new_n1385_), .S0(new_n1960_), .Y(new_n2001_));
  MX2X1    g1359(.A(new_n801_), .B(new_n670_), .S0(new_n1969_), .Y(new_n2002_));
  INVX1    g1360(.A(new_n2002_), .Y(new_n2003_));
  MX2X1    g1361(.A(new_n1491_), .B(new_n1387_), .S0(new_n1960_), .Y(new_n2004_));
  INVX1    g1362(.A(new_n2004_), .Y(new_n2005_));
  MX2X1    g1363(.A(new_n797_), .B(new_n673_), .S0(new_n1969_), .Y(new_n2006_));
  MX2X1    g1364(.A(new_n675_), .B(new_n676_), .S0(new_n1969_), .Y(new_n2007_));
  INVX1    g1365(.A(new_n2007_), .Y(new_n2008_));
  MX2X1    g1366(.A(new_n677_), .B(new_n772_), .S0(new_n1969_), .Y(new_n2009_));
  MX2X1    g1367(.A(new_n1483_), .B(new_n1391_), .S0(new_n1960_), .Y(new_n2010_));
  INVX1    g1368(.A(new_n2010_), .Y(new_n2011_));
  MX2X1    g1369(.A(new_n767_), .B(new_n678_), .S0(new_n1969_), .Y(new_n2012_));
  MX2X1    g1370(.A(new_n1479_), .B(new_n1394_), .S0(new_n1960_), .Y(new_n2013_));
  MX2X1    g1371(.A(new_n764_), .B(new_n680_), .S0(new_n1969_), .Y(new_n2014_));
  INVX1    g1372(.A(new_n2014_), .Y(new_n2015_));
  MX2X1    g1373(.A(new_n1476_), .B(new_n1396_), .S0(new_n1960_), .Y(new_n2016_));
  INVX1    g1374(.A(new_n2016_), .Y(new_n2017_));
  MX2X1    g1375(.A(new_n760_), .B(new_n683_), .S0(new_n1969_), .Y(new_n2018_));
  MX2X1    g1376(.A(new_n1472_), .B(new_n1399_), .S0(new_n1960_), .Y(new_n2019_));
  MX2X1    g1377(.A(new_n757_), .B(new_n685_), .S0(new_n1969_), .Y(new_n2020_));
  INVX1    g1378(.A(new_n2020_), .Y(new_n2021_));
  MX2X1    g1379(.A(new_n1469_), .B(new_n1401_), .S0(new_n1960_), .Y(new_n2022_));
  INVX1    g1380(.A(new_n2022_), .Y(new_n2023_));
  MX2X1    g1381(.A(new_n753_), .B(new_n688_), .S0(new_n1969_), .Y(new_n2024_));
  MX2X1    g1382(.A(new_n1465_), .B(new_n1404_), .S0(new_n1960_), .Y(new_n2025_));
  MX2X1    g1383(.A(new_n750_), .B(new_n690_), .S0(new_n1969_), .Y(new_n2026_));
  INVX1    g1384(.A(new_n2026_), .Y(new_n2027_));
  MX2X1    g1385(.A(new_n776_), .B(new_n777_), .S0(new_n1969_), .Y(new_n2028_));
  MX2X1    g1386(.A(new_n778_), .B(new_n693_), .S0(new_n1969_), .Y(new_n2029_));
  INVX1    g1387(.A(new_n2029_), .Y(new_n2030_));
  MX2X1    g1388(.A(new_n1443_), .B(new_n1409_), .S0(new_n1960_), .Y(new_n2031_));
  MX2X1    g1389(.A(new_n733_), .B(new_n694_), .S0(new_n1969_), .Y(new_n2032_));
  INVX1    g1390(.A(new_n2032_), .Y(new_n2033_));
  MX2X1    g1391(.A(new_n729_), .B(new_n697_), .S0(new_n1969_), .Y(new_n2034_));
  MX2X1    g1392(.A(new_n1440_), .B(new_n1411_), .S0(new_n1960_), .Y(new_n2035_));
  INVX1    g1393(.A(new_n2035_), .Y(new_n2036_));
  MX2X1    g1394(.A(new_n699_), .B(new_n700_), .S0(new_n1969_), .Y(new_n2037_));
  INVX1    g1395(.A(new_n2037_), .Y(new_n2038_));
  MX2X1    g1396(.A(new_n1450_), .B(new_n1451_), .S0(new_n1960_), .Y(new_n2039_));
  INVX1    g1397(.A(new_n2039_), .Y(new_n2040_));
  MX2X1    g1398(.A(new_n701_), .B(new_n717_), .S0(new_n1969_), .Y(new_n2041_));
  INVX1    g1399(.A(new_n2041_), .Y(new_n2042_));
  MX2X1    g1400(.A(new_n1452_), .B(new_n1414_), .S0(new_n1960_), .Y(new_n2043_));
  MX2X1    g1401(.A(\in1[3] ), .B(\in0[3] ), .S0(new_n1960_), .Y(new_n2044_));
  MX2X1    g1402(.A(new_n712_), .B(new_n702_), .S0(new_n1969_), .Y(new_n2045_));
  OR2X1    g1403(.A(new_n2045_), .B(new_n2044_), .Y(new_n2046_));
  MX2X1    g1404(.A(new_n719_), .B(new_n705_), .S0(new_n1969_), .Y(new_n2047_));
  MX2X1    g1405(.A(new_n1418_), .B(new_n1429_), .S0(new_n1960_), .Y(new_n2048_));
  NOR3X1   g1406(.A(new_n2048_), .B(new_n1354_), .C(new_n1292_), .Y(new_n2049_));
  MX2X1    g1407(.A(\in1[1] ), .B(\in0[1] ), .S0(new_n1960_), .Y(new_n2050_));
  AOI21X1  g1408(.A0(new_n2049_), .A1(new_n2047_), .B0(new_n2050_), .Y(new_n2051_));
  MX2X1    g1409(.A(new_n1421_), .B(new_n1417_), .S0(new_n1960_), .Y(new_n2052_));
  MX2X1    g1410(.A(\in3[2] ), .B(\in2[2] ), .S0(new_n1969_), .Y(new_n2053_));
  MX2X1    g1411(.A(\in1[2] ), .B(\in0[2] ), .S0(new_n1960_), .Y(new_n2054_));
  MX2X1    g1412(.A(new_n704_), .B(new_n709_), .S0(new_n1969_), .Y(new_n2055_));
  OAI22X1  g1413(.A0(new_n2055_), .A1(new_n2054_), .B0(new_n2049_), .B1(new_n2047_), .Y(new_n2056_));
  OAI22X1  g1414(.A0(new_n2056_), .A1(new_n2051_), .B0(new_n2053_), .B1(new_n2052_), .Y(new_n2057_));
  AND2X1   g1415(.A(new_n2045_), .B(new_n2044_), .Y(new_n2058_));
  AOI21X1  g1416(.A0(new_n2057_), .A1(new_n2046_), .B0(new_n2058_), .Y(new_n2059_));
  AOI21X1  g1417(.A0(new_n2059_), .A1(new_n2043_), .B0(new_n2042_), .Y(new_n2060_));
  INVX1    g1418(.A(new_n2043_), .Y(new_n2061_));
  NOR2X1   g1419(.A(new_n2045_), .B(new_n2044_), .Y(new_n2062_));
  MX2X1    g1420(.A(\in3[1] ), .B(\in2[1] ), .S0(new_n1969_), .Y(new_n2063_));
  NAND3X1  g1421(.A(new_n1353_), .B(new_n1352_), .C(\in3[0] ), .Y(new_n2064_));
  OAI21X1  g1422(.A0(new_n1291_), .A1(new_n1289_), .B0(\in2[0] ), .Y(new_n2065_));
  NAND3X1  g1423(.A(new_n1961_), .B(new_n2065_), .C(new_n2064_), .Y(new_n2066_));
  MX2X1    g1424(.A(new_n1419_), .B(new_n1430_), .S0(new_n1960_), .Y(new_n2067_));
  OAI21X1  g1425(.A0(new_n2066_), .A1(new_n2063_), .B0(new_n2067_), .Y(new_n2068_));
  AOI22X1  g1426(.A0(new_n2053_), .A1(new_n2052_), .B0(new_n2066_), .B1(new_n2063_), .Y(new_n2069_));
  AOI22X1  g1427(.A0(new_n2069_), .A1(new_n2068_), .B0(new_n2055_), .B1(new_n2054_), .Y(new_n2070_));
  NAND2X1  g1428(.A(new_n2045_), .B(new_n2044_), .Y(new_n2071_));
  OAI21X1  g1429(.A0(new_n2070_), .A1(new_n2062_), .B0(new_n2071_), .Y(new_n2072_));
  AND2X1   g1430(.A(new_n2072_), .B(new_n2061_), .Y(new_n2073_));
  NOR3X1   g1431(.A(new_n2073_), .B(new_n2060_), .C(new_n2040_), .Y(new_n2074_));
  OAI21X1  g1432(.A0(new_n2073_), .A1(new_n2060_), .B0(new_n2040_), .Y(new_n2075_));
  OAI21X1  g1433(.A0(new_n2074_), .A1(new_n2038_), .B0(new_n2075_), .Y(new_n2076_));
  OAI21X1  g1434(.A0(new_n2076_), .A1(new_n2036_), .B0(new_n2034_), .Y(new_n2077_));
  NAND2X1  g1435(.A(new_n2076_), .B(new_n2036_), .Y(new_n2078_));
  AOI22X1  g1436(.A0(new_n2078_), .A1(new_n2077_), .B0(new_n2033_), .B1(new_n2031_), .Y(new_n2079_));
  INVX1    g1437(.A(new_n2031_), .Y(new_n2080_));
  AND2X1   g1438(.A(new_n2032_), .B(new_n2080_), .Y(new_n2081_));
  MX2X1    g1439(.A(new_n1408_), .B(new_n1448_), .S0(new_n1960_), .Y(new_n2082_));
  INVX1    g1440(.A(new_n2082_), .Y(new_n2083_));
  NOR3X1   g1441(.A(new_n2083_), .B(new_n2081_), .C(new_n2079_), .Y(new_n2084_));
  OAI21X1  g1442(.A0(new_n2081_), .A1(new_n2079_), .B0(new_n2083_), .Y(new_n2085_));
  OAI21X1  g1443(.A0(new_n2084_), .A1(new_n2030_), .B0(new_n2085_), .Y(new_n2086_));
  MX2X1    g1444(.A(new_n1406_), .B(new_n1407_), .S0(new_n1960_), .Y(new_n2087_));
  INVX1    g1445(.A(new_n2087_), .Y(new_n2088_));
  OAI21X1  g1446(.A0(new_n2088_), .A1(new_n2086_), .B0(new_n2028_), .Y(new_n2089_));
  NAND2X1  g1447(.A(new_n2088_), .B(new_n2086_), .Y(new_n2090_));
  AOI22X1  g1448(.A0(new_n2090_), .A1(new_n2089_), .B0(new_n2027_), .B1(new_n2025_), .Y(new_n2091_));
  INVX1    g1449(.A(new_n2025_), .Y(new_n2092_));
  AND2X1   g1450(.A(new_n2026_), .B(new_n2092_), .Y(new_n2093_));
  OAI22X1  g1451(.A0(new_n2093_), .A1(new_n2091_), .B0(new_n2024_), .B1(new_n2023_), .Y(new_n2094_));
  AND2X1   g1452(.A(new_n2024_), .B(new_n2023_), .Y(new_n2095_));
  INVX1    g1453(.A(new_n2095_), .Y(new_n2096_));
  AOI22X1  g1454(.A0(new_n2096_), .A1(new_n2094_), .B0(new_n2021_), .B1(new_n2019_), .Y(new_n2097_));
  INVX1    g1455(.A(new_n2019_), .Y(new_n2098_));
  AND2X1   g1456(.A(new_n2020_), .B(new_n2098_), .Y(new_n2099_));
  OAI22X1  g1457(.A0(new_n2099_), .A1(new_n2097_), .B0(new_n2018_), .B1(new_n2017_), .Y(new_n2100_));
  AND2X1   g1458(.A(new_n2018_), .B(new_n2017_), .Y(new_n2101_));
  INVX1    g1459(.A(new_n2101_), .Y(new_n2102_));
  AOI22X1  g1460(.A0(new_n2102_), .A1(new_n2100_), .B0(new_n2015_), .B1(new_n2013_), .Y(new_n2103_));
  INVX1    g1461(.A(new_n2013_), .Y(new_n2104_));
  AND2X1   g1462(.A(new_n2014_), .B(new_n2104_), .Y(new_n2105_));
  OAI22X1  g1463(.A0(new_n2105_), .A1(new_n2103_), .B0(new_n2012_), .B1(new_n2011_), .Y(new_n2106_));
  AND2X1   g1464(.A(new_n2012_), .B(new_n2011_), .Y(new_n2107_));
  INVX1    g1465(.A(new_n2107_), .Y(new_n2108_));
  MX2X1    g1466(.A(\in1[16] ), .B(\in0[16] ), .S0(new_n1960_), .Y(new_n2109_));
  INVX1    g1467(.A(new_n2109_), .Y(new_n2110_));
  NAND3X1  g1468(.A(new_n2110_), .B(new_n2108_), .C(new_n2106_), .Y(new_n2111_));
  AOI21X1  g1469(.A0(new_n2108_), .A1(new_n2106_), .B0(new_n2110_), .Y(new_n2112_));
  AOI21X1  g1470(.A0(new_n2111_), .A1(new_n2009_), .B0(new_n2112_), .Y(new_n2113_));
  MX2X1    g1471(.A(\in1[17] ), .B(\in0[17] ), .S0(new_n1960_), .Y(new_n2114_));
  INVX1    g1472(.A(new_n2114_), .Y(new_n2115_));
  AOI21X1  g1473(.A0(new_n2115_), .A1(new_n2113_), .B0(new_n2008_), .Y(new_n2116_));
  NOR2X1   g1474(.A(new_n2115_), .B(new_n2113_), .Y(new_n2117_));
  OAI22X1  g1475(.A0(new_n2117_), .A1(new_n2116_), .B0(new_n2006_), .B1(new_n2005_), .Y(new_n2118_));
  AND2X1   g1476(.A(new_n2006_), .B(new_n2005_), .Y(new_n2119_));
  INVX1    g1477(.A(new_n2119_), .Y(new_n2120_));
  AOI22X1  g1478(.A0(new_n2120_), .A1(new_n2118_), .B0(new_n2003_), .B1(new_n2001_), .Y(new_n2121_));
  INVX1    g1479(.A(new_n2001_), .Y(new_n2122_));
  AND2X1   g1480(.A(new_n2002_), .B(new_n2122_), .Y(new_n2123_));
  OAI22X1  g1481(.A0(new_n2123_), .A1(new_n2121_), .B0(new_n2000_), .B1(new_n1999_), .Y(new_n2124_));
  AND2X1   g1482(.A(new_n2000_), .B(new_n1999_), .Y(new_n2125_));
  INVX1    g1483(.A(new_n2125_), .Y(new_n2126_));
  AOI22X1  g1484(.A0(new_n2126_), .A1(new_n2124_), .B0(new_n1997_), .B1(new_n1995_), .Y(new_n2127_));
  INVX1    g1485(.A(new_n1995_), .Y(new_n2128_));
  AND2X1   g1486(.A(new_n1996_), .B(new_n2128_), .Y(new_n2129_));
  OAI22X1  g1487(.A0(new_n2129_), .A1(new_n2127_), .B0(new_n1994_), .B1(new_n1993_), .Y(new_n2130_));
  AND2X1   g1488(.A(new_n1994_), .B(new_n1993_), .Y(new_n2131_));
  INVX1    g1489(.A(new_n2131_), .Y(new_n2132_));
  AOI22X1  g1490(.A0(new_n2132_), .A1(new_n2130_), .B0(new_n1991_), .B1(new_n1989_), .Y(new_n2133_));
  INVX1    g1491(.A(new_n1989_), .Y(new_n2134_));
  AND2X1   g1492(.A(new_n1990_), .B(new_n2134_), .Y(new_n2135_));
  MX2X1    g1493(.A(\in1[24] ), .B(\in0[24] ), .S0(new_n1960_), .Y(new_n2136_));
  NOR3X1   g1494(.A(new_n2136_), .B(new_n2135_), .C(new_n2133_), .Y(new_n2137_));
  OAI21X1  g1495(.A0(new_n2135_), .A1(new_n2133_), .B0(new_n2136_), .Y(new_n2138_));
  OAI21X1  g1496(.A0(new_n2137_), .A1(new_n1988_), .B0(new_n2138_), .Y(new_n2139_));
  MX2X1    g1497(.A(new_n1372_), .B(new_n1373_), .S0(new_n1960_), .Y(new_n2140_));
  INVX1    g1498(.A(new_n2140_), .Y(new_n2141_));
  OAI21X1  g1499(.A0(new_n2141_), .A1(new_n2139_), .B0(new_n1986_), .Y(new_n2142_));
  NAND2X1  g1500(.A(new_n2141_), .B(new_n2139_), .Y(new_n2143_));
  AOI22X1  g1501(.A0(new_n2143_), .A1(new_n2142_), .B0(new_n1985_), .B1(new_n1983_), .Y(new_n2144_));
  INVX1    g1502(.A(new_n1983_), .Y(new_n2145_));
  AND2X1   g1503(.A(new_n1984_), .B(new_n2145_), .Y(new_n2146_));
  OAI22X1  g1504(.A0(new_n2146_), .A1(new_n2144_), .B0(new_n1982_), .B1(new_n1981_), .Y(new_n2147_));
  AND2X1   g1505(.A(new_n1982_), .B(new_n1981_), .Y(new_n2148_));
  INVX1    g1506(.A(new_n2148_), .Y(new_n2149_));
  AOI22X1  g1507(.A0(new_n2149_), .A1(new_n2147_), .B0(new_n1979_), .B1(new_n1977_), .Y(new_n2150_));
  INVX1    g1508(.A(new_n1977_), .Y(new_n2151_));
  AND2X1   g1509(.A(new_n1978_), .B(new_n2151_), .Y(new_n2152_));
  OAI22X1  g1510(.A0(new_n2152_), .A1(new_n2150_), .B0(new_n1976_), .B1(new_n1975_), .Y(new_n2153_));
  AND2X1   g1511(.A(new_n1976_), .B(new_n1975_), .Y(new_n2154_));
  INVX1    g1512(.A(new_n2154_), .Y(new_n2155_));
  AOI22X1  g1513(.A0(new_n2155_), .A1(new_n2153_), .B0(new_n1973_), .B1(new_n1971_), .Y(new_n2156_));
  INVX1    g1514(.A(new_n1971_), .Y(new_n2157_));
  AND2X1   g1515(.A(new_n1972_), .B(new_n2157_), .Y(new_n2158_));
  OAI22X1  g1516(.A0(new_n2158_), .A1(new_n2156_), .B0(new_n1970_), .B1(new_n1968_), .Y(new_n2159_));
  AND2X1   g1517(.A(new_n1970_), .B(new_n1968_), .Y(new_n2160_));
  INVX1    g1518(.A(new_n2160_), .Y(new_n2161_));
  MX2X1    g1519(.A(new_n879_), .B(new_n868_), .S0(new_n1969_), .Y(new_n2162_));
  MX2X1    g1520(.A(\in1[34] ), .B(\in0[34] ), .S0(new_n1960_), .Y(new_n2163_));
  NOR2X1   g1521(.A(new_n2163_), .B(new_n2162_), .Y(new_n2164_));
  MX2X1    g1522(.A(new_n1550_), .B(new_n1556_), .S0(new_n1960_), .Y(new_n2165_));
  INVX1    g1523(.A(new_n2165_), .Y(new_n2166_));
  INVX1    g1524(.A(\in2[33] ), .Y(new_n2167_));
  MX2X1    g1525(.A(new_n873_), .B(new_n2167_), .S0(new_n1969_), .Y(new_n2168_));
  MX2X1    g1526(.A(\in1[35] ), .B(\in0[35] ), .S0(new_n1960_), .Y(new_n2169_));
  MX2X1    g1527(.A(\in3[35] ), .B(\in2[35] ), .S0(new_n1969_), .Y(new_n2170_));
  INVX1    g1528(.A(new_n2170_), .Y(new_n2171_));
  OAI22X1  g1529(.A0(new_n2171_), .A1(new_n2169_), .B0(new_n2168_), .B1(new_n2166_), .Y(new_n2172_));
  NOR2X1   g1530(.A(new_n2172_), .B(new_n2164_), .Y(new_n2173_));
  INVX1    g1531(.A(new_n2173_), .Y(new_n2174_));
  INVX1    g1532(.A(\in2[32] ), .Y(new_n2175_));
  MX2X1    g1533(.A(new_n872_), .B(new_n2175_), .S0(new_n1969_), .Y(new_n2176_));
  MX2X1    g1534(.A(new_n1549_), .B(new_n1555_), .S0(new_n1960_), .Y(new_n2177_));
  INVX1    g1535(.A(new_n2177_), .Y(new_n2178_));
  NOR2X1   g1536(.A(new_n2178_), .B(new_n2176_), .Y(new_n2179_));
  MX2X1    g1537(.A(\in1[39] ), .B(\in0[39] ), .S0(new_n1960_), .Y(new_n2180_));
  MX2X1    g1538(.A(new_n888_), .B(new_n862_), .S0(new_n1969_), .Y(new_n2181_));
  NOR2X1   g1539(.A(new_n2181_), .B(new_n2180_), .Y(new_n2182_));
  MX2X1    g1540(.A(\in3[38] ), .B(\in2[38] ), .S0(new_n1969_), .Y(new_n2183_));
  MX2X1    g1541(.A(\in1[38] ), .B(\in0[38] ), .S0(new_n1960_), .Y(new_n2184_));
  INVX1    g1542(.A(new_n2184_), .Y(new_n2185_));
  AOI21X1  g1543(.A0(new_n2185_), .A1(new_n2183_), .B0(new_n2182_), .Y(new_n2186_));
  INVX1    g1544(.A(new_n2186_), .Y(new_n2187_));
  MX2X1    g1545(.A(new_n1542_), .B(new_n1563_), .S0(new_n1960_), .Y(new_n2188_));
  INVX1    g1546(.A(new_n2188_), .Y(new_n2189_));
  MX2X1    g1547(.A(new_n865_), .B(new_n883_), .S0(new_n1969_), .Y(new_n2190_));
  MX2X1    g1548(.A(\in1[37] ), .B(\in0[37] ), .S0(new_n1960_), .Y(new_n2191_));
  MX2X1    g1549(.A(new_n866_), .B(new_n884_), .S0(new_n1969_), .Y(new_n2192_));
  OAI22X1  g1550(.A0(new_n2192_), .A1(new_n2191_), .B0(new_n2190_), .B1(new_n2189_), .Y(new_n2193_));
  NOR4X1   g1551(.A(new_n2193_), .B(new_n2187_), .C(new_n2179_), .D(new_n2174_), .Y(new_n2194_));
  INVX1    g1552(.A(new_n2194_), .Y(new_n2195_));
  AOI21X1  g1553(.A0(new_n2161_), .A1(new_n2159_), .B0(new_n2195_), .Y(new_n2196_));
  NOR2X1   g1554(.A(new_n2193_), .B(new_n2187_), .Y(new_n2197_));
  AOI22X1  g1555(.A0(new_n2178_), .A1(new_n2176_), .B0(new_n2168_), .B1(new_n2166_), .Y(new_n2198_));
  AND2X1   g1556(.A(new_n2171_), .B(new_n2169_), .Y(new_n2199_));
  INVX1    g1557(.A(new_n2199_), .Y(new_n2200_));
  AND2X1   g1558(.A(new_n2163_), .B(new_n2162_), .Y(new_n2201_));
  OAI21X1  g1559(.A0(new_n2171_), .A1(new_n2169_), .B0(new_n2201_), .Y(new_n2202_));
  AND2X1   g1560(.A(new_n2202_), .B(new_n2200_), .Y(new_n2203_));
  OAI21X1  g1561(.A0(new_n2198_), .A1(new_n2174_), .B0(new_n2203_), .Y(new_n2204_));
  OR2X1    g1562(.A(new_n2192_), .B(new_n2191_), .Y(new_n2205_));
  AND2X1   g1563(.A(new_n2190_), .B(new_n2189_), .Y(new_n2206_));
  AND2X1   g1564(.A(new_n2192_), .B(new_n2191_), .Y(new_n2207_));
  AOI21X1  g1565(.A0(new_n2206_), .A1(new_n2205_), .B0(new_n2207_), .Y(new_n2208_));
  OR2X1    g1566(.A(new_n2185_), .B(new_n2183_), .Y(new_n2209_));
  NOR2X1   g1567(.A(new_n2209_), .B(new_n2182_), .Y(new_n2210_));
  AOI21X1  g1568(.A0(new_n2181_), .A1(new_n2180_), .B0(new_n2210_), .Y(new_n2211_));
  OAI21X1  g1569(.A0(new_n2208_), .A1(new_n2187_), .B0(new_n2211_), .Y(new_n2212_));
  AOI21X1  g1570(.A0(new_n2204_), .A1(new_n2197_), .B0(new_n2212_), .Y(new_n2213_));
  INVX1    g1571(.A(new_n2213_), .Y(new_n2214_));
  MX2X1    g1572(.A(\in1[47] ), .B(\in0[47] ), .S0(new_n1960_), .Y(new_n2215_));
  MX2X1    g1573(.A(new_n924_), .B(new_n897_), .S0(new_n1969_), .Y(new_n2216_));
  NOR2X1   g1574(.A(new_n2216_), .B(new_n2215_), .Y(new_n2217_));
  MX2X1    g1575(.A(\in3[46] ), .B(\in2[46] ), .S0(new_n1969_), .Y(new_n2218_));
  MX2X1    g1576(.A(\in1[46] ), .B(\in0[46] ), .S0(new_n1960_), .Y(new_n2219_));
  INVX1    g1577(.A(new_n2219_), .Y(new_n2220_));
  AND2X1   g1578(.A(new_n2220_), .B(new_n2218_), .Y(new_n2221_));
  OR2X1    g1579(.A(new_n2221_), .B(new_n2217_), .Y(new_n2222_));
  MX2X1    g1580(.A(\in1[44] ), .B(\in0[44] ), .S0(new_n1960_), .Y(new_n2223_));
  MX2X1    g1581(.A(new_n900_), .B(new_n919_), .S0(new_n1969_), .Y(new_n2224_));
  MX2X1    g1582(.A(\in1[45] ), .B(\in0[45] ), .S0(new_n1960_), .Y(new_n2225_));
  MX2X1    g1583(.A(new_n901_), .B(new_n920_), .S0(new_n1969_), .Y(new_n2226_));
  OAI22X1  g1584(.A0(new_n2226_), .A1(new_n2225_), .B0(new_n2224_), .B1(new_n2223_), .Y(new_n2227_));
  MX2X1    g1585(.A(\in1[43] ), .B(\in0[43] ), .S0(new_n1960_), .Y(new_n2228_));
  MX2X1    g1586(.A(\in3[43] ), .B(\in2[43] ), .S0(new_n1969_), .Y(new_n2229_));
  INVX1    g1587(.A(new_n2229_), .Y(new_n2230_));
  MX2X1    g1588(.A(new_n1592_), .B(new_n1581_), .S0(new_n1960_), .Y(new_n2231_));
  INVX1    g1589(.A(new_n2231_), .Y(new_n2232_));
  MX2X1    g1590(.A(new_n915_), .B(new_n903_), .S0(new_n1969_), .Y(new_n2233_));
  OAI22X1  g1591(.A0(new_n2233_), .A1(new_n2232_), .B0(new_n2230_), .B1(new_n2228_), .Y(new_n2234_));
  INVX1    g1592(.A(\in0[41] ), .Y(new_n2235_));
  MX2X1    g1593(.A(new_n1586_), .B(new_n2235_), .S0(new_n1960_), .Y(new_n2236_));
  INVX1    g1594(.A(new_n2236_), .Y(new_n2237_));
  INVX1    g1595(.A(\in2[41] ), .Y(new_n2238_));
  MX2X1    g1596(.A(new_n908_), .B(new_n2238_), .S0(new_n1969_), .Y(new_n2239_));
  INVX1    g1597(.A(\in0[40] ), .Y(new_n2240_));
  MX2X1    g1598(.A(new_n1585_), .B(new_n2240_), .S0(new_n1960_), .Y(new_n2241_));
  INVX1    g1599(.A(new_n2241_), .Y(new_n2242_));
  INVX1    g1600(.A(\in2[40] ), .Y(new_n2243_));
  MX2X1    g1601(.A(new_n907_), .B(new_n2243_), .S0(new_n1969_), .Y(new_n2244_));
  OAI22X1  g1602(.A0(new_n2244_), .A1(new_n2242_), .B0(new_n2239_), .B1(new_n2237_), .Y(new_n2245_));
  NOR4X1   g1603(.A(new_n2245_), .B(new_n2234_), .C(new_n2227_), .D(new_n2222_), .Y(new_n2246_));
  OAI21X1  g1604(.A0(new_n2214_), .A1(new_n2196_), .B0(new_n2246_), .Y(new_n2247_));
  NOR3X1   g1605(.A(new_n2227_), .B(new_n2221_), .C(new_n2217_), .Y(new_n2248_));
  NAND2X1  g1606(.A(new_n2230_), .B(new_n2228_), .Y(new_n2249_));
  NOR2X1   g1607(.A(new_n2239_), .B(new_n2237_), .Y(new_n2250_));
  INVX1    g1608(.A(new_n2244_), .Y(new_n2251_));
  NOR3X1   g1609(.A(new_n2251_), .B(new_n2241_), .C(new_n2250_), .Y(new_n2252_));
  INVX1    g1610(.A(new_n2233_), .Y(new_n2253_));
  INVX1    g1611(.A(new_n2239_), .Y(new_n2254_));
  OAI22X1  g1612(.A0(new_n2254_), .A1(new_n2236_), .B0(new_n2253_), .B1(new_n2231_), .Y(new_n2255_));
  NOR2X1   g1613(.A(new_n2255_), .B(new_n2252_), .Y(new_n2256_));
  OAI21X1  g1614(.A0(new_n2256_), .A1(new_n2234_), .B0(new_n2249_), .Y(new_n2257_));
  AND2X1   g1615(.A(new_n2257_), .B(new_n2248_), .Y(new_n2258_));
  OR2X1    g1616(.A(new_n2226_), .B(new_n2225_), .Y(new_n2259_));
  NAND3X1  g1617(.A(new_n2259_), .B(new_n2224_), .C(new_n2223_), .Y(new_n2260_));
  NAND2X1  g1618(.A(new_n2226_), .B(new_n2225_), .Y(new_n2261_));
  AOI21X1  g1619(.A0(new_n2261_), .A1(new_n2260_), .B0(new_n2222_), .Y(new_n2262_));
  AND2X1   g1620(.A(new_n2216_), .B(new_n2215_), .Y(new_n2263_));
  NOR3X1   g1621(.A(new_n2220_), .B(new_n2218_), .C(new_n2217_), .Y(new_n2264_));
  NOR4X1   g1622(.A(new_n2264_), .B(new_n2263_), .C(new_n2262_), .D(new_n2258_), .Y(new_n2265_));
  MX2X1    g1623(.A(new_n949_), .B(new_n938_), .S0(new_n1969_), .Y(new_n2266_));
  MX2X1    g1624(.A(\in1[50] ), .B(\in0[50] ), .S0(new_n1960_), .Y(new_n2267_));
  NOR2X1   g1625(.A(new_n2267_), .B(new_n2266_), .Y(new_n2268_));
  MX2X1    g1626(.A(new_n1621_), .B(new_n1627_), .S0(new_n1960_), .Y(new_n2269_));
  INVX1    g1627(.A(new_n2269_), .Y(new_n2270_));
  INVX1    g1628(.A(\in2[49] ), .Y(new_n2271_));
  MX2X1    g1629(.A(new_n943_), .B(new_n2271_), .S0(new_n1969_), .Y(new_n2272_));
  MX2X1    g1630(.A(\in1[51] ), .B(\in0[51] ), .S0(new_n1960_), .Y(new_n2273_));
  MX2X1    g1631(.A(\in3[51] ), .B(\in2[51] ), .S0(new_n1969_), .Y(new_n2274_));
  INVX1    g1632(.A(new_n2274_), .Y(new_n2275_));
  OAI22X1  g1633(.A0(new_n2275_), .A1(new_n2273_), .B0(new_n2272_), .B1(new_n2270_), .Y(new_n2276_));
  NOR2X1   g1634(.A(new_n2276_), .B(new_n2268_), .Y(new_n2277_));
  INVX1    g1635(.A(new_n2277_), .Y(new_n2278_));
  INVX1    g1636(.A(\in2[48] ), .Y(new_n2279_));
  MX2X1    g1637(.A(new_n942_), .B(new_n2279_), .S0(new_n1969_), .Y(new_n2280_));
  MX2X1    g1638(.A(new_n1620_), .B(new_n1626_), .S0(new_n1960_), .Y(new_n2281_));
  INVX1    g1639(.A(new_n2281_), .Y(new_n2282_));
  NOR2X1   g1640(.A(new_n2282_), .B(new_n2280_), .Y(new_n2283_));
  MX2X1    g1641(.A(\in1[55] ), .B(\in0[55] ), .S0(new_n1960_), .Y(new_n2284_));
  INVX1    g1642(.A(new_n2284_), .Y(new_n2285_));
  MX2X1    g1643(.A(\in3[55] ), .B(\in2[55] ), .S0(new_n1969_), .Y(new_n2286_));
  MX2X1    g1644(.A(new_n955_), .B(new_n931_), .S0(new_n1969_), .Y(new_n2287_));
  INVX1    g1645(.A(new_n2287_), .Y(new_n2288_));
  MX2X1    g1646(.A(new_n1635_), .B(new_n1609_), .S0(new_n1960_), .Y(new_n2289_));
  AOI22X1  g1647(.A0(new_n2289_), .A1(new_n2288_), .B0(new_n2286_), .B1(new_n2285_), .Y(new_n2290_));
  INVX1    g1648(.A(new_n2290_), .Y(new_n2291_));
  INVX1    g1649(.A(\in0[53] ), .Y(new_n2292_));
  MX2X1    g1650(.A(new_n1614_), .B(new_n2292_), .S0(new_n1960_), .Y(new_n2293_));
  INVX1    g1651(.A(new_n2293_), .Y(new_n2294_));
  INVX1    g1652(.A(\in2[53] ), .Y(new_n2295_));
  MX2X1    g1653(.A(new_n936_), .B(new_n2295_), .S0(new_n1969_), .Y(new_n2296_));
  INVX1    g1654(.A(\in2[52] ), .Y(new_n2297_));
  MX2X1    g1655(.A(new_n935_), .B(new_n2297_), .S0(new_n1969_), .Y(new_n2298_));
  INVX1    g1656(.A(\in0[52] ), .Y(new_n2299_));
  MX2X1    g1657(.A(new_n1613_), .B(new_n2299_), .S0(new_n1960_), .Y(new_n2300_));
  INVX1    g1658(.A(new_n2300_), .Y(new_n2301_));
  OAI22X1  g1659(.A0(new_n2301_), .A1(new_n2298_), .B0(new_n2296_), .B1(new_n2294_), .Y(new_n2302_));
  NOR4X1   g1660(.A(new_n2302_), .B(new_n2291_), .C(new_n2283_), .D(new_n2278_), .Y(new_n2303_));
  INVX1    g1661(.A(new_n2303_), .Y(new_n2304_));
  AOI21X1  g1662(.A0(new_n2265_), .A1(new_n2247_), .B0(new_n2304_), .Y(new_n2305_));
  NOR2X1   g1663(.A(new_n2302_), .B(new_n2291_), .Y(new_n2306_));
  AOI22X1  g1664(.A0(new_n2282_), .A1(new_n2280_), .B0(new_n2272_), .B1(new_n2270_), .Y(new_n2307_));
  AND2X1   g1665(.A(new_n2275_), .B(new_n2273_), .Y(new_n2308_));
  INVX1    g1666(.A(new_n2308_), .Y(new_n2309_));
  AND2X1   g1667(.A(new_n2267_), .B(new_n2266_), .Y(new_n2310_));
  OAI21X1  g1668(.A0(new_n2275_), .A1(new_n2273_), .B0(new_n2310_), .Y(new_n2311_));
  AND2X1   g1669(.A(new_n2311_), .B(new_n2309_), .Y(new_n2312_));
  OAI21X1  g1670(.A0(new_n2307_), .A1(new_n2278_), .B0(new_n2312_), .Y(new_n2313_));
  NOR2X1   g1671(.A(new_n2286_), .B(new_n2285_), .Y(new_n2314_));
  NOR2X1   g1672(.A(new_n2296_), .B(new_n2294_), .Y(new_n2315_));
  NAND2X1  g1673(.A(new_n2301_), .B(new_n2298_), .Y(new_n2316_));
  INVX1    g1674(.A(new_n2289_), .Y(new_n2317_));
  AOI22X1  g1675(.A0(new_n2296_), .A1(new_n2294_), .B0(new_n2317_), .B1(new_n2287_), .Y(new_n2318_));
  OAI21X1  g1676(.A0(new_n2316_), .A1(new_n2315_), .B0(new_n2318_), .Y(new_n2319_));
  AOI21X1  g1677(.A0(new_n2319_), .A1(new_n2290_), .B0(new_n2314_), .Y(new_n2320_));
  INVX1    g1678(.A(new_n2320_), .Y(new_n2321_));
  AOI21X1  g1679(.A0(new_n2313_), .A1(new_n2306_), .B0(new_n2321_), .Y(new_n2322_));
  INVX1    g1680(.A(new_n2322_), .Y(new_n2323_));
  MX2X1    g1681(.A(\in1[63] ), .B(\in0[63] ), .S0(new_n1960_), .Y(new_n2324_));
  MX2X1    g1682(.A(new_n990_), .B(new_n963_), .S0(new_n1969_), .Y(new_n2325_));
  NOR2X1   g1683(.A(new_n2325_), .B(new_n2324_), .Y(new_n2326_));
  MX2X1    g1684(.A(\in3[62] ), .B(\in2[62] ), .S0(new_n1969_), .Y(new_n2327_));
  MX2X1    g1685(.A(\in1[62] ), .B(\in0[62] ), .S0(new_n1960_), .Y(new_n2328_));
  INVX1    g1686(.A(new_n2328_), .Y(new_n2329_));
  AND2X1   g1687(.A(new_n2329_), .B(new_n2327_), .Y(new_n2330_));
  OR2X1    g1688(.A(new_n2330_), .B(new_n2326_), .Y(new_n2331_));
  MX2X1    g1689(.A(\in1[60] ), .B(\in0[60] ), .S0(new_n1960_), .Y(new_n2332_));
  MX2X1    g1690(.A(new_n966_), .B(new_n985_), .S0(new_n1969_), .Y(new_n2333_));
  MX2X1    g1691(.A(\in1[61] ), .B(\in0[61] ), .S0(new_n1960_), .Y(new_n2334_));
  MX2X1    g1692(.A(new_n967_), .B(new_n986_), .S0(new_n1969_), .Y(new_n2335_));
  OAI22X1  g1693(.A0(new_n2335_), .A1(new_n2334_), .B0(new_n2333_), .B1(new_n2332_), .Y(new_n2336_));
  MX2X1    g1694(.A(\in1[59] ), .B(\in0[59] ), .S0(new_n1960_), .Y(new_n2337_));
  MX2X1    g1695(.A(\in3[59] ), .B(\in2[59] ), .S0(new_n1969_), .Y(new_n2338_));
  INVX1    g1696(.A(new_n2338_), .Y(new_n2339_));
  MX2X1    g1697(.A(new_n1659_), .B(new_n1648_), .S0(new_n1960_), .Y(new_n2340_));
  INVX1    g1698(.A(new_n2340_), .Y(new_n2341_));
  MX2X1    g1699(.A(new_n981_), .B(new_n969_), .S0(new_n1969_), .Y(new_n2342_));
  OAI22X1  g1700(.A0(new_n2342_), .A1(new_n2341_), .B0(new_n2339_), .B1(new_n2337_), .Y(new_n2343_));
  INVX1    g1701(.A(\in0[57] ), .Y(new_n2344_));
  MX2X1    g1702(.A(new_n1653_), .B(new_n2344_), .S0(new_n1960_), .Y(new_n2345_));
  INVX1    g1703(.A(new_n2345_), .Y(new_n2346_));
  INVX1    g1704(.A(\in2[57] ), .Y(new_n2347_));
  MX2X1    g1705(.A(new_n974_), .B(new_n2347_), .S0(new_n1969_), .Y(new_n2348_));
  INVX1    g1706(.A(\in0[56] ), .Y(new_n2349_));
  MX2X1    g1707(.A(new_n1652_), .B(new_n2349_), .S0(new_n1960_), .Y(new_n2350_));
  INVX1    g1708(.A(new_n2350_), .Y(new_n2351_));
  INVX1    g1709(.A(\in2[56] ), .Y(new_n2352_));
  MX2X1    g1710(.A(new_n973_), .B(new_n2352_), .S0(new_n1969_), .Y(new_n2353_));
  OAI22X1  g1711(.A0(new_n2353_), .A1(new_n2351_), .B0(new_n2348_), .B1(new_n2346_), .Y(new_n2354_));
  NOR4X1   g1712(.A(new_n2354_), .B(new_n2343_), .C(new_n2336_), .D(new_n2331_), .Y(new_n2355_));
  OAI21X1  g1713(.A0(new_n2323_), .A1(new_n2305_), .B0(new_n2355_), .Y(new_n2356_));
  NOR3X1   g1714(.A(new_n2336_), .B(new_n2330_), .C(new_n2326_), .Y(new_n2357_));
  NAND2X1  g1715(.A(new_n2339_), .B(new_n2337_), .Y(new_n2358_));
  NOR2X1   g1716(.A(new_n2348_), .B(new_n2346_), .Y(new_n2359_));
  INVX1    g1717(.A(new_n2353_), .Y(new_n2360_));
  NOR3X1   g1718(.A(new_n2360_), .B(new_n2350_), .C(new_n2359_), .Y(new_n2361_));
  INVX1    g1719(.A(new_n2342_), .Y(new_n2362_));
  INVX1    g1720(.A(new_n2348_), .Y(new_n2363_));
  OAI22X1  g1721(.A0(new_n2363_), .A1(new_n2345_), .B0(new_n2362_), .B1(new_n2340_), .Y(new_n2364_));
  NOR2X1   g1722(.A(new_n2364_), .B(new_n2361_), .Y(new_n2365_));
  OAI21X1  g1723(.A0(new_n2365_), .A1(new_n2343_), .B0(new_n2358_), .Y(new_n2366_));
  AND2X1   g1724(.A(new_n2366_), .B(new_n2357_), .Y(new_n2367_));
  OR2X1    g1725(.A(new_n2335_), .B(new_n2334_), .Y(new_n2368_));
  NAND3X1  g1726(.A(new_n2368_), .B(new_n2333_), .C(new_n2332_), .Y(new_n2369_));
  NAND2X1  g1727(.A(new_n2335_), .B(new_n2334_), .Y(new_n2370_));
  AOI21X1  g1728(.A0(new_n2370_), .A1(new_n2369_), .B0(new_n2331_), .Y(new_n2371_));
  AND2X1   g1729(.A(new_n2325_), .B(new_n2324_), .Y(new_n2372_));
  NOR3X1   g1730(.A(new_n2329_), .B(new_n2327_), .C(new_n2326_), .Y(new_n2373_));
  NOR4X1   g1731(.A(new_n2373_), .B(new_n2372_), .C(new_n2371_), .D(new_n2367_), .Y(new_n2374_));
  MX2X1    g1732(.A(\in1[67] ), .B(\in0[67] ), .S0(new_n1960_), .Y(new_n2375_));
  INVX1    g1733(.A(new_n2375_), .Y(new_n2376_));
  MX2X1    g1734(.A(\in3[67] ), .B(\in2[67] ), .S0(new_n1969_), .Y(new_n2377_));
  MX2X1    g1735(.A(new_n1008_), .B(new_n997_), .S0(new_n1969_), .Y(new_n2378_));
  INVX1    g1736(.A(new_n2378_), .Y(new_n2379_));
  MX2X1    g1737(.A(new_n1688_), .B(new_n1676_), .S0(new_n1960_), .Y(new_n2380_));
  AOI22X1  g1738(.A0(new_n2380_), .A1(new_n2379_), .B0(new_n2377_), .B1(new_n2376_), .Y(new_n2381_));
  MX2X1    g1739(.A(\in3[64] ), .B(\in2[64] ), .S0(new_n1969_), .Y(new_n2382_));
  MX2X1    g1740(.A(\in1[64] ), .B(\in0[64] ), .S0(new_n1960_), .Y(new_n2383_));
  INVX1    g1741(.A(new_n2383_), .Y(new_n2384_));
  MX2X1    g1742(.A(new_n1687_), .B(new_n1680_), .S0(new_n1960_), .Y(new_n2385_));
  INVX1    g1743(.A(new_n2385_), .Y(new_n2386_));
  MX2X1    g1744(.A(new_n1007_), .B(new_n1001_), .S0(new_n1969_), .Y(new_n2387_));
  NOR2X1   g1745(.A(new_n2387_), .B(new_n2386_), .Y(new_n2388_));
  AOI21X1  g1746(.A0(new_n2384_), .A1(new_n2382_), .B0(new_n2388_), .Y(new_n2389_));
  AND2X1   g1747(.A(new_n2389_), .B(new_n2381_), .Y(new_n2390_));
  INVX1    g1748(.A(new_n2390_), .Y(new_n2391_));
  AOI21X1  g1749(.A0(new_n2374_), .A1(new_n2356_), .B0(new_n2391_), .Y(new_n2392_));
  NOR2X1   g1750(.A(new_n2377_), .B(new_n2376_), .Y(new_n2393_));
  OR2X1    g1751(.A(new_n2384_), .B(new_n2382_), .Y(new_n2394_));
  INVX1    g1752(.A(new_n2380_), .Y(new_n2395_));
  AOI22X1  g1753(.A0(new_n2387_), .A1(new_n2386_), .B0(new_n2395_), .B1(new_n2378_), .Y(new_n2396_));
  OAI21X1  g1754(.A0(new_n2394_), .A1(new_n2388_), .B0(new_n2396_), .Y(new_n2397_));
  AOI21X1  g1755(.A0(new_n2397_), .A1(new_n2381_), .B0(new_n2393_), .Y(new_n2398_));
  INVX1    g1756(.A(new_n2398_), .Y(new_n2399_));
  MX2X1    g1757(.A(\in1[71] ), .B(\in0[71] ), .S0(new_n1960_), .Y(new_n2400_));
  MX2X1    g1758(.A(new_n1028_), .B(new_n1016_), .S0(new_n1969_), .Y(new_n2401_));
  NOR2X1   g1759(.A(new_n2401_), .B(new_n2400_), .Y(new_n2402_));
  MX2X1    g1760(.A(\in3[70] ), .B(\in2[70] ), .S0(new_n1969_), .Y(new_n2403_));
  MX2X1    g1761(.A(\in1[70] ), .B(\in0[70] ), .S0(new_n1960_), .Y(new_n2404_));
  INVX1    g1762(.A(new_n2404_), .Y(new_n2405_));
  AND2X1   g1763(.A(new_n2405_), .B(new_n2403_), .Y(new_n2406_));
  MX2X1    g1764(.A(\in1[69] ), .B(\in0[69] ), .S0(new_n1960_), .Y(new_n2407_));
  MX2X1    g1765(.A(new_n1025_), .B(new_n1019_), .S0(new_n1969_), .Y(new_n2408_));
  NOR2X1   g1766(.A(new_n2408_), .B(new_n2407_), .Y(new_n2409_));
  MX2X1    g1767(.A(\in1[68] ), .B(\in0[68] ), .S0(new_n1960_), .Y(new_n2410_));
  INVX1    g1768(.A(new_n2410_), .Y(new_n2411_));
  MX2X1    g1769(.A(\in3[68] ), .B(\in2[68] ), .S0(new_n1969_), .Y(new_n2412_));
  AND2X1   g1770(.A(new_n2412_), .B(new_n2411_), .Y(new_n2413_));
  NOR4X1   g1771(.A(new_n2413_), .B(new_n2409_), .C(new_n2406_), .D(new_n2402_), .Y(new_n2414_));
  OAI21X1  g1772(.A0(new_n2399_), .A1(new_n2392_), .B0(new_n2414_), .Y(new_n2415_));
  OR2X1    g1773(.A(new_n2412_), .B(new_n2411_), .Y(new_n2416_));
  NOR2X1   g1774(.A(new_n2416_), .B(new_n2409_), .Y(new_n2417_));
  AOI21X1  g1775(.A0(new_n2408_), .A1(new_n2407_), .B0(new_n2417_), .Y(new_n2418_));
  NOR3X1   g1776(.A(new_n2418_), .B(new_n2406_), .C(new_n2402_), .Y(new_n2419_));
  AND2X1   g1777(.A(new_n2401_), .B(new_n2400_), .Y(new_n2420_));
  OR2X1    g1778(.A(new_n2405_), .B(new_n2403_), .Y(new_n2421_));
  NOR2X1   g1779(.A(new_n2421_), .B(new_n2402_), .Y(new_n2422_));
  NOR3X1   g1780(.A(new_n2422_), .B(new_n2420_), .C(new_n2419_), .Y(new_n2423_));
  MX2X1    g1781(.A(\in1[75] ), .B(\in0[75] ), .S0(new_n1960_), .Y(new_n2424_));
  INVX1    g1782(.A(new_n2424_), .Y(new_n2425_));
  MX2X1    g1783(.A(\in3[75] ), .B(\in2[75] ), .S0(new_n1969_), .Y(new_n2426_));
  MX2X1    g1784(.A(new_n1045_), .B(new_n1034_), .S0(new_n1969_), .Y(new_n2427_));
  INVX1    g1785(.A(new_n2427_), .Y(new_n2428_));
  MX2X1    g1786(.A(new_n1724_), .B(new_n1712_), .S0(new_n1960_), .Y(new_n2429_));
  AOI22X1  g1787(.A0(new_n2429_), .A1(new_n2428_), .B0(new_n2426_), .B1(new_n2425_), .Y(new_n2430_));
  MX2X1    g1788(.A(new_n1723_), .B(new_n1716_), .S0(new_n1960_), .Y(new_n2431_));
  INVX1    g1789(.A(new_n2431_), .Y(new_n2432_));
  MX2X1    g1790(.A(new_n1044_), .B(new_n1038_), .S0(new_n1969_), .Y(new_n2433_));
  NOR2X1   g1791(.A(new_n2433_), .B(new_n2432_), .Y(new_n2434_));
  MX2X1    g1792(.A(\in3[72] ), .B(\in2[72] ), .S0(new_n1969_), .Y(new_n2435_));
  MX2X1    g1793(.A(\in1[72] ), .B(\in0[72] ), .S0(new_n1960_), .Y(new_n2436_));
  INVX1    g1794(.A(new_n2436_), .Y(new_n2437_));
  AOI21X1  g1795(.A0(new_n2437_), .A1(new_n2435_), .B0(new_n2434_), .Y(new_n2438_));
  AND2X1   g1796(.A(new_n2438_), .B(new_n2430_), .Y(new_n2439_));
  INVX1    g1797(.A(new_n2439_), .Y(new_n2440_));
  AOI21X1  g1798(.A0(new_n2423_), .A1(new_n2415_), .B0(new_n2440_), .Y(new_n2441_));
  NOR2X1   g1799(.A(new_n2426_), .B(new_n2425_), .Y(new_n2442_));
  OR2X1    g1800(.A(new_n2437_), .B(new_n2435_), .Y(new_n2443_));
  INVX1    g1801(.A(new_n2429_), .Y(new_n2444_));
  AOI22X1  g1802(.A0(new_n2433_), .A1(new_n2432_), .B0(new_n2444_), .B1(new_n2427_), .Y(new_n2445_));
  OAI21X1  g1803(.A0(new_n2443_), .A1(new_n2434_), .B0(new_n2445_), .Y(new_n2446_));
  AOI21X1  g1804(.A0(new_n2446_), .A1(new_n2430_), .B0(new_n2442_), .Y(new_n2447_));
  INVX1    g1805(.A(new_n2447_), .Y(new_n2448_));
  MX2X1    g1806(.A(\in1[79] ), .B(\in0[79] ), .S0(new_n1960_), .Y(new_n2449_));
  MX2X1    g1807(.A(new_n1065_), .B(new_n1053_), .S0(new_n1969_), .Y(new_n2450_));
  NOR2X1   g1808(.A(new_n2450_), .B(new_n2449_), .Y(new_n2451_));
  MX2X1    g1809(.A(\in3[78] ), .B(\in2[78] ), .S0(new_n1969_), .Y(new_n2452_));
  MX2X1    g1810(.A(\in1[78] ), .B(\in0[78] ), .S0(new_n1960_), .Y(new_n2453_));
  INVX1    g1811(.A(new_n2453_), .Y(new_n2454_));
  AND2X1   g1812(.A(new_n2454_), .B(new_n2452_), .Y(new_n2455_));
  MX2X1    g1813(.A(\in1[77] ), .B(\in0[77] ), .S0(new_n1960_), .Y(new_n2456_));
  MX2X1    g1814(.A(new_n1062_), .B(new_n1056_), .S0(new_n1969_), .Y(new_n2457_));
  NOR2X1   g1815(.A(new_n2457_), .B(new_n2456_), .Y(new_n2458_));
  MX2X1    g1816(.A(\in1[76] ), .B(\in0[76] ), .S0(new_n1960_), .Y(new_n2459_));
  INVX1    g1817(.A(new_n2459_), .Y(new_n2460_));
  MX2X1    g1818(.A(\in3[76] ), .B(\in2[76] ), .S0(new_n1969_), .Y(new_n2461_));
  AND2X1   g1819(.A(new_n2461_), .B(new_n2460_), .Y(new_n2462_));
  NOR4X1   g1820(.A(new_n2462_), .B(new_n2458_), .C(new_n2455_), .D(new_n2451_), .Y(new_n2463_));
  OAI21X1  g1821(.A0(new_n2448_), .A1(new_n2441_), .B0(new_n2463_), .Y(new_n2464_));
  OR2X1    g1822(.A(new_n2461_), .B(new_n2460_), .Y(new_n2465_));
  NOR2X1   g1823(.A(new_n2465_), .B(new_n2458_), .Y(new_n2466_));
  AOI21X1  g1824(.A0(new_n2457_), .A1(new_n2456_), .B0(new_n2466_), .Y(new_n2467_));
  NOR3X1   g1825(.A(new_n2467_), .B(new_n2455_), .C(new_n2451_), .Y(new_n2468_));
  AND2X1   g1826(.A(new_n2450_), .B(new_n2449_), .Y(new_n2469_));
  OR2X1    g1827(.A(new_n2454_), .B(new_n2452_), .Y(new_n2470_));
  NOR2X1   g1828(.A(new_n2470_), .B(new_n2451_), .Y(new_n2471_));
  NOR3X1   g1829(.A(new_n2471_), .B(new_n2469_), .C(new_n2468_), .Y(new_n2472_));
  MX2X1    g1830(.A(\in1[83] ), .B(\in0[83] ), .S0(new_n1960_), .Y(new_n2473_));
  INVX1    g1831(.A(new_n2473_), .Y(new_n2474_));
  MX2X1    g1832(.A(\in3[83] ), .B(\in2[83] ), .S0(new_n1969_), .Y(new_n2475_));
  MX2X1    g1833(.A(new_n1082_), .B(new_n1071_), .S0(new_n1969_), .Y(new_n2476_));
  INVX1    g1834(.A(new_n2476_), .Y(new_n2477_));
  MX2X1    g1835(.A(new_n1760_), .B(new_n1748_), .S0(new_n1960_), .Y(new_n2478_));
  AOI22X1  g1836(.A0(new_n2478_), .A1(new_n2477_), .B0(new_n2475_), .B1(new_n2474_), .Y(new_n2479_));
  MX2X1    g1837(.A(\in3[80] ), .B(\in2[80] ), .S0(new_n1969_), .Y(new_n2480_));
  MX2X1    g1838(.A(\in1[80] ), .B(\in0[80] ), .S0(new_n1960_), .Y(new_n2481_));
  INVX1    g1839(.A(new_n2481_), .Y(new_n2482_));
  MX2X1    g1840(.A(new_n1759_), .B(new_n1752_), .S0(new_n1960_), .Y(new_n2483_));
  INVX1    g1841(.A(new_n2483_), .Y(new_n2484_));
  MX2X1    g1842(.A(new_n1081_), .B(new_n1075_), .S0(new_n1969_), .Y(new_n2485_));
  NOR2X1   g1843(.A(new_n2485_), .B(new_n2484_), .Y(new_n2486_));
  AOI21X1  g1844(.A0(new_n2482_), .A1(new_n2480_), .B0(new_n2486_), .Y(new_n2487_));
  AND2X1   g1845(.A(new_n2487_), .B(new_n2479_), .Y(new_n2488_));
  INVX1    g1846(.A(new_n2488_), .Y(new_n2489_));
  AOI21X1  g1847(.A0(new_n2472_), .A1(new_n2464_), .B0(new_n2489_), .Y(new_n2490_));
  NOR2X1   g1848(.A(new_n2475_), .B(new_n2474_), .Y(new_n2491_));
  OR2X1    g1849(.A(new_n2482_), .B(new_n2480_), .Y(new_n2492_));
  INVX1    g1850(.A(new_n2478_), .Y(new_n2493_));
  AOI22X1  g1851(.A0(new_n2485_), .A1(new_n2484_), .B0(new_n2493_), .B1(new_n2476_), .Y(new_n2494_));
  OAI21X1  g1852(.A0(new_n2492_), .A1(new_n2486_), .B0(new_n2494_), .Y(new_n2495_));
  AOI21X1  g1853(.A0(new_n2495_), .A1(new_n2479_), .B0(new_n2491_), .Y(new_n2496_));
  INVX1    g1854(.A(new_n2496_), .Y(new_n2497_));
  MX2X1    g1855(.A(\in1[87] ), .B(\in0[87] ), .S0(new_n1960_), .Y(new_n2498_));
  MX2X1    g1856(.A(new_n1102_), .B(new_n1090_), .S0(new_n1969_), .Y(new_n2499_));
  NOR2X1   g1857(.A(new_n2499_), .B(new_n2498_), .Y(new_n2500_));
  MX2X1    g1858(.A(\in3[86] ), .B(\in2[86] ), .S0(new_n1969_), .Y(new_n2501_));
  MX2X1    g1859(.A(\in1[86] ), .B(\in0[86] ), .S0(new_n1960_), .Y(new_n2502_));
  INVX1    g1860(.A(new_n2502_), .Y(new_n2503_));
  AND2X1   g1861(.A(new_n2503_), .B(new_n2501_), .Y(new_n2504_));
  MX2X1    g1862(.A(\in1[85] ), .B(\in0[85] ), .S0(new_n1960_), .Y(new_n2505_));
  MX2X1    g1863(.A(new_n1099_), .B(new_n1093_), .S0(new_n1969_), .Y(new_n2506_));
  NOR2X1   g1864(.A(new_n2506_), .B(new_n2505_), .Y(new_n2507_));
  MX2X1    g1865(.A(\in1[84] ), .B(\in0[84] ), .S0(new_n1960_), .Y(new_n2508_));
  INVX1    g1866(.A(new_n2508_), .Y(new_n2509_));
  MX2X1    g1867(.A(\in3[84] ), .B(\in2[84] ), .S0(new_n1969_), .Y(new_n2510_));
  AND2X1   g1868(.A(new_n2510_), .B(new_n2509_), .Y(new_n2511_));
  NOR4X1   g1869(.A(new_n2511_), .B(new_n2507_), .C(new_n2504_), .D(new_n2500_), .Y(new_n2512_));
  OAI21X1  g1870(.A0(new_n2497_), .A1(new_n2490_), .B0(new_n2512_), .Y(new_n2513_));
  OR2X1    g1871(.A(new_n2510_), .B(new_n2509_), .Y(new_n2514_));
  NOR2X1   g1872(.A(new_n2514_), .B(new_n2507_), .Y(new_n2515_));
  AOI21X1  g1873(.A0(new_n2506_), .A1(new_n2505_), .B0(new_n2515_), .Y(new_n2516_));
  NOR3X1   g1874(.A(new_n2516_), .B(new_n2504_), .C(new_n2500_), .Y(new_n2517_));
  AND2X1   g1875(.A(new_n2499_), .B(new_n2498_), .Y(new_n2518_));
  OR2X1    g1876(.A(new_n2503_), .B(new_n2501_), .Y(new_n2519_));
  NOR2X1   g1877(.A(new_n2519_), .B(new_n2500_), .Y(new_n2520_));
  NOR3X1   g1878(.A(new_n2520_), .B(new_n2518_), .C(new_n2517_), .Y(new_n2521_));
  MX2X1    g1879(.A(\in1[91] ), .B(\in0[91] ), .S0(new_n1960_), .Y(new_n2522_));
  INVX1    g1880(.A(new_n2522_), .Y(new_n2523_));
  MX2X1    g1881(.A(\in3[91] ), .B(\in2[91] ), .S0(new_n1969_), .Y(new_n2524_));
  MX2X1    g1882(.A(new_n1119_), .B(new_n1108_), .S0(new_n1969_), .Y(new_n2525_));
  INVX1    g1883(.A(new_n2525_), .Y(new_n2526_));
  MX2X1    g1884(.A(new_n1796_), .B(new_n1784_), .S0(new_n1960_), .Y(new_n2527_));
  AOI22X1  g1885(.A0(new_n2527_), .A1(new_n2526_), .B0(new_n2524_), .B1(new_n2523_), .Y(new_n2528_));
  MX2X1    g1886(.A(new_n1795_), .B(new_n1788_), .S0(new_n1960_), .Y(new_n2529_));
  INVX1    g1887(.A(new_n2529_), .Y(new_n2530_));
  MX2X1    g1888(.A(new_n1118_), .B(new_n1112_), .S0(new_n1969_), .Y(new_n2531_));
  NOR2X1   g1889(.A(new_n2531_), .B(new_n2530_), .Y(new_n2532_));
  MX2X1    g1890(.A(\in3[88] ), .B(\in2[88] ), .S0(new_n1969_), .Y(new_n2533_));
  MX2X1    g1891(.A(\in1[88] ), .B(\in0[88] ), .S0(new_n1960_), .Y(new_n2534_));
  INVX1    g1892(.A(new_n2534_), .Y(new_n2535_));
  AOI21X1  g1893(.A0(new_n2535_), .A1(new_n2533_), .B0(new_n2532_), .Y(new_n2536_));
  AND2X1   g1894(.A(new_n2536_), .B(new_n2528_), .Y(new_n2537_));
  INVX1    g1895(.A(new_n2537_), .Y(new_n2538_));
  AOI21X1  g1896(.A0(new_n2521_), .A1(new_n2513_), .B0(new_n2538_), .Y(new_n2539_));
  NOR2X1   g1897(.A(new_n2524_), .B(new_n2523_), .Y(new_n2540_));
  OR2X1    g1898(.A(new_n2535_), .B(new_n2533_), .Y(new_n2541_));
  INVX1    g1899(.A(new_n2527_), .Y(new_n2542_));
  AOI22X1  g1900(.A0(new_n2531_), .A1(new_n2530_), .B0(new_n2542_), .B1(new_n2525_), .Y(new_n2543_));
  OAI21X1  g1901(.A0(new_n2541_), .A1(new_n2532_), .B0(new_n2543_), .Y(new_n2544_));
  AOI21X1  g1902(.A0(new_n2544_), .A1(new_n2528_), .B0(new_n2540_), .Y(new_n2545_));
  INVX1    g1903(.A(new_n2545_), .Y(new_n2546_));
  MX2X1    g1904(.A(\in1[95] ), .B(\in0[95] ), .S0(new_n1960_), .Y(new_n2547_));
  MX2X1    g1905(.A(new_n1139_), .B(new_n1127_), .S0(new_n1969_), .Y(new_n2548_));
  NOR2X1   g1906(.A(new_n2548_), .B(new_n2547_), .Y(new_n2549_));
  MX2X1    g1907(.A(\in3[94] ), .B(\in2[94] ), .S0(new_n1969_), .Y(new_n2550_));
  MX2X1    g1908(.A(\in1[94] ), .B(\in0[94] ), .S0(new_n1960_), .Y(new_n2551_));
  INVX1    g1909(.A(new_n2551_), .Y(new_n2552_));
  AND2X1   g1910(.A(new_n2552_), .B(new_n2550_), .Y(new_n2553_));
  MX2X1    g1911(.A(\in1[93] ), .B(\in0[93] ), .S0(new_n1960_), .Y(new_n2554_));
  MX2X1    g1912(.A(new_n1136_), .B(new_n1130_), .S0(new_n1969_), .Y(new_n2555_));
  NOR2X1   g1913(.A(new_n2555_), .B(new_n2554_), .Y(new_n2556_));
  MX2X1    g1914(.A(\in1[92] ), .B(\in0[92] ), .S0(new_n1960_), .Y(new_n2557_));
  INVX1    g1915(.A(new_n2557_), .Y(new_n2558_));
  MX2X1    g1916(.A(\in3[92] ), .B(\in2[92] ), .S0(new_n1969_), .Y(new_n2559_));
  AND2X1   g1917(.A(new_n2559_), .B(new_n2558_), .Y(new_n2560_));
  NOR4X1   g1918(.A(new_n2560_), .B(new_n2556_), .C(new_n2553_), .D(new_n2549_), .Y(new_n2561_));
  OAI21X1  g1919(.A0(new_n2546_), .A1(new_n2539_), .B0(new_n2561_), .Y(new_n2562_));
  OR2X1    g1920(.A(new_n2559_), .B(new_n2558_), .Y(new_n2563_));
  NOR2X1   g1921(.A(new_n2563_), .B(new_n2556_), .Y(new_n2564_));
  AOI21X1  g1922(.A0(new_n2555_), .A1(new_n2554_), .B0(new_n2564_), .Y(new_n2565_));
  NOR3X1   g1923(.A(new_n2565_), .B(new_n2553_), .C(new_n2549_), .Y(new_n2566_));
  AND2X1   g1924(.A(new_n2548_), .B(new_n2547_), .Y(new_n2567_));
  OR2X1    g1925(.A(new_n2552_), .B(new_n2550_), .Y(new_n2568_));
  NOR2X1   g1926(.A(new_n2568_), .B(new_n2549_), .Y(new_n2569_));
  NOR3X1   g1927(.A(new_n2569_), .B(new_n2567_), .C(new_n2566_), .Y(new_n2570_));
  MX2X1    g1928(.A(\in1[99] ), .B(\in0[99] ), .S0(new_n1960_), .Y(new_n2571_));
  INVX1    g1929(.A(new_n2571_), .Y(new_n2572_));
  MX2X1    g1930(.A(\in3[99] ), .B(\in2[99] ), .S0(new_n1969_), .Y(new_n2573_));
  MX2X1    g1931(.A(new_n1156_), .B(new_n1145_), .S0(new_n1969_), .Y(new_n2574_));
  INVX1    g1932(.A(new_n2574_), .Y(new_n2575_));
  MX2X1    g1933(.A(new_n1832_), .B(new_n1820_), .S0(new_n1960_), .Y(new_n2576_));
  AOI22X1  g1934(.A0(new_n2576_), .A1(new_n2575_), .B0(new_n2573_), .B1(new_n2572_), .Y(new_n2577_));
  MX2X1    g1935(.A(\in3[96] ), .B(\in2[96] ), .S0(new_n1969_), .Y(new_n2578_));
  MX2X1    g1936(.A(\in1[96] ), .B(\in0[96] ), .S0(new_n1960_), .Y(new_n2579_));
  INVX1    g1937(.A(new_n2579_), .Y(new_n2580_));
  MX2X1    g1938(.A(new_n1831_), .B(new_n1824_), .S0(new_n1960_), .Y(new_n2581_));
  INVX1    g1939(.A(new_n2581_), .Y(new_n2582_));
  MX2X1    g1940(.A(new_n1155_), .B(new_n1149_), .S0(new_n1969_), .Y(new_n2583_));
  NOR2X1   g1941(.A(new_n2583_), .B(new_n2582_), .Y(new_n2584_));
  AOI21X1  g1942(.A0(new_n2580_), .A1(new_n2578_), .B0(new_n2584_), .Y(new_n2585_));
  AND2X1   g1943(.A(new_n2585_), .B(new_n2577_), .Y(new_n2586_));
  INVX1    g1944(.A(new_n2586_), .Y(new_n2587_));
  AOI21X1  g1945(.A0(new_n2570_), .A1(new_n2562_), .B0(new_n2587_), .Y(new_n2588_));
  NOR2X1   g1946(.A(new_n2573_), .B(new_n2572_), .Y(new_n2589_));
  OR2X1    g1947(.A(new_n2580_), .B(new_n2578_), .Y(new_n2590_));
  INVX1    g1948(.A(new_n2576_), .Y(new_n2591_));
  AOI22X1  g1949(.A0(new_n2583_), .A1(new_n2582_), .B0(new_n2591_), .B1(new_n2574_), .Y(new_n2592_));
  OAI21X1  g1950(.A0(new_n2590_), .A1(new_n2584_), .B0(new_n2592_), .Y(new_n2593_));
  AOI21X1  g1951(.A0(new_n2593_), .A1(new_n2577_), .B0(new_n2589_), .Y(new_n2594_));
  INVX1    g1952(.A(new_n2594_), .Y(new_n2595_));
  MX2X1    g1953(.A(\in1[103] ), .B(\in0[103] ), .S0(new_n1960_), .Y(new_n2596_));
  MX2X1    g1954(.A(new_n1176_), .B(new_n1164_), .S0(new_n1969_), .Y(new_n2597_));
  NOR2X1   g1955(.A(new_n2597_), .B(new_n2596_), .Y(new_n2598_));
  MX2X1    g1956(.A(\in3[102] ), .B(\in2[102] ), .S0(new_n1969_), .Y(new_n2599_));
  MX2X1    g1957(.A(\in1[102] ), .B(\in0[102] ), .S0(new_n1960_), .Y(new_n2600_));
  INVX1    g1958(.A(new_n2600_), .Y(new_n2601_));
  AND2X1   g1959(.A(new_n2601_), .B(new_n2599_), .Y(new_n2602_));
  MX2X1    g1960(.A(\in1[101] ), .B(\in0[101] ), .S0(new_n1960_), .Y(new_n2603_));
  MX2X1    g1961(.A(new_n1173_), .B(new_n1167_), .S0(new_n1969_), .Y(new_n2604_));
  NOR2X1   g1962(.A(new_n2604_), .B(new_n2603_), .Y(new_n2605_));
  MX2X1    g1963(.A(\in1[100] ), .B(\in0[100] ), .S0(new_n1960_), .Y(new_n2606_));
  INVX1    g1964(.A(new_n2606_), .Y(new_n2607_));
  MX2X1    g1965(.A(\in3[100] ), .B(\in2[100] ), .S0(new_n1969_), .Y(new_n2608_));
  AND2X1   g1966(.A(new_n2608_), .B(new_n2607_), .Y(new_n2609_));
  NOR4X1   g1967(.A(new_n2609_), .B(new_n2605_), .C(new_n2602_), .D(new_n2598_), .Y(new_n2610_));
  OAI21X1  g1968(.A0(new_n2595_), .A1(new_n2588_), .B0(new_n2610_), .Y(new_n2611_));
  OR2X1    g1969(.A(new_n2608_), .B(new_n2607_), .Y(new_n2612_));
  NOR2X1   g1970(.A(new_n2612_), .B(new_n2605_), .Y(new_n2613_));
  AOI21X1  g1971(.A0(new_n2604_), .A1(new_n2603_), .B0(new_n2613_), .Y(new_n2614_));
  NOR3X1   g1972(.A(new_n2614_), .B(new_n2602_), .C(new_n2598_), .Y(new_n2615_));
  AND2X1   g1973(.A(new_n2597_), .B(new_n2596_), .Y(new_n2616_));
  OR2X1    g1974(.A(new_n2601_), .B(new_n2599_), .Y(new_n2617_));
  NOR2X1   g1975(.A(new_n2617_), .B(new_n2598_), .Y(new_n2618_));
  NOR3X1   g1976(.A(new_n2618_), .B(new_n2616_), .C(new_n2615_), .Y(new_n2619_));
  MX2X1    g1977(.A(\in1[107] ), .B(\in0[107] ), .S0(new_n1960_), .Y(new_n2620_));
  INVX1    g1978(.A(new_n2620_), .Y(new_n2621_));
  MX2X1    g1979(.A(\in3[107] ), .B(\in2[107] ), .S0(new_n1969_), .Y(new_n2622_));
  MX2X1    g1980(.A(new_n1193_), .B(new_n1182_), .S0(new_n1969_), .Y(new_n2623_));
  INVX1    g1981(.A(new_n2623_), .Y(new_n2624_));
  MX2X1    g1982(.A(new_n1868_), .B(new_n1856_), .S0(new_n1960_), .Y(new_n2625_));
  AOI22X1  g1983(.A0(new_n2625_), .A1(new_n2624_), .B0(new_n2622_), .B1(new_n2621_), .Y(new_n2626_));
  MX2X1    g1984(.A(new_n1867_), .B(new_n1860_), .S0(new_n1960_), .Y(new_n2627_));
  INVX1    g1985(.A(new_n2627_), .Y(new_n2628_));
  MX2X1    g1986(.A(new_n1192_), .B(new_n1186_), .S0(new_n1969_), .Y(new_n2629_));
  NOR2X1   g1987(.A(new_n2629_), .B(new_n2628_), .Y(new_n2630_));
  MX2X1    g1988(.A(\in3[104] ), .B(\in2[104] ), .S0(new_n1969_), .Y(new_n2631_));
  MX2X1    g1989(.A(\in1[104] ), .B(\in0[104] ), .S0(new_n1960_), .Y(new_n2632_));
  INVX1    g1990(.A(new_n2632_), .Y(new_n2633_));
  AOI21X1  g1991(.A0(new_n2633_), .A1(new_n2631_), .B0(new_n2630_), .Y(new_n2634_));
  AND2X1   g1992(.A(new_n2634_), .B(new_n2626_), .Y(new_n2635_));
  INVX1    g1993(.A(new_n2635_), .Y(new_n2636_));
  AOI21X1  g1994(.A0(new_n2619_), .A1(new_n2611_), .B0(new_n2636_), .Y(new_n2637_));
  NOR2X1   g1995(.A(new_n2622_), .B(new_n2621_), .Y(new_n2638_));
  OR2X1    g1996(.A(new_n2633_), .B(new_n2631_), .Y(new_n2639_));
  INVX1    g1997(.A(new_n2625_), .Y(new_n2640_));
  AOI22X1  g1998(.A0(new_n2629_), .A1(new_n2628_), .B0(new_n2640_), .B1(new_n2623_), .Y(new_n2641_));
  OAI21X1  g1999(.A0(new_n2639_), .A1(new_n2630_), .B0(new_n2641_), .Y(new_n2642_));
  AOI21X1  g2000(.A0(new_n2642_), .A1(new_n2626_), .B0(new_n2638_), .Y(new_n2643_));
  INVX1    g2001(.A(new_n2643_), .Y(new_n2644_));
  MX2X1    g2002(.A(\in1[111] ), .B(\in0[111] ), .S0(new_n1960_), .Y(new_n2645_));
  MX2X1    g2003(.A(new_n1213_), .B(new_n1201_), .S0(new_n1969_), .Y(new_n2646_));
  NOR2X1   g2004(.A(new_n2646_), .B(new_n2645_), .Y(new_n2647_));
  MX2X1    g2005(.A(\in3[110] ), .B(\in2[110] ), .S0(new_n1969_), .Y(new_n2648_));
  MX2X1    g2006(.A(\in1[110] ), .B(\in0[110] ), .S0(new_n1960_), .Y(new_n2649_));
  INVX1    g2007(.A(new_n2649_), .Y(new_n2650_));
  AND2X1   g2008(.A(new_n2650_), .B(new_n2648_), .Y(new_n2651_));
  MX2X1    g2009(.A(\in1[109] ), .B(\in0[109] ), .S0(new_n1960_), .Y(new_n2652_));
  MX2X1    g2010(.A(new_n1210_), .B(new_n1204_), .S0(new_n1969_), .Y(new_n2653_));
  NOR2X1   g2011(.A(new_n2653_), .B(new_n2652_), .Y(new_n2654_));
  MX2X1    g2012(.A(\in1[108] ), .B(\in0[108] ), .S0(new_n1960_), .Y(new_n2655_));
  INVX1    g2013(.A(new_n2655_), .Y(new_n2656_));
  MX2X1    g2014(.A(\in3[108] ), .B(\in2[108] ), .S0(new_n1969_), .Y(new_n2657_));
  AND2X1   g2015(.A(new_n2657_), .B(new_n2656_), .Y(new_n2658_));
  NOR4X1   g2016(.A(new_n2658_), .B(new_n2654_), .C(new_n2651_), .D(new_n2647_), .Y(new_n2659_));
  OAI21X1  g2017(.A0(new_n2644_), .A1(new_n2637_), .B0(new_n2659_), .Y(new_n2660_));
  OR2X1    g2018(.A(new_n2657_), .B(new_n2656_), .Y(new_n2661_));
  NOR2X1   g2019(.A(new_n2661_), .B(new_n2654_), .Y(new_n2662_));
  AOI21X1  g2020(.A0(new_n2653_), .A1(new_n2652_), .B0(new_n2662_), .Y(new_n2663_));
  NOR3X1   g2021(.A(new_n2663_), .B(new_n2651_), .C(new_n2647_), .Y(new_n2664_));
  AND2X1   g2022(.A(new_n2646_), .B(new_n2645_), .Y(new_n2665_));
  OR2X1    g2023(.A(new_n2650_), .B(new_n2648_), .Y(new_n2666_));
  NOR2X1   g2024(.A(new_n2666_), .B(new_n2647_), .Y(new_n2667_));
  NOR3X1   g2025(.A(new_n2667_), .B(new_n2665_), .C(new_n2664_), .Y(new_n2668_));
  MX2X1    g2026(.A(\in1[115] ), .B(\in0[115] ), .S0(new_n1960_), .Y(new_n2669_));
  INVX1    g2027(.A(new_n2669_), .Y(new_n2670_));
  MX2X1    g2028(.A(\in3[115] ), .B(\in2[115] ), .S0(new_n1969_), .Y(new_n2671_));
  MX2X1    g2029(.A(new_n1230_), .B(new_n1219_), .S0(new_n1969_), .Y(new_n2672_));
  INVX1    g2030(.A(new_n2672_), .Y(new_n2673_));
  MX2X1    g2031(.A(new_n1904_), .B(new_n1892_), .S0(new_n1960_), .Y(new_n2674_));
  AOI22X1  g2032(.A0(new_n2674_), .A1(new_n2673_), .B0(new_n2671_), .B1(new_n2670_), .Y(new_n2675_));
  MX2X1    g2033(.A(\in3[112] ), .B(\in2[112] ), .S0(new_n1969_), .Y(new_n2676_));
  MX2X1    g2034(.A(\in1[112] ), .B(\in0[112] ), .S0(new_n1960_), .Y(new_n2677_));
  INVX1    g2035(.A(new_n2677_), .Y(new_n2678_));
  MX2X1    g2036(.A(new_n1903_), .B(new_n1896_), .S0(new_n1960_), .Y(new_n2679_));
  INVX1    g2037(.A(new_n2679_), .Y(new_n2680_));
  MX2X1    g2038(.A(new_n1229_), .B(new_n1223_), .S0(new_n1969_), .Y(new_n2681_));
  NOR2X1   g2039(.A(new_n2681_), .B(new_n2680_), .Y(new_n2682_));
  AOI21X1  g2040(.A0(new_n2678_), .A1(new_n2676_), .B0(new_n2682_), .Y(new_n2683_));
  AND2X1   g2041(.A(new_n2683_), .B(new_n2675_), .Y(new_n2684_));
  INVX1    g2042(.A(new_n2684_), .Y(new_n2685_));
  AOI21X1  g2043(.A0(new_n2668_), .A1(new_n2660_), .B0(new_n2685_), .Y(new_n2686_));
  NOR2X1   g2044(.A(new_n2671_), .B(new_n2670_), .Y(new_n2687_));
  OR2X1    g2045(.A(new_n2678_), .B(new_n2676_), .Y(new_n2688_));
  INVX1    g2046(.A(new_n2674_), .Y(new_n2689_));
  AOI22X1  g2047(.A0(new_n2681_), .A1(new_n2680_), .B0(new_n2689_), .B1(new_n2672_), .Y(new_n2690_));
  OAI21X1  g2048(.A0(new_n2688_), .A1(new_n2682_), .B0(new_n2690_), .Y(new_n2691_));
  AOI21X1  g2049(.A0(new_n2691_), .A1(new_n2675_), .B0(new_n2687_), .Y(new_n2692_));
  INVX1    g2050(.A(new_n2692_), .Y(new_n2693_));
  MX2X1    g2051(.A(\in1[119] ), .B(\in0[119] ), .S0(new_n1960_), .Y(new_n2694_));
  MX2X1    g2052(.A(new_n1250_), .B(new_n1238_), .S0(new_n1969_), .Y(new_n2695_));
  NOR2X1   g2053(.A(new_n2695_), .B(new_n2694_), .Y(new_n2696_));
  MX2X1    g2054(.A(\in3[118] ), .B(\in2[118] ), .S0(new_n1969_), .Y(new_n2697_));
  MX2X1    g2055(.A(\in1[118] ), .B(\in0[118] ), .S0(new_n1960_), .Y(new_n2698_));
  INVX1    g2056(.A(new_n2698_), .Y(new_n2699_));
  AND2X1   g2057(.A(new_n2699_), .B(new_n2697_), .Y(new_n2700_));
  MX2X1    g2058(.A(\in1[117] ), .B(\in0[117] ), .S0(new_n1960_), .Y(new_n2701_));
  MX2X1    g2059(.A(new_n1247_), .B(new_n1241_), .S0(new_n1969_), .Y(new_n2702_));
  NOR2X1   g2060(.A(new_n2702_), .B(new_n2701_), .Y(new_n2703_));
  MX2X1    g2061(.A(\in1[116] ), .B(\in0[116] ), .S0(new_n1960_), .Y(new_n2704_));
  INVX1    g2062(.A(new_n2704_), .Y(new_n2705_));
  MX2X1    g2063(.A(\in3[116] ), .B(\in2[116] ), .S0(new_n1969_), .Y(new_n2706_));
  AND2X1   g2064(.A(new_n2706_), .B(new_n2705_), .Y(new_n2707_));
  NOR4X1   g2065(.A(new_n2707_), .B(new_n2703_), .C(new_n2700_), .D(new_n2696_), .Y(new_n2708_));
  OAI21X1  g2066(.A0(new_n2693_), .A1(new_n2686_), .B0(new_n2708_), .Y(new_n2709_));
  OR2X1    g2067(.A(new_n2706_), .B(new_n2705_), .Y(new_n2710_));
  NOR2X1   g2068(.A(new_n2710_), .B(new_n2703_), .Y(new_n2711_));
  AOI21X1  g2069(.A0(new_n2702_), .A1(new_n2701_), .B0(new_n2711_), .Y(new_n2712_));
  NOR3X1   g2070(.A(new_n2712_), .B(new_n2700_), .C(new_n2696_), .Y(new_n2713_));
  AND2X1   g2071(.A(new_n2695_), .B(new_n2694_), .Y(new_n2714_));
  OR2X1    g2072(.A(new_n2699_), .B(new_n2697_), .Y(new_n2715_));
  NOR2X1   g2073(.A(new_n2715_), .B(new_n2696_), .Y(new_n2716_));
  NOR3X1   g2074(.A(new_n2716_), .B(new_n2714_), .C(new_n2713_), .Y(new_n2717_));
  MX2X1    g2075(.A(\in1[123] ), .B(\in0[123] ), .S0(new_n1960_), .Y(new_n2718_));
  INVX1    g2076(.A(new_n2718_), .Y(new_n2719_));
  MX2X1    g2077(.A(\in3[123] ), .B(\in2[123] ), .S0(new_n1969_), .Y(new_n2720_));
  MX2X1    g2078(.A(new_n1267_), .B(new_n1256_), .S0(new_n1969_), .Y(new_n2721_));
  INVX1    g2079(.A(new_n2721_), .Y(new_n2722_));
  MX2X1    g2080(.A(new_n1940_), .B(new_n1928_), .S0(new_n1960_), .Y(new_n2723_));
  AOI22X1  g2081(.A0(new_n2723_), .A1(new_n2722_), .B0(new_n2720_), .B1(new_n2719_), .Y(new_n2724_));
  MX2X1    g2082(.A(new_n1939_), .B(new_n1932_), .S0(new_n1960_), .Y(new_n2725_));
  INVX1    g2083(.A(new_n2725_), .Y(new_n2726_));
  MX2X1    g2084(.A(new_n1266_), .B(new_n1260_), .S0(new_n1969_), .Y(new_n2727_));
  NOR2X1   g2085(.A(new_n2727_), .B(new_n2726_), .Y(new_n2728_));
  MX2X1    g2086(.A(\in3[120] ), .B(\in2[120] ), .S0(new_n1969_), .Y(new_n2729_));
  MX2X1    g2087(.A(\in1[120] ), .B(\in0[120] ), .S0(new_n1960_), .Y(new_n2730_));
  INVX1    g2088(.A(new_n2730_), .Y(new_n2731_));
  AOI21X1  g2089(.A0(new_n2731_), .A1(new_n2729_), .B0(new_n2728_), .Y(new_n2732_));
  AND2X1   g2090(.A(new_n2732_), .B(new_n2724_), .Y(new_n2733_));
  INVX1    g2091(.A(new_n2733_), .Y(new_n2734_));
  AOI21X1  g2092(.A0(new_n2717_), .A1(new_n2709_), .B0(new_n2734_), .Y(new_n2735_));
  NOR2X1   g2093(.A(new_n2720_), .B(new_n2719_), .Y(new_n2736_));
  OR2X1    g2094(.A(new_n2731_), .B(new_n2729_), .Y(new_n2737_));
  INVX1    g2095(.A(new_n2723_), .Y(new_n2738_));
  AOI22X1  g2096(.A0(new_n2727_), .A1(new_n2726_), .B0(new_n2738_), .B1(new_n2721_), .Y(new_n2739_));
  OAI21X1  g2097(.A0(new_n2737_), .A1(new_n2728_), .B0(new_n2739_), .Y(new_n2740_));
  AOI21X1  g2098(.A0(new_n2740_), .A1(new_n2724_), .B0(new_n2736_), .Y(new_n2741_));
  INVX1    g2099(.A(new_n2741_), .Y(new_n2742_));
  MX2X1    g2100(.A(new_n1952_), .B(new_n1947_), .S0(new_n1960_), .Y(new_n2743_));
  INVX1    g2101(.A(new_n2743_), .Y(new_n2744_));
  MX2X1    g2102(.A(new_n1283_), .B(new_n1277_), .S0(new_n1969_), .Y(new_n2745_));
  NOR2X1   g2103(.A(new_n2745_), .B(new_n2744_), .Y(new_n2746_));
  MX2X1    g2104(.A(new_n1954_), .B(new_n1946_), .S0(new_n1960_), .Y(new_n2747_));
  INVX1    g2105(.A(new_n2747_), .Y(new_n2748_));
  MX2X1    g2106(.A(new_n1285_), .B(new_n1276_), .S0(new_n1969_), .Y(new_n2749_));
  NOR2X1   g2107(.A(new_n2749_), .B(new_n2748_), .Y(new_n2750_));
  MX2X1    g2108(.A(new_n1953_), .B(new_n1949_), .S0(new_n1960_), .Y(new_n2751_));
  INVX1    g2109(.A(new_n2751_), .Y(new_n2752_));
  MX2X1    g2110(.A(new_n1284_), .B(new_n1279_), .S0(new_n1969_), .Y(new_n2753_));
  OAI22X1  g2111(.A0(new_n2753_), .A1(new_n2752_), .B0(new_n1964_), .B1(new_n1962_), .Y(new_n2754_));
  NOR3X1   g2112(.A(new_n2754_), .B(new_n2750_), .C(new_n2746_), .Y(new_n2755_));
  OAI21X1  g2113(.A0(new_n2742_), .A1(new_n2735_), .B0(new_n2755_), .Y(new_n2756_));
  NOR2X1   g2114(.A(new_n1964_), .B(new_n1962_), .Y(new_n2757_));
  NOR2X1   g2115(.A(new_n2750_), .B(new_n2746_), .Y(new_n2758_));
  INVX1    g2116(.A(new_n2749_), .Y(new_n2759_));
  INVX1    g2117(.A(new_n2753_), .Y(new_n2760_));
  OAI22X1  g2118(.A0(new_n2760_), .A1(new_n2751_), .B0(new_n2759_), .B1(new_n2747_), .Y(new_n2761_));
  AOI22X1  g2119(.A0(new_n2761_), .A1(new_n2758_), .B0(new_n2745_), .B1(new_n2744_), .Y(new_n2762_));
  NOR2X1   g2120(.A(new_n2762_), .B(new_n2757_), .Y(new_n2763_));
  INVX1    g2121(.A(new_n2763_), .Y(new_n2764_));
  NAND3X1  g2122(.A(new_n2764_), .B(new_n2756_), .C(new_n1966_), .Y(new_n2765_));
  MX2X1    g2123(.A(new_n1355_), .B(new_n1961_), .S0(new_n2765_), .Y(\result[0] ));
  MX2X1    g2124(.A(new_n2063_), .B(new_n2050_), .S0(new_n2765_), .Y(\result[1] ));
  MX2X1    g2125(.A(new_n2053_), .B(new_n2054_), .S0(new_n2765_), .Y(\result[2] ));
  INVX1    g2126(.A(new_n2045_), .Y(new_n2769_));
  MX2X1    g2127(.A(new_n2769_), .B(new_n2044_), .S0(new_n2765_), .Y(\result[3] ));
  MX2X1    g2128(.A(new_n2042_), .B(new_n2061_), .S0(new_n2765_), .Y(\result[4] ));
  MX2X1    g2129(.A(new_n2038_), .B(new_n2040_), .S0(new_n2765_), .Y(\result[5] ));
  INVX1    g2130(.A(new_n2034_), .Y(new_n2773_));
  MX2X1    g2131(.A(new_n2773_), .B(new_n2036_), .S0(new_n2765_), .Y(\result[6] ));
  MX2X1    g2132(.A(new_n2033_), .B(new_n2080_), .S0(new_n2765_), .Y(\result[7] ));
  MX2X1    g2133(.A(new_n2030_), .B(new_n2083_), .S0(new_n2765_), .Y(\result[8] ));
  INVX1    g2134(.A(new_n2028_), .Y(new_n2777_));
  MX2X1    g2135(.A(new_n2777_), .B(new_n2088_), .S0(new_n2765_), .Y(\result[9] ));
  MX2X1    g2136(.A(new_n2027_), .B(new_n2092_), .S0(new_n2765_), .Y(\result[10] ));
  INVX1    g2137(.A(new_n2024_), .Y(new_n2780_));
  MX2X1    g2138(.A(new_n2780_), .B(new_n2023_), .S0(new_n2765_), .Y(\result[11] ));
  MX2X1    g2139(.A(new_n2021_), .B(new_n2098_), .S0(new_n2765_), .Y(\result[12] ));
  INVX1    g2140(.A(new_n2018_), .Y(new_n2783_));
  MX2X1    g2141(.A(new_n2783_), .B(new_n2017_), .S0(new_n2765_), .Y(\result[13] ));
  MX2X1    g2142(.A(new_n2015_), .B(new_n2104_), .S0(new_n2765_), .Y(\result[14] ));
  INVX1    g2143(.A(new_n2012_), .Y(new_n2786_));
  MX2X1    g2144(.A(new_n2786_), .B(new_n2011_), .S0(new_n2765_), .Y(\result[15] ));
  INVX1    g2145(.A(new_n2009_), .Y(new_n2788_));
  MX2X1    g2146(.A(new_n2788_), .B(new_n2109_), .S0(new_n2765_), .Y(\result[16] ));
  MX2X1    g2147(.A(new_n2008_), .B(new_n2114_), .S0(new_n2765_), .Y(\result[17] ));
  INVX1    g2148(.A(new_n2006_), .Y(new_n2791_));
  MX2X1    g2149(.A(new_n2791_), .B(new_n2005_), .S0(new_n2765_), .Y(\result[18] ));
  MX2X1    g2150(.A(new_n2003_), .B(new_n2122_), .S0(new_n2765_), .Y(\result[19] ));
  INVX1    g2151(.A(new_n2000_), .Y(new_n2794_));
  MX2X1    g2152(.A(new_n2794_), .B(new_n1999_), .S0(new_n2765_), .Y(\result[20] ));
  MX2X1    g2153(.A(new_n1997_), .B(new_n2128_), .S0(new_n2765_), .Y(\result[21] ));
  INVX1    g2154(.A(new_n1994_), .Y(new_n2797_));
  MX2X1    g2155(.A(new_n2797_), .B(new_n1993_), .S0(new_n2765_), .Y(\result[22] ));
  MX2X1    g2156(.A(new_n1991_), .B(new_n2134_), .S0(new_n2765_), .Y(\result[23] ));
  MX2X1    g2157(.A(new_n1988_), .B(new_n2136_), .S0(new_n2765_), .Y(\result[24] ));
  INVX1    g2158(.A(new_n1986_), .Y(new_n2801_));
  MX2X1    g2159(.A(new_n2801_), .B(new_n2141_), .S0(new_n2765_), .Y(\result[25] ));
  MX2X1    g2160(.A(new_n1985_), .B(new_n2145_), .S0(new_n2765_), .Y(\result[26] ));
  INVX1    g2161(.A(new_n1982_), .Y(new_n2804_));
  MX2X1    g2162(.A(new_n2804_), .B(new_n1981_), .S0(new_n2765_), .Y(\result[27] ));
  MX2X1    g2163(.A(new_n1979_), .B(new_n2151_), .S0(new_n2765_), .Y(\result[28] ));
  INVX1    g2164(.A(new_n1976_), .Y(new_n2807_));
  MX2X1    g2165(.A(new_n2807_), .B(new_n1975_), .S0(new_n2765_), .Y(\result[29] ));
  MX2X1    g2166(.A(new_n1973_), .B(new_n2157_), .S0(new_n2765_), .Y(\result[30] ));
  INVX1    g2167(.A(new_n1970_), .Y(new_n2810_));
  MX2X1    g2168(.A(new_n2810_), .B(new_n1968_), .S0(new_n2765_), .Y(\result[31] ));
  INVX1    g2169(.A(new_n2176_), .Y(new_n2812_));
  MX2X1    g2170(.A(new_n2812_), .B(new_n2178_), .S0(new_n2765_), .Y(\result[32] ));
  INVX1    g2171(.A(new_n2168_), .Y(new_n2814_));
  MX2X1    g2172(.A(new_n2814_), .B(new_n2166_), .S0(new_n2765_), .Y(\result[33] ));
  INVX1    g2173(.A(new_n2162_), .Y(new_n2816_));
  MX2X1    g2174(.A(new_n2816_), .B(new_n2163_), .S0(new_n2765_), .Y(\result[34] ));
  MX2X1    g2175(.A(new_n2170_), .B(new_n2169_), .S0(new_n2765_), .Y(\result[35] ));
  INVX1    g2176(.A(new_n2190_), .Y(new_n2819_));
  MX2X1    g2177(.A(new_n2819_), .B(new_n2189_), .S0(new_n2765_), .Y(\result[36] ));
  INVX1    g2178(.A(new_n2192_), .Y(new_n2821_));
  MX2X1    g2179(.A(new_n2821_), .B(new_n2191_), .S0(new_n2765_), .Y(\result[37] ));
  MX2X1    g2180(.A(new_n2183_), .B(new_n2184_), .S0(new_n2765_), .Y(\result[38] ));
  INVX1    g2181(.A(new_n2181_), .Y(new_n2824_));
  MX2X1    g2182(.A(new_n2824_), .B(new_n2180_), .S0(new_n2765_), .Y(\result[39] ));
  MX2X1    g2183(.A(new_n2251_), .B(new_n2242_), .S0(new_n2765_), .Y(\result[40] ));
  MX2X1    g2184(.A(new_n2254_), .B(new_n2237_), .S0(new_n2765_), .Y(\result[41] ));
  MX2X1    g2185(.A(new_n2253_), .B(new_n2232_), .S0(new_n2765_), .Y(\result[42] ));
  MX2X1    g2186(.A(new_n2229_), .B(new_n2228_), .S0(new_n2765_), .Y(\result[43] ));
  INVX1    g2187(.A(new_n2224_), .Y(new_n2830_));
  MX2X1    g2188(.A(new_n2830_), .B(new_n2223_), .S0(new_n2765_), .Y(\result[44] ));
  INVX1    g2189(.A(new_n2226_), .Y(new_n2832_));
  MX2X1    g2190(.A(new_n2832_), .B(new_n2225_), .S0(new_n2765_), .Y(\result[45] ));
  MX2X1    g2191(.A(new_n2218_), .B(new_n2219_), .S0(new_n2765_), .Y(\result[46] ));
  INVX1    g2192(.A(new_n2216_), .Y(new_n2835_));
  MX2X1    g2193(.A(new_n2835_), .B(new_n2215_), .S0(new_n2765_), .Y(\result[47] ));
  INVX1    g2194(.A(new_n2280_), .Y(new_n2837_));
  MX2X1    g2195(.A(new_n2837_), .B(new_n2282_), .S0(new_n2765_), .Y(\result[48] ));
  INVX1    g2196(.A(new_n2272_), .Y(new_n2839_));
  MX2X1    g2197(.A(new_n2839_), .B(new_n2270_), .S0(new_n2765_), .Y(\result[49] ));
  INVX1    g2198(.A(new_n2266_), .Y(new_n2841_));
  MX2X1    g2199(.A(new_n2841_), .B(new_n2267_), .S0(new_n2765_), .Y(\result[50] ));
  MX2X1    g2200(.A(new_n2274_), .B(new_n2273_), .S0(new_n2765_), .Y(\result[51] ));
  INVX1    g2201(.A(new_n2298_), .Y(new_n2844_));
  MX2X1    g2202(.A(new_n2844_), .B(new_n2301_), .S0(new_n2765_), .Y(\result[52] ));
  INVX1    g2203(.A(new_n2296_), .Y(new_n2846_));
  MX2X1    g2204(.A(new_n2846_), .B(new_n2294_), .S0(new_n2765_), .Y(\result[53] ));
  MX2X1    g2205(.A(new_n2288_), .B(new_n2317_), .S0(new_n2765_), .Y(\result[54] ));
  MX2X1    g2206(.A(new_n2286_), .B(new_n2284_), .S0(new_n2765_), .Y(\result[55] ));
  MX2X1    g2207(.A(new_n2360_), .B(new_n2351_), .S0(new_n2765_), .Y(\result[56] ));
  MX2X1    g2208(.A(new_n2363_), .B(new_n2346_), .S0(new_n2765_), .Y(\result[57] ));
  MX2X1    g2209(.A(new_n2362_), .B(new_n2341_), .S0(new_n2765_), .Y(\result[58] ));
  MX2X1    g2210(.A(new_n2338_), .B(new_n2337_), .S0(new_n2765_), .Y(\result[59] ));
  INVX1    g2211(.A(new_n2333_), .Y(new_n2854_));
  MX2X1    g2212(.A(new_n2854_), .B(new_n2332_), .S0(new_n2765_), .Y(\result[60] ));
  INVX1    g2213(.A(new_n2335_), .Y(new_n2856_));
  MX2X1    g2214(.A(new_n2856_), .B(new_n2334_), .S0(new_n2765_), .Y(\result[61] ));
  MX2X1    g2215(.A(new_n2327_), .B(new_n2328_), .S0(new_n2765_), .Y(\result[62] ));
  INVX1    g2216(.A(new_n2325_), .Y(new_n2859_));
  MX2X1    g2217(.A(new_n2859_), .B(new_n2324_), .S0(new_n2765_), .Y(\result[63] ));
  MX2X1    g2218(.A(new_n2382_), .B(new_n2383_), .S0(new_n2765_), .Y(\result[64] ));
  INVX1    g2219(.A(new_n2387_), .Y(new_n2862_));
  MX2X1    g2220(.A(new_n2862_), .B(new_n2386_), .S0(new_n2765_), .Y(\result[65] ));
  MX2X1    g2221(.A(new_n2379_), .B(new_n2395_), .S0(new_n2765_), .Y(\result[66] ));
  MX2X1    g2222(.A(new_n2377_), .B(new_n2375_), .S0(new_n2765_), .Y(\result[67] ));
  MX2X1    g2223(.A(new_n2412_), .B(new_n2410_), .S0(new_n2765_), .Y(\result[68] ));
  INVX1    g2224(.A(new_n2408_), .Y(new_n2867_));
  MX2X1    g2225(.A(new_n2867_), .B(new_n2407_), .S0(new_n2765_), .Y(\result[69] ));
  MX2X1    g2226(.A(new_n2403_), .B(new_n2404_), .S0(new_n2765_), .Y(\result[70] ));
  INVX1    g2227(.A(new_n2401_), .Y(new_n2870_));
  MX2X1    g2228(.A(new_n2870_), .B(new_n2400_), .S0(new_n2765_), .Y(\result[71] ));
  MX2X1    g2229(.A(new_n2435_), .B(new_n2436_), .S0(new_n2765_), .Y(\result[72] ));
  INVX1    g2230(.A(new_n2433_), .Y(new_n2873_));
  MX2X1    g2231(.A(new_n2873_), .B(new_n2432_), .S0(new_n2765_), .Y(\result[73] ));
  MX2X1    g2232(.A(new_n2428_), .B(new_n2444_), .S0(new_n2765_), .Y(\result[74] ));
  MX2X1    g2233(.A(new_n2426_), .B(new_n2424_), .S0(new_n2765_), .Y(\result[75] ));
  MX2X1    g2234(.A(new_n2461_), .B(new_n2459_), .S0(new_n2765_), .Y(\result[76] ));
  INVX1    g2235(.A(new_n2457_), .Y(new_n2878_));
  MX2X1    g2236(.A(new_n2878_), .B(new_n2456_), .S0(new_n2765_), .Y(\result[77] ));
  MX2X1    g2237(.A(new_n2452_), .B(new_n2453_), .S0(new_n2765_), .Y(\result[78] ));
  INVX1    g2238(.A(new_n2450_), .Y(new_n2881_));
  MX2X1    g2239(.A(new_n2881_), .B(new_n2449_), .S0(new_n2765_), .Y(\result[79] ));
  MX2X1    g2240(.A(new_n2480_), .B(new_n2481_), .S0(new_n2765_), .Y(\result[80] ));
  INVX1    g2241(.A(new_n2485_), .Y(new_n2884_));
  MX2X1    g2242(.A(new_n2884_), .B(new_n2484_), .S0(new_n2765_), .Y(\result[81] ));
  MX2X1    g2243(.A(new_n2477_), .B(new_n2493_), .S0(new_n2765_), .Y(\result[82] ));
  MX2X1    g2244(.A(new_n2475_), .B(new_n2473_), .S0(new_n2765_), .Y(\result[83] ));
  MX2X1    g2245(.A(new_n2510_), .B(new_n2508_), .S0(new_n2765_), .Y(\result[84] ));
  INVX1    g2246(.A(new_n2506_), .Y(new_n2889_));
  MX2X1    g2247(.A(new_n2889_), .B(new_n2505_), .S0(new_n2765_), .Y(\result[85] ));
  MX2X1    g2248(.A(new_n2501_), .B(new_n2502_), .S0(new_n2765_), .Y(\result[86] ));
  INVX1    g2249(.A(new_n2499_), .Y(new_n2892_));
  MX2X1    g2250(.A(new_n2892_), .B(new_n2498_), .S0(new_n2765_), .Y(\result[87] ));
  MX2X1    g2251(.A(new_n2533_), .B(new_n2534_), .S0(new_n2765_), .Y(\result[88] ));
  INVX1    g2252(.A(new_n2531_), .Y(new_n2895_));
  MX2X1    g2253(.A(new_n2895_), .B(new_n2530_), .S0(new_n2765_), .Y(\result[89] ));
  MX2X1    g2254(.A(new_n2526_), .B(new_n2542_), .S0(new_n2765_), .Y(\result[90] ));
  MX2X1    g2255(.A(new_n2524_), .B(new_n2522_), .S0(new_n2765_), .Y(\result[91] ));
  MX2X1    g2256(.A(new_n2559_), .B(new_n2557_), .S0(new_n2765_), .Y(\result[92] ));
  INVX1    g2257(.A(new_n2555_), .Y(new_n2900_));
  MX2X1    g2258(.A(new_n2900_), .B(new_n2554_), .S0(new_n2765_), .Y(\result[93] ));
  MX2X1    g2259(.A(new_n2550_), .B(new_n2551_), .S0(new_n2765_), .Y(\result[94] ));
  INVX1    g2260(.A(new_n2548_), .Y(new_n2903_));
  MX2X1    g2261(.A(new_n2903_), .B(new_n2547_), .S0(new_n2765_), .Y(\result[95] ));
  MX2X1    g2262(.A(new_n2578_), .B(new_n2579_), .S0(new_n2765_), .Y(\result[96] ));
  INVX1    g2263(.A(new_n2583_), .Y(new_n2906_));
  MX2X1    g2264(.A(new_n2906_), .B(new_n2582_), .S0(new_n2765_), .Y(\result[97] ));
  MX2X1    g2265(.A(new_n2575_), .B(new_n2591_), .S0(new_n2765_), .Y(\result[98] ));
  MX2X1    g2266(.A(new_n2573_), .B(new_n2571_), .S0(new_n2765_), .Y(\result[99] ));
  MX2X1    g2267(.A(new_n2608_), .B(new_n2606_), .S0(new_n2765_), .Y(\result[100] ));
  INVX1    g2268(.A(new_n2604_), .Y(new_n2911_));
  MX2X1    g2269(.A(new_n2911_), .B(new_n2603_), .S0(new_n2765_), .Y(\result[101] ));
  MX2X1    g2270(.A(new_n2599_), .B(new_n2600_), .S0(new_n2765_), .Y(\result[102] ));
  INVX1    g2271(.A(new_n2597_), .Y(new_n2914_));
  MX2X1    g2272(.A(new_n2914_), .B(new_n2596_), .S0(new_n2765_), .Y(\result[103] ));
  MX2X1    g2273(.A(new_n2631_), .B(new_n2632_), .S0(new_n2765_), .Y(\result[104] ));
  INVX1    g2274(.A(new_n2629_), .Y(new_n2917_));
  MX2X1    g2275(.A(new_n2917_), .B(new_n2628_), .S0(new_n2765_), .Y(\result[105] ));
  MX2X1    g2276(.A(new_n2624_), .B(new_n2640_), .S0(new_n2765_), .Y(\result[106] ));
  MX2X1    g2277(.A(new_n2622_), .B(new_n2620_), .S0(new_n2765_), .Y(\result[107] ));
  MX2X1    g2278(.A(new_n2657_), .B(new_n2655_), .S0(new_n2765_), .Y(\result[108] ));
  INVX1    g2279(.A(new_n2653_), .Y(new_n2922_));
  MX2X1    g2280(.A(new_n2922_), .B(new_n2652_), .S0(new_n2765_), .Y(\result[109] ));
  MX2X1    g2281(.A(new_n2648_), .B(new_n2649_), .S0(new_n2765_), .Y(\result[110] ));
  INVX1    g2282(.A(new_n2646_), .Y(new_n2925_));
  MX2X1    g2283(.A(new_n2925_), .B(new_n2645_), .S0(new_n2765_), .Y(\result[111] ));
  MX2X1    g2284(.A(new_n2676_), .B(new_n2677_), .S0(new_n2765_), .Y(\result[112] ));
  INVX1    g2285(.A(new_n2681_), .Y(new_n2928_));
  MX2X1    g2286(.A(new_n2928_), .B(new_n2680_), .S0(new_n2765_), .Y(\result[113] ));
  MX2X1    g2287(.A(new_n2673_), .B(new_n2689_), .S0(new_n2765_), .Y(\result[114] ));
  MX2X1    g2288(.A(new_n2671_), .B(new_n2669_), .S0(new_n2765_), .Y(\result[115] ));
  MX2X1    g2289(.A(new_n2706_), .B(new_n2704_), .S0(new_n2765_), .Y(\result[116] ));
  INVX1    g2290(.A(new_n2702_), .Y(new_n2933_));
  MX2X1    g2291(.A(new_n2933_), .B(new_n2701_), .S0(new_n2765_), .Y(\result[117] ));
  MX2X1    g2292(.A(new_n2697_), .B(new_n2698_), .S0(new_n2765_), .Y(\result[118] ));
  INVX1    g2293(.A(new_n2695_), .Y(new_n2936_));
  MX2X1    g2294(.A(new_n2936_), .B(new_n2694_), .S0(new_n2765_), .Y(\result[119] ));
  MX2X1    g2295(.A(new_n2729_), .B(new_n2730_), .S0(new_n2765_), .Y(\result[120] ));
  INVX1    g2296(.A(new_n2727_), .Y(new_n2939_));
  MX2X1    g2297(.A(new_n2939_), .B(new_n2726_), .S0(new_n2765_), .Y(\result[121] ));
  MX2X1    g2298(.A(new_n2722_), .B(new_n2738_), .S0(new_n2765_), .Y(\result[122] ));
  MX2X1    g2299(.A(new_n2720_), .B(new_n2718_), .S0(new_n2765_), .Y(\result[123] ));
  MX2X1    g2300(.A(new_n2760_), .B(new_n2752_), .S0(new_n2765_), .Y(\result[124] ));
  MX2X1    g2301(.A(new_n2759_), .B(new_n2748_), .S0(new_n2765_), .Y(\result[125] ));
  INVX1    g2302(.A(new_n2745_), .Y(new_n2945_));
  MX2X1    g2303(.A(new_n2945_), .B(new_n2744_), .S0(new_n2765_), .Y(\result[126] ));
  INVX1    g2304(.A(new_n1962_), .Y(new_n2947_));
  AOI21X1  g2305(.A0(new_n2756_), .A1(new_n2947_), .B0(new_n1964_), .Y(\result[127] ));
  INVX1    g2306(.A(new_n1969_), .Y(new_n2949_));
  INVX1    g2307(.A(new_n1960_), .Y(new_n2950_));
  MX2X1    g2308(.A(new_n2949_), .B(new_n2950_), .S0(new_n2765_), .Y(\address[0] ));
  AND2X1   g2309(.A(new_n2764_), .B(new_n2756_), .Y(new_n2952_));
  AND2X1   g2310(.A(new_n2952_), .B(new_n1966_), .Y(\address[1] ));
endmodule


