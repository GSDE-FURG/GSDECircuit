// Benchmark "top" written by ABC on Mon Sep 21 04:01:57 2020

module top ( 
    \count[0] , \count[1] , \count[2] , \count[3] , \count[4] , \count[5] ,
    \count[6] , \count[7] ,
    \selectp1[0] , \selectp1[1] , \selectp1[2] , \selectp1[3] ,
    \selectp1[4] , \selectp1[5] , \selectp1[6] , \selectp1[7] ,
    \selectp1[8] , \selectp1[9] , \selectp1[10] , \selectp1[11] ,
    \selectp1[12] , \selectp1[13] , \selectp1[14] , \selectp1[15] ,
    \selectp1[16] , \selectp1[17] , \selectp1[18] , \selectp1[19] ,
    \selectp1[20] , \selectp1[21] , \selectp1[22] , \selectp1[23] ,
    \selectp1[24] , \selectp1[25] , \selectp1[26] , \selectp1[27] ,
    \selectp1[28] , \selectp1[29] , \selectp1[30] , \selectp1[31] ,
    \selectp1[32] , \selectp1[33] , \selectp1[34] , \selectp1[35] ,
    \selectp1[36] , \selectp1[37] , \selectp1[38] , \selectp1[39] ,
    \selectp1[40] , \selectp1[41] , \selectp1[42] , \selectp1[43] ,
    \selectp1[44] , \selectp1[45] , \selectp1[46] , \selectp1[47] ,
    \selectp1[48] , \selectp1[49] , \selectp1[50] , \selectp1[51] ,
    \selectp1[52] , \selectp1[53] , \selectp1[54] , \selectp1[55] ,
    \selectp1[56] , \selectp1[57] , \selectp1[58] , \selectp1[59] ,
    \selectp1[60] , \selectp1[61] , \selectp1[62] , \selectp1[63] ,
    \selectp1[64] , \selectp1[65] , \selectp1[66] , \selectp1[67] ,
    \selectp1[68] , \selectp1[69] , \selectp1[70] , \selectp1[71] ,
    \selectp1[72] , \selectp1[73] , \selectp1[74] , \selectp1[75] ,
    \selectp1[76] , \selectp1[77] , \selectp1[78] , \selectp1[79] ,
    \selectp1[80] , \selectp1[81] , \selectp1[82] , \selectp1[83] ,
    \selectp1[84] , \selectp1[85] , \selectp1[86] , \selectp1[87] ,
    \selectp1[88] , \selectp1[89] , \selectp1[90] , \selectp1[91] ,
    \selectp1[92] , \selectp1[93] , \selectp1[94] , \selectp1[95] ,
    \selectp1[96] , \selectp1[97] , \selectp1[98] , \selectp1[99] ,
    \selectp1[100] , \selectp1[101] , \selectp1[102] , \selectp1[103] ,
    \selectp1[104] , \selectp1[105] , \selectp1[106] , \selectp1[107] ,
    \selectp1[108] , \selectp1[109] , \selectp1[110] , \selectp1[111] ,
    \selectp1[112] , \selectp1[113] , \selectp1[114] , \selectp1[115] ,
    \selectp1[116] , \selectp1[117] , \selectp1[118] , \selectp1[119] ,
    \selectp1[120] , \selectp1[121] , \selectp1[122] , \selectp1[123] ,
    \selectp1[124] , \selectp1[125] , \selectp1[126] , \selectp1[127] ,
    \selectp2[0] , \selectp2[1] , \selectp2[2] , \selectp2[3] ,
    \selectp2[4] , \selectp2[5] , \selectp2[6] , \selectp2[7] ,
    \selectp2[8] , \selectp2[9] , \selectp2[10] , \selectp2[11] ,
    \selectp2[12] , \selectp2[13] , \selectp2[14] , \selectp2[15] ,
    \selectp2[16] , \selectp2[17] , \selectp2[18] , \selectp2[19] ,
    \selectp2[20] , \selectp2[21] , \selectp2[22] , \selectp2[23] ,
    \selectp2[24] , \selectp2[25] , \selectp2[26] , \selectp2[27] ,
    \selectp2[28] , \selectp2[29] , \selectp2[30] , \selectp2[31] ,
    \selectp2[32] , \selectp2[33] , \selectp2[34] , \selectp2[35] ,
    \selectp2[36] , \selectp2[37] , \selectp2[38] , \selectp2[39] ,
    \selectp2[40] , \selectp2[41] , \selectp2[42] , \selectp2[43] ,
    \selectp2[44] , \selectp2[45] , \selectp2[46] , \selectp2[47] ,
    \selectp2[48] , \selectp2[49] , \selectp2[50] , \selectp2[51] ,
    \selectp2[52] , \selectp2[53] , \selectp2[54] , \selectp2[55] ,
    \selectp2[56] , \selectp2[57] , \selectp2[58] , \selectp2[59] ,
    \selectp2[60] , \selectp2[61] , \selectp2[62] , \selectp2[63] ,
    \selectp2[64] , \selectp2[65] , \selectp2[66] , \selectp2[67] ,
    \selectp2[68] , \selectp2[69] , \selectp2[70] , \selectp2[71] ,
    \selectp2[72] , \selectp2[73] , \selectp2[74] , \selectp2[75] ,
    \selectp2[76] , \selectp2[77] , \selectp2[78] , \selectp2[79] ,
    \selectp2[80] , \selectp2[81] , \selectp2[82] , \selectp2[83] ,
    \selectp2[84] , \selectp2[85] , \selectp2[86] , \selectp2[87] ,
    \selectp2[88] , \selectp2[89] , \selectp2[90] , \selectp2[91] ,
    \selectp2[92] , \selectp2[93] , \selectp2[94] , \selectp2[95] ,
    \selectp2[96] , \selectp2[97] , \selectp2[98] , \selectp2[99] ,
    \selectp2[100] , \selectp2[101] , \selectp2[102] , \selectp2[103] ,
    \selectp2[104] , \selectp2[105] , \selectp2[106] , \selectp2[107] ,
    \selectp2[108] , \selectp2[109] , \selectp2[110] , \selectp2[111] ,
    \selectp2[112] , \selectp2[113] , \selectp2[114] , \selectp2[115] ,
    \selectp2[116] , \selectp2[117] , \selectp2[118] , \selectp2[119] ,
    \selectp2[120] , \selectp2[121] , \selectp2[122] , \selectp2[123] ,
    \selectp2[124] , \selectp2[125] , \selectp2[126] , \selectp2[127]   );
  input  \count[0] , \count[1] , \count[2] , \count[3] , \count[4] ,
    \count[5] , \count[6] , \count[7] ;
  output \selectp1[0] , \selectp1[1] , \selectp1[2] , \selectp1[3] ,
    \selectp1[4] , \selectp1[5] , \selectp1[6] , \selectp1[7] ,
    \selectp1[8] , \selectp1[9] , \selectp1[10] , \selectp1[11] ,
    \selectp1[12] , \selectp1[13] , \selectp1[14] , \selectp1[15] ,
    \selectp1[16] , \selectp1[17] , \selectp1[18] , \selectp1[19] ,
    \selectp1[20] , \selectp1[21] , \selectp1[22] , \selectp1[23] ,
    \selectp1[24] , \selectp1[25] , \selectp1[26] , \selectp1[27] ,
    \selectp1[28] , \selectp1[29] , \selectp1[30] , \selectp1[31] ,
    \selectp1[32] , \selectp1[33] , \selectp1[34] , \selectp1[35] ,
    \selectp1[36] , \selectp1[37] , \selectp1[38] , \selectp1[39] ,
    \selectp1[40] , \selectp1[41] , \selectp1[42] , \selectp1[43] ,
    \selectp1[44] , \selectp1[45] , \selectp1[46] , \selectp1[47] ,
    \selectp1[48] , \selectp1[49] , \selectp1[50] , \selectp1[51] ,
    \selectp1[52] , \selectp1[53] , \selectp1[54] , \selectp1[55] ,
    \selectp1[56] , \selectp1[57] , \selectp1[58] , \selectp1[59] ,
    \selectp1[60] , \selectp1[61] , \selectp1[62] , \selectp1[63] ,
    \selectp1[64] , \selectp1[65] , \selectp1[66] , \selectp1[67] ,
    \selectp1[68] , \selectp1[69] , \selectp1[70] , \selectp1[71] ,
    \selectp1[72] , \selectp1[73] , \selectp1[74] , \selectp1[75] ,
    \selectp1[76] , \selectp1[77] , \selectp1[78] , \selectp1[79] ,
    \selectp1[80] , \selectp1[81] , \selectp1[82] , \selectp1[83] ,
    \selectp1[84] , \selectp1[85] , \selectp1[86] , \selectp1[87] ,
    \selectp1[88] , \selectp1[89] , \selectp1[90] , \selectp1[91] ,
    \selectp1[92] , \selectp1[93] , \selectp1[94] , \selectp1[95] ,
    \selectp1[96] , \selectp1[97] , \selectp1[98] , \selectp1[99] ,
    \selectp1[100] , \selectp1[101] , \selectp1[102] , \selectp1[103] ,
    \selectp1[104] , \selectp1[105] , \selectp1[106] , \selectp1[107] ,
    \selectp1[108] , \selectp1[109] , \selectp1[110] , \selectp1[111] ,
    \selectp1[112] , \selectp1[113] , \selectp1[114] , \selectp1[115] ,
    \selectp1[116] , \selectp1[117] , \selectp1[118] , \selectp1[119] ,
    \selectp1[120] , \selectp1[121] , \selectp1[122] , \selectp1[123] ,
    \selectp1[124] , \selectp1[125] , \selectp1[126] , \selectp1[127] ,
    \selectp2[0] , \selectp2[1] , \selectp2[2] , \selectp2[3] ,
    \selectp2[4] , \selectp2[5] , \selectp2[6] , \selectp2[7] ,
    \selectp2[8] , \selectp2[9] , \selectp2[10] , \selectp2[11] ,
    \selectp2[12] , \selectp2[13] , \selectp2[14] , \selectp2[15] ,
    \selectp2[16] , \selectp2[17] , \selectp2[18] , \selectp2[19] ,
    \selectp2[20] , \selectp2[21] , \selectp2[22] , \selectp2[23] ,
    \selectp2[24] , \selectp2[25] , \selectp2[26] , \selectp2[27] ,
    \selectp2[28] , \selectp2[29] , \selectp2[30] , \selectp2[31] ,
    \selectp2[32] , \selectp2[33] , \selectp2[34] , \selectp2[35] ,
    \selectp2[36] , \selectp2[37] , \selectp2[38] , \selectp2[39] ,
    \selectp2[40] , \selectp2[41] , \selectp2[42] , \selectp2[43] ,
    \selectp2[44] , \selectp2[45] , \selectp2[46] , \selectp2[47] ,
    \selectp2[48] , \selectp2[49] , \selectp2[50] , \selectp2[51] ,
    \selectp2[52] , \selectp2[53] , \selectp2[54] , \selectp2[55] ,
    \selectp2[56] , \selectp2[57] , \selectp2[58] , \selectp2[59] ,
    \selectp2[60] , \selectp2[61] , \selectp2[62] , \selectp2[63] ,
    \selectp2[64] , \selectp2[65] , \selectp2[66] , \selectp2[67] ,
    \selectp2[68] , \selectp2[69] , \selectp2[70] , \selectp2[71] ,
    \selectp2[72] , \selectp2[73] , \selectp2[74] , \selectp2[75] ,
    \selectp2[76] , \selectp2[77] , \selectp2[78] , \selectp2[79] ,
    \selectp2[80] , \selectp2[81] , \selectp2[82] , \selectp2[83] ,
    \selectp2[84] , \selectp2[85] , \selectp2[86] , \selectp2[87] ,
    \selectp2[88] , \selectp2[89] , \selectp2[90] , \selectp2[91] ,
    \selectp2[92] , \selectp2[93] , \selectp2[94] , \selectp2[95] ,
    \selectp2[96] , \selectp2[97] , \selectp2[98] , \selectp2[99] ,
    \selectp2[100] , \selectp2[101] , \selectp2[102] , \selectp2[103] ,
    \selectp2[104] , \selectp2[105] , \selectp2[106] , \selectp2[107] ,
    \selectp2[108] , \selectp2[109] , \selectp2[110] , \selectp2[111] ,
    \selectp2[112] , \selectp2[113] , \selectp2[114] , \selectp2[115] ,
    \selectp2[116] , \selectp2[117] , \selectp2[118] , \selectp2[119] ,
    \selectp2[120] , \selectp2[121] , \selectp2[122] , \selectp2[123] ,
    \selectp2[124] , \selectp2[125] , \selectp2[126] , \selectp2[127] ;
  wire new_n265_, new_n266_, new_n267_, new_n269_, new_n270_, new_n272_,
    new_n273_, new_n275_, new_n277_, new_n278_, new_n280_, new_n282_,
    new_n284_, new_n286_, new_n287_, new_n289_, new_n291_, new_n293_,
    new_n295_, new_n297_, new_n299_, new_n301_, new_n303_, new_n304_,
    new_n321_, new_n322_, new_n339_, new_n356_, new_n357_, new_n374_,
    new_n391_, new_n408_, new_n425_, new_n442_, new_n459_, new_n476_,
    new_n493_, new_n510_, new_n527_, new_n544_;
  INVX1    g000(.A(\count[7] ), .Y(new_n265_));
  NOR4X1   g001(.A(new_n265_), .B(\count[6] ), .C(\count[5] ), .D(\count[4] ), .Y(new_n266_));
  NOR4X1   g002(.A(\count[3] ), .B(\count[2] ), .C(\count[1] ), .D(\count[0] ), .Y(new_n267_));
  AND2X1   g003(.A(new_n267_), .B(new_n266_), .Y(\selectp1[0] ));
  INVX1    g004(.A(\count[0] ), .Y(new_n269_));
  NOR4X1   g005(.A(\count[3] ), .B(\count[2] ), .C(\count[1] ), .D(new_n269_), .Y(new_n270_));
  AND2X1   g006(.A(new_n270_), .B(new_n266_), .Y(\selectp1[1] ));
  INVX1    g007(.A(\count[1] ), .Y(new_n272_));
  NOR4X1   g008(.A(\count[3] ), .B(\count[2] ), .C(new_n272_), .D(\count[0] ), .Y(new_n273_));
  AND2X1   g009(.A(new_n273_), .B(new_n266_), .Y(\selectp1[2] ));
  NOR4X1   g010(.A(\count[3] ), .B(\count[2] ), .C(new_n272_), .D(new_n269_), .Y(new_n275_));
  AND2X1   g011(.A(new_n275_), .B(new_n266_), .Y(\selectp1[3] ));
  INVX1    g012(.A(\count[2] ), .Y(new_n277_));
  NOR4X1   g013(.A(\count[3] ), .B(new_n277_), .C(\count[1] ), .D(\count[0] ), .Y(new_n278_));
  AND2X1   g014(.A(new_n278_), .B(new_n266_), .Y(\selectp1[4] ));
  NOR4X1   g015(.A(\count[3] ), .B(new_n277_), .C(\count[1] ), .D(new_n269_), .Y(new_n280_));
  AND2X1   g016(.A(new_n280_), .B(new_n266_), .Y(\selectp1[5] ));
  NOR4X1   g017(.A(\count[3] ), .B(new_n277_), .C(new_n272_), .D(\count[0] ), .Y(new_n282_));
  AND2X1   g018(.A(new_n282_), .B(new_n266_), .Y(\selectp1[6] ));
  NOR4X1   g019(.A(\count[3] ), .B(new_n277_), .C(new_n272_), .D(new_n269_), .Y(new_n284_));
  AND2X1   g020(.A(new_n284_), .B(new_n266_), .Y(\selectp1[7] ));
  INVX1    g021(.A(\count[3] ), .Y(new_n286_));
  NOR4X1   g022(.A(new_n286_), .B(\count[2] ), .C(\count[1] ), .D(\count[0] ), .Y(new_n287_));
  AND2X1   g023(.A(new_n287_), .B(new_n266_), .Y(\selectp1[8] ));
  NOR4X1   g024(.A(new_n286_), .B(\count[2] ), .C(\count[1] ), .D(new_n269_), .Y(new_n289_));
  AND2X1   g025(.A(new_n289_), .B(new_n266_), .Y(\selectp1[9] ));
  NOR4X1   g026(.A(new_n286_), .B(\count[2] ), .C(new_n272_), .D(\count[0] ), .Y(new_n291_));
  AND2X1   g027(.A(new_n291_), .B(new_n266_), .Y(\selectp1[10] ));
  NOR4X1   g028(.A(new_n286_), .B(\count[2] ), .C(new_n272_), .D(new_n269_), .Y(new_n293_));
  AND2X1   g029(.A(new_n293_), .B(new_n266_), .Y(\selectp1[11] ));
  NOR4X1   g030(.A(new_n286_), .B(new_n277_), .C(\count[1] ), .D(\count[0] ), .Y(new_n295_));
  AND2X1   g031(.A(new_n295_), .B(new_n266_), .Y(\selectp1[12] ));
  NOR4X1   g032(.A(new_n286_), .B(new_n277_), .C(\count[1] ), .D(new_n269_), .Y(new_n297_));
  AND2X1   g033(.A(new_n297_), .B(new_n266_), .Y(\selectp1[13] ));
  NOR4X1   g034(.A(new_n286_), .B(new_n277_), .C(new_n272_), .D(\count[0] ), .Y(new_n299_));
  AND2X1   g035(.A(new_n299_), .B(new_n266_), .Y(\selectp1[14] ));
  NOR4X1   g036(.A(new_n286_), .B(new_n277_), .C(new_n272_), .D(new_n269_), .Y(new_n301_));
  AND2X1   g037(.A(new_n301_), .B(new_n266_), .Y(\selectp1[15] ));
  INVX1    g038(.A(\count[4] ), .Y(new_n303_));
  NOR4X1   g039(.A(new_n265_), .B(\count[6] ), .C(\count[5] ), .D(new_n303_), .Y(new_n304_));
  AND2X1   g040(.A(new_n304_), .B(new_n267_), .Y(\selectp1[16] ));
  AND2X1   g041(.A(new_n304_), .B(new_n270_), .Y(\selectp1[17] ));
  AND2X1   g042(.A(new_n304_), .B(new_n273_), .Y(\selectp1[18] ));
  AND2X1   g043(.A(new_n304_), .B(new_n275_), .Y(\selectp1[19] ));
  AND2X1   g044(.A(new_n304_), .B(new_n278_), .Y(\selectp1[20] ));
  AND2X1   g045(.A(new_n304_), .B(new_n280_), .Y(\selectp1[21] ));
  AND2X1   g046(.A(new_n304_), .B(new_n282_), .Y(\selectp1[22] ));
  AND2X1   g047(.A(new_n304_), .B(new_n284_), .Y(\selectp1[23] ));
  AND2X1   g048(.A(new_n304_), .B(new_n287_), .Y(\selectp1[24] ));
  AND2X1   g049(.A(new_n304_), .B(new_n289_), .Y(\selectp1[25] ));
  AND2X1   g050(.A(new_n304_), .B(new_n291_), .Y(\selectp1[26] ));
  AND2X1   g051(.A(new_n304_), .B(new_n293_), .Y(\selectp1[27] ));
  AND2X1   g052(.A(new_n304_), .B(new_n295_), .Y(\selectp1[28] ));
  AND2X1   g053(.A(new_n304_), .B(new_n297_), .Y(\selectp1[29] ));
  AND2X1   g054(.A(new_n304_), .B(new_n299_), .Y(\selectp1[30] ));
  AND2X1   g055(.A(new_n304_), .B(new_n301_), .Y(\selectp1[31] ));
  INVX1    g056(.A(\count[5] ), .Y(new_n321_));
  NOR4X1   g057(.A(new_n265_), .B(\count[6] ), .C(new_n321_), .D(\count[4] ), .Y(new_n322_));
  AND2X1   g058(.A(new_n322_), .B(new_n267_), .Y(\selectp1[32] ));
  AND2X1   g059(.A(new_n322_), .B(new_n270_), .Y(\selectp1[33] ));
  AND2X1   g060(.A(new_n322_), .B(new_n273_), .Y(\selectp1[34] ));
  AND2X1   g061(.A(new_n322_), .B(new_n275_), .Y(\selectp1[35] ));
  AND2X1   g062(.A(new_n322_), .B(new_n278_), .Y(\selectp1[36] ));
  AND2X1   g063(.A(new_n322_), .B(new_n280_), .Y(\selectp1[37] ));
  AND2X1   g064(.A(new_n322_), .B(new_n282_), .Y(\selectp1[38] ));
  AND2X1   g065(.A(new_n322_), .B(new_n284_), .Y(\selectp1[39] ));
  AND2X1   g066(.A(new_n322_), .B(new_n287_), .Y(\selectp1[40] ));
  AND2X1   g067(.A(new_n322_), .B(new_n289_), .Y(\selectp1[41] ));
  AND2X1   g068(.A(new_n322_), .B(new_n291_), .Y(\selectp1[42] ));
  AND2X1   g069(.A(new_n322_), .B(new_n293_), .Y(\selectp1[43] ));
  AND2X1   g070(.A(new_n322_), .B(new_n295_), .Y(\selectp1[44] ));
  AND2X1   g071(.A(new_n322_), .B(new_n297_), .Y(\selectp1[45] ));
  AND2X1   g072(.A(new_n322_), .B(new_n299_), .Y(\selectp1[46] ));
  AND2X1   g073(.A(new_n322_), .B(new_n301_), .Y(\selectp1[47] ));
  NOR4X1   g074(.A(new_n265_), .B(\count[6] ), .C(new_n321_), .D(new_n303_), .Y(new_n339_));
  AND2X1   g075(.A(new_n339_), .B(new_n267_), .Y(\selectp1[48] ));
  AND2X1   g076(.A(new_n339_), .B(new_n270_), .Y(\selectp1[49] ));
  AND2X1   g077(.A(new_n339_), .B(new_n273_), .Y(\selectp1[50] ));
  AND2X1   g078(.A(new_n339_), .B(new_n275_), .Y(\selectp1[51] ));
  AND2X1   g079(.A(new_n339_), .B(new_n278_), .Y(\selectp1[52] ));
  AND2X1   g080(.A(new_n339_), .B(new_n280_), .Y(\selectp1[53] ));
  AND2X1   g081(.A(new_n339_), .B(new_n282_), .Y(\selectp1[54] ));
  AND2X1   g082(.A(new_n339_), .B(new_n284_), .Y(\selectp1[55] ));
  AND2X1   g083(.A(new_n339_), .B(new_n287_), .Y(\selectp1[56] ));
  AND2X1   g084(.A(new_n339_), .B(new_n289_), .Y(\selectp1[57] ));
  AND2X1   g085(.A(new_n339_), .B(new_n291_), .Y(\selectp1[58] ));
  AND2X1   g086(.A(new_n339_), .B(new_n293_), .Y(\selectp1[59] ));
  AND2X1   g087(.A(new_n339_), .B(new_n295_), .Y(\selectp1[60] ));
  AND2X1   g088(.A(new_n339_), .B(new_n297_), .Y(\selectp1[61] ));
  AND2X1   g089(.A(new_n339_), .B(new_n299_), .Y(\selectp1[62] ));
  AND2X1   g090(.A(new_n339_), .B(new_n301_), .Y(\selectp1[63] ));
  INVX1    g091(.A(\count[6] ), .Y(new_n356_));
  NOR4X1   g092(.A(new_n265_), .B(new_n356_), .C(\count[5] ), .D(\count[4] ), .Y(new_n357_));
  AND2X1   g093(.A(new_n357_), .B(new_n267_), .Y(\selectp1[64] ));
  AND2X1   g094(.A(new_n357_), .B(new_n270_), .Y(\selectp1[65] ));
  AND2X1   g095(.A(new_n357_), .B(new_n273_), .Y(\selectp1[66] ));
  AND2X1   g096(.A(new_n357_), .B(new_n275_), .Y(\selectp1[67] ));
  AND2X1   g097(.A(new_n357_), .B(new_n278_), .Y(\selectp1[68] ));
  AND2X1   g098(.A(new_n357_), .B(new_n280_), .Y(\selectp1[69] ));
  AND2X1   g099(.A(new_n357_), .B(new_n282_), .Y(\selectp1[70] ));
  AND2X1   g100(.A(new_n357_), .B(new_n284_), .Y(\selectp1[71] ));
  AND2X1   g101(.A(new_n357_), .B(new_n287_), .Y(\selectp1[72] ));
  AND2X1   g102(.A(new_n357_), .B(new_n289_), .Y(\selectp1[73] ));
  AND2X1   g103(.A(new_n357_), .B(new_n291_), .Y(\selectp1[74] ));
  AND2X1   g104(.A(new_n357_), .B(new_n293_), .Y(\selectp1[75] ));
  AND2X1   g105(.A(new_n357_), .B(new_n295_), .Y(\selectp1[76] ));
  AND2X1   g106(.A(new_n357_), .B(new_n297_), .Y(\selectp1[77] ));
  AND2X1   g107(.A(new_n357_), .B(new_n299_), .Y(\selectp1[78] ));
  AND2X1   g108(.A(new_n357_), .B(new_n301_), .Y(\selectp1[79] ));
  NOR4X1   g109(.A(new_n265_), .B(new_n356_), .C(\count[5] ), .D(new_n303_), .Y(new_n374_));
  AND2X1   g110(.A(new_n374_), .B(new_n267_), .Y(\selectp1[80] ));
  AND2X1   g111(.A(new_n374_), .B(new_n270_), .Y(\selectp1[81] ));
  AND2X1   g112(.A(new_n374_), .B(new_n273_), .Y(\selectp1[82] ));
  AND2X1   g113(.A(new_n374_), .B(new_n275_), .Y(\selectp1[83] ));
  AND2X1   g114(.A(new_n374_), .B(new_n278_), .Y(\selectp1[84] ));
  AND2X1   g115(.A(new_n374_), .B(new_n280_), .Y(\selectp1[85] ));
  AND2X1   g116(.A(new_n374_), .B(new_n282_), .Y(\selectp1[86] ));
  AND2X1   g117(.A(new_n374_), .B(new_n284_), .Y(\selectp1[87] ));
  AND2X1   g118(.A(new_n374_), .B(new_n287_), .Y(\selectp1[88] ));
  AND2X1   g119(.A(new_n374_), .B(new_n289_), .Y(\selectp1[89] ));
  AND2X1   g120(.A(new_n374_), .B(new_n291_), .Y(\selectp1[90] ));
  AND2X1   g121(.A(new_n374_), .B(new_n293_), .Y(\selectp1[91] ));
  AND2X1   g122(.A(new_n374_), .B(new_n295_), .Y(\selectp1[92] ));
  AND2X1   g123(.A(new_n374_), .B(new_n297_), .Y(\selectp1[93] ));
  AND2X1   g124(.A(new_n374_), .B(new_n299_), .Y(\selectp1[94] ));
  AND2X1   g125(.A(new_n374_), .B(new_n301_), .Y(\selectp1[95] ));
  NOR4X1   g126(.A(new_n265_), .B(new_n356_), .C(new_n321_), .D(\count[4] ), .Y(new_n391_));
  AND2X1   g127(.A(new_n391_), .B(new_n267_), .Y(\selectp1[96] ));
  AND2X1   g128(.A(new_n391_), .B(new_n270_), .Y(\selectp1[97] ));
  AND2X1   g129(.A(new_n391_), .B(new_n273_), .Y(\selectp1[98] ));
  AND2X1   g130(.A(new_n391_), .B(new_n275_), .Y(\selectp1[99] ));
  AND2X1   g131(.A(new_n391_), .B(new_n278_), .Y(\selectp1[100] ));
  AND2X1   g132(.A(new_n391_), .B(new_n280_), .Y(\selectp1[101] ));
  AND2X1   g133(.A(new_n391_), .B(new_n282_), .Y(\selectp1[102] ));
  AND2X1   g134(.A(new_n391_), .B(new_n284_), .Y(\selectp1[103] ));
  AND2X1   g135(.A(new_n391_), .B(new_n287_), .Y(\selectp1[104] ));
  AND2X1   g136(.A(new_n391_), .B(new_n289_), .Y(\selectp1[105] ));
  AND2X1   g137(.A(new_n391_), .B(new_n291_), .Y(\selectp1[106] ));
  AND2X1   g138(.A(new_n391_), .B(new_n293_), .Y(\selectp1[107] ));
  AND2X1   g139(.A(new_n391_), .B(new_n295_), .Y(\selectp1[108] ));
  AND2X1   g140(.A(new_n391_), .B(new_n297_), .Y(\selectp1[109] ));
  AND2X1   g141(.A(new_n391_), .B(new_n299_), .Y(\selectp1[110] ));
  AND2X1   g142(.A(new_n391_), .B(new_n301_), .Y(\selectp1[111] ));
  NOR4X1   g143(.A(new_n265_), .B(new_n356_), .C(new_n321_), .D(new_n303_), .Y(new_n408_));
  AND2X1   g144(.A(new_n408_), .B(new_n267_), .Y(\selectp1[112] ));
  AND2X1   g145(.A(new_n408_), .B(new_n270_), .Y(\selectp1[113] ));
  AND2X1   g146(.A(new_n408_), .B(new_n273_), .Y(\selectp1[114] ));
  AND2X1   g147(.A(new_n408_), .B(new_n275_), .Y(\selectp1[115] ));
  AND2X1   g148(.A(new_n408_), .B(new_n278_), .Y(\selectp1[116] ));
  AND2X1   g149(.A(new_n408_), .B(new_n280_), .Y(\selectp1[117] ));
  AND2X1   g150(.A(new_n408_), .B(new_n282_), .Y(\selectp1[118] ));
  AND2X1   g151(.A(new_n408_), .B(new_n284_), .Y(\selectp1[119] ));
  AND2X1   g152(.A(new_n408_), .B(new_n287_), .Y(\selectp1[120] ));
  AND2X1   g153(.A(new_n408_), .B(new_n289_), .Y(\selectp1[121] ));
  AND2X1   g154(.A(new_n408_), .B(new_n291_), .Y(\selectp1[122] ));
  AND2X1   g155(.A(new_n408_), .B(new_n293_), .Y(\selectp1[123] ));
  AND2X1   g156(.A(new_n408_), .B(new_n295_), .Y(\selectp1[124] ));
  AND2X1   g157(.A(new_n408_), .B(new_n297_), .Y(\selectp1[125] ));
  AND2X1   g158(.A(new_n408_), .B(new_n299_), .Y(\selectp1[126] ));
  AND2X1   g159(.A(new_n408_), .B(new_n301_), .Y(\selectp1[127] ));
  NOR4X1   g160(.A(\count[7] ), .B(\count[6] ), .C(\count[5] ), .D(\count[4] ), .Y(new_n425_));
  AND2X1   g161(.A(new_n425_), .B(new_n267_), .Y(\selectp2[0] ));
  AND2X1   g162(.A(new_n425_), .B(new_n270_), .Y(\selectp2[1] ));
  AND2X1   g163(.A(new_n425_), .B(new_n273_), .Y(\selectp2[2] ));
  AND2X1   g164(.A(new_n425_), .B(new_n275_), .Y(\selectp2[3] ));
  AND2X1   g165(.A(new_n425_), .B(new_n278_), .Y(\selectp2[4] ));
  AND2X1   g166(.A(new_n425_), .B(new_n280_), .Y(\selectp2[5] ));
  AND2X1   g167(.A(new_n425_), .B(new_n282_), .Y(\selectp2[6] ));
  AND2X1   g168(.A(new_n425_), .B(new_n284_), .Y(\selectp2[7] ));
  AND2X1   g169(.A(new_n425_), .B(new_n287_), .Y(\selectp2[8] ));
  AND2X1   g170(.A(new_n425_), .B(new_n289_), .Y(\selectp2[9] ));
  AND2X1   g171(.A(new_n425_), .B(new_n291_), .Y(\selectp2[10] ));
  AND2X1   g172(.A(new_n425_), .B(new_n293_), .Y(\selectp2[11] ));
  AND2X1   g173(.A(new_n425_), .B(new_n295_), .Y(\selectp2[12] ));
  AND2X1   g174(.A(new_n425_), .B(new_n297_), .Y(\selectp2[13] ));
  AND2X1   g175(.A(new_n425_), .B(new_n299_), .Y(\selectp2[14] ));
  AND2X1   g176(.A(new_n425_), .B(new_n301_), .Y(\selectp2[15] ));
  NOR4X1   g177(.A(\count[7] ), .B(\count[6] ), .C(\count[5] ), .D(new_n303_), .Y(new_n442_));
  AND2X1   g178(.A(new_n442_), .B(new_n267_), .Y(\selectp2[16] ));
  AND2X1   g179(.A(new_n442_), .B(new_n270_), .Y(\selectp2[17] ));
  AND2X1   g180(.A(new_n442_), .B(new_n273_), .Y(\selectp2[18] ));
  AND2X1   g181(.A(new_n442_), .B(new_n275_), .Y(\selectp2[19] ));
  AND2X1   g182(.A(new_n442_), .B(new_n278_), .Y(\selectp2[20] ));
  AND2X1   g183(.A(new_n442_), .B(new_n280_), .Y(\selectp2[21] ));
  AND2X1   g184(.A(new_n442_), .B(new_n282_), .Y(\selectp2[22] ));
  AND2X1   g185(.A(new_n442_), .B(new_n284_), .Y(\selectp2[23] ));
  AND2X1   g186(.A(new_n442_), .B(new_n287_), .Y(\selectp2[24] ));
  AND2X1   g187(.A(new_n442_), .B(new_n289_), .Y(\selectp2[25] ));
  AND2X1   g188(.A(new_n442_), .B(new_n291_), .Y(\selectp2[26] ));
  AND2X1   g189(.A(new_n442_), .B(new_n293_), .Y(\selectp2[27] ));
  AND2X1   g190(.A(new_n442_), .B(new_n295_), .Y(\selectp2[28] ));
  AND2X1   g191(.A(new_n442_), .B(new_n297_), .Y(\selectp2[29] ));
  AND2X1   g192(.A(new_n442_), .B(new_n299_), .Y(\selectp2[30] ));
  AND2X1   g193(.A(new_n442_), .B(new_n301_), .Y(\selectp2[31] ));
  NOR4X1   g194(.A(\count[7] ), .B(\count[6] ), .C(new_n321_), .D(\count[4] ), .Y(new_n459_));
  AND2X1   g195(.A(new_n459_), .B(new_n267_), .Y(\selectp2[32] ));
  AND2X1   g196(.A(new_n459_), .B(new_n270_), .Y(\selectp2[33] ));
  AND2X1   g197(.A(new_n459_), .B(new_n273_), .Y(\selectp2[34] ));
  AND2X1   g198(.A(new_n459_), .B(new_n275_), .Y(\selectp2[35] ));
  AND2X1   g199(.A(new_n459_), .B(new_n278_), .Y(\selectp2[36] ));
  AND2X1   g200(.A(new_n459_), .B(new_n280_), .Y(\selectp2[37] ));
  AND2X1   g201(.A(new_n459_), .B(new_n282_), .Y(\selectp2[38] ));
  AND2X1   g202(.A(new_n459_), .B(new_n284_), .Y(\selectp2[39] ));
  AND2X1   g203(.A(new_n459_), .B(new_n287_), .Y(\selectp2[40] ));
  AND2X1   g204(.A(new_n459_), .B(new_n289_), .Y(\selectp2[41] ));
  AND2X1   g205(.A(new_n459_), .B(new_n291_), .Y(\selectp2[42] ));
  AND2X1   g206(.A(new_n459_), .B(new_n293_), .Y(\selectp2[43] ));
  AND2X1   g207(.A(new_n459_), .B(new_n295_), .Y(\selectp2[44] ));
  AND2X1   g208(.A(new_n459_), .B(new_n297_), .Y(\selectp2[45] ));
  AND2X1   g209(.A(new_n459_), .B(new_n299_), .Y(\selectp2[46] ));
  AND2X1   g210(.A(new_n459_), .B(new_n301_), .Y(\selectp2[47] ));
  NOR4X1   g211(.A(\count[7] ), .B(\count[6] ), .C(new_n321_), .D(new_n303_), .Y(new_n476_));
  AND2X1   g212(.A(new_n476_), .B(new_n267_), .Y(\selectp2[48] ));
  AND2X1   g213(.A(new_n476_), .B(new_n270_), .Y(\selectp2[49] ));
  AND2X1   g214(.A(new_n476_), .B(new_n273_), .Y(\selectp2[50] ));
  AND2X1   g215(.A(new_n476_), .B(new_n275_), .Y(\selectp2[51] ));
  AND2X1   g216(.A(new_n476_), .B(new_n278_), .Y(\selectp2[52] ));
  AND2X1   g217(.A(new_n476_), .B(new_n280_), .Y(\selectp2[53] ));
  AND2X1   g218(.A(new_n476_), .B(new_n282_), .Y(\selectp2[54] ));
  AND2X1   g219(.A(new_n476_), .B(new_n284_), .Y(\selectp2[55] ));
  AND2X1   g220(.A(new_n476_), .B(new_n287_), .Y(\selectp2[56] ));
  AND2X1   g221(.A(new_n476_), .B(new_n289_), .Y(\selectp2[57] ));
  AND2X1   g222(.A(new_n476_), .B(new_n291_), .Y(\selectp2[58] ));
  AND2X1   g223(.A(new_n476_), .B(new_n293_), .Y(\selectp2[59] ));
  AND2X1   g224(.A(new_n476_), .B(new_n295_), .Y(\selectp2[60] ));
  AND2X1   g225(.A(new_n476_), .B(new_n297_), .Y(\selectp2[61] ));
  AND2X1   g226(.A(new_n476_), .B(new_n299_), .Y(\selectp2[62] ));
  AND2X1   g227(.A(new_n476_), .B(new_n301_), .Y(\selectp2[63] ));
  NOR4X1   g228(.A(\count[7] ), .B(new_n356_), .C(\count[5] ), .D(\count[4] ), .Y(new_n493_));
  AND2X1   g229(.A(new_n493_), .B(new_n267_), .Y(\selectp2[64] ));
  AND2X1   g230(.A(new_n493_), .B(new_n270_), .Y(\selectp2[65] ));
  AND2X1   g231(.A(new_n493_), .B(new_n273_), .Y(\selectp2[66] ));
  AND2X1   g232(.A(new_n493_), .B(new_n275_), .Y(\selectp2[67] ));
  AND2X1   g233(.A(new_n493_), .B(new_n278_), .Y(\selectp2[68] ));
  AND2X1   g234(.A(new_n493_), .B(new_n280_), .Y(\selectp2[69] ));
  AND2X1   g235(.A(new_n493_), .B(new_n282_), .Y(\selectp2[70] ));
  AND2X1   g236(.A(new_n493_), .B(new_n284_), .Y(\selectp2[71] ));
  AND2X1   g237(.A(new_n493_), .B(new_n287_), .Y(\selectp2[72] ));
  AND2X1   g238(.A(new_n493_), .B(new_n289_), .Y(\selectp2[73] ));
  AND2X1   g239(.A(new_n493_), .B(new_n291_), .Y(\selectp2[74] ));
  AND2X1   g240(.A(new_n493_), .B(new_n293_), .Y(\selectp2[75] ));
  AND2X1   g241(.A(new_n493_), .B(new_n295_), .Y(\selectp2[76] ));
  AND2X1   g242(.A(new_n493_), .B(new_n297_), .Y(\selectp2[77] ));
  AND2X1   g243(.A(new_n493_), .B(new_n299_), .Y(\selectp2[78] ));
  AND2X1   g244(.A(new_n493_), .B(new_n301_), .Y(\selectp2[79] ));
  NOR4X1   g245(.A(\count[7] ), .B(new_n356_), .C(\count[5] ), .D(new_n303_), .Y(new_n510_));
  AND2X1   g246(.A(new_n510_), .B(new_n267_), .Y(\selectp2[80] ));
  AND2X1   g247(.A(new_n510_), .B(new_n270_), .Y(\selectp2[81] ));
  AND2X1   g248(.A(new_n510_), .B(new_n273_), .Y(\selectp2[82] ));
  AND2X1   g249(.A(new_n510_), .B(new_n275_), .Y(\selectp2[83] ));
  AND2X1   g250(.A(new_n510_), .B(new_n278_), .Y(\selectp2[84] ));
  AND2X1   g251(.A(new_n510_), .B(new_n280_), .Y(\selectp2[85] ));
  AND2X1   g252(.A(new_n510_), .B(new_n282_), .Y(\selectp2[86] ));
  AND2X1   g253(.A(new_n510_), .B(new_n284_), .Y(\selectp2[87] ));
  AND2X1   g254(.A(new_n510_), .B(new_n287_), .Y(\selectp2[88] ));
  AND2X1   g255(.A(new_n510_), .B(new_n289_), .Y(\selectp2[89] ));
  AND2X1   g256(.A(new_n510_), .B(new_n291_), .Y(\selectp2[90] ));
  AND2X1   g257(.A(new_n510_), .B(new_n293_), .Y(\selectp2[91] ));
  AND2X1   g258(.A(new_n510_), .B(new_n295_), .Y(\selectp2[92] ));
  AND2X1   g259(.A(new_n510_), .B(new_n297_), .Y(\selectp2[93] ));
  AND2X1   g260(.A(new_n510_), .B(new_n299_), .Y(\selectp2[94] ));
  AND2X1   g261(.A(new_n510_), .B(new_n301_), .Y(\selectp2[95] ));
  NOR4X1   g262(.A(\count[7] ), .B(new_n356_), .C(new_n321_), .D(\count[4] ), .Y(new_n527_));
  AND2X1   g263(.A(new_n527_), .B(new_n267_), .Y(\selectp2[96] ));
  AND2X1   g264(.A(new_n527_), .B(new_n270_), .Y(\selectp2[97] ));
  AND2X1   g265(.A(new_n527_), .B(new_n273_), .Y(\selectp2[98] ));
  AND2X1   g266(.A(new_n527_), .B(new_n275_), .Y(\selectp2[99] ));
  AND2X1   g267(.A(new_n527_), .B(new_n278_), .Y(\selectp2[100] ));
  AND2X1   g268(.A(new_n527_), .B(new_n280_), .Y(\selectp2[101] ));
  AND2X1   g269(.A(new_n527_), .B(new_n282_), .Y(\selectp2[102] ));
  AND2X1   g270(.A(new_n527_), .B(new_n284_), .Y(\selectp2[103] ));
  AND2X1   g271(.A(new_n527_), .B(new_n287_), .Y(\selectp2[104] ));
  AND2X1   g272(.A(new_n527_), .B(new_n289_), .Y(\selectp2[105] ));
  AND2X1   g273(.A(new_n527_), .B(new_n291_), .Y(\selectp2[106] ));
  AND2X1   g274(.A(new_n527_), .B(new_n293_), .Y(\selectp2[107] ));
  AND2X1   g275(.A(new_n527_), .B(new_n295_), .Y(\selectp2[108] ));
  AND2X1   g276(.A(new_n527_), .B(new_n297_), .Y(\selectp2[109] ));
  AND2X1   g277(.A(new_n527_), .B(new_n299_), .Y(\selectp2[110] ));
  AND2X1   g278(.A(new_n527_), .B(new_n301_), .Y(\selectp2[111] ));
  NOR4X1   g279(.A(\count[7] ), .B(new_n356_), .C(new_n321_), .D(new_n303_), .Y(new_n544_));
  AND2X1   g280(.A(new_n544_), .B(new_n267_), .Y(\selectp2[112] ));
  AND2X1   g281(.A(new_n544_), .B(new_n270_), .Y(\selectp2[113] ));
  AND2X1   g282(.A(new_n544_), .B(new_n273_), .Y(\selectp2[114] ));
  AND2X1   g283(.A(new_n544_), .B(new_n275_), .Y(\selectp2[115] ));
  AND2X1   g284(.A(new_n544_), .B(new_n278_), .Y(\selectp2[116] ));
  AND2X1   g285(.A(new_n544_), .B(new_n280_), .Y(\selectp2[117] ));
  AND2X1   g286(.A(new_n544_), .B(new_n282_), .Y(\selectp2[118] ));
  AND2X1   g287(.A(new_n544_), .B(new_n284_), .Y(\selectp2[119] ));
  AND2X1   g288(.A(new_n544_), .B(new_n287_), .Y(\selectp2[120] ));
  AND2X1   g289(.A(new_n544_), .B(new_n289_), .Y(\selectp2[121] ));
  AND2X1   g290(.A(new_n544_), .B(new_n291_), .Y(\selectp2[122] ));
  AND2X1   g291(.A(new_n544_), .B(new_n293_), .Y(\selectp2[123] ));
  AND2X1   g292(.A(new_n544_), .B(new_n295_), .Y(\selectp2[124] ));
  AND2X1   g293(.A(new_n544_), .B(new_n297_), .Y(\selectp2[125] ));
  AND2X1   g294(.A(new_n544_), .B(new_n299_), .Y(\selectp2[126] ));
  AND2X1   g295(.A(new_n544_), .B(new_n301_), .Y(\selectp2[127] ));
endmodule


