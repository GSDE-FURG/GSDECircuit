//Converted to Combinational (Partial output: n3119gat) , Module name: s5378_n3119gat , Timestamp: 2018-12-03T15:51:03.229508 
module s5378_n3119gat ( n3095gat, n3086gat, n3087gat, n160gat, n553gat, n957gat, n816gat, n1294gat, n1241gat, n1298gat, n1068gat, n861gat, n865gat, n1080gat, n1148gat, n3083gat, n3084gat, n3085gat, n3088gat, n3093gat, n3119gat );
input n3095gat, n3086gat, n3087gat, n160gat, n553gat, n957gat, n816gat, n1294gat, n1241gat, n1298gat, n1068gat, n861gat, n865gat, n1080gat, n1148gat, n3083gat, n3084gat, n3085gat, n3088gat, n3093gat;
output n3119gat;
wire n343, n722, n784_1, n812, n808, n810, n811, n721, n780, n783, n809_1, n798, n806, n789_1, n807, n797, n719_1, n720, n715, n748, n779_1, n714_1, n709_1, n781, n782, n707, n805, n801, n803, n804_1, n788, n785, n786, n787, n796, n792, n794_1, n795, n718, n650, n622, n703, n704_1, n706, n713, n708, n705, n799_1, n800, n802, n701, n741, n790, n791, n793;
OAI21X1  g193(.A0(n784_1), .A1(n722), .B0(n343), .Y(n3119gat));
NAND4X1  g192(.A(n811), .B(n810), .C(n808), .D(n812), .Y(n343));
INVX1    g101(.A(n721), .Y(n722));
AND2X1   g163(.A(n783), .B(n780), .Y(n784_1));
NAND3X1  g191(.A(n806), .B(n798), .C(n809_1), .Y(n812));
NAND3X1  g187(.A(n807), .B(n798), .C(n789_1), .Y(n808));
NAND3X1  g189(.A(n807), .B(n797), .C(n809_1), .Y(n810));
NAND3X1  g190(.A(n806), .B(n797), .C(n789_1), .Y(n811));
NOR2X1   g100(.A(n720), .B(n719_1), .Y(n721));
AOI22X1  g159(.A0(n714_1), .A1(n779_1), .B0(n748), .B1(n715), .Y(n780));
AOI22X1  g162(.A0(n707), .A1(n782), .B0(n781), .B1(n709_1), .Y(n783));
INVX1    g188(.A(n789_1), .Y(n809_1));
INVX1    g177(.A(n797), .Y(n798));
NOR4X1   g185(.A(n804_1), .B(n803), .C(n801), .D(n805), .Y(n806));
NOR4X1   g168(.A(n787), .B(n786), .C(n785), .D(n788), .Y(n789_1));
INVX1    g186(.A(n806), .Y(n807));
NOR4X1   g176(.A(n795), .B(n794_1), .C(n792), .D(n796), .Y(n797));
OAI21X1  g098(.A0(n622), .A1(n650), .B0(n718), .Y(n719_1));
OAI21X1  g099(.A0(n3087gat), .A1(n3086gat), .B0(n3095gat), .Y(n720));
NOR3X1   g094(.A(n706), .B(n704_1), .C(n703), .Y(n715));
INVX1    g127(.A(n160gat), .Y(n748));
INVX1    g158(.A(n553gat), .Y(n779_1));
NOR3X1   g093(.A(n706), .B(n704_1), .C(n713), .Y(n714_1));
NOR3X1   g088(.A(n708), .B(n704_1), .C(n703), .Y(n709_1));
INVX1    g160(.A(n957gat), .Y(n781));
INVX1    g161(.A(n816gat), .Y(n782));
NOR3X1   g086(.A(n706), .B(n705), .C(n703), .Y(n707));
NOR3X1   g184(.A(n1298gat), .B(n1241gat), .C(n1294gat), .Y(n805));
NOR3X1   g180(.A(n1298gat), .B(n800), .C(n799_1), .Y(n801));
NOR3X1   g182(.A(n802), .B(n800), .C(n1294gat), .Y(n803));
NOR3X1   g183(.A(n802), .B(n1241gat), .C(n799_1), .Y(n804_1));
NOR3X1   g167(.A(n861gat), .B(n957gat), .C(n1068gat), .Y(n788));
NOR3X1   g164(.A(n861gat), .B(n781), .C(n701), .Y(n785));
NOR3X1   g165(.A(n741), .B(n781), .C(n1068gat), .Y(n786));
NOR3X1   g166(.A(n741), .B(n957gat), .C(n701), .Y(n787));
NOR3X1   g175(.A(n1148gat), .B(n1080gat), .C(n865gat), .Y(n796));
NOR3X1   g171(.A(n1148gat), .B(n791), .C(n790), .Y(n792));
NOR3X1   g173(.A(n793), .B(n791), .C(n865gat), .Y(n794_1));
NOR3X1   g174(.A(n793), .B(n1080gat), .C(n790), .Y(n795));
OAI21X1  g097(.A0(n3084gat), .A1(n3083gat), .B0(n3095gat), .Y(n718));
INVX1    g029(.A(n3085gat), .Y(n650));
INVX1    g001(.A(n3095gat), .Y(n622));
AOI22X1  g082(.A0(n3093gat), .A1(n3087gat), .B0(n3088gat), .B1(n3095gat), .Y(n703));
AOI22X1  g083(.A0(n3093gat), .A1(n3086gat), .B0(n3087gat), .B1(n3095gat), .Y(n704_1));
AOI22X1  g085(.A0(n3093gat), .A1(n3085gat), .B0(n3086gat), .B1(n3095gat), .Y(n706));
INVX1    g092(.A(n703), .Y(n713));
INVX1    g087(.A(n706), .Y(n708));
INVX1    g084(.A(n704_1), .Y(n705));
INVX1    g178(.A(n1294gat), .Y(n799_1));
INVX1    g179(.A(n1241gat), .Y(n800));
INVX1    g181(.A(n1298gat), .Y(n802));
INVX1    g080(.A(n1068gat), .Y(n701));
INVX1    g120(.A(n861gat), .Y(n741));
INVX1    g169(.A(n865gat), .Y(n790));
INVX1    g170(.A(n1080gat), .Y(n791));
INVX1    g172(.A(n1148gat), .Y(n793));

endmodule
