//Converted to Combinational (Partial output: n1146) , Module name: s9234_n1146 , Timestamp: 2018-12-03T15:51:03.594285 
module s9234_n1146 ( g94, g102, g89, g98, g152, g107, g114, g123, g188, g157, g139, g128, g131, g135, g179, g161, g143, g170, n1146 );
input g94, g102, g89, g98, g152, g107, g114, g123, g188, g157, g139, g128, g131, g135, g179, g161, g143, g170;
output n1146;
wire n1160, n1156_1, n1790, n1159, n1140, n788, n1157, n1078, n1132, n1155, n1136_1, n1789, n1786, n1158, n1128, n784, n1129, n1131_1, n1151_1, n1154, n1135, n1788, n783, n780, n1127, n708, n1130, n1149, n1150, n1152, n1143, n1153, n1134, n1787, n1318, n781_1, n782, n1126_1, n1138, n1142, n1141_1, n1144, n1133, n1612;
OAI21X1  g1081(.A0(n1790), .A1(n1156_1), .B0(n1160), .Y(n1146));
OR4X1    g0451(.A(n1157), .B(n788), .C(n1140), .D(n1159), .Y(n1160));
OAI21X1  g0447(.A0(n1155), .A1(n1132), .B0(n1078), .Y(n1156_1));
MX2X1    g1080(.A(n1786), .B(n1789), .S0(n1136_1), .Y(n1790));
INVX1    g0450(.A(n1158), .Y(n1159));
NOR3X1   g0431(.A(g102), .B(n1128), .C(g94), .Y(n1140));
NOR4X1   g0080(.A(g98), .B(g94), .C(g89), .D(g102), .Y(n788));
OR2X1    g0448(.A(n1155), .B(n1132), .Y(n1157));
INVX1    g0369(.A(n788), .Y(n1078));
OAI21X1  g0423(.A0(n1131_1), .A1(n1129), .B0(n784), .Y(n1132));
NOR2X1   g0446(.A(n1154), .B(n1151_1), .Y(n1155));
NAND2X1  g0427(.A(n1135), .B(n1132), .Y(n1136_1));
XOR2X1   g1079(.A(n1788), .B(g152), .Y(n1789));
INVX1    g1076(.A(g152), .Y(n1786));
AOI21X1  g0449(.A0(n1128), .A1(g94), .B0(n1131_1), .Y(n1158));
INVX1    g0419(.A(g98), .Y(n1128));
INVX1    g0076(.A(n783), .Y(n784));
AOI21X1  g0420(.A0(n1128), .A1(n1127), .B0(n780), .Y(n1129));
NOR3X1   g0422(.A(g107), .B(n1130), .C(n708), .Y(n1131_1));
NOR2X1   g0442(.A(n1150), .B(n1149), .Y(n1151_1));
NOR3X1   g0445(.A(n1153), .B(n1143), .C(n1152), .Y(n1154));
OAI21X1  g0426(.A0(n1134), .A1(g107), .B0(n784), .Y(n1135));
MX2X1    g1078(.A(n1318), .B(n1787), .S0(n1135), .Y(n1788));
NAND3X1  g0075(.A(n782), .B(g114), .C(n781_1), .Y(n783));
INVX1    g0072(.A(g123), .Y(n780));
INVX1    g0418(.A(g94), .Y(n1127));
INVX1    g0000(.A(g89), .Y(n708));
INVX1    g0421(.A(g102), .Y(n1130));
NAND2X1  g0440(.A(n1138), .B(n1126_1), .Y(n1149));
OR4X1    g0441(.A(n1141_1), .B(n1140), .C(g188), .D(n1142), .Y(n1150));
INVX1    g0443(.A(g188), .Y(n1152));
NOR3X1   g0434(.A(n1142), .B(n1141_1), .C(n1140), .Y(n1143));
OR2X1    g0444(.A(n1144), .B(n1126_1), .Y(n1153));
NOR4X1   g0425(.A(g107), .B(n1130), .C(g94), .D(n1133), .Y(n1134));
XOR2X1   g1077(.A(n1143), .B(n1612), .Y(n1787));
INVX1    g0609(.A(g157), .Y(n1318));
INVX1    g0073(.A(g139), .Y(n781_1));
NOR3X1   g0074(.A(g135), .B(g131), .C(g128), .Y(n782));
INVX1    g0417(.A(g179), .Y(n1126_1));
NOR4X1   g0429(.A(g152), .B(g170), .C(g143), .D(g161), .Y(n1138));
NOR3X1   g0433(.A(g102), .B(g98), .C(n1127), .Y(n1142));
NOR2X1   g0432(.A(n1130), .B(g94), .Y(n1141_1));
NAND4X1  g0435(.A(g152), .B(g170), .C(g143), .D(g161), .Y(n1144));
OR2X1    g0424(.A(g98), .B(g89), .Y(n1133));
INVX1    g0902(.A(g143), .Y(n1612));

endmodule
