//Converted to Combinational , Module name: s344 , Timestamp: 2018-12-03T15:51:01.401054 
module s344 ( START, B0, B1, B2, B3, A0, A1, A2, A3, CT2, CT1, CT0, ACVQN3, ACVQN2, ACVQN1, ACVQN0, MRVQN3, MRVQN2, MRVQN1, MRVQN0, AX3, AX2, AX1, AX0, P4, P5, P6, P7, P0, P1, P2, P3, CNTVCON2, CNTVCO2, READY, n41, n46, n51, n56, n61, n66, n71, n76, n81, n86, n91, n96, n101, n106, n111 );
input START, B0, B1, B2, B3, A0, A1, A2, A3, CT2, CT1, CT0, ACVQN3, ACVQN2, ACVQN1, ACVQN0, MRVQN3, MRVQN2, MRVQN1, MRVQN0, AX3, AX2, AX1, AX0;
output P4, P5, P6, P7, P0, P1, P2, P3, CNTVCON2, CNTVCO2, READY, n41, n46, n51, n56, n61, n66, n71, n76, n81, n86, n91, n96, n101, n106, n111;
wire n73, n74, n75, n79, n81_1, n82, n83, n86_1, n87, n88, n89, n90, n91_1, n92, n93, n94, n95, n96_1, n97, n98, n99, n101_1, n102, n103, n105, n106_1, n107, n108, n109, n110, n111_1, n112, n113, n114, n115, n116, n118, n119, n120, n122, n123, n124, n125, n127, n128, n130, n131, n133, n134;
INVX1    g00(.A(ACVQN0), .Y(P4));
INVX1    g01(.A(ACVQN1), .Y(P5));
INVX1    g02(.A(ACVQN2), .Y(P6));
INVX1    g03(.A(ACVQN3), .Y(P7));
INVX1    g04(.A(MRVQN0), .Y(P0));
INVX1    g05(.A(MRVQN1), .Y(P1));
INVX1    g06(.A(MRVQN2), .Y(P2));
INVX1    g07(.A(MRVQN3), .Y(P3));
INVX1    g08(.A(CT2), .Y(n73));
INVX1    g09(.A(CT1), .Y(n74));
INVX1    g10(.A(CT0), .Y(n75));
NOR3X1   g11(.A(n75), .B(n74), .C(n73), .Y(CNTVCO2));
INVX1    g12(.A(CNTVCO2), .Y(CNTVCON2));
NOR3X1   g13(.A(n75), .B(CT1), .C(n73), .Y(READY));
AOI21X1  g14(.A0(CT0), .A1(CT1), .B0(CT2), .Y(n79));
NOR3X1   g15(.A(n79), .B(CNTVCO2), .C(START), .Y(n41));
OAI21X1  g16(.A0(CT1), .A1(n73), .B0(CT0), .Y(n81_1));
INVX1    g17(.A(START), .Y(n82));
OAI21X1  g18(.A0(n81_1), .A1(n74), .B0(n82), .Y(n83));
AOI21X1  g19(.A0(n81_1), .A1(n74), .B0(n83), .Y(n46));
AND2X1   g20(.A(n81_1), .B(n82), .Y(n51));
NOR3X1   g21(.A(CT0), .B(CT1), .C(CT2), .Y(n86_1));
NOR2X1   g22(.A(n86_1), .B(READY), .Y(n87));
NAND3X1  g23(.A(AX0), .B(P0), .C(P4), .Y(n88));
AOI21X1  g24(.A0(AX1), .A1(P0), .B0(P5), .Y(n89));
NAND3X1  g25(.A(AX1), .B(P0), .C(P5), .Y(n90));
OAI21X1  g26(.A0(n89), .A1(n88), .B0(n90), .Y(n91_1));
INVX1    g27(.A(AX2), .Y(n92));
OAI21X1  g28(.A0(n92), .A1(MRVQN0), .B0(ACVQN2), .Y(n93));
NOR3X1   g29(.A(n92), .B(MRVQN0), .C(ACVQN2), .Y(n94));
AOI21X1  g30(.A0(n93), .A1(n91_1), .B0(n94), .Y(n95));
AOI21X1  g31(.A0(AX3), .A1(P0), .B0(P7), .Y(n96_1));
NAND3X1  g32(.A(AX3), .B(P0), .C(P7), .Y(n97));
OAI21X1  g33(.A0(n96_1), .A1(n95), .B0(n97), .Y(n98));
MX2X1    g34(.A(P7), .B(n98), .S0(n87), .Y(n99));
NAND2X1  g35(.A(n99), .B(n82), .Y(n56));
AND2X1   g36(.A(n96_1), .B(n95), .Y(n101_1));
OAI22X1  g37(.A0(n98), .A1(n101_1), .B0(n97), .B1(n95), .Y(n102));
MX2X1    g38(.A(P6), .B(n102), .S0(n87), .Y(n103));
NAND2X1  g39(.A(n103), .B(n82), .Y(n61));
INVX1    g40(.A(AX0), .Y(n105));
NOR3X1   g41(.A(n105), .B(MRVQN0), .C(ACVQN0), .Y(n106_1));
INVX1    g42(.A(AX1), .Y(n107));
OAI21X1  g43(.A0(n107), .A1(MRVQN0), .B0(ACVQN1), .Y(n108));
NOR3X1   g44(.A(n107), .B(MRVQN0), .C(ACVQN1), .Y(n109));
AOI21X1  g45(.A0(n108), .A1(n106_1), .B0(n109), .Y(n110));
INVX1    g46(.A(n94), .Y(n111_1));
INVX1    g47(.A(n93), .Y(n112));
OAI21X1  g48(.A0(n112), .A1(n110), .B0(n111_1), .Y(n113));
NOR2X1   g49(.A(n93), .B(n91_1), .Y(n114));
OAI22X1  g50(.A0(n113), .A1(n114), .B0(n111_1), .B1(n110), .Y(n115));
MX2X1    g51(.A(P5), .B(n115), .S0(n87), .Y(n116));
NAND2X1  g52(.A(n116), .B(n82), .Y(n66));
NOR2X1   g53(.A(n108), .B(n106_1), .Y(n118));
OAI22X1  g54(.A0(n91_1), .A1(n118), .B0(n90), .B1(n88), .Y(n119));
MX2X1    g55(.A(P4), .B(n119), .S0(n87), .Y(n120));
NAND2X1  g56(.A(n120), .B(n82), .Y(n71));
INVX1    g57(.A(B3), .Y(n122));
MX2X1    g58(.A(n122), .B(MRVQN3), .S0(READY), .Y(n123));
NOR2X1   g59(.A(n105), .B(MRVQN0), .Y(n124));
XOR2X1   g60(.A(n124), .B(ACVQN0), .Y(n125));
MX2X1    g61(.A(n123), .B(n125), .S0(n87), .Y(n76));
INVX1    g62(.A(B2), .Y(n127));
MX2X1    g63(.A(n127), .B(MRVQN2), .S0(READY), .Y(n128));
MX2X1    g64(.A(n128), .B(MRVQN3), .S0(n87), .Y(n81));
INVX1    g65(.A(B1), .Y(n130));
MX2X1    g66(.A(n130), .B(MRVQN1), .S0(READY), .Y(n131));
MX2X1    g67(.A(n131), .B(MRVQN2), .S0(n87), .Y(n86));
INVX1    g68(.A(B0), .Y(n133));
MX2X1    g69(.A(n133), .B(MRVQN0), .S0(READY), .Y(n134));
MX2X1    g70(.A(n134), .B(MRVQN1), .S0(n87), .Y(n91));
MX2X1    g71(.A(AX3), .B(A3), .S0(n86_1), .Y(n96));
MX2X1    g72(.A(AX2), .B(A2), .S0(n86_1), .Y(n101));
MX2X1    g73(.A(AX1), .B(A1), .S0(n86_1), .Y(n106));
MX2X1    g74(.A(AX0), .B(A0), .S0(n86_1), .Y(n111));
endmodule
