//Converted to Combinational , Module name: s713 , Timestamp: 2018-12-03T15:51:01.939971 
module s713 ( G1, G2, G3, G4, G5, G6, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G64, G65, G66, G67, G68, G69, G70, G71, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G103BF, G104BF, G105BF, G106BF, G107, G83, G84, G85, G86BF, G87BF, G88BF, G89BF, G90, G91, G92, G94, G95BF, G96BF, G97BF, G98BF, G99BF, G100BF, G101BF, n117, n122, n127, n132, n137, n142, n147, n152, n157, n162, n167, n172, n177, n182, n187, n192, n197, n202, n207 );
input G1, G2, G3, G4, G5, G6, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G64, G65, G66, G67, G68, G69, G70, G71, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82;
output G103BF, G104BF, G105BF, G106BF, G107, G83, G84, G85, G86BF, G87BF, G88BF, G89BF, G90, G91, G92, G94, G95BF, G96BF, G97BF, G98BF, G99BF, G100BF, G101BF, n117, n122, n127, n132, n137, n142, n147, n152, n157, n162, n167, n172, n177, n182, n187, n192, n197, n202, n207;
wire n115, n116, n117_1, n118, n119, n120, n121, n122_1, n123, n124, n125, n126, n127_1, n128, n129, n130, n131, n132_1, n133, n134, n135, n136, n137_1, n138, n139, n140, n141, n142_1, n143, n147_1, n151, n153, n155, n157_1, n159, n164, n165, n166, n167_1, n168, n169, n170, n171, n172_1, n173, n174, n175, n176, n177_1, n178, n179, n180, n181, n182_1, n183, n184, n185, n187_1, n188, n190, n203, n208, n209, n210, n211, n213, n214, n215, n216, n218, n219, n220, n222, n223, n224;
INVX1    g000(.A(G3), .Y(n115));
INVX1    g001(.A(G75), .Y(n116));
INVX1    g002(.A(G77), .Y(n117_1));
INVX1    g003(.A(G78), .Y(n118));
INVX1    g004(.A(G13), .Y(n119));
NAND4X1  g005(.A(G10), .B(G9), .C(n115), .D(n119), .Y(n120));
INVX1    g006(.A(G25), .Y(n121));
NOR2X1   g007(.A(G11), .B(G3), .Y(n122_1));
NOR3X1   g008(.A(n122_1), .B(G67), .C(n121), .Y(n123));
AOI21X1  g009(.A0(n123), .A1(n120), .B0(G3), .Y(n124));
OR2X1    g010(.A(n124), .B(n118), .Y(n125));
INVX1    g011(.A(G2), .Y(n126));
AND2X1   g012(.A(G66), .B(n126), .Y(n127_1));
OAI21X1  g013(.A0(n124), .A1(n118), .B0(n127_1), .Y(n128));
INVX1    g014(.A(G9), .Y(n129));
NOR4X1   g015(.A(G10), .B(n129), .C(G3), .D(G13), .Y(n130));
OAI21X1  g016(.A0(G11), .A1(G3), .B0(G24), .Y(n131));
NOR2X1   g017(.A(n131), .B(n130), .Y(n132_1));
AOI21X1  g018(.A0(n132_1), .A1(n128), .B0(G3), .Y(n133));
OAI21X1  g019(.A0(n133), .A1(n117_1), .B0(n125), .Y(n134));
INVX1    g020(.A(G23), .Y(n135));
INVX1    g021(.A(G10), .Y(n136));
NOR4X1   g022(.A(n136), .B(G9), .C(G3), .D(G13), .Y(n137_1));
NOR4X1   g023(.A(n122_1), .B(G65), .C(n135), .D(n137_1), .Y(n138));
OAI21X1  g024(.A0(n138), .A1(G3), .B0(G76), .Y(n139));
NAND3X1  g025(.A(n139), .B(G64), .C(n126), .Y(n140));
NOR4X1   g026(.A(G10), .B(G9), .C(G3), .D(G13), .Y(n141));
OAI21X1  g027(.A0(G11), .A1(G3), .B0(G22), .Y(n142_1));
NOR2X1   g028(.A(n142_1), .B(n141), .Y(n143));
OAI21X1  g029(.A0(n140), .A1(n134), .B0(n143), .Y(G86BF));
AOI21X1  g030(.A0(G86BF), .A1(n115), .B0(n116), .Y(n117));
NAND2X1  g031(.A(n117), .B(G14), .Y(G103BF));
INVX1    g032(.A(n139), .Y(n147_1));
NAND2X1  g033(.A(n147_1), .B(G15), .Y(G104BF));
NOR2X1   g034(.A(n133), .B(n117_1), .Y(n127));
NAND2X1  g035(.A(n127), .B(G16), .Y(G105BF));
INVX1    g036(.A(n125), .Y(n151));
NAND2X1  g037(.A(n151), .B(G17), .Y(G106BF));
NAND2X1  g038(.A(G79), .B(G18), .Y(n153));
NOR2X1   g039(.A(n153), .B(G4), .Y(G107));
NAND2X1  g040(.A(G80), .B(G19), .Y(n155));
NOR2X1   g041(.A(n155), .B(G4), .Y(G83));
NAND2X1  g042(.A(G81), .B(G20), .Y(n157_1));
NOR2X1   g043(.A(n157_1), .B(G4), .Y(G84));
NAND2X1  g044(.A(G82), .B(G21), .Y(n159));
NOR2X1   g045(.A(n159), .B(G4), .Y(G85));
INVX1    g046(.A(n138), .Y(G87BF));
NAND2X1  g047(.A(n132_1), .B(n128), .Y(G88BF));
NAND2X1  g048(.A(n123), .B(n120), .Y(G89BF));
INVX1    g049(.A(G74), .Y(n164));
INVX1    g050(.A(G4), .Y(n165));
AND2X1   g051(.A(G73), .B(n165), .Y(n166));
NAND4X1  g052(.A(n119), .B(n136), .C(n129), .D(n166), .Y(n167_1));
NOR3X1   g053(.A(n167_1), .B(G86BF), .C(n164), .Y(n168));
NAND3X1  g054(.A(n132_1), .B(n128), .C(G70), .Y(n169));
INVX1    g055(.A(G72), .Y(n170));
NAND3X1  g056(.A(n123), .B(n120), .C(G68), .Y(n171));
NAND2X1  g057(.A(G71), .B(n165), .Y(n172_1));
NOR2X1   g058(.A(n172_1), .B(G11), .Y(n173));
NAND2X1  g059(.A(G69), .B(n165), .Y(n174));
INVX1    g060(.A(n174), .Y(n175));
NAND3X1  g061(.A(n175), .B(n173), .C(n166), .Y(n176));
OR4X1    g062(.A(n171), .B(G87BF), .C(n170), .D(n176), .Y(n177_1));
NOR4X1   g063(.A(n169), .B(G86BF), .C(n164), .D(n177_1), .Y(n178));
OR4X1    g064(.A(G13), .B(G10), .C(n129), .D(n174), .Y(n179));
AND2X1   g065(.A(n138), .B(G72), .Y(n180));
NOR4X1   g066(.A(G13), .B(n136), .C(G9), .D(n172_1), .Y(n181));
OR4X1    g067(.A(G13), .B(n136), .C(n129), .D(n171), .Y(n182_1));
NAND3X1  g068(.A(n182_1), .B(G26), .C(G12), .Y(n183));
AOI21X1  g069(.A0(n181), .A1(n180), .B0(n183), .Y(n184));
OAI21X1  g070(.A0(n179), .A1(n169), .B0(n184), .Y(n185));
NOR3X1   g071(.A(n185), .B(n178), .C(n168), .Y(G90));
NAND2X1  g072(.A(G28), .B(G12), .Y(n187_1));
NAND2X1  g073(.A(G13), .B(G11), .Y(n188));
NOR2X1   g074(.A(n188), .B(n187_1), .Y(G92));
OR2X1    g075(.A(n140), .B(n134), .Y(n190));
NAND4X1  g076(.A(n190), .B(G74), .C(G30), .D(n143), .Y(G95BF));
NAND3X1  g077(.A(G73), .B(G31), .C(n165), .Y(G96BF));
NAND3X1  g078(.A(n138), .B(G72), .C(G32), .Y(G97BF));
NAND3X1  g079(.A(G71), .B(G33), .C(n165), .Y(G98BF));
NAND4X1  g080(.A(n128), .B(G70), .C(G34), .D(n132_1), .Y(G99BF));
NAND3X1  g081(.A(G69), .B(G35), .C(n165), .Y(G100BF));
NAND4X1  g082(.A(n120), .B(G68), .C(G36), .D(n123), .Y(G101BF));
NOR4X1   g083(.A(n127), .B(n151), .C(G2), .D(n139), .Y(n122));
NOR3X1   g084(.A(n124), .B(n118), .C(G2), .Y(n132));
NOR2X1   g085(.A(n171), .B(G89BF), .Y(n137));
MX2X1    g086(.A(G70), .B(n175), .S0(G88BF), .Y(n142));
OAI21X1  g087(.A0(n169), .A1(G88BF), .B0(n175), .Y(n147));
INVX1    g088(.A(n172_1), .Y(n203));
MX2X1    g089(.A(n203), .B(G72), .S0(n138), .Y(n152));
OAI21X1  g090(.A0(G87BF), .A1(n170), .B0(n203), .Y(n157));
MX2X1    g091(.A(G74), .B(n166), .S0(G86BF), .Y(n162));
OAI21X1  g092(.A0(G86BF), .A1(n164), .B0(n166), .Y(n167));
NAND2X1  g093(.A(n117), .B(n126), .Y(n208));
NAND4X1  g094(.A(n139), .B(n125), .C(G8), .D(n166), .Y(n209));
NOR4X1   g095(.A(G86BF), .B(n127), .C(n164), .D(n209), .Y(n210));
AOI21X1  g096(.A0(n117), .A1(G8), .B0(n210), .Y(n211));
NAND2X1  g097(.A(n211), .B(n208), .Y(n172));
NAND4X1  g098(.A(n138), .B(G72), .C(G5), .D(n203), .Y(n213));
NOR2X1   g099(.A(n213), .B(n151), .Y(n214));
OAI21X1  g100(.A0(n133), .A1(n117_1), .B0(n214), .Y(n215));
OAI21X1  g101(.A0(G5), .A1(n126), .B0(n147_1), .Y(n216));
OAI21X1  g102(.A0(n215), .A1(n117), .B0(n216), .Y(n177));
NAND4X1  g103(.A(n139), .B(n125), .C(G6), .D(n175), .Y(n218));
OR2X1    g104(.A(n218), .B(n169), .Y(n219));
OAI21X1  g105(.A0(G6), .A1(n126), .B0(n127), .Y(n220));
OAI21X1  g106(.A0(n219), .A1(n117), .B0(n220), .Y(n182));
INVX1    g107(.A(G1), .Y(n222));
OR4X1    g108(.A(n147_1), .B(n127), .C(n222), .D(n171), .Y(n223));
OAI21X1  g109(.A0(n126), .A1(G1), .B0(n151), .Y(n224));
OAI21X1  g110(.A0(n223), .A1(n117), .B0(n224), .Y(n187));
NOR3X1   g111(.A(n208), .B(n147_1), .C(n134), .Y(n192));
NOR4X1   g112(.A(n151), .B(n117_1), .C(G2), .D(n133), .Y(n202));
BUFX1    g113(.A(G27), .Y(G91));
BUFX1    g114(.A(G29), .Y(G94));
NOR4X1   g115(.A(n127), .B(n151), .C(G2), .D(n139), .Y(n197));
NOR3X1   g116(.A(n124), .B(n118), .C(G2), .Y(n207));
endmodule
