//Converted to Combinational (Partial output: n7440) , Module name: s38417_n7440 , Timestamp: 2018-12-03T15:51:14.854831 
module s38417_n7440 ( g2625, g2682, g2619, g2679, g2685, g2624, g185, g2616, g2993, g3006, g3010, g3032, g3036, g2598, g2670, g2676, g2673, g2998, g3024, g3002, g3013, g3018, g3028, g2656, g2655, g2657, g2659, g2658, g2660, g2650, g2649, g2651, g2661, g2667, g2664, g2639, g2564, g2641, g2454, g2400, g2412, g2458, g2456, g2406, g2424, g2428, g2426, g2653, g2652, g2654, g2439, g2443, g2441, g2469, g2399, g2471, g2643, g2647, g2645, n7440 );
input g2625, g2682, g2619, g2679, g2685, g2624, g185, g2616, g2993, g3006, g3010, g3032, g3036, g2598, g2670, g2676, g2673, g2998, g3024, g3002, g3013, g3018, g3028, g2656, g2655, g2657, g2659, g2658, g2660, g2650, g2649, g2651, g2661, g2667, g2664, g2639, g2564, g2641, g2454, g2400, g2412, g2458, g2456, g2406, g2424, g2428, g2426, g2653, g2652, g2654, g2439, g2443, g2441, g2469, g2399, g2471, g2643, g2647, g2645;
output n7440;
wire n9164, n5982, n9044, n9163, n9161, n5981_1, n9042, n9043, n9135, n9162, n9154, n9089, n5976_1, n5980, n9134, n9119, n9125, n9130, n9151, n9079, n9088, n9084, n9085, n5971_1, n5975, n5979, n9116, n9131, n9133, n9132, n9118, n9105, n9113, n9115, n9124, n9120, n9122, n9123, n9129, n9126, n9127, n9128, n9142, n9146, n9150, n9078, n9074, n9075, n9086, n9087, n7285, n5970, n5974, n5972, n5973, n5977, n5978, n9104, n9097, n9013, n9014, n9017, n9019, n9020, n9027, n9107, n9117, n9094, n9098, n9101, n9112, n7480, n9069, n9114, n9030, n9111, n7475, n7490, n9121, n9025, n9026, n9141, n9137, n9139, n9140, n9143, n9144, n9145, n9147, n9148, n9149, n9076, n9077, n7130, n9000, n9001, n9102, n9103, n9095, n9096, n5326, n8978, n9003, n9015, n9016, n9099, n9100, n9108, n9109, n9110, n9021, n7485, n9136, n9138, n9054, n8982, n8983;
MX2X1    g4120(.A(g2682), .B(n9164), .S0(g2625), .Y(n7440));
AOI22X1  g4118(.A0(n9161), .A1(n9163), .B0(n9044), .B1(n5982), .Y(n9164));
INVX1    g0939(.A(n5981_1), .Y(n5982));
AND2X1   g3998(.A(n9043), .B(n9042), .Y(n9044));
AOI21X1  g4117(.A0(n9162), .A1(n9135), .B0(n5982), .Y(n9163));
NAND3X1  g4115(.A(n9135), .B(n9089), .C(n9154), .Y(n9161));
NOR2X1   g0938(.A(n5980), .B(n5976_1), .Y(n5981_1));
NAND2X1  g3996(.A(g2679), .B(g2619), .Y(n9042));
AOI22X1  g3997(.A0(g2682), .A1(g2625), .B0(g2624), .B1(g2685), .Y(n9043));
NOR4X1   g4089(.A(n9130), .B(n9125), .C(n9119), .D(n9134), .Y(n9135));
NOR2X1   g4116(.A(n9151), .B(n9154), .Y(n9162));
INVX1    g4108(.A(n9079), .Y(n9154));
AOI21X1  g4043(.A0(n9085), .A1(n9084), .B0(n9088), .Y(n9089));
NAND2X1  g0933(.A(n5975), .B(n5971_1), .Y(n5976_1));
INVX1    g0937(.A(n5979), .Y(n5980));
OAI22X1  g4088(.A0(n9132), .A1(n9133), .B0(n9131), .B1(n9116), .Y(n9134));
NAND4X1  g4073(.A(n9115), .B(n9113), .C(n9105), .D(n9118), .Y(n9119));
NAND4X1  g4079(.A(n9123), .B(n9122), .C(n9120), .D(n9124), .Y(n9125));
NAND4X1  g4084(.A(n9128), .B(n9127), .C(n9126), .D(n9129), .Y(n9130));
NOR3X1   g4105(.A(n9150), .B(n9146), .C(n9142), .Y(n9151));
AOI21X1  g4033(.A0(n9075), .A1(n9074), .B0(n9078), .Y(n9079));
NAND2X1  g4042(.A(n9087), .B(n9086), .Y(n9088));
INVX1    g4038(.A(n7285), .Y(n9084));
AND2X1   g4039(.A(g2616), .B(g185), .Y(n9085));
NOR3X1   g0928(.A(g3006), .B(n5970), .C(g2993), .Y(n5971_1));
NOR4X1   g0932(.A(g3010), .B(n5973), .C(n5972), .D(n5974), .Y(n5975));
NOR4X1   g0936(.A(g3036), .B(n5978), .C(n5977), .D(g3032), .Y(n5979));
INVX1    g4070(.A(n9104), .Y(n9116));
OR4X1    g4085(.A(n9017), .B(n9014), .C(n9013), .D(n9097), .Y(n9131));
OR4X1    g4087(.A(n9027), .B(n9020), .C(n9019), .D(n9104), .Y(n9133));
OR2X1    g4086(.A(n9107), .B(n9097), .Y(n9132));
NAND3X1  g4072(.A(n9117), .B(n9116), .C(n9107), .Y(n9118));
OR4X1    g4059(.A(n9101), .B(n9098), .C(n9094), .D(n9104), .Y(n9105));
OR4X1    g4067(.A(n9097), .B(n9017), .C(n7480), .D(n9112), .Y(n9113));
NAND3X1  g4069(.A(n9114), .B(n9107), .C(n9069), .Y(n9115));
OR4X1    g4078(.A(n9107), .B(n9027), .C(n9030), .D(n9104), .Y(n9124));
OR4X1    g4074(.A(n9097), .B(n7490), .C(n7475), .D(n9111), .Y(n9120));
NAND3X1  g4076(.A(n9121), .B(n7490), .C(n9017), .Y(n9122));
NAND4X1  g4077(.A(n9097), .B(n7490), .C(n7475), .D(n9111), .Y(n9123));
OR4X1    g4083(.A(n9026), .B(n9025), .C(n9030), .D(n9111), .Y(n9129));
OR4X1    g4080(.A(n9097), .B(n9027), .C(n9030), .D(n9107), .Y(n9126));
OAI21X1  g4081(.A0(n9020), .A1(n9019), .B0(n9114), .Y(n9127));
OR4X1    g4082(.A(n9101), .B(n9097), .C(n9017), .D(n9116), .Y(n9128));
OR4X1    g4096(.A(n9140), .B(n9139), .C(n9137), .D(n9141), .Y(n9142));
NAND3X1  g4100(.A(n9145), .B(n9144), .C(n9143), .Y(n9146));
NAND3X1  g4104(.A(n9149), .B(n9148), .C(n9147), .Y(n9150));
NAND2X1  g4032(.A(n9077), .B(n9076), .Y(n9078));
INVX1    g4028(.A(n7130), .Y(n9074));
AND2X1   g4029(.A(g2598), .B(g185), .Y(n9075));
NAND2X1  g4040(.A(g2670), .B(g2619), .Y(n9086));
AOI22X1  g4041(.A0(g2673), .A1(g2625), .B0(g2624), .B1(g2676), .Y(n9087));
AND2X1   g3956(.A(n9001), .B(n9000), .Y(n7285));
INVX1    g0927(.A(g2998), .Y(n5970));
INVX1    g0931(.A(g3024), .Y(n5974));
INVX1    g0929(.A(g3002), .Y(n5972));
INVX1    g0930(.A(g3013), .Y(n5973));
INVX1    g0934(.A(g3018), .Y(n5977));
INVX1    g0935(.A(g3028), .Y(n5978));
AND2X1   g4058(.A(n9103), .B(n9102), .Y(n9104));
AND2X1   g4051(.A(n9096), .B(n9095), .Y(n9097));
NOR2X1   g3967(.A(g2656), .B(n5326), .Y(n9013));
OAI22X1  g3968(.A0(g2657), .A1(n9003), .B0(n8978), .B1(g2655), .Y(n9014));
NOR2X1   g3971(.A(n9016), .B(n9015), .Y(n9017));
NOR2X1   g3973(.A(g2659), .B(n5326), .Y(n9019));
OAI22X1  g3974(.A0(g2660), .A1(n9003), .B0(n8978), .B1(g2658), .Y(n9020));
NOR2X1   g3981(.A(n9026), .B(n9025), .Y(n9027));
INVX1    g4061(.A(n9101), .Y(n9107));
NOR4X1   g4071(.A(n9026), .B(n9025), .C(n9030), .D(n9097), .Y(n9117));
OR4X1    g4048(.A(n9025), .B(n9016), .C(n9015), .D(n9026), .Y(n9094));
INVX1    g4052(.A(n9097), .Y(n9098));
AND2X1   g4055(.A(n9100), .B(n9099), .Y(n9101));
NAND2X1  g4066(.A(n9111), .B(n9107), .Y(n9112));
INVX1    g4060(.A(n9030), .Y(n7480));
NOR4X1   g4023(.A(n9015), .B(n9014), .C(n9013), .D(n9016), .Y(n9069));
AND2X1   g4068(.A(n9104), .B(n9097), .Y(n9114));
NOR2X1   g3984(.A(n9014), .B(n9013), .Y(n9030));
NAND3X1  g4065(.A(n9110), .B(n9109), .C(n9108), .Y(n9111));
INVX1    g3978(.A(n9021), .Y(n7475));
INVX1    g4015(.A(n9027), .Y(n7490));
AND2X1   g4075(.A(n9101), .B(n9097), .Y(n9121));
NOR2X1   g3979(.A(g2650), .B(n5326), .Y(n9025));
OAI22X1  g3980(.A0(g2651), .A1(n9003), .B0(n8978), .B1(g2649), .Y(n9026));
NOR4X1   g4095(.A(n9098), .B(n9027), .C(n9030), .D(n9112), .Y(n9141));
NOR3X1   g4091(.A(n9136), .B(n9027), .C(n7485), .Y(n9137));
NOR2X1   g4093(.A(n9138), .B(n9094), .Y(n9139));
NOR4X1   g4094(.A(n9097), .B(n9094), .C(n7475), .D(n9116), .Y(n9140));
NAND4X1  g4097(.A(n9101), .B(n9027), .C(n7485), .D(n9116), .Y(n9143));
OR4X1    g4098(.A(n9101), .B(n9097), .C(n9021), .D(n9104), .Y(n9144));
OR4X1    g4099(.A(n9098), .B(n9027), .C(n9017), .D(n9116), .Y(n9145));
NAND2X1  g4101(.A(n9117), .B(n9101), .Y(n9147));
NAND2X1  g4102(.A(n9121), .B(n9054), .Y(n9148));
OR4X1    g4103(.A(n9027), .B(n7485), .C(n7480), .D(n9111), .Y(n9149));
NAND2X1  g4030(.A(g2661), .B(g2619), .Y(n9076));
AOI22X1  g4031(.A0(g2664), .A1(g2625), .B0(g2624), .B1(g2667), .Y(n9077));
AND2X1   g3938(.A(n8983), .B(n8982), .Y(n7130));
NAND2X1  g3954(.A(g2639), .B(g2619), .Y(n9000));
AOI22X1  g3955(.A0(g2641), .A1(g2625), .B0(g2624), .B1(g2564), .Y(n9001));
NAND2X1  g4056(.A(g2400), .B(g2454), .Y(n9102));
AOI22X1  g4057(.A0(g2406), .A1(g2456), .B0(g2458), .B1(g2412), .Y(n9103));
NAND2X1  g4049(.A(g2400), .B(g2424), .Y(n9095));
AOI22X1  g4050(.A0(g2406), .A1(g2426), .B0(g2428), .B1(g2412), .Y(n9096));
INVX1    g0284(.A(g2619), .Y(n5326));
INVX1    g3932(.A(g2624), .Y(n8978));
INVX1    g3957(.A(g2625), .Y(n9003));
NOR2X1   g3969(.A(g2653), .B(n5326), .Y(n9015));
OAI22X1  g3970(.A0(g2654), .A1(n9003), .B0(n8978), .B1(g2652), .Y(n9016));
NAND2X1  g4053(.A(g2400), .B(g2439), .Y(n9099));
AOI22X1  g4054(.A0(g2406), .A1(g2441), .B0(g2443), .B1(g2412), .Y(n9100));
NAND2X1  g4062(.A(g2400), .B(g2469), .Y(n9108));
NAND2X1  g4063(.A(g2412), .B(g2399), .Y(n9109));
NAND2X1  g4064(.A(g2406), .B(g2471), .Y(n9110));
NOR2X1   g3975(.A(n9020), .B(n9019), .Y(n9021));
INVX1    g3977(.A(n9017), .Y(n7485));
NAND4X1  g4090(.A(n9107), .B(n9097), .C(n9021), .D(n9116), .Y(n9136));
NAND4X1  g4092(.A(n9107), .B(n9098), .C(n9030), .D(n9111), .Y(n9138));
NOR3X1   g4008(.A(n9017), .B(n9014), .C(n9013), .Y(n9054));
NAND2X1  g3936(.A(g2643), .B(g2619), .Y(n8982));
AOI22X1  g3937(.A0(g2645), .A1(g2625), .B0(g2624), .B1(g2647), .Y(n8983));

endmodule
