// Benchmark "top" written by ABC on Wed Sep 23 03:15:56 2020

module top ( 
    \in0[0] , \in0[1] , \in0[2] , \in0[3] , \in0[4] , \in0[5] , \in0[6] ,
    \in0[7] , \in0[8] , \in0[9] , \in0[10] , \in0[11] , \in0[12] ,
    \in0[13] , \in0[14] , \in0[15] , \in0[16] , \in0[17] , \in0[18] ,
    \in0[19] , \in0[20] , \in0[21] , \in0[22] , \in0[23] , \in0[24] ,
    \in0[25] , \in0[26] , \in0[27] , \in0[28] , \in0[29] , \in0[30] ,
    \in0[31] , \in0[32] , \in0[33] , \in0[34] , \in0[35] , \in0[36] ,
    \in0[37] , \in0[38] , \in0[39] , \in0[40] , \in0[41] , \in0[42] ,
    \in0[43] , \in0[44] , \in0[45] , \in0[46] , \in0[47] , \in0[48] ,
    \in0[49] , \in0[50] , \in0[51] , \in0[52] , \in0[53] , \in0[54] ,
    \in0[55] , \in0[56] , \in0[57] , \in0[58] , \in0[59] , \in0[60] ,
    \in0[61] , \in0[62] , \in0[63] , \in0[64] , \in0[65] , \in0[66] ,
    \in0[67] , \in0[68] , \in0[69] , \in0[70] , \in0[71] , \in0[72] ,
    \in0[73] , \in0[74] , \in0[75] , \in0[76] , \in0[77] , \in0[78] ,
    \in0[79] , \in0[80] , \in0[81] , \in0[82] , \in0[83] , \in0[84] ,
    \in0[85] , \in0[86] , \in0[87] , \in0[88] , \in0[89] , \in0[90] ,
    \in0[91] , \in0[92] , \in0[93] , \in0[94] , \in0[95] , \in0[96] ,
    \in0[97] , \in0[98] , \in0[99] , \in0[100] , \in0[101] , \in0[102] ,
    \in0[103] , \in0[104] , \in0[105] , \in0[106] , \in0[107] , \in0[108] ,
    \in0[109] , \in0[110] , \in0[111] , \in0[112] , \in0[113] , \in0[114] ,
    \in0[115] , \in0[116] , \in0[117] , \in0[118] , \in0[119] , \in0[120] ,
    \in0[121] , \in0[122] , \in0[123] , \in0[124] , \in0[125] , \in0[126] ,
    \in0[127] , \in1[0] , \in1[1] , \in1[2] , \in1[3] , \in1[4] , \in1[5] ,
    \in1[6] , \in1[7] , \in1[8] , \in1[9] , \in1[10] , \in1[11] ,
    \in1[12] , \in1[13] , \in1[14] , \in1[15] , \in1[16] , \in1[17] ,
    \in1[18] , \in1[19] , \in1[20] , \in1[21] , \in1[22] , \in1[23] ,
    \in1[24] , \in1[25] , \in1[26] , \in1[27] , \in1[28] , \in1[29] ,
    \in1[30] , \in1[31] , \in1[32] , \in1[33] , \in1[34] , \in1[35] ,
    \in1[36] , \in1[37] , \in1[38] , \in1[39] , \in1[40] , \in1[41] ,
    \in1[42] , \in1[43] , \in1[44] , \in1[45] , \in1[46] , \in1[47] ,
    \in1[48] , \in1[49] , \in1[50] , \in1[51] , \in1[52] , \in1[53] ,
    \in1[54] , \in1[55] , \in1[56] , \in1[57] , \in1[58] , \in1[59] ,
    \in1[60] , \in1[61] , \in1[62] , \in1[63] , \in1[64] , \in1[65] ,
    \in1[66] , \in1[67] , \in1[68] , \in1[69] , \in1[70] , \in1[71] ,
    \in1[72] , \in1[73] , \in1[74] , \in1[75] , \in1[76] , \in1[77] ,
    \in1[78] , \in1[79] , \in1[80] , \in1[81] , \in1[82] , \in1[83] ,
    \in1[84] , \in1[85] , \in1[86] , \in1[87] , \in1[88] , \in1[89] ,
    \in1[90] , \in1[91] , \in1[92] , \in1[93] , \in1[94] , \in1[95] ,
    \in1[96] , \in1[97] , \in1[98] , \in1[99] , \in1[100] , \in1[101] ,
    \in1[102] , \in1[103] , \in1[104] , \in1[105] , \in1[106] , \in1[107] ,
    \in1[108] , \in1[109] , \in1[110] , \in1[111] , \in1[112] , \in1[113] ,
    \in1[114] , \in1[115] , \in1[116] , \in1[117] , \in1[118] , \in1[119] ,
    \in1[120] , \in1[121] , \in1[122] , \in1[123] , \in1[124] , \in1[125] ,
    \in1[126] , \in1[127] , \in2[0] , \in2[1] , \in2[2] , \in2[3] ,
    \in2[4] , \in2[5] , \in2[6] , \in2[7] , \in2[8] , \in2[9] , \in2[10] ,
    \in2[11] , \in2[12] , \in2[13] , \in2[14] , \in2[15] , \in2[16] ,
    \in2[17] , \in2[18] , \in2[19] , \in2[20] , \in2[21] , \in2[22] ,
    \in2[23] , \in2[24] , \in2[25] , \in2[26] , \in2[27] , \in2[28] ,
    \in2[29] , \in2[30] , \in2[31] , \in2[32] , \in2[33] , \in2[34] ,
    \in2[35] , \in2[36] , \in2[37] , \in2[38] , \in2[39] , \in2[40] ,
    \in2[41] , \in2[42] , \in2[43] , \in2[44] , \in2[45] , \in2[46] ,
    \in2[47] , \in2[48] , \in2[49] , \in2[50] , \in2[51] , \in2[52] ,
    \in2[53] , \in2[54] , \in2[55] , \in2[56] , \in2[57] , \in2[58] ,
    \in2[59] , \in2[60] , \in2[61] , \in2[62] , \in2[63] , \in2[64] ,
    \in2[65] , \in2[66] , \in2[67] , \in2[68] , \in2[69] , \in2[70] ,
    \in2[71] , \in2[72] , \in2[73] , \in2[74] , \in2[75] , \in2[76] ,
    \in2[77] , \in2[78] , \in2[79] , \in2[80] , \in2[81] , \in2[82] ,
    \in2[83] , \in2[84] , \in2[85] , \in2[86] , \in2[87] , \in2[88] ,
    \in2[89] , \in2[90] , \in2[91] , \in2[92] , \in2[93] , \in2[94] ,
    \in2[95] , \in2[96] , \in2[97] , \in2[98] , \in2[99] , \in2[100] ,
    \in2[101] , \in2[102] , \in2[103] , \in2[104] , \in2[105] , \in2[106] ,
    \in2[107] , \in2[108] , \in2[109] , \in2[110] , \in2[111] , \in2[112] ,
    \in2[113] , \in2[114] , \in2[115] , \in2[116] , \in2[117] , \in2[118] ,
    \in2[119] , \in2[120] , \in2[121] , \in2[122] , \in2[123] , \in2[124] ,
    \in2[125] , \in2[126] , \in2[127] , \in3[0] , \in3[1] , \in3[2] ,
    \in3[3] , \in3[4] , \in3[5] , \in3[6] , \in3[7] , \in3[8] , \in3[9] ,
    \in3[10] , \in3[11] , \in3[12] , \in3[13] , \in3[14] , \in3[15] ,
    \in3[16] , \in3[17] , \in3[18] , \in3[19] , \in3[20] , \in3[21] ,
    \in3[22] , \in3[23] , \in3[24] , \in3[25] , \in3[26] , \in3[27] ,
    \in3[28] , \in3[29] , \in3[30] , \in3[31] , \in3[32] , \in3[33] ,
    \in3[34] , \in3[35] , \in3[36] , \in3[37] , \in3[38] , \in3[39] ,
    \in3[40] , \in3[41] , \in3[42] , \in3[43] , \in3[44] , \in3[45] ,
    \in3[46] , \in3[47] , \in3[48] , \in3[49] , \in3[50] , \in3[51] ,
    \in3[52] , \in3[53] , \in3[54] , \in3[55] , \in3[56] , \in3[57] ,
    \in3[58] , \in3[59] , \in3[60] , \in3[61] , \in3[62] , \in3[63] ,
    \in3[64] , \in3[65] , \in3[66] , \in3[67] , \in3[68] , \in3[69] ,
    \in3[70] , \in3[71] , \in3[72] , \in3[73] , \in3[74] , \in3[75] ,
    \in3[76] , \in3[77] , \in3[78] , \in3[79] , \in3[80] , \in3[81] ,
    \in3[82] , \in3[83] , \in3[84] , \in3[85] , \in3[86] , \in3[87] ,
    \in3[88] , \in3[89] , \in3[90] , \in3[91] , \in3[92] , \in3[93] ,
    \in3[94] , \in3[95] , \in3[96] , \in3[97] , \in3[98] , \in3[99] ,
    \in3[100] , \in3[101] , \in3[102] , \in3[103] , \in3[104] , \in3[105] ,
    \in3[106] , \in3[107] , \in3[108] , \in3[109] , \in3[110] , \in3[111] ,
    \in3[112] , \in3[113] , \in3[114] , \in3[115] , \in3[116] , \in3[117] ,
    \in3[118] , \in3[119] , \in3[120] , \in3[121] , \in3[122] , \in3[123] ,
    \in3[124] , \in3[125] , \in3[126] , \in3[127] ,
    \result[0] , \result[1] , \result[2] , \result[3] , \result[4] ,
    \result[5] , \result[6] , \result[7] , \result[8] , \result[9] ,
    \result[10] , \result[11] , \result[12] , \result[13] , \result[14] ,
    \result[15] , \result[16] , \result[17] , \result[18] , \result[19] ,
    \result[20] , \result[21] , \result[22] , \result[23] , \result[24] ,
    \result[25] , \result[26] , \result[27] , \result[28] , \result[29] ,
    \result[30] , \result[31] , \result[32] , \result[33] , \result[34] ,
    \result[35] , \result[36] , \result[37] , \result[38] , \result[39] ,
    \result[40] , \result[41] , \result[42] , \result[43] , \result[44] ,
    \result[45] , \result[46] , \result[47] , \result[48] , \result[49] ,
    \result[50] , \result[51] , \result[52] , \result[53] , \result[54] ,
    \result[55] , \result[56] , \result[57] , \result[58] , \result[59] ,
    \result[60] , \result[61] , \result[62] , \result[63] , \result[64] ,
    \result[65] , \result[66] , \result[67] , \result[68] , \result[69] ,
    \result[70] , \result[71] , \result[72] , \result[73] , \result[74] ,
    \result[75] , \result[76] , \result[77] , \result[78] , \result[79] ,
    \result[80] , \result[81] , \result[82] , \result[83] , \result[84] ,
    \result[85] , \result[86] , \result[87] , \result[88] , \result[89] ,
    \result[90] , \result[91] , \result[92] , \result[93] , \result[94] ,
    \result[95] , \result[96] , \result[97] , \result[98] , \result[99] ,
    \result[100] , \result[101] , \result[102] , \result[103] ,
    \result[104] , \result[105] , \result[106] , \result[107] ,
    \result[108] , \result[109] , \result[110] , \result[111] ,
    \result[112] , \result[113] , \result[114] , \result[115] ,
    \result[116] , \result[117] , \result[118] , \result[119] ,
    \result[120] , \result[121] , \result[122] , \result[123] ,
    \result[124] , \result[125] , \result[126] , \result[127] ,
    \address[0] , \address[1]   );
  input  \in0[0] , \in0[1] , \in0[2] , \in0[3] , \in0[4] , \in0[5] ,
    \in0[6] , \in0[7] , \in0[8] , \in0[9] , \in0[10] , \in0[11] ,
    \in0[12] , \in0[13] , \in0[14] , \in0[15] , \in0[16] , \in0[17] ,
    \in0[18] , \in0[19] , \in0[20] , \in0[21] , \in0[22] , \in0[23] ,
    \in0[24] , \in0[25] , \in0[26] , \in0[27] , \in0[28] , \in0[29] ,
    \in0[30] , \in0[31] , \in0[32] , \in0[33] , \in0[34] , \in0[35] ,
    \in0[36] , \in0[37] , \in0[38] , \in0[39] , \in0[40] , \in0[41] ,
    \in0[42] , \in0[43] , \in0[44] , \in0[45] , \in0[46] , \in0[47] ,
    \in0[48] , \in0[49] , \in0[50] , \in0[51] , \in0[52] , \in0[53] ,
    \in0[54] , \in0[55] , \in0[56] , \in0[57] , \in0[58] , \in0[59] ,
    \in0[60] , \in0[61] , \in0[62] , \in0[63] , \in0[64] , \in0[65] ,
    \in0[66] , \in0[67] , \in0[68] , \in0[69] , \in0[70] , \in0[71] ,
    \in0[72] , \in0[73] , \in0[74] , \in0[75] , \in0[76] , \in0[77] ,
    \in0[78] , \in0[79] , \in0[80] , \in0[81] , \in0[82] , \in0[83] ,
    \in0[84] , \in0[85] , \in0[86] , \in0[87] , \in0[88] , \in0[89] ,
    \in0[90] , \in0[91] , \in0[92] , \in0[93] , \in0[94] , \in0[95] ,
    \in0[96] , \in0[97] , \in0[98] , \in0[99] , \in0[100] , \in0[101] ,
    \in0[102] , \in0[103] , \in0[104] , \in0[105] , \in0[106] , \in0[107] ,
    \in0[108] , \in0[109] , \in0[110] , \in0[111] , \in0[112] , \in0[113] ,
    \in0[114] , \in0[115] , \in0[116] , \in0[117] , \in0[118] , \in0[119] ,
    \in0[120] , \in0[121] , \in0[122] , \in0[123] , \in0[124] , \in0[125] ,
    \in0[126] , \in0[127] , \in1[0] , \in1[1] , \in1[2] , \in1[3] ,
    \in1[4] , \in1[5] , \in1[6] , \in1[7] , \in1[8] , \in1[9] , \in1[10] ,
    \in1[11] , \in1[12] , \in1[13] , \in1[14] , \in1[15] , \in1[16] ,
    \in1[17] , \in1[18] , \in1[19] , \in1[20] , \in1[21] , \in1[22] ,
    \in1[23] , \in1[24] , \in1[25] , \in1[26] , \in1[27] , \in1[28] ,
    \in1[29] , \in1[30] , \in1[31] , \in1[32] , \in1[33] , \in1[34] ,
    \in1[35] , \in1[36] , \in1[37] , \in1[38] , \in1[39] , \in1[40] ,
    \in1[41] , \in1[42] , \in1[43] , \in1[44] , \in1[45] , \in1[46] ,
    \in1[47] , \in1[48] , \in1[49] , \in1[50] , \in1[51] , \in1[52] ,
    \in1[53] , \in1[54] , \in1[55] , \in1[56] , \in1[57] , \in1[58] ,
    \in1[59] , \in1[60] , \in1[61] , \in1[62] , \in1[63] , \in1[64] ,
    \in1[65] , \in1[66] , \in1[67] , \in1[68] , \in1[69] , \in1[70] ,
    \in1[71] , \in1[72] , \in1[73] , \in1[74] , \in1[75] , \in1[76] ,
    \in1[77] , \in1[78] , \in1[79] , \in1[80] , \in1[81] , \in1[82] ,
    \in1[83] , \in1[84] , \in1[85] , \in1[86] , \in1[87] , \in1[88] ,
    \in1[89] , \in1[90] , \in1[91] , \in1[92] , \in1[93] , \in1[94] ,
    \in1[95] , \in1[96] , \in1[97] , \in1[98] , \in1[99] , \in1[100] ,
    \in1[101] , \in1[102] , \in1[103] , \in1[104] , \in1[105] , \in1[106] ,
    \in1[107] , \in1[108] , \in1[109] , \in1[110] , \in1[111] , \in1[112] ,
    \in1[113] , \in1[114] , \in1[115] , \in1[116] , \in1[117] , \in1[118] ,
    \in1[119] , \in1[120] , \in1[121] , \in1[122] , \in1[123] , \in1[124] ,
    \in1[125] , \in1[126] , \in1[127] , \in2[0] , \in2[1] , \in2[2] ,
    \in2[3] , \in2[4] , \in2[5] , \in2[6] , \in2[7] , \in2[8] , \in2[9] ,
    \in2[10] , \in2[11] , \in2[12] , \in2[13] , \in2[14] , \in2[15] ,
    \in2[16] , \in2[17] , \in2[18] , \in2[19] , \in2[20] , \in2[21] ,
    \in2[22] , \in2[23] , \in2[24] , \in2[25] , \in2[26] , \in2[27] ,
    \in2[28] , \in2[29] , \in2[30] , \in2[31] , \in2[32] , \in2[33] ,
    \in2[34] , \in2[35] , \in2[36] , \in2[37] , \in2[38] , \in2[39] ,
    \in2[40] , \in2[41] , \in2[42] , \in2[43] , \in2[44] , \in2[45] ,
    \in2[46] , \in2[47] , \in2[48] , \in2[49] , \in2[50] , \in2[51] ,
    \in2[52] , \in2[53] , \in2[54] , \in2[55] , \in2[56] , \in2[57] ,
    \in2[58] , \in2[59] , \in2[60] , \in2[61] , \in2[62] , \in2[63] ,
    \in2[64] , \in2[65] , \in2[66] , \in2[67] , \in2[68] , \in2[69] ,
    \in2[70] , \in2[71] , \in2[72] , \in2[73] , \in2[74] , \in2[75] ,
    \in2[76] , \in2[77] , \in2[78] , \in2[79] , \in2[80] , \in2[81] ,
    \in2[82] , \in2[83] , \in2[84] , \in2[85] , \in2[86] , \in2[87] ,
    \in2[88] , \in2[89] , \in2[90] , \in2[91] , \in2[92] , \in2[93] ,
    \in2[94] , \in2[95] , \in2[96] , \in2[97] , \in2[98] , \in2[99] ,
    \in2[100] , \in2[101] , \in2[102] , \in2[103] , \in2[104] , \in2[105] ,
    \in2[106] , \in2[107] , \in2[108] , \in2[109] , \in2[110] , \in2[111] ,
    \in2[112] , \in2[113] , \in2[114] , \in2[115] , \in2[116] , \in2[117] ,
    \in2[118] , \in2[119] , \in2[120] , \in2[121] , \in2[122] , \in2[123] ,
    \in2[124] , \in2[125] , \in2[126] , \in2[127] , \in3[0] , \in3[1] ,
    \in3[2] , \in3[3] , \in3[4] , \in3[5] , \in3[6] , \in3[7] , \in3[8] ,
    \in3[9] , \in3[10] , \in3[11] , \in3[12] , \in3[13] , \in3[14] ,
    \in3[15] , \in3[16] , \in3[17] , \in3[18] , \in3[19] , \in3[20] ,
    \in3[21] , \in3[22] , \in3[23] , \in3[24] , \in3[25] , \in3[26] ,
    \in3[27] , \in3[28] , \in3[29] , \in3[30] , \in3[31] , \in3[32] ,
    \in3[33] , \in3[34] , \in3[35] , \in3[36] , \in3[37] , \in3[38] ,
    \in3[39] , \in3[40] , \in3[41] , \in3[42] , \in3[43] , \in3[44] ,
    \in3[45] , \in3[46] , \in3[47] , \in3[48] , \in3[49] , \in3[50] ,
    \in3[51] , \in3[52] , \in3[53] , \in3[54] , \in3[55] , \in3[56] ,
    \in3[57] , \in3[58] , \in3[59] , \in3[60] , \in3[61] , \in3[62] ,
    \in3[63] , \in3[64] , \in3[65] , \in3[66] , \in3[67] , \in3[68] ,
    \in3[69] , \in3[70] , \in3[71] , \in3[72] , \in3[73] , \in3[74] ,
    \in3[75] , \in3[76] , \in3[77] , \in3[78] , \in3[79] , \in3[80] ,
    \in3[81] , \in3[82] , \in3[83] , \in3[84] , \in3[85] , \in3[86] ,
    \in3[87] , \in3[88] , \in3[89] , \in3[90] , \in3[91] , \in3[92] ,
    \in3[93] , \in3[94] , \in3[95] , \in3[96] , \in3[97] , \in3[98] ,
    \in3[99] , \in3[100] , \in3[101] , \in3[102] , \in3[103] , \in3[104] ,
    \in3[105] , \in3[106] , \in3[107] , \in3[108] , \in3[109] , \in3[110] ,
    \in3[111] , \in3[112] , \in3[113] , \in3[114] , \in3[115] , \in3[116] ,
    \in3[117] , \in3[118] , \in3[119] , \in3[120] , \in3[121] , \in3[122] ,
    \in3[123] , \in3[124] , \in3[125] , \in3[126] , \in3[127] ;
  output \result[0] , \result[1] , \result[2] , \result[3] , \result[4] ,
    \result[5] , \result[6] , \result[7] , \result[8] , \result[9] ,
    \result[10] , \result[11] , \result[12] , \result[13] , \result[14] ,
    \result[15] , \result[16] , \result[17] , \result[18] , \result[19] ,
    \result[20] , \result[21] , \result[22] , \result[23] , \result[24] ,
    \result[25] , \result[26] , \result[27] , \result[28] , \result[29] ,
    \result[30] , \result[31] , \result[32] , \result[33] , \result[34] ,
    \result[35] , \result[36] , \result[37] , \result[38] , \result[39] ,
    \result[40] , \result[41] , \result[42] , \result[43] , \result[44] ,
    \result[45] , \result[46] , \result[47] , \result[48] , \result[49] ,
    \result[50] , \result[51] , \result[52] , \result[53] , \result[54] ,
    \result[55] , \result[56] , \result[57] , \result[58] , \result[59] ,
    \result[60] , \result[61] , \result[62] , \result[63] , \result[64] ,
    \result[65] , \result[66] , \result[67] , \result[68] , \result[69] ,
    \result[70] , \result[71] , \result[72] , \result[73] , \result[74] ,
    \result[75] , \result[76] , \result[77] , \result[78] , \result[79] ,
    \result[80] , \result[81] , \result[82] , \result[83] , \result[84] ,
    \result[85] , \result[86] , \result[87] , \result[88] , \result[89] ,
    \result[90] , \result[91] , \result[92] , \result[93] , \result[94] ,
    \result[95] , \result[96] , \result[97] , \result[98] , \result[99] ,
    \result[100] , \result[101] , \result[102] , \result[103] ,
    \result[104] , \result[105] , \result[106] , \result[107] ,
    \result[108] , \result[109] , \result[110] , \result[111] ,
    \result[112] , \result[113] , \result[114] , \result[115] ,
    \result[116] , \result[117] , \result[118] , \result[119] ,
    \result[120] , \result[121] , \result[122] , \result[123] ,
    \result[124] , \result[125] , \result[126] , \result[127] ,
    \address[0] , \address[1] ;
  wire new_n643_, new_n644_, new_n645_, new_n646_, new_n647_, new_n648_,
    new_n649_, new_n650_, new_n651_, new_n652_, new_n653_, new_n654_,
    new_n655_, new_n656_, new_n657_, new_n658_, new_n659_, new_n660_,
    new_n661_, new_n662_, new_n663_, new_n664_, new_n665_, new_n666_,
    new_n667_, new_n668_, new_n669_, new_n670_, new_n671_, new_n672_,
    new_n673_, new_n674_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n687_, new_n688_, new_n689_, new_n690_,
    new_n691_, new_n692_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n817_, new_n818_, new_n819_, new_n820_, new_n821_, new_n822_,
    new_n823_, new_n824_, new_n825_, new_n826_, new_n827_, new_n828_,
    new_n829_, new_n830_, new_n831_, new_n832_, new_n833_, new_n834_,
    new_n835_, new_n836_, new_n837_, new_n838_, new_n839_, new_n840_,
    new_n841_, new_n842_, new_n843_, new_n844_, new_n845_, new_n846_,
    new_n847_, new_n848_, new_n849_, new_n850_, new_n851_, new_n852_,
    new_n853_, new_n854_, new_n855_, new_n856_, new_n857_, new_n858_,
    new_n859_, new_n860_, new_n861_, new_n862_, new_n863_, new_n864_,
    new_n865_, new_n866_, new_n867_, new_n868_, new_n869_, new_n870_,
    new_n871_, new_n872_, new_n873_, new_n874_, new_n875_, new_n876_,
    new_n877_, new_n878_, new_n879_, new_n880_, new_n881_, new_n882_,
    new_n883_, new_n884_, new_n885_, new_n886_, new_n887_, new_n888_,
    new_n889_, new_n890_, new_n891_, new_n892_, new_n893_, new_n894_,
    new_n895_, new_n896_, new_n897_, new_n898_, new_n899_, new_n900_,
    new_n901_, new_n902_, new_n903_, new_n904_, new_n905_, new_n906_,
    new_n907_, new_n908_, new_n909_, new_n910_, new_n911_, new_n912_,
    new_n913_, new_n914_, new_n915_, new_n916_, new_n917_, new_n918_,
    new_n919_, new_n920_, new_n921_, new_n922_, new_n923_, new_n924_,
    new_n925_, new_n926_, new_n927_, new_n928_, new_n929_, new_n930_,
    new_n931_, new_n932_, new_n933_, new_n934_, new_n935_, new_n936_,
    new_n937_, new_n938_, new_n939_, new_n940_, new_n941_, new_n942_,
    new_n943_, new_n944_, new_n945_, new_n946_, new_n947_, new_n948_,
    new_n949_, new_n950_, new_n951_, new_n952_, new_n953_, new_n954_,
    new_n955_, new_n956_, new_n957_, new_n958_, new_n959_, new_n960_,
    new_n961_, new_n962_, new_n963_, new_n964_, new_n965_, new_n966_,
    new_n967_, new_n968_, new_n969_, new_n970_, new_n971_, new_n972_,
    new_n973_, new_n974_, new_n975_, new_n976_, new_n977_, new_n978_,
    new_n979_, new_n980_, new_n981_, new_n982_, new_n983_, new_n984_,
    new_n985_, new_n986_, new_n987_, new_n988_, new_n989_, new_n990_,
    new_n991_, new_n992_, new_n993_, new_n994_, new_n995_, new_n996_,
    new_n997_, new_n998_, new_n999_, new_n1000_, new_n1001_, new_n1002_,
    new_n1003_, new_n1004_, new_n1005_, new_n1006_, new_n1007_, new_n1008_,
    new_n1009_, new_n1010_, new_n1011_, new_n1012_, new_n1013_, new_n1014_,
    new_n1015_, new_n1016_, new_n1017_, new_n1018_, new_n1019_, new_n1020_,
    new_n1021_, new_n1022_, new_n1023_, new_n1024_, new_n1025_, new_n1026_,
    new_n1027_, new_n1028_, new_n1029_, new_n1030_, new_n1031_, new_n1032_,
    new_n1033_, new_n1034_, new_n1035_, new_n1036_, new_n1037_, new_n1038_,
    new_n1039_, new_n1040_, new_n1041_, new_n1042_, new_n1043_, new_n1044_,
    new_n1045_, new_n1046_, new_n1047_, new_n1048_, new_n1049_, new_n1050_,
    new_n1051_, new_n1052_, new_n1053_, new_n1054_, new_n1055_, new_n1056_,
    new_n1057_, new_n1058_, new_n1059_, new_n1060_, new_n1061_, new_n1062_,
    new_n1063_, new_n1064_, new_n1065_, new_n1066_, new_n1067_, new_n1068_,
    new_n1069_, new_n1070_, new_n1071_, new_n1072_, new_n1073_, new_n1074_,
    new_n1075_, new_n1076_, new_n1077_, new_n1078_, new_n1079_, new_n1080_,
    new_n1081_, new_n1082_, new_n1083_, new_n1084_, new_n1085_, new_n1086_,
    new_n1087_, new_n1088_, new_n1089_, new_n1090_, new_n1091_, new_n1092_,
    new_n1093_, new_n1094_, new_n1095_, new_n1096_, new_n1097_, new_n1098_,
    new_n1099_, new_n1100_, new_n1101_, new_n1102_, new_n1103_, new_n1104_,
    new_n1105_, new_n1106_, new_n1107_, new_n1108_, new_n1109_, new_n1110_,
    new_n1111_, new_n1112_, new_n1113_, new_n1114_, new_n1115_, new_n1116_,
    new_n1117_, new_n1118_, new_n1119_, new_n1120_, new_n1121_, new_n1122_,
    new_n1123_, new_n1124_, new_n1125_, new_n1126_, new_n1127_, new_n1128_,
    new_n1129_, new_n1130_, new_n1131_, new_n1132_, new_n1133_, new_n1134_,
    new_n1135_, new_n1136_, new_n1137_, new_n1138_, new_n1139_, new_n1140_,
    new_n1141_, new_n1142_, new_n1143_, new_n1144_, new_n1145_, new_n1146_,
    new_n1147_, new_n1148_, new_n1149_, new_n1150_, new_n1151_, new_n1152_,
    new_n1153_, new_n1154_, new_n1155_, new_n1156_, new_n1157_, new_n1158_,
    new_n1159_, new_n1160_, new_n1161_, new_n1162_, new_n1163_, new_n1164_,
    new_n1165_, new_n1166_, new_n1167_, new_n1168_, new_n1169_, new_n1170_,
    new_n1171_, new_n1172_, new_n1173_, new_n1174_, new_n1175_, new_n1176_,
    new_n1177_, new_n1178_, new_n1179_, new_n1180_, new_n1181_, new_n1182_,
    new_n1183_, new_n1184_, new_n1185_, new_n1186_, new_n1187_, new_n1188_,
    new_n1189_, new_n1190_, new_n1191_, new_n1192_, new_n1193_, new_n1194_,
    new_n1195_, new_n1196_, new_n1197_, new_n1198_, new_n1199_, new_n1200_,
    new_n1201_, new_n1202_, new_n1203_, new_n1204_, new_n1205_, new_n1206_,
    new_n1207_, new_n1208_, new_n1209_, new_n1210_, new_n1211_, new_n1212_,
    new_n1213_, new_n1214_, new_n1215_, new_n1216_, new_n1217_, new_n1218_,
    new_n1219_, new_n1220_, new_n1221_, new_n1222_, new_n1223_, new_n1224_,
    new_n1225_, new_n1226_, new_n1227_, new_n1228_, new_n1229_, new_n1230_,
    new_n1231_, new_n1232_, new_n1233_, new_n1234_, new_n1235_, new_n1236_,
    new_n1237_, new_n1238_, new_n1239_, new_n1240_, new_n1241_, new_n1242_,
    new_n1243_, new_n1244_, new_n1245_, new_n1246_, new_n1247_, new_n1248_,
    new_n1249_, new_n1250_, new_n1251_, new_n1252_, new_n1253_, new_n1254_,
    new_n1255_, new_n1256_, new_n1257_, new_n1258_, new_n1259_, new_n1260_,
    new_n1261_, new_n1262_, new_n1263_, new_n1264_, new_n1265_, new_n1266_,
    new_n1267_, new_n1268_, new_n1269_, new_n1270_, new_n1271_, new_n1272_,
    new_n1273_, new_n1274_, new_n1275_, new_n1276_, new_n1277_, new_n1278_,
    new_n1279_, new_n1280_, new_n1281_, new_n1282_, new_n1283_, new_n1284_,
    new_n1285_, new_n1286_, new_n1287_, new_n1288_, new_n1289_, new_n1290_,
    new_n1291_, new_n1292_, new_n1293_, new_n1294_, new_n1295_, new_n1296_,
    new_n1297_, new_n1298_, new_n1299_, new_n1300_, new_n1301_, new_n1302_,
    new_n1303_, new_n1304_, new_n1305_, new_n1306_, new_n1307_, new_n1308_,
    new_n1309_, new_n1310_, new_n1311_, new_n1312_, new_n1313_, new_n1314_,
    new_n1315_, new_n1316_, new_n1317_, new_n1318_, new_n1319_, new_n1320_,
    new_n1321_, new_n1322_, new_n1323_, new_n1324_, new_n1325_, new_n1326_,
    new_n1327_, new_n1328_, new_n1329_, new_n1330_, new_n1331_, new_n1332_,
    new_n1333_, new_n1334_, new_n1335_, new_n1336_, new_n1337_, new_n1338_,
    new_n1339_, new_n1340_, new_n1341_, new_n1342_, new_n1343_, new_n1344_,
    new_n1345_, new_n1346_, new_n1347_, new_n1348_, new_n1349_, new_n1350_,
    new_n1351_, new_n1352_, new_n1353_, new_n1354_, new_n1355_, new_n1356_,
    new_n1357_, new_n1358_, new_n1359_, new_n1360_, new_n1361_, new_n1362_,
    new_n1363_, new_n1364_, new_n1365_, new_n1366_, new_n1367_, new_n1368_,
    new_n1369_, new_n1370_, new_n1371_, new_n1372_, new_n1373_, new_n1374_,
    new_n1375_, new_n1376_, new_n1377_, new_n1378_, new_n1379_, new_n1380_,
    new_n1381_, new_n1382_, new_n1383_, new_n1384_, new_n1385_, new_n1386_,
    new_n1387_, new_n1388_, new_n1389_, new_n1390_, new_n1391_, new_n1392_,
    new_n1393_, new_n1394_, new_n1395_, new_n1396_, new_n1397_, new_n1398_,
    new_n1399_, new_n1400_, new_n1401_, new_n1402_, new_n1403_, new_n1404_,
    new_n1405_, new_n1406_, new_n1407_, new_n1408_, new_n1409_, new_n1410_,
    new_n1411_, new_n1412_, new_n1413_, new_n1414_, new_n1415_, new_n1416_,
    new_n1417_, new_n1418_, new_n1419_, new_n1420_, new_n1421_, new_n1422_,
    new_n1423_, new_n1424_, new_n1425_, new_n1426_, new_n1427_, new_n1428_,
    new_n1429_, new_n1430_, new_n1431_, new_n1432_, new_n1433_, new_n1434_,
    new_n1435_, new_n1436_, new_n1437_, new_n1438_, new_n1439_, new_n1440_,
    new_n1441_, new_n1442_, new_n1443_, new_n1444_, new_n1445_, new_n1446_,
    new_n1447_, new_n1448_, new_n1449_, new_n1450_, new_n1451_, new_n1452_,
    new_n1453_, new_n1454_, new_n1455_, new_n1456_, new_n1457_, new_n1458_,
    new_n1459_, new_n1460_, new_n1461_, new_n1462_, new_n1463_, new_n1464_,
    new_n1465_, new_n1466_, new_n1467_, new_n1468_, new_n1469_, new_n1470_,
    new_n1471_, new_n1472_, new_n1473_, new_n1474_, new_n1475_, new_n1476_,
    new_n1477_, new_n1478_, new_n1479_, new_n1480_, new_n1481_, new_n1482_,
    new_n1483_, new_n1484_, new_n1485_, new_n1486_, new_n1487_, new_n1488_,
    new_n1489_, new_n1490_, new_n1491_, new_n1492_, new_n1493_, new_n1494_,
    new_n1495_, new_n1496_, new_n1497_, new_n1498_, new_n1499_, new_n1500_,
    new_n1501_, new_n1502_, new_n1503_, new_n1504_, new_n1505_, new_n1506_,
    new_n1507_, new_n1508_, new_n1509_, new_n1510_, new_n1511_, new_n1512_,
    new_n1513_, new_n1514_, new_n1515_, new_n1516_, new_n1517_, new_n1518_,
    new_n1519_, new_n1520_, new_n1521_, new_n1522_, new_n1523_, new_n1524_,
    new_n1525_, new_n1526_, new_n1527_, new_n1528_, new_n1529_, new_n1530_,
    new_n1531_, new_n1532_, new_n1533_, new_n1534_, new_n1535_, new_n1536_,
    new_n1537_, new_n1538_, new_n1539_, new_n1540_, new_n1541_, new_n1542_,
    new_n1543_, new_n1544_, new_n1545_, new_n1546_, new_n1547_, new_n1548_,
    new_n1549_, new_n1550_, new_n1551_, new_n1552_, new_n1553_, new_n1554_,
    new_n1555_, new_n1556_, new_n1557_, new_n1558_, new_n1559_, new_n1560_,
    new_n1561_, new_n1562_, new_n1563_, new_n1564_, new_n1565_, new_n1566_,
    new_n1567_, new_n1568_, new_n1569_, new_n1570_, new_n1571_, new_n1572_,
    new_n1573_, new_n1574_, new_n1575_, new_n1576_, new_n1577_, new_n1578_,
    new_n1579_, new_n1580_, new_n1581_, new_n1582_, new_n1583_, new_n1584_,
    new_n1585_, new_n1586_, new_n1587_, new_n1588_, new_n1589_, new_n1590_,
    new_n1591_, new_n1592_, new_n1593_, new_n1594_, new_n1595_, new_n1596_,
    new_n1597_, new_n1598_, new_n1599_, new_n1600_, new_n1601_, new_n1602_,
    new_n1603_, new_n1604_, new_n1605_, new_n1606_, new_n1607_, new_n1608_,
    new_n1609_, new_n1610_, new_n1611_, new_n1612_, new_n1613_, new_n1614_,
    new_n1615_, new_n1616_, new_n1617_, new_n1618_, new_n1619_, new_n1620_,
    new_n1621_, new_n1622_, new_n1623_, new_n1624_, new_n1625_, new_n1626_,
    new_n1627_, new_n1628_, new_n1629_, new_n1630_, new_n1631_, new_n1632_,
    new_n1633_, new_n1634_, new_n1635_, new_n1636_, new_n1637_, new_n1638_,
    new_n1639_, new_n1640_, new_n1641_, new_n1642_, new_n1643_, new_n1644_,
    new_n1645_, new_n1646_, new_n1647_, new_n1648_, new_n1649_, new_n1650_,
    new_n1651_, new_n1652_, new_n1653_, new_n1654_, new_n1655_, new_n1656_,
    new_n1657_, new_n1658_, new_n1659_, new_n1660_, new_n1661_, new_n1662_,
    new_n1663_, new_n1664_, new_n1665_, new_n1666_, new_n1667_, new_n1668_,
    new_n1669_, new_n1670_, new_n1671_, new_n1672_, new_n1673_, new_n1674_,
    new_n1675_, new_n1676_, new_n1677_, new_n1678_, new_n1679_, new_n1680_,
    new_n1681_, new_n1682_, new_n1683_, new_n1684_, new_n1685_, new_n1686_,
    new_n1687_, new_n1688_, new_n1689_, new_n1690_, new_n1691_, new_n1692_,
    new_n1693_, new_n1694_, new_n1695_, new_n1696_, new_n1697_, new_n1698_,
    new_n1699_, new_n1700_, new_n1701_, new_n1702_, new_n1703_, new_n1704_,
    new_n1705_, new_n1706_, new_n1707_, new_n1708_, new_n1709_, new_n1710_,
    new_n1711_, new_n1712_, new_n1713_, new_n1714_, new_n1715_, new_n1716_,
    new_n1717_, new_n1718_, new_n1719_, new_n1720_, new_n1721_, new_n1722_,
    new_n1723_, new_n1724_, new_n1725_, new_n1726_, new_n1727_, new_n1728_,
    new_n1729_, new_n1730_, new_n1731_, new_n1732_, new_n1733_, new_n1734_,
    new_n1735_, new_n1736_, new_n1737_, new_n1738_, new_n1739_, new_n1740_,
    new_n1741_, new_n1742_, new_n1743_, new_n1744_, new_n1745_, new_n1746_,
    new_n1747_, new_n1748_, new_n1749_, new_n1750_, new_n1751_, new_n1752_,
    new_n1753_, new_n1754_, new_n1755_, new_n1756_, new_n1757_, new_n1758_,
    new_n1759_, new_n1760_, new_n1761_, new_n1762_, new_n1763_, new_n1764_,
    new_n1765_, new_n1766_, new_n1767_, new_n1768_, new_n1769_, new_n1770_,
    new_n1771_, new_n1772_, new_n1773_, new_n1774_, new_n1775_, new_n1776_,
    new_n1777_, new_n1778_, new_n1779_, new_n1780_, new_n1781_, new_n1782_,
    new_n1783_, new_n1784_, new_n1785_, new_n1786_, new_n1787_, new_n1788_,
    new_n1789_, new_n1790_, new_n1791_, new_n1792_, new_n1793_, new_n1794_,
    new_n1795_, new_n1796_, new_n1797_, new_n1798_, new_n1799_, new_n1800_,
    new_n1801_, new_n1802_, new_n1803_, new_n1804_, new_n1805_, new_n1806_,
    new_n1807_, new_n1808_, new_n1809_, new_n1810_, new_n1811_, new_n1812_,
    new_n1813_, new_n1814_, new_n1815_, new_n1816_, new_n1817_, new_n1818_,
    new_n1819_, new_n1820_, new_n1821_, new_n1822_, new_n1823_, new_n1824_,
    new_n1825_, new_n1826_, new_n1827_, new_n1828_, new_n1829_, new_n1830_,
    new_n1831_, new_n1832_, new_n1833_, new_n1834_, new_n1835_, new_n1836_,
    new_n1837_, new_n1838_, new_n1839_, new_n1840_, new_n1841_, new_n1842_,
    new_n1843_, new_n1844_, new_n1845_, new_n1846_, new_n1847_, new_n1848_,
    new_n1849_, new_n1850_, new_n1851_, new_n1852_, new_n1853_, new_n1854_,
    new_n1855_, new_n1856_, new_n1857_, new_n1858_, new_n1859_, new_n1860_,
    new_n1861_, new_n1862_, new_n1863_, new_n1864_, new_n1865_, new_n1866_,
    new_n1867_, new_n1868_, new_n1869_, new_n1870_, new_n1871_, new_n1872_,
    new_n1873_, new_n1874_, new_n1875_, new_n1876_, new_n1877_, new_n1878_,
    new_n1879_, new_n1880_, new_n1881_, new_n1882_, new_n1883_, new_n1884_,
    new_n1885_, new_n1886_, new_n1887_, new_n1888_, new_n1889_, new_n1890_,
    new_n1891_, new_n1892_, new_n1893_, new_n1894_, new_n1895_, new_n1896_,
    new_n1897_, new_n1898_, new_n1899_, new_n1900_, new_n1901_, new_n1902_,
    new_n1903_, new_n1904_, new_n1905_, new_n1906_, new_n1907_, new_n1908_,
    new_n1909_, new_n1910_, new_n1911_, new_n1912_, new_n1913_, new_n1914_,
    new_n1915_, new_n1916_, new_n1917_, new_n1918_, new_n1919_, new_n1920_,
    new_n1921_, new_n1922_, new_n1923_, new_n1924_, new_n1925_, new_n1926_,
    new_n1927_, new_n1928_, new_n1929_, new_n1930_, new_n1931_, new_n1932_,
    new_n1933_, new_n1934_, new_n1935_, new_n1936_, new_n1937_, new_n1938_,
    new_n1939_, new_n1940_, new_n1941_, new_n1942_, new_n1943_, new_n1944_,
    new_n1945_, new_n1946_, new_n1947_, new_n1948_, new_n1949_, new_n1950_,
    new_n1951_, new_n1952_, new_n1953_, new_n1954_, new_n1955_, new_n1956_,
    new_n1957_, new_n1958_, new_n1959_, new_n1960_, new_n1961_, new_n1962_,
    new_n1963_, new_n1964_, new_n1965_, new_n1966_, new_n1967_, new_n1968_,
    new_n1969_, new_n1970_, new_n1971_, new_n1972_, new_n1973_, new_n1974_,
    new_n1975_, new_n1976_, new_n1977_, new_n1978_, new_n1979_, new_n1980_,
    new_n1981_, new_n1982_, new_n1983_, new_n1984_, new_n1985_, new_n1986_,
    new_n1987_, new_n1988_, new_n1989_, new_n1990_, new_n1991_, new_n1992_,
    new_n1993_, new_n1994_, new_n1995_, new_n1996_, new_n1997_, new_n1998_,
    new_n1999_, new_n2000_, new_n2001_, new_n2002_, new_n2003_, new_n2004_,
    new_n2005_, new_n2006_, new_n2007_, new_n2008_, new_n2009_, new_n2010_,
    new_n2011_, new_n2012_, new_n2013_, new_n2014_, new_n2015_, new_n2016_,
    new_n2017_, new_n2018_, new_n2019_, new_n2020_, new_n2021_, new_n2022_,
    new_n2023_, new_n2024_, new_n2025_, new_n2026_, new_n2027_, new_n2028_,
    new_n2029_, new_n2030_, new_n2031_, new_n2032_, new_n2033_, new_n2034_,
    new_n2035_, new_n2036_, new_n2037_, new_n2038_, new_n2039_, new_n2040_,
    new_n2041_, new_n2042_, new_n2043_, new_n2044_, new_n2045_, new_n2046_,
    new_n2047_, new_n2048_, new_n2049_, new_n2050_, new_n2051_, new_n2052_,
    new_n2053_, new_n2054_, new_n2055_, new_n2056_, new_n2057_, new_n2058_,
    new_n2059_, new_n2060_, new_n2061_, new_n2062_, new_n2063_, new_n2064_,
    new_n2065_, new_n2066_, new_n2067_, new_n2068_, new_n2069_, new_n2070_,
    new_n2071_, new_n2072_, new_n2073_, new_n2074_, new_n2075_, new_n2076_,
    new_n2077_, new_n2078_, new_n2079_, new_n2080_, new_n2081_, new_n2082_,
    new_n2083_, new_n2084_, new_n2085_, new_n2086_, new_n2087_, new_n2088_,
    new_n2089_, new_n2090_, new_n2091_, new_n2092_, new_n2093_, new_n2094_,
    new_n2095_, new_n2096_, new_n2097_, new_n2098_, new_n2099_, new_n2100_,
    new_n2101_, new_n2102_, new_n2103_, new_n2104_, new_n2105_, new_n2106_,
    new_n2107_, new_n2108_, new_n2109_, new_n2110_, new_n2111_, new_n2112_,
    new_n2113_, new_n2114_, new_n2115_, new_n2116_, new_n2117_, new_n2118_,
    new_n2119_, new_n2120_, new_n2121_, new_n2122_, new_n2123_, new_n2124_,
    new_n2125_, new_n2126_, new_n2127_, new_n2128_, new_n2129_, new_n2130_,
    new_n2131_, new_n2132_, new_n2133_, new_n2134_, new_n2135_, new_n2136_,
    new_n2137_, new_n2138_, new_n2139_, new_n2140_, new_n2141_, new_n2142_,
    new_n2143_, new_n2144_, new_n2145_, new_n2146_, new_n2147_, new_n2148_,
    new_n2149_, new_n2150_, new_n2151_, new_n2152_, new_n2153_, new_n2154_,
    new_n2155_, new_n2156_, new_n2157_, new_n2158_, new_n2159_, new_n2160_,
    new_n2161_, new_n2162_, new_n2163_, new_n2164_, new_n2165_, new_n2166_,
    new_n2167_, new_n2168_, new_n2169_, new_n2170_, new_n2171_, new_n2172_,
    new_n2173_, new_n2174_, new_n2175_, new_n2176_, new_n2177_, new_n2178_,
    new_n2179_, new_n2180_, new_n2181_, new_n2182_, new_n2183_, new_n2184_,
    new_n2185_, new_n2186_, new_n2187_, new_n2188_, new_n2189_, new_n2190_,
    new_n2191_, new_n2192_, new_n2193_, new_n2194_, new_n2195_, new_n2196_,
    new_n2197_, new_n2198_, new_n2199_, new_n2200_, new_n2201_, new_n2202_,
    new_n2203_, new_n2204_, new_n2205_, new_n2206_, new_n2207_, new_n2208_,
    new_n2209_, new_n2210_, new_n2211_, new_n2212_, new_n2213_, new_n2214_,
    new_n2215_, new_n2216_, new_n2217_, new_n2218_, new_n2219_, new_n2220_,
    new_n2221_, new_n2222_, new_n2223_, new_n2224_, new_n2225_, new_n2226_,
    new_n2227_, new_n2228_, new_n2229_, new_n2230_, new_n2231_, new_n2232_,
    new_n2233_, new_n2234_, new_n2235_, new_n2236_, new_n2237_, new_n2238_,
    new_n2239_, new_n2240_, new_n2241_, new_n2242_, new_n2243_, new_n2244_,
    new_n2245_, new_n2246_, new_n2247_, new_n2248_, new_n2249_, new_n2250_,
    new_n2251_, new_n2252_, new_n2253_, new_n2254_, new_n2255_, new_n2256_,
    new_n2257_, new_n2258_, new_n2259_, new_n2260_, new_n2261_, new_n2262_,
    new_n2263_, new_n2264_, new_n2265_, new_n2266_, new_n2267_, new_n2268_,
    new_n2269_, new_n2270_, new_n2271_, new_n2272_, new_n2273_, new_n2274_,
    new_n2275_, new_n2276_, new_n2277_, new_n2278_, new_n2279_, new_n2280_,
    new_n2281_, new_n2282_, new_n2283_, new_n2284_, new_n2285_, new_n2286_,
    new_n2287_, new_n2288_, new_n2289_, new_n2290_, new_n2291_, new_n2292_,
    new_n2293_, new_n2294_, new_n2295_, new_n2296_, new_n2297_, new_n2298_,
    new_n2299_, new_n2300_, new_n2301_, new_n2302_, new_n2303_, new_n2304_,
    new_n2305_, new_n2306_, new_n2307_, new_n2308_, new_n2309_, new_n2310_,
    new_n2311_, new_n2312_, new_n2313_, new_n2314_, new_n2315_, new_n2316_,
    new_n2317_, new_n2318_, new_n2319_, new_n2320_, new_n2321_, new_n2322_,
    new_n2323_, new_n2324_, new_n2325_, new_n2326_, new_n2327_, new_n2328_,
    new_n2329_, new_n2330_, new_n2331_, new_n2332_, new_n2333_, new_n2334_,
    new_n2335_, new_n2336_, new_n2337_, new_n2338_, new_n2339_, new_n2340_,
    new_n2341_, new_n2342_, new_n2343_, new_n2344_, new_n2345_, new_n2346_,
    new_n2347_, new_n2348_, new_n2349_, new_n2350_, new_n2351_, new_n2352_,
    new_n2353_, new_n2354_, new_n2355_, new_n2356_, new_n2357_, new_n2358_,
    new_n2359_, new_n2360_, new_n2361_, new_n2362_, new_n2363_, new_n2364_,
    new_n2365_, new_n2366_, new_n2367_, new_n2368_, new_n2369_, new_n2370_,
    new_n2371_, new_n2372_, new_n2373_, new_n2374_, new_n2375_, new_n2376_,
    new_n2377_, new_n2378_, new_n2379_, new_n2380_, new_n2381_, new_n2382_,
    new_n2383_, new_n2384_, new_n2385_, new_n2386_, new_n2387_, new_n2388_,
    new_n2389_, new_n2390_, new_n2391_, new_n2392_, new_n2393_, new_n2394_,
    new_n2395_, new_n2396_, new_n2397_, new_n2398_, new_n2399_, new_n2400_,
    new_n2401_, new_n2402_, new_n2403_, new_n2404_, new_n2405_, new_n2406_,
    new_n2407_, new_n2408_, new_n2409_, new_n2410_, new_n2411_, new_n2412_,
    new_n2413_, new_n2414_, new_n2415_, new_n2416_, new_n2417_, new_n2418_,
    new_n2419_, new_n2420_, new_n2421_, new_n2422_, new_n2423_, new_n2424_,
    new_n2425_, new_n2426_, new_n2427_, new_n2428_, new_n2429_, new_n2430_,
    new_n2431_, new_n2432_, new_n2433_, new_n2434_, new_n2435_, new_n2436_,
    new_n2437_, new_n2438_, new_n2439_, new_n2440_, new_n2441_, new_n2442_,
    new_n2443_, new_n2444_, new_n2445_, new_n2446_, new_n2447_, new_n2448_,
    new_n2449_, new_n2450_, new_n2451_, new_n2452_, new_n2453_, new_n2454_,
    new_n2455_, new_n2456_, new_n2457_, new_n2458_, new_n2459_, new_n2460_,
    new_n2461_, new_n2462_, new_n2463_, new_n2464_, new_n2465_, new_n2466_,
    new_n2467_, new_n2468_, new_n2469_, new_n2470_, new_n2471_, new_n2472_,
    new_n2473_, new_n2474_, new_n2475_, new_n2476_, new_n2477_, new_n2478_,
    new_n2479_, new_n2480_, new_n2481_, new_n2482_, new_n2483_, new_n2484_,
    new_n2485_, new_n2486_, new_n2487_, new_n2488_, new_n2489_, new_n2490_,
    new_n2491_, new_n2492_, new_n2493_, new_n2494_, new_n2495_, new_n2496_,
    new_n2497_, new_n2498_, new_n2499_, new_n2500_, new_n2501_, new_n2502_,
    new_n2503_, new_n2504_, new_n2505_, new_n2506_, new_n2507_, new_n2508_,
    new_n2509_, new_n2510_, new_n2511_, new_n2512_, new_n2513_, new_n2514_,
    new_n2515_, new_n2516_, new_n2517_, new_n2518_, new_n2519_, new_n2520_,
    new_n2521_, new_n2522_, new_n2523_, new_n2524_, new_n2525_, new_n2526_,
    new_n2527_, new_n2528_, new_n2529_, new_n2530_, new_n2531_, new_n2532_,
    new_n2533_, new_n2534_, new_n2535_, new_n2536_, new_n2537_, new_n2538_,
    new_n2539_, new_n2540_, new_n2541_, new_n2542_, new_n2543_, new_n2544_,
    new_n2545_, new_n2546_, new_n2547_, new_n2548_, new_n2549_, new_n2550_,
    new_n2551_, new_n2552_, new_n2553_, new_n2554_, new_n2555_, new_n2556_,
    new_n2557_, new_n2558_, new_n2559_, new_n2560_, new_n2561_, new_n2562_,
    new_n2563_, new_n2564_, new_n2565_, new_n2566_, new_n2567_, new_n2568_,
    new_n2569_, new_n2570_, new_n2571_, new_n2572_, new_n2573_, new_n2574_,
    new_n2575_, new_n2576_, new_n2577_, new_n2578_, new_n2579_, new_n2580_,
    new_n2581_, new_n2582_, new_n2583_, new_n2584_, new_n2585_, new_n2586_,
    new_n2587_, new_n2588_, new_n2589_, new_n2590_, new_n2591_, new_n2592_,
    new_n2593_, new_n2594_, new_n2595_, new_n2596_, new_n2597_, new_n2598_,
    new_n2599_, new_n2600_, new_n2601_, new_n2602_, new_n2603_, new_n2604_,
    new_n2605_, new_n2606_, new_n2607_, new_n2608_, new_n2609_, new_n2610_,
    new_n2611_, new_n2612_, new_n2613_, new_n2614_, new_n2615_, new_n2616_,
    new_n2617_, new_n2618_, new_n2619_, new_n2620_, new_n2621_, new_n2622_,
    new_n2623_, new_n2624_, new_n2625_, new_n2626_, new_n2627_, new_n2628_,
    new_n2629_, new_n2630_, new_n2631_, new_n2632_, new_n2633_, new_n2634_,
    new_n2635_, new_n2636_, new_n2637_, new_n2638_, new_n2639_, new_n2640_,
    new_n2641_, new_n2642_, new_n2643_, new_n2644_, new_n2645_, new_n2646_,
    new_n2647_, new_n2648_, new_n2649_, new_n2650_, new_n2651_, new_n2652_,
    new_n2653_, new_n2654_, new_n2655_, new_n2656_, new_n2657_, new_n2658_,
    new_n2659_, new_n2660_, new_n2661_, new_n2662_, new_n2663_, new_n2664_,
    new_n2665_, new_n2666_, new_n2667_, new_n2668_, new_n2669_, new_n2670_,
    new_n2671_, new_n2672_, new_n2673_, new_n2674_, new_n2675_, new_n2676_,
    new_n2677_, new_n2678_, new_n2679_, new_n2680_, new_n2681_, new_n2682_,
    new_n2683_, new_n2684_, new_n2685_, new_n2686_, new_n2687_, new_n2688_,
    new_n2689_, new_n2690_, new_n2691_, new_n2692_, new_n2693_, new_n2694_,
    new_n2695_, new_n2696_, new_n2697_, new_n2698_, new_n2699_, new_n2700_,
    new_n2701_, new_n2702_, new_n2703_, new_n2704_, new_n2705_, new_n2706_,
    new_n2707_, new_n2708_, new_n2709_, new_n2710_, new_n2711_, new_n2712_,
    new_n2713_, new_n2714_, new_n2715_, new_n2716_, new_n2717_, new_n2718_,
    new_n2719_, new_n2720_, new_n2721_, new_n2722_, new_n2723_, new_n2724_,
    new_n2725_, new_n2726_, new_n2727_, new_n2728_, new_n2729_, new_n2730_,
    new_n2731_, new_n2732_, new_n2733_, new_n2734_, new_n2735_, new_n2736_,
    new_n2737_, new_n2738_, new_n2739_, new_n2740_, new_n2741_, new_n2742_,
    new_n2743_, new_n2744_, new_n2745_, new_n2746_, new_n2747_, new_n2748_,
    new_n2749_, new_n2750_, new_n2751_, new_n2752_, new_n2753_, new_n2754_,
    new_n2755_, new_n2756_, new_n2757_, new_n2758_, new_n2759_, new_n2760_,
    new_n2761_, new_n2762_, new_n2763_, new_n2764_, new_n2765_, new_n2766_,
    new_n2767_, new_n2768_, new_n2769_, new_n2770_, new_n2771_, new_n2772_,
    new_n2773_, new_n2774_, new_n2775_, new_n2776_, new_n2777_, new_n2778_,
    new_n2779_, new_n2780_, new_n2781_, new_n2782_, new_n2783_, new_n2784_,
    new_n2785_, new_n2786_, new_n2787_, new_n2788_, new_n2789_, new_n2790_,
    new_n2791_, new_n2792_, new_n2793_, new_n2794_, new_n2795_, new_n2796_,
    new_n2797_, new_n2798_, new_n2799_, new_n2800_, new_n2801_, new_n2802_,
    new_n2803_, new_n2804_, new_n2805_, new_n2806_, new_n2807_, new_n2808_,
    new_n2809_, new_n2810_, new_n2811_, new_n2812_, new_n2813_, new_n2814_,
    new_n2815_, new_n2816_, new_n2817_, new_n2818_, new_n2819_, new_n2820_,
    new_n2821_, new_n2822_, new_n2823_, new_n2824_, new_n2825_, new_n2826_,
    new_n2827_, new_n2828_, new_n2829_, new_n2830_, new_n2831_, new_n2832_,
    new_n2833_, new_n2834_, new_n2835_, new_n2836_, new_n2837_, new_n2838_,
    new_n2839_, new_n2840_, new_n2841_, new_n2842_, new_n2843_, new_n2844_,
    new_n2845_, new_n2846_, new_n2847_, new_n2848_, new_n2849_, new_n2850_,
    new_n2851_, new_n2852_, new_n2853_, new_n2854_, new_n2855_, new_n2856_,
    new_n2857_, new_n2858_, new_n2859_, new_n2860_, new_n2861_, new_n2862_,
    new_n2863_, new_n2864_, new_n2865_, new_n2866_, new_n2867_, new_n2868_,
    new_n2869_, new_n2870_, new_n2871_, new_n2872_, new_n2873_, new_n2874_,
    new_n2875_, new_n2876_, new_n2877_, new_n2878_, new_n2879_, new_n2880_,
    new_n2881_, new_n2882_, new_n2883_, new_n2884_, new_n2885_, new_n2886_,
    new_n2887_, new_n2888_, new_n2889_, new_n2890_, new_n2891_, new_n2892_,
    new_n2893_, new_n2894_, new_n2895_, new_n2896_, new_n2897_, new_n2898_,
    new_n2899_, new_n2900_, new_n2901_, new_n2902_, new_n2903_, new_n2904_,
    new_n2905_, new_n2906_, new_n2907_, new_n2908_, new_n2909_, new_n2910_,
    new_n2911_, new_n2912_, new_n2913_, new_n2914_, new_n2915_, new_n2916_,
    new_n2917_, new_n2918_, new_n2919_, new_n2920_, new_n2921_, new_n2922_,
    new_n2923_, new_n2924_, new_n2925_, new_n2926_, new_n2927_, new_n2928_,
    new_n2929_, new_n2930_, new_n2931_, new_n2932_, new_n2933_, new_n2934_,
    new_n2935_, new_n2936_, new_n2937_, new_n2938_, new_n2939_, new_n2940_,
    new_n2941_, new_n2942_, new_n2943_, new_n2944_, new_n2945_, new_n2946_,
    new_n2947_, new_n2948_, new_n2949_, new_n2950_, new_n2951_, new_n2952_,
    new_n2953_, new_n2954_, new_n2955_, new_n2956_, new_n2957_, new_n2958_,
    new_n2959_, new_n2960_, new_n2961_, new_n2962_, new_n2963_, new_n2964_,
    new_n2965_, new_n2966_, new_n2967_, new_n2968_, new_n2969_, new_n2970_,
    new_n2971_, new_n2972_, new_n2973_, new_n2974_, new_n2975_, new_n2976_,
    new_n2977_, new_n2978_, new_n2979_, new_n2980_, new_n2981_, new_n2982_,
    new_n2983_, new_n2984_, new_n2985_, new_n2986_, new_n2987_, new_n2988_,
    new_n2989_, new_n2990_, new_n2991_, new_n2992_, new_n2993_, new_n2994_,
    new_n2995_, new_n2996_, new_n2997_, new_n2998_, new_n2999_, new_n3000_,
    new_n3001_, new_n3002_, new_n3003_, new_n3004_, new_n3005_, new_n3006_,
    new_n3007_, new_n3008_, new_n3009_, new_n3010_, new_n3011_, new_n3012_,
    new_n3013_, new_n3014_, new_n3015_, new_n3016_, new_n3017_, new_n3018_,
    new_n3019_, new_n3020_, new_n3021_, new_n3022_, new_n3023_, new_n3024_,
    new_n3025_, new_n3026_, new_n3027_, new_n3028_, new_n3029_, new_n3030_,
    new_n3031_, new_n3032_, new_n3033_, new_n3034_, new_n3035_, new_n3036_,
    new_n3037_, new_n3038_, new_n3039_, new_n3040_, new_n3041_, new_n3042_,
    new_n3043_, new_n3044_, new_n3045_, new_n3046_, new_n3047_, new_n3048_,
    new_n3049_, new_n3050_, new_n3051_, new_n3052_, new_n3053_, new_n3054_,
    new_n3055_, new_n3056_, new_n3057_, new_n3058_, new_n3059_, new_n3060_,
    new_n3061_, new_n3062_, new_n3063_, new_n3064_, new_n3065_, new_n3066_,
    new_n3067_, new_n3068_, new_n3069_, new_n3070_, new_n3071_, new_n3072_,
    new_n3073_, new_n3074_, new_n3075_, new_n3076_, new_n3077_, new_n3078_,
    new_n3079_, new_n3080_, new_n3081_, new_n3082_, new_n3083_, new_n3084_,
    new_n3085_, new_n3086_, new_n3087_, new_n3088_, new_n3089_, new_n3090_,
    new_n3091_, new_n3092_, new_n3093_, new_n3094_, new_n3095_, new_n3096_,
    new_n3097_, new_n3098_, new_n3099_, new_n3100_, new_n3101_, new_n3102_,
    new_n3103_, new_n3104_, new_n3105_, new_n3106_, new_n3107_, new_n3108_,
    new_n3109_, new_n3110_, new_n3111_, new_n3112_, new_n3113_, new_n3114_,
    new_n3115_, new_n3116_, new_n3117_, new_n3118_, new_n3119_, new_n3120_,
    new_n3121_, new_n3122_, new_n3123_, new_n3124_, new_n3125_, new_n3126_,
    new_n3127_, new_n3128_, new_n3129_, new_n3130_, new_n3131_, new_n3132_,
    new_n3133_, new_n3134_, new_n3135_, new_n3136_, new_n3137_, new_n3138_,
    new_n3139_, new_n3140_, new_n3141_, new_n3142_, new_n3143_, new_n3144_,
    new_n3145_, new_n3146_, new_n3147_, new_n3148_, new_n3149_, new_n3150_,
    new_n3151_, new_n3152_, new_n3153_, new_n3154_, new_n3155_, new_n3156_,
    new_n3157_, new_n3158_, new_n3159_, new_n3160_, new_n3161_, new_n3162_,
    new_n3163_, new_n3164_, new_n3165_, new_n3166_, new_n3167_, new_n3168_,
    new_n3169_, new_n3171_, new_n3172_, new_n3174_, new_n3176_, new_n3178_,
    new_n3179_, new_n3181_, new_n3183_, new_n3185_, new_n3187_, new_n3189_,
    new_n3191_, new_n3193_, new_n3195_, new_n3197_, new_n3199_, new_n3201_,
    new_n3203_, new_n3205_, new_n3207_, new_n3209_, new_n3211_, new_n3212_,
    new_n3214_, new_n3216_, new_n3217_, new_n3219_, new_n3221_, new_n3222_,
    new_n3224_, new_n3226_, new_n3228_, new_n3230_, new_n3232_, new_n3234_,
    new_n3236_, new_n3238_, new_n3240_, new_n3242_, new_n3244_, new_n3246_,
    new_n3248_, new_n3250_, new_n3252_, new_n3254_, new_n3256_, new_n3258_,
    new_n3259_, new_n3261_, new_n3263_, new_n3265_, new_n3267_, new_n3269_,
    new_n3271_, new_n3273_, new_n3275_, new_n3277_, new_n3279_, new_n3281_,
    new_n3283_, new_n3285_, new_n3287_, new_n3289_, new_n3291_, new_n3292_,
    new_n3294_, new_n3296_, new_n3298_, new_n3300_, new_n3302_, new_n3304_,
    new_n3306_, new_n3308_, new_n3310_, new_n3312_, new_n3314_, new_n3316_,
    new_n3318_, new_n3320_, new_n3322_, new_n3324_, new_n3326_, new_n3328_,
    new_n3330_, new_n3332_, new_n3334_, new_n3336_, new_n3338_, new_n3340_,
    new_n3342_, new_n3344_, new_n3346_, new_n3348_, new_n3350_, new_n3352_,
    new_n3354_, new_n3356_, new_n3358_, new_n3360_, new_n3362_, new_n3364_,
    new_n3366_, new_n3368_, new_n3370_, new_n3372_, new_n3374_, new_n3376_,
    new_n3378_, new_n3380_, new_n3382_, new_n3384_, new_n3386_, new_n3388_,
    new_n3390_, new_n3392_, new_n3394_, new_n3396_, new_n3398_, new_n3400_,
    new_n3402_, new_n3404_, new_n3406_, new_n3408_, new_n3410_, new_n3412_,
    new_n3414_, new_n3416_, new_n3418_, new_n3420_, new_n3422_, new_n3424_,
    new_n3426_, new_n3428_, new_n3430_, new_n3432_, new_n3434_;
  INVX1    g0000(.A(\in1[0] ), .Y(new_n643_));
  INVX1    g0001(.A(\in0[31] ), .Y(new_n644_));
  AND2X1   g0002(.A(\in1[31] ), .B(new_n644_), .Y(new_n645_));
  INVX1    g0003(.A(\in0[30] ), .Y(new_n646_));
  AND2X1   g0004(.A(\in1[30] ), .B(new_n646_), .Y(new_n647_));
  INVX1    g0005(.A(new_n647_), .Y(new_n648_));
  INVX1    g0006(.A(\in0[29] ), .Y(new_n649_));
  AND2X1   g0007(.A(\in1[29] ), .B(new_n649_), .Y(new_n650_));
  INVX1    g0008(.A(\in0[28] ), .Y(new_n651_));
  AND2X1   g0009(.A(\in1[28] ), .B(new_n651_), .Y(new_n652_));
  INVX1    g0010(.A(new_n652_), .Y(new_n653_));
  INVX1    g0011(.A(\in0[27] ), .Y(new_n654_));
  AND2X1   g0012(.A(\in1[27] ), .B(new_n654_), .Y(new_n655_));
  INVX1    g0013(.A(\in0[26] ), .Y(new_n656_));
  AND2X1   g0014(.A(\in1[26] ), .B(new_n656_), .Y(new_n657_));
  INVX1    g0015(.A(new_n657_), .Y(new_n658_));
  INVX1    g0016(.A(\in0[24] ), .Y(new_n659_));
  INVX1    g0017(.A(\in0[23] ), .Y(new_n660_));
  AND2X1   g0018(.A(\in1[23] ), .B(new_n660_), .Y(new_n661_));
  INVX1    g0019(.A(new_n661_), .Y(new_n662_));
  INVX1    g0020(.A(\in0[22] ), .Y(new_n663_));
  AND2X1   g0021(.A(\in1[22] ), .B(new_n663_), .Y(new_n664_));
  INVX1    g0022(.A(\in0[21] ), .Y(new_n665_));
  AND2X1   g0023(.A(\in1[21] ), .B(new_n665_), .Y(new_n666_));
  INVX1    g0024(.A(new_n666_), .Y(new_n667_));
  INVX1    g0025(.A(\in0[20] ), .Y(new_n668_));
  AND2X1   g0026(.A(\in1[20] ), .B(new_n668_), .Y(new_n669_));
  INVX1    g0027(.A(\in0[19] ), .Y(new_n670_));
  AND2X1   g0028(.A(\in1[19] ), .B(new_n670_), .Y(new_n671_));
  INVX1    g0029(.A(new_n671_), .Y(new_n672_));
  INVX1    g0030(.A(\in0[18] ), .Y(new_n673_));
  AND2X1   g0031(.A(\in1[18] ), .B(new_n673_), .Y(new_n674_));
  INVX1    g0032(.A(\in1[17] ), .Y(new_n675_));
  INVX1    g0033(.A(\in0[17] ), .Y(new_n676_));
  INVX1    g0034(.A(\in1[16] ), .Y(new_n677_));
  INVX1    g0035(.A(\in0[15] ), .Y(new_n678_));
  AND2X1   g0036(.A(\in1[15] ), .B(new_n678_), .Y(new_n679_));
  INVX1    g0037(.A(\in0[14] ), .Y(new_n680_));
  AND2X1   g0038(.A(\in1[14] ), .B(new_n680_), .Y(new_n681_));
  INVX1    g0039(.A(new_n681_), .Y(new_n682_));
  INVX1    g0040(.A(\in0[13] ), .Y(new_n683_));
  AND2X1   g0041(.A(\in1[13] ), .B(new_n683_), .Y(new_n684_));
  INVX1    g0042(.A(\in0[12] ), .Y(new_n685_));
  AND2X1   g0043(.A(\in1[12] ), .B(new_n685_), .Y(new_n686_));
  INVX1    g0044(.A(new_n686_), .Y(new_n687_));
  INVX1    g0045(.A(\in0[11] ), .Y(new_n688_));
  AND2X1   g0046(.A(\in1[11] ), .B(new_n688_), .Y(new_n689_));
  INVX1    g0047(.A(\in0[10] ), .Y(new_n690_));
  AND2X1   g0048(.A(\in1[10] ), .B(new_n690_), .Y(new_n691_));
  INVX1    g0049(.A(new_n691_), .Y(new_n692_));
  INVX1    g0050(.A(\in0[8] ), .Y(new_n693_));
  INVX1    g0051(.A(\in0[7] ), .Y(new_n694_));
  AND2X1   g0052(.A(\in1[7] ), .B(new_n694_), .Y(new_n695_));
  INVX1    g0053(.A(new_n695_), .Y(new_n696_));
  INVX1    g0054(.A(\in0[6] ), .Y(new_n697_));
  AND2X1   g0055(.A(\in1[6] ), .B(new_n697_), .Y(new_n698_));
  INVX1    g0056(.A(\in1[5] ), .Y(new_n699_));
  INVX1    g0057(.A(\in0[5] ), .Y(new_n700_));
  INVX1    g0058(.A(\in1[4] ), .Y(new_n701_));
  INVX1    g0059(.A(\in0[3] ), .Y(new_n702_));
  AND2X1   g0060(.A(\in1[3] ), .B(new_n702_), .Y(new_n703_));
  INVX1    g0061(.A(\in1[2] ), .Y(new_n704_));
  INVX1    g0062(.A(\in0[0] ), .Y(new_n705_));
  INVX1    g0063(.A(\in0[1] ), .Y(new_n706_));
  OAI22X1  g0064(.A0(\in1[1] ), .A1(new_n706_), .B0(\in1[0] ), .B1(new_n705_), .Y(new_n707_));
  INVX1    g0065(.A(\in0[2] ), .Y(new_n708_));
  AOI22X1  g0066(.A0(\in1[2] ), .A1(new_n708_), .B0(\in1[1] ), .B1(new_n706_), .Y(new_n709_));
  AOI22X1  g0067(.A0(new_n709_), .A1(new_n707_), .B0(new_n704_), .B1(\in0[2] ), .Y(new_n710_));
  OR2X1    g0068(.A(\in1[3] ), .B(new_n702_), .Y(new_n711_));
  OAI21X1  g0069(.A0(new_n710_), .A1(new_n703_), .B0(new_n711_), .Y(new_n712_));
  OAI21X1  g0070(.A0(new_n712_), .A1(\in0[4] ), .B0(new_n701_), .Y(new_n713_));
  INVX1    g0071(.A(\in0[4] ), .Y(new_n714_));
  INVX1    g0072(.A(\in1[3] ), .Y(new_n715_));
  OR2X1    g0073(.A(new_n715_), .B(\in0[3] ), .Y(new_n716_));
  INVX1    g0074(.A(\in1[1] ), .Y(new_n717_));
  AOI22X1  g0075(.A0(new_n717_), .A1(\in0[1] ), .B0(new_n643_), .B1(\in0[0] ), .Y(new_n718_));
  OAI22X1  g0076(.A0(new_n704_), .A1(\in0[2] ), .B0(new_n717_), .B1(\in0[1] ), .Y(new_n719_));
  OAI22X1  g0077(.A0(new_n719_), .A1(new_n718_), .B0(\in1[2] ), .B1(new_n708_), .Y(new_n720_));
  AND2X1   g0078(.A(new_n715_), .B(\in0[3] ), .Y(new_n721_));
  AOI21X1  g0079(.A0(new_n720_), .A1(new_n716_), .B0(new_n721_), .Y(new_n722_));
  OR2X1    g0080(.A(new_n722_), .B(new_n714_), .Y(new_n723_));
  NAND3X1  g0081(.A(new_n723_), .B(new_n713_), .C(new_n700_), .Y(new_n724_));
  AOI21X1  g0082(.A0(new_n723_), .A1(new_n713_), .B0(new_n700_), .Y(new_n725_));
  AOI21X1  g0083(.A0(new_n724_), .A1(new_n699_), .B0(new_n725_), .Y(new_n726_));
  INVX1    g0084(.A(\in1[6] ), .Y(new_n727_));
  AND2X1   g0085(.A(new_n727_), .B(\in0[6] ), .Y(new_n728_));
  INVX1    g0086(.A(new_n728_), .Y(new_n729_));
  OAI21X1  g0087(.A0(new_n726_), .A1(new_n698_), .B0(new_n729_), .Y(new_n730_));
  INVX1    g0088(.A(\in1[7] ), .Y(new_n731_));
  AND2X1   g0089(.A(new_n731_), .B(\in0[7] ), .Y(new_n732_));
  AOI21X1  g0090(.A0(new_n730_), .A1(new_n696_), .B0(new_n732_), .Y(new_n733_));
  AOI21X1  g0091(.A0(new_n733_), .A1(new_n693_), .B0(\in1[8] ), .Y(new_n734_));
  INVX1    g0092(.A(new_n698_), .Y(new_n735_));
  AOI21X1  g0093(.A0(new_n722_), .A1(new_n714_), .B0(\in1[4] ), .Y(new_n736_));
  AND2X1   g0094(.A(new_n712_), .B(\in0[4] ), .Y(new_n737_));
  NOR3X1   g0095(.A(new_n737_), .B(new_n736_), .C(\in0[5] ), .Y(new_n738_));
  OAI21X1  g0096(.A0(new_n737_), .A1(new_n736_), .B0(\in0[5] ), .Y(new_n739_));
  OAI21X1  g0097(.A0(new_n738_), .A1(\in1[5] ), .B0(new_n739_), .Y(new_n740_));
  AOI21X1  g0098(.A0(new_n740_), .A1(new_n735_), .B0(new_n728_), .Y(new_n741_));
  INVX1    g0099(.A(new_n732_), .Y(new_n742_));
  OAI21X1  g0100(.A0(new_n741_), .A1(new_n695_), .B0(new_n742_), .Y(new_n743_));
  AND2X1   g0101(.A(new_n743_), .B(\in0[8] ), .Y(new_n744_));
  NOR3X1   g0102(.A(new_n744_), .B(new_n734_), .C(\in0[9] ), .Y(new_n745_));
  OAI21X1  g0103(.A0(new_n744_), .A1(new_n734_), .B0(\in0[9] ), .Y(new_n746_));
  OAI21X1  g0104(.A0(new_n745_), .A1(\in1[9] ), .B0(new_n746_), .Y(new_n747_));
  INVX1    g0105(.A(\in1[10] ), .Y(new_n748_));
  AND2X1   g0106(.A(new_n748_), .B(\in0[10] ), .Y(new_n749_));
  AOI21X1  g0107(.A0(new_n747_), .A1(new_n692_), .B0(new_n749_), .Y(new_n750_));
  INVX1    g0108(.A(\in1[11] ), .Y(new_n751_));
  AND2X1   g0109(.A(new_n751_), .B(\in0[11] ), .Y(new_n752_));
  INVX1    g0110(.A(new_n752_), .Y(new_n753_));
  OAI21X1  g0111(.A0(new_n750_), .A1(new_n689_), .B0(new_n753_), .Y(new_n754_));
  INVX1    g0112(.A(\in1[12] ), .Y(new_n755_));
  AND2X1   g0113(.A(new_n755_), .B(\in0[12] ), .Y(new_n756_));
  AOI21X1  g0114(.A0(new_n754_), .A1(new_n687_), .B0(new_n756_), .Y(new_n757_));
  INVX1    g0115(.A(\in1[13] ), .Y(new_n758_));
  AND2X1   g0116(.A(new_n758_), .B(\in0[13] ), .Y(new_n759_));
  INVX1    g0117(.A(new_n759_), .Y(new_n760_));
  OAI21X1  g0118(.A0(new_n757_), .A1(new_n684_), .B0(new_n760_), .Y(new_n761_));
  INVX1    g0119(.A(\in1[14] ), .Y(new_n762_));
  AND2X1   g0120(.A(new_n762_), .B(\in0[14] ), .Y(new_n763_));
  AOI21X1  g0121(.A0(new_n761_), .A1(new_n682_), .B0(new_n763_), .Y(new_n764_));
  INVX1    g0122(.A(\in1[15] ), .Y(new_n765_));
  AND2X1   g0123(.A(new_n765_), .B(\in0[15] ), .Y(new_n766_));
  INVX1    g0124(.A(new_n766_), .Y(new_n767_));
  OAI21X1  g0125(.A0(new_n764_), .A1(new_n679_), .B0(new_n767_), .Y(new_n768_));
  OAI21X1  g0126(.A0(new_n768_), .A1(\in0[16] ), .B0(new_n677_), .Y(new_n769_));
  INVX1    g0127(.A(\in0[16] ), .Y(new_n770_));
  INVX1    g0128(.A(new_n679_), .Y(new_n771_));
  INVX1    g0129(.A(new_n684_), .Y(new_n772_));
  INVX1    g0130(.A(new_n689_), .Y(new_n773_));
  INVX1    g0131(.A(\in1[9] ), .Y(new_n774_));
  INVX1    g0132(.A(\in0[9] ), .Y(new_n775_));
  INVX1    g0133(.A(\in1[8] ), .Y(new_n776_));
  OAI21X1  g0134(.A0(new_n743_), .A1(\in0[8] ), .B0(new_n776_), .Y(new_n777_));
  OR2X1    g0135(.A(new_n733_), .B(new_n693_), .Y(new_n778_));
  NAND3X1  g0136(.A(new_n778_), .B(new_n777_), .C(new_n775_), .Y(new_n779_));
  AOI21X1  g0137(.A0(new_n778_), .A1(new_n777_), .B0(new_n775_), .Y(new_n780_));
  AOI21X1  g0138(.A0(new_n779_), .A1(new_n774_), .B0(new_n780_), .Y(new_n781_));
  INVX1    g0139(.A(new_n749_), .Y(new_n782_));
  OAI21X1  g0140(.A0(new_n781_), .A1(new_n691_), .B0(new_n782_), .Y(new_n783_));
  AOI21X1  g0141(.A0(new_n783_), .A1(new_n773_), .B0(new_n752_), .Y(new_n784_));
  INVX1    g0142(.A(new_n756_), .Y(new_n785_));
  OAI21X1  g0143(.A0(new_n784_), .A1(new_n686_), .B0(new_n785_), .Y(new_n786_));
  AOI21X1  g0144(.A0(new_n786_), .A1(new_n772_), .B0(new_n759_), .Y(new_n787_));
  INVX1    g0145(.A(new_n763_), .Y(new_n788_));
  OAI21X1  g0146(.A0(new_n787_), .A1(new_n681_), .B0(new_n788_), .Y(new_n789_));
  AOI21X1  g0147(.A0(new_n789_), .A1(new_n771_), .B0(new_n766_), .Y(new_n790_));
  OR2X1    g0148(.A(new_n790_), .B(new_n770_), .Y(new_n791_));
  NAND3X1  g0149(.A(new_n791_), .B(new_n769_), .C(new_n676_), .Y(new_n792_));
  AOI21X1  g0150(.A0(new_n791_), .A1(new_n769_), .B0(new_n676_), .Y(new_n793_));
  AOI21X1  g0151(.A0(new_n792_), .A1(new_n675_), .B0(new_n793_), .Y(new_n794_));
  INVX1    g0152(.A(\in1[18] ), .Y(new_n795_));
  AND2X1   g0153(.A(new_n795_), .B(\in0[18] ), .Y(new_n796_));
  INVX1    g0154(.A(new_n796_), .Y(new_n797_));
  OAI21X1  g0155(.A0(new_n794_), .A1(new_n674_), .B0(new_n797_), .Y(new_n798_));
  INVX1    g0156(.A(\in1[19] ), .Y(new_n799_));
  AND2X1   g0157(.A(new_n799_), .B(\in0[19] ), .Y(new_n800_));
  AOI21X1  g0158(.A0(new_n798_), .A1(new_n672_), .B0(new_n800_), .Y(new_n801_));
  INVX1    g0159(.A(\in1[20] ), .Y(new_n802_));
  AND2X1   g0160(.A(new_n802_), .B(\in0[20] ), .Y(new_n803_));
  INVX1    g0161(.A(new_n803_), .Y(new_n804_));
  OAI21X1  g0162(.A0(new_n801_), .A1(new_n669_), .B0(new_n804_), .Y(new_n805_));
  INVX1    g0163(.A(\in1[21] ), .Y(new_n806_));
  AND2X1   g0164(.A(new_n806_), .B(\in0[21] ), .Y(new_n807_));
  AOI21X1  g0165(.A0(new_n805_), .A1(new_n667_), .B0(new_n807_), .Y(new_n808_));
  INVX1    g0166(.A(\in1[22] ), .Y(new_n809_));
  AND2X1   g0167(.A(new_n809_), .B(\in0[22] ), .Y(new_n810_));
  INVX1    g0168(.A(new_n810_), .Y(new_n811_));
  OAI21X1  g0169(.A0(new_n808_), .A1(new_n664_), .B0(new_n811_), .Y(new_n812_));
  INVX1    g0170(.A(\in1[23] ), .Y(new_n813_));
  AND2X1   g0171(.A(new_n813_), .B(\in0[23] ), .Y(new_n814_));
  AOI21X1  g0172(.A0(new_n812_), .A1(new_n662_), .B0(new_n814_), .Y(new_n815_));
  AOI21X1  g0173(.A0(new_n815_), .A1(new_n659_), .B0(\in1[24] ), .Y(new_n816_));
  INVX1    g0174(.A(new_n664_), .Y(new_n817_));
  INVX1    g0175(.A(new_n669_), .Y(new_n818_));
  INVX1    g0176(.A(new_n674_), .Y(new_n819_));
  AOI21X1  g0177(.A0(new_n790_), .A1(new_n770_), .B0(\in1[16] ), .Y(new_n820_));
  AND2X1   g0178(.A(new_n768_), .B(\in0[16] ), .Y(new_n821_));
  NOR3X1   g0179(.A(new_n821_), .B(new_n820_), .C(\in0[17] ), .Y(new_n822_));
  OAI21X1  g0180(.A0(new_n821_), .A1(new_n820_), .B0(\in0[17] ), .Y(new_n823_));
  OAI21X1  g0181(.A0(new_n822_), .A1(\in1[17] ), .B0(new_n823_), .Y(new_n824_));
  AOI21X1  g0182(.A0(new_n824_), .A1(new_n819_), .B0(new_n796_), .Y(new_n825_));
  INVX1    g0183(.A(new_n800_), .Y(new_n826_));
  OAI21X1  g0184(.A0(new_n825_), .A1(new_n671_), .B0(new_n826_), .Y(new_n827_));
  AOI21X1  g0185(.A0(new_n827_), .A1(new_n818_), .B0(new_n803_), .Y(new_n828_));
  INVX1    g0186(.A(new_n807_), .Y(new_n829_));
  OAI21X1  g0187(.A0(new_n828_), .A1(new_n666_), .B0(new_n829_), .Y(new_n830_));
  AOI21X1  g0188(.A0(new_n830_), .A1(new_n817_), .B0(new_n810_), .Y(new_n831_));
  INVX1    g0189(.A(new_n814_), .Y(new_n832_));
  OAI21X1  g0190(.A0(new_n831_), .A1(new_n661_), .B0(new_n832_), .Y(new_n833_));
  AND2X1   g0191(.A(new_n833_), .B(\in0[24] ), .Y(new_n834_));
  NOR3X1   g0192(.A(new_n834_), .B(new_n816_), .C(\in0[25] ), .Y(new_n835_));
  OAI21X1  g0193(.A0(new_n834_), .A1(new_n816_), .B0(\in0[25] ), .Y(new_n836_));
  OAI21X1  g0194(.A0(new_n835_), .A1(\in1[25] ), .B0(new_n836_), .Y(new_n837_));
  INVX1    g0195(.A(\in1[26] ), .Y(new_n838_));
  AND2X1   g0196(.A(new_n838_), .B(\in0[26] ), .Y(new_n839_));
  AOI21X1  g0197(.A0(new_n837_), .A1(new_n658_), .B0(new_n839_), .Y(new_n840_));
  INVX1    g0198(.A(\in1[27] ), .Y(new_n841_));
  AND2X1   g0199(.A(new_n841_), .B(\in0[27] ), .Y(new_n842_));
  INVX1    g0200(.A(new_n842_), .Y(new_n843_));
  OAI21X1  g0201(.A0(new_n840_), .A1(new_n655_), .B0(new_n843_), .Y(new_n844_));
  INVX1    g0202(.A(\in1[28] ), .Y(new_n845_));
  AND2X1   g0203(.A(new_n845_), .B(\in0[28] ), .Y(new_n846_));
  AOI21X1  g0204(.A0(new_n844_), .A1(new_n653_), .B0(new_n846_), .Y(new_n847_));
  INVX1    g0205(.A(\in1[29] ), .Y(new_n848_));
  AND2X1   g0206(.A(new_n848_), .B(\in0[29] ), .Y(new_n849_));
  INVX1    g0207(.A(new_n849_), .Y(new_n850_));
  OAI21X1  g0208(.A0(new_n847_), .A1(new_n650_), .B0(new_n850_), .Y(new_n851_));
  INVX1    g0209(.A(\in1[30] ), .Y(new_n852_));
  AND2X1   g0210(.A(new_n852_), .B(\in0[30] ), .Y(new_n853_));
  AOI21X1  g0211(.A0(new_n851_), .A1(new_n648_), .B0(new_n853_), .Y(new_n854_));
  INVX1    g0212(.A(\in1[31] ), .Y(new_n855_));
  AND2X1   g0213(.A(new_n855_), .B(\in0[31] ), .Y(new_n856_));
  INVX1    g0214(.A(new_n856_), .Y(new_n857_));
  OAI21X1  g0215(.A0(new_n854_), .A1(new_n645_), .B0(new_n857_), .Y(new_n858_));
  INVX1    g0216(.A(\in0[38] ), .Y(new_n859_));
  INVX1    g0217(.A(\in0[39] ), .Y(new_n860_));
  AOI22X1  g0218(.A0(\in1[39] ), .A1(new_n860_), .B0(\in1[38] ), .B1(new_n859_), .Y(new_n861_));
  INVX1    g0219(.A(new_n861_), .Y(new_n862_));
  INVX1    g0220(.A(\in1[36] ), .Y(new_n863_));
  INVX1    g0221(.A(\in1[37] ), .Y(new_n864_));
  OAI22X1  g0222(.A0(new_n864_), .A1(\in0[37] ), .B0(new_n863_), .B1(\in0[36] ), .Y(new_n865_));
  INVX1    g0223(.A(\in0[34] ), .Y(new_n866_));
  INVX1    g0224(.A(\in0[35] ), .Y(new_n867_));
  AOI22X1  g0225(.A0(\in1[35] ), .A1(new_n867_), .B0(\in1[34] ), .B1(new_n866_), .Y(new_n868_));
  INVX1    g0226(.A(new_n868_), .Y(new_n869_));
  INVX1    g0227(.A(\in1[32] ), .Y(new_n870_));
  INVX1    g0228(.A(\in1[33] ), .Y(new_n871_));
  OAI22X1  g0229(.A0(new_n871_), .A1(\in0[33] ), .B0(new_n870_), .B1(\in0[32] ), .Y(new_n872_));
  NOR4X1   g0230(.A(new_n872_), .B(new_n869_), .C(new_n865_), .D(new_n862_), .Y(new_n873_));
  NOR2X1   g0231(.A(new_n865_), .B(new_n862_), .Y(new_n874_));
  AND2X1   g0232(.A(new_n870_), .B(\in0[32] ), .Y(new_n875_));
  OAI21X1  g0233(.A0(new_n871_), .A1(\in0[33] ), .B0(new_n875_), .Y(new_n876_));
  INVX1    g0234(.A(\in1[34] ), .Y(new_n877_));
  AOI22X1  g0235(.A0(new_n877_), .A1(\in0[34] ), .B0(new_n871_), .B1(\in0[33] ), .Y(new_n878_));
  AND2X1   g0236(.A(new_n878_), .B(new_n876_), .Y(new_n879_));
  OAI22X1  g0237(.A0(new_n879_), .A1(new_n869_), .B0(\in1[35] ), .B1(new_n867_), .Y(new_n880_));
  INVX1    g0238(.A(\in0[36] ), .Y(new_n881_));
  INVX1    g0239(.A(\in0[37] ), .Y(new_n882_));
  AND2X1   g0240(.A(\in1[37] ), .B(new_n882_), .Y(new_n883_));
  NOR3X1   g0241(.A(new_n883_), .B(\in1[36] ), .C(new_n881_), .Y(new_n884_));
  AOI21X1  g0242(.A0(new_n864_), .A1(\in0[37] ), .B0(new_n884_), .Y(new_n885_));
  INVX1    g0243(.A(\in1[39] ), .Y(new_n886_));
  AND2X1   g0244(.A(\in1[39] ), .B(new_n860_), .Y(new_n887_));
  NOR3X1   g0245(.A(new_n887_), .B(\in1[38] ), .C(new_n859_), .Y(new_n888_));
  AOI21X1  g0246(.A0(new_n886_), .A1(\in0[39] ), .B0(new_n888_), .Y(new_n889_));
  OAI21X1  g0247(.A0(new_n885_), .A1(new_n862_), .B0(new_n889_), .Y(new_n890_));
  AOI21X1  g0248(.A0(new_n880_), .A1(new_n874_), .B0(new_n890_), .Y(new_n891_));
  INVX1    g0249(.A(new_n891_), .Y(new_n892_));
  AOI21X1  g0250(.A0(new_n873_), .A1(new_n858_), .B0(new_n892_), .Y(new_n893_));
  INVX1    g0251(.A(\in0[46] ), .Y(new_n894_));
  INVX1    g0252(.A(\in0[47] ), .Y(new_n895_));
  AOI22X1  g0253(.A0(\in1[47] ), .A1(new_n895_), .B0(\in1[46] ), .B1(new_n894_), .Y(new_n896_));
  INVX1    g0254(.A(new_n896_), .Y(new_n897_));
  INVX1    g0255(.A(\in1[44] ), .Y(new_n898_));
  INVX1    g0256(.A(\in1[45] ), .Y(new_n899_));
  OAI22X1  g0257(.A0(new_n899_), .A1(\in0[45] ), .B0(new_n898_), .B1(\in0[44] ), .Y(new_n900_));
  INVX1    g0258(.A(\in0[42] ), .Y(new_n901_));
  INVX1    g0259(.A(\in0[43] ), .Y(new_n902_));
  AOI22X1  g0260(.A0(\in1[43] ), .A1(new_n902_), .B0(\in1[42] ), .B1(new_n901_), .Y(new_n903_));
  INVX1    g0261(.A(new_n903_), .Y(new_n904_));
  INVX1    g0262(.A(\in1[40] ), .Y(new_n905_));
  INVX1    g0263(.A(\in1[41] ), .Y(new_n906_));
  OAI22X1  g0264(.A0(new_n906_), .A1(\in0[41] ), .B0(new_n905_), .B1(\in0[40] ), .Y(new_n907_));
  NOR4X1   g0265(.A(new_n907_), .B(new_n904_), .C(new_n900_), .D(new_n897_), .Y(new_n908_));
  INVX1    g0266(.A(new_n908_), .Y(new_n909_));
  NOR2X1   g0267(.A(new_n900_), .B(new_n897_), .Y(new_n910_));
  AND2X1   g0268(.A(new_n905_), .B(\in0[40] ), .Y(new_n911_));
  OAI21X1  g0269(.A0(new_n906_), .A1(\in0[41] ), .B0(new_n911_), .Y(new_n912_));
  INVX1    g0270(.A(\in1[42] ), .Y(new_n913_));
  AOI22X1  g0271(.A0(new_n913_), .A1(\in0[42] ), .B0(new_n906_), .B1(\in0[41] ), .Y(new_n914_));
  AND2X1   g0272(.A(new_n914_), .B(new_n912_), .Y(new_n915_));
  OAI22X1  g0273(.A0(new_n915_), .A1(new_n904_), .B0(\in1[43] ), .B1(new_n902_), .Y(new_n916_));
  INVX1    g0274(.A(\in0[44] ), .Y(new_n917_));
  INVX1    g0275(.A(\in0[45] ), .Y(new_n918_));
  AND2X1   g0276(.A(\in1[45] ), .B(new_n918_), .Y(new_n919_));
  NOR3X1   g0277(.A(new_n919_), .B(\in1[44] ), .C(new_n917_), .Y(new_n920_));
  AOI21X1  g0278(.A0(new_n899_), .A1(\in0[45] ), .B0(new_n920_), .Y(new_n921_));
  INVX1    g0279(.A(\in1[47] ), .Y(new_n922_));
  AND2X1   g0280(.A(\in1[47] ), .B(new_n895_), .Y(new_n923_));
  NOR3X1   g0281(.A(new_n923_), .B(\in1[46] ), .C(new_n894_), .Y(new_n924_));
  AOI21X1  g0282(.A0(new_n922_), .A1(\in0[47] ), .B0(new_n924_), .Y(new_n925_));
  OAI21X1  g0283(.A0(new_n921_), .A1(new_n897_), .B0(new_n925_), .Y(new_n926_));
  AOI21X1  g0284(.A0(new_n916_), .A1(new_n910_), .B0(new_n926_), .Y(new_n927_));
  OAI21X1  g0285(.A0(new_n909_), .A1(new_n893_), .B0(new_n927_), .Y(new_n928_));
  INVX1    g0286(.A(\in0[54] ), .Y(new_n929_));
  INVX1    g0287(.A(\in0[55] ), .Y(new_n930_));
  AOI22X1  g0288(.A0(\in1[55] ), .A1(new_n930_), .B0(\in1[54] ), .B1(new_n929_), .Y(new_n931_));
  INVX1    g0289(.A(new_n931_), .Y(new_n932_));
  INVX1    g0290(.A(\in1[52] ), .Y(new_n933_));
  INVX1    g0291(.A(\in1[53] ), .Y(new_n934_));
  OAI22X1  g0292(.A0(new_n934_), .A1(\in0[53] ), .B0(new_n933_), .B1(\in0[52] ), .Y(new_n935_));
  INVX1    g0293(.A(\in0[50] ), .Y(new_n936_));
  INVX1    g0294(.A(\in0[51] ), .Y(new_n937_));
  AOI22X1  g0295(.A0(\in1[51] ), .A1(new_n937_), .B0(\in1[50] ), .B1(new_n936_), .Y(new_n938_));
  INVX1    g0296(.A(new_n938_), .Y(new_n939_));
  INVX1    g0297(.A(\in1[48] ), .Y(new_n940_));
  INVX1    g0298(.A(\in1[49] ), .Y(new_n941_));
  OAI22X1  g0299(.A0(new_n941_), .A1(\in0[49] ), .B0(new_n940_), .B1(\in0[48] ), .Y(new_n942_));
  NOR4X1   g0300(.A(new_n942_), .B(new_n939_), .C(new_n935_), .D(new_n932_), .Y(new_n943_));
  NOR2X1   g0301(.A(new_n935_), .B(new_n932_), .Y(new_n944_));
  AND2X1   g0302(.A(new_n940_), .B(\in0[48] ), .Y(new_n945_));
  OAI21X1  g0303(.A0(new_n941_), .A1(\in0[49] ), .B0(new_n945_), .Y(new_n946_));
  INVX1    g0304(.A(\in1[50] ), .Y(new_n947_));
  AOI22X1  g0305(.A0(new_n947_), .A1(\in0[50] ), .B0(new_n941_), .B1(\in0[49] ), .Y(new_n948_));
  AND2X1   g0306(.A(new_n948_), .B(new_n946_), .Y(new_n949_));
  OAI22X1  g0307(.A0(new_n949_), .A1(new_n939_), .B0(\in1[51] ), .B1(new_n937_), .Y(new_n950_));
  AND2X1   g0308(.A(new_n933_), .B(\in0[52] ), .Y(new_n951_));
  OAI21X1  g0309(.A0(new_n934_), .A1(\in0[53] ), .B0(new_n951_), .Y(new_n952_));
  INVX1    g0310(.A(\in1[54] ), .Y(new_n953_));
  AOI22X1  g0311(.A0(new_n953_), .A1(\in0[54] ), .B0(new_n934_), .B1(\in0[53] ), .Y(new_n954_));
  AND2X1   g0312(.A(new_n954_), .B(new_n952_), .Y(new_n955_));
  OAI22X1  g0313(.A0(new_n955_), .A1(new_n932_), .B0(\in1[55] ), .B1(new_n930_), .Y(new_n956_));
  AOI21X1  g0314(.A0(new_n950_), .A1(new_n944_), .B0(new_n956_), .Y(new_n957_));
  INVX1    g0315(.A(new_n957_), .Y(new_n958_));
  AOI21X1  g0316(.A0(new_n943_), .A1(new_n928_), .B0(new_n958_), .Y(new_n959_));
  INVX1    g0317(.A(\in0[62] ), .Y(new_n960_));
  INVX1    g0318(.A(\in0[63] ), .Y(new_n961_));
  AOI22X1  g0319(.A0(\in1[63] ), .A1(new_n961_), .B0(\in1[62] ), .B1(new_n960_), .Y(new_n962_));
  INVX1    g0320(.A(new_n962_), .Y(new_n963_));
  INVX1    g0321(.A(\in1[60] ), .Y(new_n964_));
  INVX1    g0322(.A(\in1[61] ), .Y(new_n965_));
  OAI22X1  g0323(.A0(new_n965_), .A1(\in0[61] ), .B0(new_n964_), .B1(\in0[60] ), .Y(new_n966_));
  INVX1    g0324(.A(\in0[58] ), .Y(new_n967_));
  INVX1    g0325(.A(\in0[59] ), .Y(new_n968_));
  AOI22X1  g0326(.A0(\in1[59] ), .A1(new_n968_), .B0(\in1[58] ), .B1(new_n967_), .Y(new_n969_));
  INVX1    g0327(.A(new_n969_), .Y(new_n970_));
  INVX1    g0328(.A(\in1[56] ), .Y(new_n971_));
  INVX1    g0329(.A(\in1[57] ), .Y(new_n972_));
  OAI22X1  g0330(.A0(new_n972_), .A1(\in0[57] ), .B0(new_n971_), .B1(\in0[56] ), .Y(new_n973_));
  NOR4X1   g0331(.A(new_n973_), .B(new_n970_), .C(new_n966_), .D(new_n963_), .Y(new_n974_));
  INVX1    g0332(.A(new_n974_), .Y(new_n975_));
  NOR2X1   g0333(.A(new_n966_), .B(new_n963_), .Y(new_n976_));
  AND2X1   g0334(.A(new_n971_), .B(\in0[56] ), .Y(new_n977_));
  OAI21X1  g0335(.A0(new_n972_), .A1(\in0[57] ), .B0(new_n977_), .Y(new_n978_));
  INVX1    g0336(.A(\in1[58] ), .Y(new_n979_));
  AOI22X1  g0337(.A0(new_n979_), .A1(\in0[58] ), .B0(new_n972_), .B1(\in0[57] ), .Y(new_n980_));
  AND2X1   g0338(.A(new_n980_), .B(new_n978_), .Y(new_n981_));
  OAI22X1  g0339(.A0(new_n981_), .A1(new_n970_), .B0(\in1[59] ), .B1(new_n968_), .Y(new_n982_));
  INVX1    g0340(.A(\in0[60] ), .Y(new_n983_));
  INVX1    g0341(.A(\in0[61] ), .Y(new_n984_));
  AND2X1   g0342(.A(\in1[61] ), .B(new_n984_), .Y(new_n985_));
  NOR3X1   g0343(.A(new_n985_), .B(\in1[60] ), .C(new_n983_), .Y(new_n986_));
  AOI21X1  g0344(.A0(new_n965_), .A1(\in0[61] ), .B0(new_n986_), .Y(new_n987_));
  INVX1    g0345(.A(\in1[63] ), .Y(new_n988_));
  AND2X1   g0346(.A(\in1[63] ), .B(new_n961_), .Y(new_n989_));
  NOR3X1   g0347(.A(new_n989_), .B(\in1[62] ), .C(new_n960_), .Y(new_n990_));
  AOI21X1  g0348(.A0(new_n988_), .A1(\in0[63] ), .B0(new_n990_), .Y(new_n991_));
  OAI21X1  g0349(.A0(new_n987_), .A1(new_n963_), .B0(new_n991_), .Y(new_n992_));
  AOI21X1  g0350(.A0(new_n982_), .A1(new_n976_), .B0(new_n992_), .Y(new_n993_));
  OAI21X1  g0351(.A0(new_n975_), .A1(new_n959_), .B0(new_n993_), .Y(new_n994_));
  INVX1    g0352(.A(\in0[66] ), .Y(new_n995_));
  INVX1    g0353(.A(\in0[67] ), .Y(new_n996_));
  AOI22X1  g0354(.A0(\in1[67] ), .A1(new_n996_), .B0(\in1[66] ), .B1(new_n995_), .Y(new_n997_));
  INVX1    g0355(.A(\in0[64] ), .Y(new_n998_));
  INVX1    g0356(.A(\in0[65] ), .Y(new_n999_));
  AOI22X1  g0357(.A0(\in1[65] ), .A1(new_n999_), .B0(\in1[64] ), .B1(new_n998_), .Y(new_n1000_));
  AND2X1   g0358(.A(new_n1000_), .B(new_n997_), .Y(new_n1001_));
  OR2X1    g0359(.A(\in1[67] ), .B(new_n996_), .Y(new_n1002_));
  AND2X1   g0360(.A(\in1[65] ), .B(new_n999_), .Y(new_n1003_));
  NOR3X1   g0361(.A(new_n1003_), .B(\in1[64] ), .C(new_n998_), .Y(new_n1004_));
  INVX1    g0362(.A(\in1[65] ), .Y(new_n1005_));
  INVX1    g0363(.A(\in1[66] ), .Y(new_n1006_));
  AOI22X1  g0364(.A0(new_n1006_), .A1(\in0[66] ), .B0(new_n1005_), .B1(\in0[65] ), .Y(new_n1007_));
  INVX1    g0365(.A(new_n1007_), .Y(new_n1008_));
  OAI21X1  g0366(.A0(new_n1008_), .A1(new_n1004_), .B0(new_n997_), .Y(new_n1009_));
  AND2X1   g0367(.A(new_n1009_), .B(new_n1002_), .Y(new_n1010_));
  INVX1    g0368(.A(new_n1010_), .Y(new_n1011_));
  AOI21X1  g0369(.A0(new_n1001_), .A1(new_n994_), .B0(new_n1011_), .Y(new_n1012_));
  INVX1    g0370(.A(\in0[70] ), .Y(new_n1013_));
  INVX1    g0371(.A(\in0[71] ), .Y(new_n1014_));
  AOI22X1  g0372(.A0(\in1[71] ), .A1(new_n1014_), .B0(\in1[70] ), .B1(new_n1013_), .Y(new_n1015_));
  INVX1    g0373(.A(\in0[68] ), .Y(new_n1016_));
  INVX1    g0374(.A(\in0[69] ), .Y(new_n1017_));
  AOI22X1  g0375(.A0(\in1[69] ), .A1(new_n1017_), .B0(\in1[68] ), .B1(new_n1016_), .Y(new_n1018_));
  AND2X1   g0376(.A(new_n1018_), .B(new_n1015_), .Y(new_n1019_));
  INVX1    g0377(.A(new_n1019_), .Y(new_n1020_));
  AND2X1   g0378(.A(\in1[69] ), .B(new_n1017_), .Y(new_n1021_));
  NOR3X1   g0379(.A(new_n1021_), .B(\in1[68] ), .C(new_n1016_), .Y(new_n1022_));
  INVX1    g0380(.A(\in1[69] ), .Y(new_n1023_));
  AND2X1   g0381(.A(new_n1023_), .B(\in0[69] ), .Y(new_n1024_));
  OAI21X1  g0382(.A0(new_n1024_), .A1(new_n1022_), .B0(new_n1015_), .Y(new_n1025_));
  INVX1    g0383(.A(\in1[71] ), .Y(new_n1026_));
  AND2X1   g0384(.A(\in1[71] ), .B(new_n1014_), .Y(new_n1027_));
  NOR3X1   g0385(.A(new_n1027_), .B(\in1[70] ), .C(new_n1013_), .Y(new_n1028_));
  AOI21X1  g0386(.A0(new_n1026_), .A1(\in0[71] ), .B0(new_n1028_), .Y(new_n1029_));
  AND2X1   g0387(.A(new_n1029_), .B(new_n1025_), .Y(new_n1030_));
  OAI21X1  g0388(.A0(new_n1020_), .A1(new_n1012_), .B0(new_n1030_), .Y(new_n1031_));
  INVX1    g0389(.A(\in0[74] ), .Y(new_n1032_));
  INVX1    g0390(.A(\in0[75] ), .Y(new_n1033_));
  AOI22X1  g0391(.A0(\in1[75] ), .A1(new_n1033_), .B0(\in1[74] ), .B1(new_n1032_), .Y(new_n1034_));
  INVX1    g0392(.A(\in0[72] ), .Y(new_n1035_));
  INVX1    g0393(.A(\in0[73] ), .Y(new_n1036_));
  AOI22X1  g0394(.A0(\in1[73] ), .A1(new_n1036_), .B0(\in1[72] ), .B1(new_n1035_), .Y(new_n1037_));
  AND2X1   g0395(.A(new_n1037_), .B(new_n1034_), .Y(new_n1038_));
  OR2X1    g0396(.A(\in1[75] ), .B(new_n1033_), .Y(new_n1039_));
  AND2X1   g0397(.A(\in1[73] ), .B(new_n1036_), .Y(new_n1040_));
  NOR3X1   g0398(.A(new_n1040_), .B(\in1[72] ), .C(new_n1035_), .Y(new_n1041_));
  INVX1    g0399(.A(\in1[73] ), .Y(new_n1042_));
  INVX1    g0400(.A(\in1[74] ), .Y(new_n1043_));
  AOI22X1  g0401(.A0(new_n1043_), .A1(\in0[74] ), .B0(new_n1042_), .B1(\in0[73] ), .Y(new_n1044_));
  INVX1    g0402(.A(new_n1044_), .Y(new_n1045_));
  OAI21X1  g0403(.A0(new_n1045_), .A1(new_n1041_), .B0(new_n1034_), .Y(new_n1046_));
  AND2X1   g0404(.A(new_n1046_), .B(new_n1039_), .Y(new_n1047_));
  INVX1    g0405(.A(new_n1047_), .Y(new_n1048_));
  AOI21X1  g0406(.A0(new_n1038_), .A1(new_n1031_), .B0(new_n1048_), .Y(new_n1049_));
  INVX1    g0407(.A(\in0[78] ), .Y(new_n1050_));
  INVX1    g0408(.A(\in0[79] ), .Y(new_n1051_));
  AOI22X1  g0409(.A0(\in1[79] ), .A1(new_n1051_), .B0(\in1[78] ), .B1(new_n1050_), .Y(new_n1052_));
  INVX1    g0410(.A(\in0[76] ), .Y(new_n1053_));
  INVX1    g0411(.A(\in0[77] ), .Y(new_n1054_));
  AOI22X1  g0412(.A0(\in1[77] ), .A1(new_n1054_), .B0(\in1[76] ), .B1(new_n1053_), .Y(new_n1055_));
  AND2X1   g0413(.A(new_n1055_), .B(new_n1052_), .Y(new_n1056_));
  INVX1    g0414(.A(new_n1056_), .Y(new_n1057_));
  AND2X1   g0415(.A(\in1[77] ), .B(new_n1054_), .Y(new_n1058_));
  NOR3X1   g0416(.A(new_n1058_), .B(\in1[76] ), .C(new_n1053_), .Y(new_n1059_));
  INVX1    g0417(.A(\in1[77] ), .Y(new_n1060_));
  AND2X1   g0418(.A(new_n1060_), .B(\in0[77] ), .Y(new_n1061_));
  OAI21X1  g0419(.A0(new_n1061_), .A1(new_n1059_), .B0(new_n1052_), .Y(new_n1062_));
  INVX1    g0420(.A(\in1[79] ), .Y(new_n1063_));
  AND2X1   g0421(.A(\in1[79] ), .B(new_n1051_), .Y(new_n1064_));
  NOR3X1   g0422(.A(new_n1064_), .B(\in1[78] ), .C(new_n1050_), .Y(new_n1065_));
  AOI21X1  g0423(.A0(new_n1063_), .A1(\in0[79] ), .B0(new_n1065_), .Y(new_n1066_));
  AND2X1   g0424(.A(new_n1066_), .B(new_n1062_), .Y(new_n1067_));
  OAI21X1  g0425(.A0(new_n1057_), .A1(new_n1049_), .B0(new_n1067_), .Y(new_n1068_));
  INVX1    g0426(.A(\in0[82] ), .Y(new_n1069_));
  INVX1    g0427(.A(\in0[83] ), .Y(new_n1070_));
  AOI22X1  g0428(.A0(\in1[83] ), .A1(new_n1070_), .B0(\in1[82] ), .B1(new_n1069_), .Y(new_n1071_));
  INVX1    g0429(.A(\in0[80] ), .Y(new_n1072_));
  INVX1    g0430(.A(\in0[81] ), .Y(new_n1073_));
  AOI22X1  g0431(.A0(\in1[81] ), .A1(new_n1073_), .B0(\in1[80] ), .B1(new_n1072_), .Y(new_n1074_));
  AND2X1   g0432(.A(new_n1074_), .B(new_n1071_), .Y(new_n1075_));
  OR2X1    g0433(.A(\in1[83] ), .B(new_n1070_), .Y(new_n1076_));
  AND2X1   g0434(.A(\in1[81] ), .B(new_n1073_), .Y(new_n1077_));
  NOR3X1   g0435(.A(new_n1077_), .B(\in1[80] ), .C(new_n1072_), .Y(new_n1078_));
  INVX1    g0436(.A(\in1[81] ), .Y(new_n1079_));
  INVX1    g0437(.A(\in1[82] ), .Y(new_n1080_));
  AOI22X1  g0438(.A0(new_n1080_), .A1(\in0[82] ), .B0(new_n1079_), .B1(\in0[81] ), .Y(new_n1081_));
  INVX1    g0439(.A(new_n1081_), .Y(new_n1082_));
  OAI21X1  g0440(.A0(new_n1082_), .A1(new_n1078_), .B0(new_n1071_), .Y(new_n1083_));
  AND2X1   g0441(.A(new_n1083_), .B(new_n1076_), .Y(new_n1084_));
  INVX1    g0442(.A(new_n1084_), .Y(new_n1085_));
  AOI21X1  g0443(.A0(new_n1075_), .A1(new_n1068_), .B0(new_n1085_), .Y(new_n1086_));
  INVX1    g0444(.A(\in0[86] ), .Y(new_n1087_));
  INVX1    g0445(.A(\in0[87] ), .Y(new_n1088_));
  AOI22X1  g0446(.A0(\in1[87] ), .A1(new_n1088_), .B0(\in1[86] ), .B1(new_n1087_), .Y(new_n1089_));
  INVX1    g0447(.A(\in0[84] ), .Y(new_n1090_));
  INVX1    g0448(.A(\in0[85] ), .Y(new_n1091_));
  AOI22X1  g0449(.A0(\in1[85] ), .A1(new_n1091_), .B0(\in1[84] ), .B1(new_n1090_), .Y(new_n1092_));
  AND2X1   g0450(.A(new_n1092_), .B(new_n1089_), .Y(new_n1093_));
  INVX1    g0451(.A(new_n1093_), .Y(new_n1094_));
  AND2X1   g0452(.A(\in1[85] ), .B(new_n1091_), .Y(new_n1095_));
  NOR3X1   g0453(.A(new_n1095_), .B(\in1[84] ), .C(new_n1090_), .Y(new_n1096_));
  INVX1    g0454(.A(\in1[85] ), .Y(new_n1097_));
  AND2X1   g0455(.A(new_n1097_), .B(\in0[85] ), .Y(new_n1098_));
  OAI21X1  g0456(.A0(new_n1098_), .A1(new_n1096_), .B0(new_n1089_), .Y(new_n1099_));
  INVX1    g0457(.A(\in1[87] ), .Y(new_n1100_));
  AND2X1   g0458(.A(\in1[87] ), .B(new_n1088_), .Y(new_n1101_));
  NOR3X1   g0459(.A(new_n1101_), .B(\in1[86] ), .C(new_n1087_), .Y(new_n1102_));
  AOI21X1  g0460(.A0(new_n1100_), .A1(\in0[87] ), .B0(new_n1102_), .Y(new_n1103_));
  AND2X1   g0461(.A(new_n1103_), .B(new_n1099_), .Y(new_n1104_));
  OAI21X1  g0462(.A0(new_n1094_), .A1(new_n1086_), .B0(new_n1104_), .Y(new_n1105_));
  INVX1    g0463(.A(\in0[90] ), .Y(new_n1106_));
  INVX1    g0464(.A(\in0[91] ), .Y(new_n1107_));
  AOI22X1  g0465(.A0(\in1[91] ), .A1(new_n1107_), .B0(\in1[90] ), .B1(new_n1106_), .Y(new_n1108_));
  INVX1    g0466(.A(\in0[88] ), .Y(new_n1109_));
  INVX1    g0467(.A(\in0[89] ), .Y(new_n1110_));
  AOI22X1  g0468(.A0(\in1[89] ), .A1(new_n1110_), .B0(\in1[88] ), .B1(new_n1109_), .Y(new_n1111_));
  AND2X1   g0469(.A(new_n1111_), .B(new_n1108_), .Y(new_n1112_));
  OR2X1    g0470(.A(\in1[91] ), .B(new_n1107_), .Y(new_n1113_));
  AND2X1   g0471(.A(\in1[89] ), .B(new_n1110_), .Y(new_n1114_));
  NOR3X1   g0472(.A(new_n1114_), .B(\in1[88] ), .C(new_n1109_), .Y(new_n1115_));
  INVX1    g0473(.A(\in1[89] ), .Y(new_n1116_));
  INVX1    g0474(.A(\in1[90] ), .Y(new_n1117_));
  AOI22X1  g0475(.A0(new_n1117_), .A1(\in0[90] ), .B0(new_n1116_), .B1(\in0[89] ), .Y(new_n1118_));
  INVX1    g0476(.A(new_n1118_), .Y(new_n1119_));
  OAI21X1  g0477(.A0(new_n1119_), .A1(new_n1115_), .B0(new_n1108_), .Y(new_n1120_));
  AND2X1   g0478(.A(new_n1120_), .B(new_n1113_), .Y(new_n1121_));
  INVX1    g0479(.A(new_n1121_), .Y(new_n1122_));
  AOI21X1  g0480(.A0(new_n1112_), .A1(new_n1105_), .B0(new_n1122_), .Y(new_n1123_));
  INVX1    g0481(.A(\in0[94] ), .Y(new_n1124_));
  INVX1    g0482(.A(\in0[95] ), .Y(new_n1125_));
  AOI22X1  g0483(.A0(\in1[95] ), .A1(new_n1125_), .B0(\in1[94] ), .B1(new_n1124_), .Y(new_n1126_));
  INVX1    g0484(.A(\in0[92] ), .Y(new_n1127_));
  INVX1    g0485(.A(\in0[93] ), .Y(new_n1128_));
  AOI22X1  g0486(.A0(\in1[93] ), .A1(new_n1128_), .B0(\in1[92] ), .B1(new_n1127_), .Y(new_n1129_));
  AND2X1   g0487(.A(new_n1129_), .B(new_n1126_), .Y(new_n1130_));
  INVX1    g0488(.A(new_n1130_), .Y(new_n1131_));
  AND2X1   g0489(.A(\in1[93] ), .B(new_n1128_), .Y(new_n1132_));
  NOR3X1   g0490(.A(new_n1132_), .B(\in1[92] ), .C(new_n1127_), .Y(new_n1133_));
  INVX1    g0491(.A(\in1[93] ), .Y(new_n1134_));
  AND2X1   g0492(.A(new_n1134_), .B(\in0[93] ), .Y(new_n1135_));
  OAI21X1  g0493(.A0(new_n1135_), .A1(new_n1133_), .B0(new_n1126_), .Y(new_n1136_));
  INVX1    g0494(.A(\in1[95] ), .Y(new_n1137_));
  AND2X1   g0495(.A(\in1[95] ), .B(new_n1125_), .Y(new_n1138_));
  NOR3X1   g0496(.A(new_n1138_), .B(\in1[94] ), .C(new_n1124_), .Y(new_n1139_));
  AOI21X1  g0497(.A0(new_n1137_), .A1(\in0[95] ), .B0(new_n1139_), .Y(new_n1140_));
  AND2X1   g0498(.A(new_n1140_), .B(new_n1136_), .Y(new_n1141_));
  OAI21X1  g0499(.A0(new_n1131_), .A1(new_n1123_), .B0(new_n1141_), .Y(new_n1142_));
  INVX1    g0500(.A(\in0[98] ), .Y(new_n1143_));
  INVX1    g0501(.A(\in0[99] ), .Y(new_n1144_));
  AOI22X1  g0502(.A0(\in1[99] ), .A1(new_n1144_), .B0(\in1[98] ), .B1(new_n1143_), .Y(new_n1145_));
  INVX1    g0503(.A(\in0[96] ), .Y(new_n1146_));
  INVX1    g0504(.A(\in0[97] ), .Y(new_n1147_));
  AOI22X1  g0505(.A0(\in1[97] ), .A1(new_n1147_), .B0(\in1[96] ), .B1(new_n1146_), .Y(new_n1148_));
  AND2X1   g0506(.A(new_n1148_), .B(new_n1145_), .Y(new_n1149_));
  OR2X1    g0507(.A(\in1[99] ), .B(new_n1144_), .Y(new_n1150_));
  AND2X1   g0508(.A(\in1[97] ), .B(new_n1147_), .Y(new_n1151_));
  NOR3X1   g0509(.A(new_n1151_), .B(\in1[96] ), .C(new_n1146_), .Y(new_n1152_));
  INVX1    g0510(.A(\in1[97] ), .Y(new_n1153_));
  INVX1    g0511(.A(\in1[98] ), .Y(new_n1154_));
  AOI22X1  g0512(.A0(new_n1154_), .A1(\in0[98] ), .B0(new_n1153_), .B1(\in0[97] ), .Y(new_n1155_));
  INVX1    g0513(.A(new_n1155_), .Y(new_n1156_));
  OAI21X1  g0514(.A0(new_n1156_), .A1(new_n1152_), .B0(new_n1145_), .Y(new_n1157_));
  AND2X1   g0515(.A(new_n1157_), .B(new_n1150_), .Y(new_n1158_));
  INVX1    g0516(.A(new_n1158_), .Y(new_n1159_));
  AOI21X1  g0517(.A0(new_n1149_), .A1(new_n1142_), .B0(new_n1159_), .Y(new_n1160_));
  INVX1    g0518(.A(\in0[102] ), .Y(new_n1161_));
  INVX1    g0519(.A(\in0[103] ), .Y(new_n1162_));
  AOI22X1  g0520(.A0(\in1[103] ), .A1(new_n1162_), .B0(\in1[102] ), .B1(new_n1161_), .Y(new_n1163_));
  INVX1    g0521(.A(\in0[100] ), .Y(new_n1164_));
  INVX1    g0522(.A(\in0[101] ), .Y(new_n1165_));
  AOI22X1  g0523(.A0(\in1[101] ), .A1(new_n1165_), .B0(\in1[100] ), .B1(new_n1164_), .Y(new_n1166_));
  AND2X1   g0524(.A(new_n1166_), .B(new_n1163_), .Y(new_n1167_));
  INVX1    g0525(.A(new_n1167_), .Y(new_n1168_));
  AND2X1   g0526(.A(\in1[101] ), .B(new_n1165_), .Y(new_n1169_));
  NOR3X1   g0527(.A(new_n1169_), .B(\in1[100] ), .C(new_n1164_), .Y(new_n1170_));
  INVX1    g0528(.A(\in1[101] ), .Y(new_n1171_));
  AND2X1   g0529(.A(new_n1171_), .B(\in0[101] ), .Y(new_n1172_));
  OAI21X1  g0530(.A0(new_n1172_), .A1(new_n1170_), .B0(new_n1163_), .Y(new_n1173_));
  INVX1    g0531(.A(\in1[103] ), .Y(new_n1174_));
  AND2X1   g0532(.A(\in1[103] ), .B(new_n1162_), .Y(new_n1175_));
  NOR3X1   g0533(.A(new_n1175_), .B(\in1[102] ), .C(new_n1161_), .Y(new_n1176_));
  AOI21X1  g0534(.A0(new_n1174_), .A1(\in0[103] ), .B0(new_n1176_), .Y(new_n1177_));
  AND2X1   g0535(.A(new_n1177_), .B(new_n1173_), .Y(new_n1178_));
  OAI21X1  g0536(.A0(new_n1168_), .A1(new_n1160_), .B0(new_n1178_), .Y(new_n1179_));
  INVX1    g0537(.A(\in0[106] ), .Y(new_n1180_));
  INVX1    g0538(.A(\in0[107] ), .Y(new_n1181_));
  AOI22X1  g0539(.A0(\in1[107] ), .A1(new_n1181_), .B0(\in1[106] ), .B1(new_n1180_), .Y(new_n1182_));
  INVX1    g0540(.A(\in0[104] ), .Y(new_n1183_));
  INVX1    g0541(.A(\in0[105] ), .Y(new_n1184_));
  AOI22X1  g0542(.A0(\in1[105] ), .A1(new_n1184_), .B0(\in1[104] ), .B1(new_n1183_), .Y(new_n1185_));
  AND2X1   g0543(.A(new_n1185_), .B(new_n1182_), .Y(new_n1186_));
  OR2X1    g0544(.A(\in1[107] ), .B(new_n1181_), .Y(new_n1187_));
  AND2X1   g0545(.A(\in1[105] ), .B(new_n1184_), .Y(new_n1188_));
  NOR3X1   g0546(.A(new_n1188_), .B(\in1[104] ), .C(new_n1183_), .Y(new_n1189_));
  INVX1    g0547(.A(\in1[105] ), .Y(new_n1190_));
  INVX1    g0548(.A(\in1[106] ), .Y(new_n1191_));
  AOI22X1  g0549(.A0(new_n1191_), .A1(\in0[106] ), .B0(new_n1190_), .B1(\in0[105] ), .Y(new_n1192_));
  INVX1    g0550(.A(new_n1192_), .Y(new_n1193_));
  OAI21X1  g0551(.A0(new_n1193_), .A1(new_n1189_), .B0(new_n1182_), .Y(new_n1194_));
  AND2X1   g0552(.A(new_n1194_), .B(new_n1187_), .Y(new_n1195_));
  INVX1    g0553(.A(new_n1195_), .Y(new_n1196_));
  AOI21X1  g0554(.A0(new_n1186_), .A1(new_n1179_), .B0(new_n1196_), .Y(new_n1197_));
  INVX1    g0555(.A(\in0[110] ), .Y(new_n1198_));
  INVX1    g0556(.A(\in0[111] ), .Y(new_n1199_));
  AOI22X1  g0557(.A0(\in1[111] ), .A1(new_n1199_), .B0(\in1[110] ), .B1(new_n1198_), .Y(new_n1200_));
  INVX1    g0558(.A(\in0[108] ), .Y(new_n1201_));
  INVX1    g0559(.A(\in0[109] ), .Y(new_n1202_));
  AOI22X1  g0560(.A0(\in1[109] ), .A1(new_n1202_), .B0(\in1[108] ), .B1(new_n1201_), .Y(new_n1203_));
  AND2X1   g0561(.A(new_n1203_), .B(new_n1200_), .Y(new_n1204_));
  INVX1    g0562(.A(new_n1204_), .Y(new_n1205_));
  AND2X1   g0563(.A(\in1[109] ), .B(new_n1202_), .Y(new_n1206_));
  NOR3X1   g0564(.A(new_n1206_), .B(\in1[108] ), .C(new_n1201_), .Y(new_n1207_));
  INVX1    g0565(.A(\in1[109] ), .Y(new_n1208_));
  AND2X1   g0566(.A(new_n1208_), .B(\in0[109] ), .Y(new_n1209_));
  OAI21X1  g0567(.A0(new_n1209_), .A1(new_n1207_), .B0(new_n1200_), .Y(new_n1210_));
  INVX1    g0568(.A(\in1[111] ), .Y(new_n1211_));
  AND2X1   g0569(.A(\in1[111] ), .B(new_n1199_), .Y(new_n1212_));
  NOR3X1   g0570(.A(new_n1212_), .B(\in1[110] ), .C(new_n1198_), .Y(new_n1213_));
  AOI21X1  g0571(.A0(new_n1211_), .A1(\in0[111] ), .B0(new_n1213_), .Y(new_n1214_));
  AND2X1   g0572(.A(new_n1214_), .B(new_n1210_), .Y(new_n1215_));
  OAI21X1  g0573(.A0(new_n1205_), .A1(new_n1197_), .B0(new_n1215_), .Y(new_n1216_));
  INVX1    g0574(.A(\in0[114] ), .Y(new_n1217_));
  INVX1    g0575(.A(\in0[115] ), .Y(new_n1218_));
  AOI22X1  g0576(.A0(\in1[115] ), .A1(new_n1218_), .B0(\in1[114] ), .B1(new_n1217_), .Y(new_n1219_));
  INVX1    g0577(.A(\in0[112] ), .Y(new_n1220_));
  INVX1    g0578(.A(\in0[113] ), .Y(new_n1221_));
  AOI22X1  g0579(.A0(\in1[113] ), .A1(new_n1221_), .B0(\in1[112] ), .B1(new_n1220_), .Y(new_n1222_));
  AND2X1   g0580(.A(new_n1222_), .B(new_n1219_), .Y(new_n1223_));
  OR2X1    g0581(.A(\in1[115] ), .B(new_n1218_), .Y(new_n1224_));
  AND2X1   g0582(.A(\in1[113] ), .B(new_n1221_), .Y(new_n1225_));
  NOR3X1   g0583(.A(new_n1225_), .B(\in1[112] ), .C(new_n1220_), .Y(new_n1226_));
  INVX1    g0584(.A(\in1[113] ), .Y(new_n1227_));
  INVX1    g0585(.A(\in1[114] ), .Y(new_n1228_));
  AOI22X1  g0586(.A0(new_n1228_), .A1(\in0[114] ), .B0(new_n1227_), .B1(\in0[113] ), .Y(new_n1229_));
  INVX1    g0587(.A(new_n1229_), .Y(new_n1230_));
  OAI21X1  g0588(.A0(new_n1230_), .A1(new_n1226_), .B0(new_n1219_), .Y(new_n1231_));
  AND2X1   g0589(.A(new_n1231_), .B(new_n1224_), .Y(new_n1232_));
  INVX1    g0590(.A(new_n1232_), .Y(new_n1233_));
  AOI21X1  g0591(.A0(new_n1223_), .A1(new_n1216_), .B0(new_n1233_), .Y(new_n1234_));
  INVX1    g0592(.A(\in0[118] ), .Y(new_n1235_));
  INVX1    g0593(.A(\in0[119] ), .Y(new_n1236_));
  AOI22X1  g0594(.A0(\in1[119] ), .A1(new_n1236_), .B0(\in1[118] ), .B1(new_n1235_), .Y(new_n1237_));
  INVX1    g0595(.A(\in0[116] ), .Y(new_n1238_));
  INVX1    g0596(.A(\in0[117] ), .Y(new_n1239_));
  AOI22X1  g0597(.A0(\in1[117] ), .A1(new_n1239_), .B0(\in1[116] ), .B1(new_n1238_), .Y(new_n1240_));
  AND2X1   g0598(.A(new_n1240_), .B(new_n1237_), .Y(new_n1241_));
  INVX1    g0599(.A(new_n1241_), .Y(new_n1242_));
  AND2X1   g0600(.A(\in1[117] ), .B(new_n1239_), .Y(new_n1243_));
  NOR3X1   g0601(.A(new_n1243_), .B(\in1[116] ), .C(new_n1238_), .Y(new_n1244_));
  INVX1    g0602(.A(\in1[117] ), .Y(new_n1245_));
  AND2X1   g0603(.A(new_n1245_), .B(\in0[117] ), .Y(new_n1246_));
  OAI21X1  g0604(.A0(new_n1246_), .A1(new_n1244_), .B0(new_n1237_), .Y(new_n1247_));
  INVX1    g0605(.A(\in1[119] ), .Y(new_n1248_));
  AND2X1   g0606(.A(\in1[119] ), .B(new_n1236_), .Y(new_n1249_));
  NOR3X1   g0607(.A(new_n1249_), .B(\in1[118] ), .C(new_n1235_), .Y(new_n1250_));
  AOI21X1  g0608(.A0(new_n1248_), .A1(\in0[119] ), .B0(new_n1250_), .Y(new_n1251_));
  AND2X1   g0609(.A(new_n1251_), .B(new_n1247_), .Y(new_n1252_));
  OAI21X1  g0610(.A0(new_n1242_), .A1(new_n1234_), .B0(new_n1252_), .Y(new_n1253_));
  INVX1    g0611(.A(\in0[122] ), .Y(new_n1254_));
  INVX1    g0612(.A(\in0[123] ), .Y(new_n1255_));
  AOI22X1  g0613(.A0(\in1[123] ), .A1(new_n1255_), .B0(\in1[122] ), .B1(new_n1254_), .Y(new_n1256_));
  INVX1    g0614(.A(\in0[120] ), .Y(new_n1257_));
  INVX1    g0615(.A(\in0[121] ), .Y(new_n1258_));
  AOI22X1  g0616(.A0(\in1[121] ), .A1(new_n1258_), .B0(\in1[120] ), .B1(new_n1257_), .Y(new_n1259_));
  AND2X1   g0617(.A(new_n1259_), .B(new_n1256_), .Y(new_n1260_));
  OR2X1    g0618(.A(\in1[123] ), .B(new_n1255_), .Y(new_n1261_));
  AND2X1   g0619(.A(\in1[121] ), .B(new_n1258_), .Y(new_n1262_));
  NOR3X1   g0620(.A(new_n1262_), .B(\in1[120] ), .C(new_n1257_), .Y(new_n1263_));
  INVX1    g0621(.A(\in1[121] ), .Y(new_n1264_));
  INVX1    g0622(.A(\in1[122] ), .Y(new_n1265_));
  AOI22X1  g0623(.A0(new_n1265_), .A1(\in0[122] ), .B0(new_n1264_), .B1(\in0[121] ), .Y(new_n1266_));
  INVX1    g0624(.A(new_n1266_), .Y(new_n1267_));
  OAI21X1  g0625(.A0(new_n1267_), .A1(new_n1263_), .B0(new_n1256_), .Y(new_n1268_));
  AND2X1   g0626(.A(new_n1268_), .B(new_n1261_), .Y(new_n1269_));
  INVX1    g0627(.A(new_n1269_), .Y(new_n1270_));
  AOI21X1  g0628(.A0(new_n1260_), .A1(new_n1253_), .B0(new_n1270_), .Y(new_n1271_));
  INVX1    g0629(.A(\in1[127] ), .Y(new_n1272_));
  AND2X1   g0630(.A(new_n1272_), .B(\in0[127] ), .Y(new_n1273_));
  INVX1    g0631(.A(\in0[125] ), .Y(new_n1274_));
  INVX1    g0632(.A(\in0[126] ), .Y(new_n1275_));
  AOI22X1  g0633(.A0(\in1[126] ), .A1(new_n1275_), .B0(\in1[125] ), .B1(new_n1274_), .Y(new_n1276_));
  INVX1    g0634(.A(\in0[124] ), .Y(new_n1277_));
  AOI22X1  g0635(.A0(new_n1272_), .A1(\in0[127] ), .B0(\in1[124] ), .B1(new_n1277_), .Y(new_n1278_));
  AND2X1   g0636(.A(new_n1278_), .B(new_n1276_), .Y(new_n1279_));
  INVX1    g0637(.A(new_n1279_), .Y(new_n1280_));
  INVX1    g0638(.A(\in1[126] ), .Y(new_n1281_));
  OAI22X1  g0639(.A0(\in1[125] ), .A1(new_n1274_), .B0(\in1[124] ), .B1(new_n1277_), .Y(new_n1282_));
  AOI22X1  g0640(.A0(new_n1282_), .A1(new_n1276_), .B0(new_n1281_), .B1(\in0[126] ), .Y(new_n1283_));
  OAI22X1  g0641(.A0(new_n1283_), .A1(new_n1273_), .B0(new_n1280_), .B1(new_n1271_), .Y(new_n1284_));
  INVX1    g0642(.A(\in0[127] ), .Y(new_n1285_));
  AND2X1   g0643(.A(\in1[127] ), .B(new_n1285_), .Y(new_n1286_));
  NOR3X1   g0644(.A(new_n1286_), .B(new_n1284_), .C(new_n643_), .Y(new_n1287_));
  INVX1    g0645(.A(new_n645_), .Y(new_n1288_));
  INVX1    g0646(.A(new_n650_), .Y(new_n1289_));
  INVX1    g0647(.A(new_n655_), .Y(new_n1290_));
  INVX1    g0648(.A(\in1[25] ), .Y(new_n1291_));
  INVX1    g0649(.A(\in0[25] ), .Y(new_n1292_));
  INVX1    g0650(.A(\in1[24] ), .Y(new_n1293_));
  OAI21X1  g0651(.A0(new_n833_), .A1(\in0[24] ), .B0(new_n1293_), .Y(new_n1294_));
  OR2X1    g0652(.A(new_n815_), .B(new_n659_), .Y(new_n1295_));
  NAND3X1  g0653(.A(new_n1295_), .B(new_n1294_), .C(new_n1292_), .Y(new_n1296_));
  AOI21X1  g0654(.A0(new_n1295_), .A1(new_n1294_), .B0(new_n1292_), .Y(new_n1297_));
  AOI21X1  g0655(.A0(new_n1296_), .A1(new_n1291_), .B0(new_n1297_), .Y(new_n1298_));
  INVX1    g0656(.A(new_n839_), .Y(new_n1299_));
  OAI21X1  g0657(.A0(new_n1298_), .A1(new_n657_), .B0(new_n1299_), .Y(new_n1300_));
  AOI21X1  g0658(.A0(new_n1300_), .A1(new_n1290_), .B0(new_n842_), .Y(new_n1301_));
  INVX1    g0659(.A(new_n846_), .Y(new_n1302_));
  OAI21X1  g0660(.A0(new_n1301_), .A1(new_n652_), .B0(new_n1302_), .Y(new_n1303_));
  AOI21X1  g0661(.A0(new_n1303_), .A1(new_n1289_), .B0(new_n849_), .Y(new_n1304_));
  INVX1    g0662(.A(new_n853_), .Y(new_n1305_));
  OAI21X1  g0663(.A0(new_n1304_), .A1(new_n647_), .B0(new_n1305_), .Y(new_n1306_));
  AOI21X1  g0664(.A0(new_n1306_), .A1(new_n1288_), .B0(new_n856_), .Y(new_n1307_));
  INVX1    g0665(.A(new_n873_), .Y(new_n1308_));
  OAI21X1  g0666(.A0(new_n1308_), .A1(new_n1307_), .B0(new_n891_), .Y(new_n1309_));
  INVX1    g0667(.A(new_n927_), .Y(new_n1310_));
  AOI21X1  g0668(.A0(new_n908_), .A1(new_n1309_), .B0(new_n1310_), .Y(new_n1311_));
  INVX1    g0669(.A(new_n943_), .Y(new_n1312_));
  OAI21X1  g0670(.A0(new_n1312_), .A1(new_n1311_), .B0(new_n957_), .Y(new_n1313_));
  INVX1    g0671(.A(new_n993_), .Y(new_n1314_));
  AOI21X1  g0672(.A0(new_n974_), .A1(new_n1313_), .B0(new_n1314_), .Y(new_n1315_));
  INVX1    g0673(.A(new_n1001_), .Y(new_n1316_));
  OAI21X1  g0674(.A0(new_n1316_), .A1(new_n1315_), .B0(new_n1010_), .Y(new_n1317_));
  INVX1    g0675(.A(new_n1030_), .Y(new_n1318_));
  AOI21X1  g0676(.A0(new_n1019_), .A1(new_n1317_), .B0(new_n1318_), .Y(new_n1319_));
  INVX1    g0677(.A(new_n1038_), .Y(new_n1320_));
  OAI21X1  g0678(.A0(new_n1320_), .A1(new_n1319_), .B0(new_n1047_), .Y(new_n1321_));
  INVX1    g0679(.A(new_n1067_), .Y(new_n1322_));
  AOI21X1  g0680(.A0(new_n1056_), .A1(new_n1321_), .B0(new_n1322_), .Y(new_n1323_));
  INVX1    g0681(.A(new_n1075_), .Y(new_n1324_));
  OAI21X1  g0682(.A0(new_n1324_), .A1(new_n1323_), .B0(new_n1084_), .Y(new_n1325_));
  INVX1    g0683(.A(new_n1104_), .Y(new_n1326_));
  AOI21X1  g0684(.A0(new_n1093_), .A1(new_n1325_), .B0(new_n1326_), .Y(new_n1327_));
  INVX1    g0685(.A(new_n1112_), .Y(new_n1328_));
  OAI21X1  g0686(.A0(new_n1328_), .A1(new_n1327_), .B0(new_n1121_), .Y(new_n1329_));
  INVX1    g0687(.A(new_n1141_), .Y(new_n1330_));
  AOI21X1  g0688(.A0(new_n1130_), .A1(new_n1329_), .B0(new_n1330_), .Y(new_n1331_));
  INVX1    g0689(.A(new_n1149_), .Y(new_n1332_));
  OAI21X1  g0690(.A0(new_n1332_), .A1(new_n1331_), .B0(new_n1158_), .Y(new_n1333_));
  INVX1    g0691(.A(new_n1178_), .Y(new_n1334_));
  AOI21X1  g0692(.A0(new_n1167_), .A1(new_n1333_), .B0(new_n1334_), .Y(new_n1335_));
  INVX1    g0693(.A(new_n1186_), .Y(new_n1336_));
  OAI21X1  g0694(.A0(new_n1336_), .A1(new_n1335_), .B0(new_n1195_), .Y(new_n1337_));
  INVX1    g0695(.A(new_n1215_), .Y(new_n1338_));
  AOI21X1  g0696(.A0(new_n1204_), .A1(new_n1337_), .B0(new_n1338_), .Y(new_n1339_));
  INVX1    g0697(.A(new_n1223_), .Y(new_n1340_));
  OAI21X1  g0698(.A0(new_n1340_), .A1(new_n1339_), .B0(new_n1232_), .Y(new_n1341_));
  INVX1    g0699(.A(new_n1252_), .Y(new_n1342_));
  AOI21X1  g0700(.A0(new_n1241_), .A1(new_n1341_), .B0(new_n1342_), .Y(new_n1343_));
  INVX1    g0701(.A(new_n1260_), .Y(new_n1344_));
  OAI21X1  g0702(.A0(new_n1344_), .A1(new_n1343_), .B0(new_n1269_), .Y(new_n1345_));
  NOR2X1   g0703(.A(new_n1283_), .B(new_n1273_), .Y(new_n1346_));
  AOI21X1  g0704(.A0(new_n1279_), .A1(new_n1345_), .B0(new_n1346_), .Y(new_n1347_));
  INVX1    g0705(.A(new_n1286_), .Y(new_n1348_));
  AOI21X1  g0706(.A0(new_n1348_), .A1(new_n1347_), .B0(new_n705_), .Y(new_n1349_));
  NOR2X1   g0707(.A(new_n1349_), .B(new_n1287_), .Y(new_n1350_));
  INVX1    g0708(.A(\in2[127] ), .Y(new_n1351_));
  INVX1    g0709(.A(\in3[127] ), .Y(new_n1352_));
  INVX1    g0710(.A(\in2[31] ), .Y(new_n1353_));
  AND2X1   g0711(.A(\in3[31] ), .B(new_n1353_), .Y(new_n1354_));
  INVX1    g0712(.A(new_n1354_), .Y(new_n1355_));
  INVX1    g0713(.A(\in2[30] ), .Y(new_n1356_));
  AND2X1   g0714(.A(\in3[30] ), .B(new_n1356_), .Y(new_n1357_));
  INVX1    g0715(.A(\in2[29] ), .Y(new_n1358_));
  AND2X1   g0716(.A(\in3[29] ), .B(new_n1358_), .Y(new_n1359_));
  INVX1    g0717(.A(new_n1359_), .Y(new_n1360_));
  INVX1    g0718(.A(\in2[28] ), .Y(new_n1361_));
  AND2X1   g0719(.A(\in3[28] ), .B(new_n1361_), .Y(new_n1362_));
  INVX1    g0720(.A(\in2[27] ), .Y(new_n1363_));
  AND2X1   g0721(.A(\in3[27] ), .B(new_n1363_), .Y(new_n1364_));
  INVX1    g0722(.A(new_n1364_), .Y(new_n1365_));
  INVX1    g0723(.A(\in2[26] ), .Y(new_n1366_));
  AND2X1   g0724(.A(\in3[26] ), .B(new_n1366_), .Y(new_n1367_));
  INVX1    g0725(.A(\in3[25] ), .Y(new_n1368_));
  INVX1    g0726(.A(\in2[25] ), .Y(new_n1369_));
  INVX1    g0727(.A(\in3[24] ), .Y(new_n1370_));
  INVX1    g0728(.A(\in2[23] ), .Y(new_n1371_));
  AND2X1   g0729(.A(\in3[23] ), .B(new_n1371_), .Y(new_n1372_));
  INVX1    g0730(.A(\in2[22] ), .Y(new_n1373_));
  AND2X1   g0731(.A(\in3[22] ), .B(new_n1373_), .Y(new_n1374_));
  INVX1    g0732(.A(new_n1374_), .Y(new_n1375_));
  INVX1    g0733(.A(\in2[21] ), .Y(new_n1376_));
  AND2X1   g0734(.A(\in3[21] ), .B(new_n1376_), .Y(new_n1377_));
  INVX1    g0735(.A(\in2[20] ), .Y(new_n1378_));
  AND2X1   g0736(.A(\in3[20] ), .B(new_n1378_), .Y(new_n1379_));
  INVX1    g0737(.A(new_n1379_), .Y(new_n1380_));
  INVX1    g0738(.A(\in2[19] ), .Y(new_n1381_));
  AND2X1   g0739(.A(\in3[19] ), .B(new_n1381_), .Y(new_n1382_));
  INVX1    g0740(.A(\in2[18] ), .Y(new_n1383_));
  AND2X1   g0741(.A(\in3[18] ), .B(new_n1383_), .Y(new_n1384_));
  INVX1    g0742(.A(new_n1384_), .Y(new_n1385_));
  INVX1    g0743(.A(\in2[16] ), .Y(new_n1386_));
  INVX1    g0744(.A(\in2[15] ), .Y(new_n1387_));
  AND2X1   g0745(.A(\in3[15] ), .B(new_n1387_), .Y(new_n1388_));
  INVX1    g0746(.A(new_n1388_), .Y(new_n1389_));
  INVX1    g0747(.A(\in2[14] ), .Y(new_n1390_));
  AND2X1   g0748(.A(\in3[14] ), .B(new_n1390_), .Y(new_n1391_));
  INVX1    g0749(.A(\in2[13] ), .Y(new_n1392_));
  AND2X1   g0750(.A(\in3[13] ), .B(new_n1392_), .Y(new_n1393_));
  INVX1    g0751(.A(new_n1393_), .Y(new_n1394_));
  INVX1    g0752(.A(\in2[12] ), .Y(new_n1395_));
  AND2X1   g0753(.A(\in3[12] ), .B(new_n1395_), .Y(new_n1396_));
  INVX1    g0754(.A(\in2[11] ), .Y(new_n1397_));
  AND2X1   g0755(.A(\in3[11] ), .B(new_n1397_), .Y(new_n1398_));
  INVX1    g0756(.A(new_n1398_), .Y(new_n1399_));
  INVX1    g0757(.A(\in2[10] ), .Y(new_n1400_));
  AND2X1   g0758(.A(\in3[10] ), .B(new_n1400_), .Y(new_n1401_));
  INVX1    g0759(.A(\in3[9] ), .Y(new_n1402_));
  INVX1    g0760(.A(\in2[9] ), .Y(new_n1403_));
  INVX1    g0761(.A(\in3[8] ), .Y(new_n1404_));
  INVX1    g0762(.A(\in2[7] ), .Y(new_n1405_));
  AND2X1   g0763(.A(\in3[7] ), .B(new_n1405_), .Y(new_n1406_));
  INVX1    g0764(.A(\in2[6] ), .Y(new_n1407_));
  AND2X1   g0765(.A(\in3[6] ), .B(new_n1407_), .Y(new_n1408_));
  INVX1    g0766(.A(new_n1408_), .Y(new_n1409_));
  INVX1    g0767(.A(\in2[4] ), .Y(new_n1410_));
  INVX1    g0768(.A(\in2[3] ), .Y(new_n1411_));
  AND2X1   g0769(.A(\in3[3] ), .B(new_n1411_), .Y(new_n1412_));
  INVX1    g0770(.A(new_n1412_), .Y(new_n1413_));
  INVX1    g0771(.A(\in2[2] ), .Y(new_n1414_));
  INVX1    g0772(.A(\in3[1] ), .Y(new_n1415_));
  INVX1    g0773(.A(\in3[0] ), .Y(new_n1416_));
  AND2X1   g0774(.A(new_n1416_), .B(\in2[0] ), .Y(new_n1417_));
  AOI21X1  g0775(.A0(new_n1417_), .A1(\in2[1] ), .B0(new_n1415_), .Y(new_n1418_));
  INVX1    g0776(.A(\in3[2] ), .Y(new_n1419_));
  OAI22X1  g0777(.A0(new_n1417_), .A1(\in2[1] ), .B0(new_n1419_), .B1(\in2[2] ), .Y(new_n1420_));
  OAI22X1  g0778(.A0(new_n1420_), .A1(new_n1418_), .B0(\in3[2] ), .B1(new_n1414_), .Y(new_n1421_));
  INVX1    g0779(.A(\in3[3] ), .Y(new_n1422_));
  AND2X1   g0780(.A(new_n1422_), .B(\in2[3] ), .Y(new_n1423_));
  AOI21X1  g0781(.A0(new_n1421_), .A1(new_n1413_), .B0(new_n1423_), .Y(new_n1424_));
  AOI21X1  g0782(.A0(new_n1424_), .A1(new_n1410_), .B0(\in3[4] ), .Y(new_n1425_));
  INVX1    g0783(.A(\in2[1] ), .Y(new_n1426_));
  INVX1    g0784(.A(\in2[0] ), .Y(new_n1427_));
  OR2X1    g0785(.A(\in3[0] ), .B(new_n1427_), .Y(new_n1428_));
  OAI21X1  g0786(.A0(new_n1428_), .A1(new_n1426_), .B0(\in3[1] ), .Y(new_n1429_));
  AOI22X1  g0787(.A0(new_n1428_), .A1(new_n1426_), .B0(\in3[2] ), .B1(new_n1414_), .Y(new_n1430_));
  AOI22X1  g0788(.A0(new_n1430_), .A1(new_n1429_), .B0(new_n1419_), .B1(\in2[2] ), .Y(new_n1431_));
  INVX1    g0789(.A(new_n1423_), .Y(new_n1432_));
  OAI21X1  g0790(.A0(new_n1431_), .A1(new_n1412_), .B0(new_n1432_), .Y(new_n1433_));
  AND2X1   g0791(.A(new_n1433_), .B(\in2[4] ), .Y(new_n1434_));
  NOR3X1   g0792(.A(new_n1434_), .B(new_n1425_), .C(\in2[5] ), .Y(new_n1435_));
  OAI21X1  g0793(.A0(new_n1434_), .A1(new_n1425_), .B0(\in2[5] ), .Y(new_n1436_));
  OAI21X1  g0794(.A0(new_n1435_), .A1(\in3[5] ), .B0(new_n1436_), .Y(new_n1437_));
  INVX1    g0795(.A(\in3[6] ), .Y(new_n1438_));
  AND2X1   g0796(.A(new_n1438_), .B(\in2[6] ), .Y(new_n1439_));
  AOI21X1  g0797(.A0(new_n1437_), .A1(new_n1409_), .B0(new_n1439_), .Y(new_n1440_));
  INVX1    g0798(.A(\in3[7] ), .Y(new_n1441_));
  AND2X1   g0799(.A(new_n1441_), .B(\in2[7] ), .Y(new_n1442_));
  INVX1    g0800(.A(new_n1442_), .Y(new_n1443_));
  OAI21X1  g0801(.A0(new_n1440_), .A1(new_n1406_), .B0(new_n1443_), .Y(new_n1444_));
  OAI21X1  g0802(.A0(new_n1444_), .A1(\in2[8] ), .B0(new_n1404_), .Y(new_n1445_));
  INVX1    g0803(.A(\in2[8] ), .Y(new_n1446_));
  INVX1    g0804(.A(new_n1406_), .Y(new_n1447_));
  INVX1    g0805(.A(\in3[5] ), .Y(new_n1448_));
  INVX1    g0806(.A(\in2[5] ), .Y(new_n1449_));
  INVX1    g0807(.A(\in3[4] ), .Y(new_n1450_));
  OAI21X1  g0808(.A0(new_n1433_), .A1(\in2[4] ), .B0(new_n1450_), .Y(new_n1451_));
  OR2X1    g0809(.A(new_n1424_), .B(new_n1410_), .Y(new_n1452_));
  NAND3X1  g0810(.A(new_n1452_), .B(new_n1451_), .C(new_n1449_), .Y(new_n1453_));
  AOI21X1  g0811(.A0(new_n1452_), .A1(new_n1451_), .B0(new_n1449_), .Y(new_n1454_));
  AOI21X1  g0812(.A0(new_n1453_), .A1(new_n1448_), .B0(new_n1454_), .Y(new_n1455_));
  INVX1    g0813(.A(new_n1439_), .Y(new_n1456_));
  OAI21X1  g0814(.A0(new_n1455_), .A1(new_n1408_), .B0(new_n1456_), .Y(new_n1457_));
  AOI21X1  g0815(.A0(new_n1457_), .A1(new_n1447_), .B0(new_n1442_), .Y(new_n1458_));
  OR2X1    g0816(.A(new_n1458_), .B(new_n1446_), .Y(new_n1459_));
  NAND3X1  g0817(.A(new_n1459_), .B(new_n1445_), .C(new_n1403_), .Y(new_n1460_));
  AOI21X1  g0818(.A0(new_n1459_), .A1(new_n1445_), .B0(new_n1403_), .Y(new_n1461_));
  AOI21X1  g0819(.A0(new_n1460_), .A1(new_n1402_), .B0(new_n1461_), .Y(new_n1462_));
  INVX1    g0820(.A(\in3[10] ), .Y(new_n1463_));
  AND2X1   g0821(.A(new_n1463_), .B(\in2[10] ), .Y(new_n1464_));
  INVX1    g0822(.A(new_n1464_), .Y(new_n1465_));
  OAI21X1  g0823(.A0(new_n1462_), .A1(new_n1401_), .B0(new_n1465_), .Y(new_n1466_));
  INVX1    g0824(.A(\in3[11] ), .Y(new_n1467_));
  AND2X1   g0825(.A(new_n1467_), .B(\in2[11] ), .Y(new_n1468_));
  AOI21X1  g0826(.A0(new_n1466_), .A1(new_n1399_), .B0(new_n1468_), .Y(new_n1469_));
  INVX1    g0827(.A(\in3[12] ), .Y(new_n1470_));
  AND2X1   g0828(.A(new_n1470_), .B(\in2[12] ), .Y(new_n1471_));
  INVX1    g0829(.A(new_n1471_), .Y(new_n1472_));
  OAI21X1  g0830(.A0(new_n1469_), .A1(new_n1396_), .B0(new_n1472_), .Y(new_n1473_));
  INVX1    g0831(.A(\in3[13] ), .Y(new_n1474_));
  AND2X1   g0832(.A(new_n1474_), .B(\in2[13] ), .Y(new_n1475_));
  AOI21X1  g0833(.A0(new_n1473_), .A1(new_n1394_), .B0(new_n1475_), .Y(new_n1476_));
  INVX1    g0834(.A(\in3[14] ), .Y(new_n1477_));
  AND2X1   g0835(.A(new_n1477_), .B(\in2[14] ), .Y(new_n1478_));
  INVX1    g0836(.A(new_n1478_), .Y(new_n1479_));
  OAI21X1  g0837(.A0(new_n1476_), .A1(new_n1391_), .B0(new_n1479_), .Y(new_n1480_));
  INVX1    g0838(.A(\in3[15] ), .Y(new_n1481_));
  AND2X1   g0839(.A(new_n1481_), .B(\in2[15] ), .Y(new_n1482_));
  AOI21X1  g0840(.A0(new_n1480_), .A1(new_n1389_), .B0(new_n1482_), .Y(new_n1483_));
  AOI21X1  g0841(.A0(new_n1483_), .A1(new_n1386_), .B0(\in3[16] ), .Y(new_n1484_));
  INVX1    g0842(.A(new_n1391_), .Y(new_n1485_));
  INVX1    g0843(.A(new_n1396_), .Y(new_n1486_));
  INVX1    g0844(.A(new_n1401_), .Y(new_n1487_));
  AOI21X1  g0845(.A0(new_n1458_), .A1(new_n1446_), .B0(\in3[8] ), .Y(new_n1488_));
  AND2X1   g0846(.A(new_n1444_), .B(\in2[8] ), .Y(new_n1489_));
  NOR3X1   g0847(.A(new_n1489_), .B(new_n1488_), .C(\in2[9] ), .Y(new_n1490_));
  OAI21X1  g0848(.A0(new_n1489_), .A1(new_n1488_), .B0(\in2[9] ), .Y(new_n1491_));
  OAI21X1  g0849(.A0(new_n1490_), .A1(\in3[9] ), .B0(new_n1491_), .Y(new_n1492_));
  AOI21X1  g0850(.A0(new_n1492_), .A1(new_n1487_), .B0(new_n1464_), .Y(new_n1493_));
  INVX1    g0851(.A(new_n1468_), .Y(new_n1494_));
  OAI21X1  g0852(.A0(new_n1493_), .A1(new_n1398_), .B0(new_n1494_), .Y(new_n1495_));
  AOI21X1  g0853(.A0(new_n1495_), .A1(new_n1486_), .B0(new_n1471_), .Y(new_n1496_));
  INVX1    g0854(.A(new_n1475_), .Y(new_n1497_));
  OAI21X1  g0855(.A0(new_n1496_), .A1(new_n1393_), .B0(new_n1497_), .Y(new_n1498_));
  AOI21X1  g0856(.A0(new_n1498_), .A1(new_n1485_), .B0(new_n1478_), .Y(new_n1499_));
  INVX1    g0857(.A(new_n1482_), .Y(new_n1500_));
  OAI21X1  g0858(.A0(new_n1499_), .A1(new_n1388_), .B0(new_n1500_), .Y(new_n1501_));
  AND2X1   g0859(.A(new_n1501_), .B(\in2[16] ), .Y(new_n1502_));
  NOR3X1   g0860(.A(new_n1502_), .B(new_n1484_), .C(\in2[17] ), .Y(new_n1503_));
  OAI21X1  g0861(.A0(new_n1502_), .A1(new_n1484_), .B0(\in2[17] ), .Y(new_n1504_));
  OAI21X1  g0862(.A0(new_n1503_), .A1(\in3[17] ), .B0(new_n1504_), .Y(new_n1505_));
  INVX1    g0863(.A(\in3[18] ), .Y(new_n1506_));
  AND2X1   g0864(.A(new_n1506_), .B(\in2[18] ), .Y(new_n1507_));
  AOI21X1  g0865(.A0(new_n1505_), .A1(new_n1385_), .B0(new_n1507_), .Y(new_n1508_));
  INVX1    g0866(.A(\in3[19] ), .Y(new_n1509_));
  AND2X1   g0867(.A(new_n1509_), .B(\in2[19] ), .Y(new_n1510_));
  INVX1    g0868(.A(new_n1510_), .Y(new_n1511_));
  OAI21X1  g0869(.A0(new_n1508_), .A1(new_n1382_), .B0(new_n1511_), .Y(new_n1512_));
  INVX1    g0870(.A(\in3[20] ), .Y(new_n1513_));
  AND2X1   g0871(.A(new_n1513_), .B(\in2[20] ), .Y(new_n1514_));
  AOI21X1  g0872(.A0(new_n1512_), .A1(new_n1380_), .B0(new_n1514_), .Y(new_n1515_));
  INVX1    g0873(.A(\in3[21] ), .Y(new_n1516_));
  AND2X1   g0874(.A(new_n1516_), .B(\in2[21] ), .Y(new_n1517_));
  INVX1    g0875(.A(new_n1517_), .Y(new_n1518_));
  OAI21X1  g0876(.A0(new_n1515_), .A1(new_n1377_), .B0(new_n1518_), .Y(new_n1519_));
  INVX1    g0877(.A(\in3[22] ), .Y(new_n1520_));
  AND2X1   g0878(.A(new_n1520_), .B(\in2[22] ), .Y(new_n1521_));
  AOI21X1  g0879(.A0(new_n1519_), .A1(new_n1375_), .B0(new_n1521_), .Y(new_n1522_));
  INVX1    g0880(.A(\in3[23] ), .Y(new_n1523_));
  AND2X1   g0881(.A(new_n1523_), .B(\in2[23] ), .Y(new_n1524_));
  INVX1    g0882(.A(new_n1524_), .Y(new_n1525_));
  OAI21X1  g0883(.A0(new_n1522_), .A1(new_n1372_), .B0(new_n1525_), .Y(new_n1526_));
  OAI21X1  g0884(.A0(new_n1526_), .A1(\in2[24] ), .B0(new_n1370_), .Y(new_n1527_));
  INVX1    g0885(.A(\in2[24] ), .Y(new_n1528_));
  INVX1    g0886(.A(new_n1372_), .Y(new_n1529_));
  INVX1    g0887(.A(new_n1377_), .Y(new_n1530_));
  INVX1    g0888(.A(new_n1382_), .Y(new_n1531_));
  INVX1    g0889(.A(\in3[17] ), .Y(new_n1532_));
  INVX1    g0890(.A(\in2[17] ), .Y(new_n1533_));
  INVX1    g0891(.A(\in3[16] ), .Y(new_n1534_));
  OAI21X1  g0892(.A0(new_n1501_), .A1(\in2[16] ), .B0(new_n1534_), .Y(new_n1535_));
  OR2X1    g0893(.A(new_n1483_), .B(new_n1386_), .Y(new_n1536_));
  NAND3X1  g0894(.A(new_n1536_), .B(new_n1535_), .C(new_n1533_), .Y(new_n1537_));
  AOI21X1  g0895(.A0(new_n1536_), .A1(new_n1535_), .B0(new_n1533_), .Y(new_n1538_));
  AOI21X1  g0896(.A0(new_n1537_), .A1(new_n1532_), .B0(new_n1538_), .Y(new_n1539_));
  INVX1    g0897(.A(new_n1507_), .Y(new_n1540_));
  OAI21X1  g0898(.A0(new_n1539_), .A1(new_n1384_), .B0(new_n1540_), .Y(new_n1541_));
  AOI21X1  g0899(.A0(new_n1541_), .A1(new_n1531_), .B0(new_n1510_), .Y(new_n1542_));
  INVX1    g0900(.A(new_n1514_), .Y(new_n1543_));
  OAI21X1  g0901(.A0(new_n1542_), .A1(new_n1379_), .B0(new_n1543_), .Y(new_n1544_));
  AOI21X1  g0902(.A0(new_n1544_), .A1(new_n1530_), .B0(new_n1517_), .Y(new_n1545_));
  INVX1    g0903(.A(new_n1521_), .Y(new_n1546_));
  OAI21X1  g0904(.A0(new_n1545_), .A1(new_n1374_), .B0(new_n1546_), .Y(new_n1547_));
  AOI21X1  g0905(.A0(new_n1547_), .A1(new_n1529_), .B0(new_n1524_), .Y(new_n1548_));
  OR2X1    g0906(.A(new_n1548_), .B(new_n1528_), .Y(new_n1549_));
  NAND3X1  g0907(.A(new_n1549_), .B(new_n1527_), .C(new_n1369_), .Y(new_n1550_));
  AOI21X1  g0908(.A0(new_n1549_), .A1(new_n1527_), .B0(new_n1369_), .Y(new_n1551_));
  AOI21X1  g0909(.A0(new_n1550_), .A1(new_n1368_), .B0(new_n1551_), .Y(new_n1552_));
  INVX1    g0910(.A(\in3[26] ), .Y(new_n1553_));
  AND2X1   g0911(.A(new_n1553_), .B(\in2[26] ), .Y(new_n1554_));
  INVX1    g0912(.A(new_n1554_), .Y(new_n1555_));
  OAI21X1  g0913(.A0(new_n1552_), .A1(new_n1367_), .B0(new_n1555_), .Y(new_n1556_));
  INVX1    g0914(.A(\in3[27] ), .Y(new_n1557_));
  AND2X1   g0915(.A(new_n1557_), .B(\in2[27] ), .Y(new_n1558_));
  AOI21X1  g0916(.A0(new_n1556_), .A1(new_n1365_), .B0(new_n1558_), .Y(new_n1559_));
  INVX1    g0917(.A(\in3[28] ), .Y(new_n1560_));
  AND2X1   g0918(.A(new_n1560_), .B(\in2[28] ), .Y(new_n1561_));
  INVX1    g0919(.A(new_n1561_), .Y(new_n1562_));
  OAI21X1  g0920(.A0(new_n1559_), .A1(new_n1362_), .B0(new_n1562_), .Y(new_n1563_));
  INVX1    g0921(.A(\in3[29] ), .Y(new_n1564_));
  AND2X1   g0922(.A(new_n1564_), .B(\in2[29] ), .Y(new_n1565_));
  AOI21X1  g0923(.A0(new_n1563_), .A1(new_n1360_), .B0(new_n1565_), .Y(new_n1566_));
  INVX1    g0924(.A(\in3[30] ), .Y(new_n1567_));
  AND2X1   g0925(.A(new_n1567_), .B(\in2[30] ), .Y(new_n1568_));
  INVX1    g0926(.A(new_n1568_), .Y(new_n1569_));
  OAI21X1  g0927(.A0(new_n1566_), .A1(new_n1357_), .B0(new_n1569_), .Y(new_n1570_));
  INVX1    g0928(.A(\in3[31] ), .Y(new_n1571_));
  AND2X1   g0929(.A(new_n1571_), .B(\in2[31] ), .Y(new_n1572_));
  AOI21X1  g0930(.A0(new_n1570_), .A1(new_n1355_), .B0(new_n1572_), .Y(new_n1573_));
  INVX1    g0931(.A(\in2[38] ), .Y(new_n1574_));
  INVX1    g0932(.A(\in2[39] ), .Y(new_n1575_));
  AOI22X1  g0933(.A0(\in3[39] ), .A1(new_n1575_), .B0(\in3[38] ), .B1(new_n1574_), .Y(new_n1576_));
  INVX1    g0934(.A(new_n1576_), .Y(new_n1577_));
  INVX1    g0935(.A(\in3[36] ), .Y(new_n1578_));
  INVX1    g0936(.A(\in3[37] ), .Y(new_n1579_));
  OAI22X1  g0937(.A0(new_n1579_), .A1(\in2[37] ), .B0(new_n1578_), .B1(\in2[36] ), .Y(new_n1580_));
  INVX1    g0938(.A(\in2[34] ), .Y(new_n1581_));
  INVX1    g0939(.A(\in2[35] ), .Y(new_n1582_));
  AOI22X1  g0940(.A0(\in3[35] ), .A1(new_n1582_), .B0(\in3[34] ), .B1(new_n1581_), .Y(new_n1583_));
  INVX1    g0941(.A(new_n1583_), .Y(new_n1584_));
  INVX1    g0942(.A(\in3[32] ), .Y(new_n1585_));
  INVX1    g0943(.A(\in3[33] ), .Y(new_n1586_));
  OAI22X1  g0944(.A0(new_n1586_), .A1(\in2[33] ), .B0(new_n1585_), .B1(\in2[32] ), .Y(new_n1587_));
  NOR4X1   g0945(.A(new_n1587_), .B(new_n1584_), .C(new_n1580_), .D(new_n1577_), .Y(new_n1588_));
  INVX1    g0946(.A(new_n1588_), .Y(new_n1589_));
  NOR2X1   g0947(.A(new_n1580_), .B(new_n1577_), .Y(new_n1590_));
  AND2X1   g0948(.A(new_n1585_), .B(\in2[32] ), .Y(new_n1591_));
  OAI21X1  g0949(.A0(new_n1586_), .A1(\in2[33] ), .B0(new_n1591_), .Y(new_n1592_));
  INVX1    g0950(.A(\in3[34] ), .Y(new_n1593_));
  AOI22X1  g0951(.A0(new_n1593_), .A1(\in2[34] ), .B0(new_n1586_), .B1(\in2[33] ), .Y(new_n1594_));
  AND2X1   g0952(.A(new_n1594_), .B(new_n1592_), .Y(new_n1595_));
  OAI22X1  g0953(.A0(new_n1595_), .A1(new_n1584_), .B0(\in3[35] ), .B1(new_n1582_), .Y(new_n1596_));
  NOR2X1   g0954(.A(new_n1579_), .B(\in2[37] ), .Y(new_n1597_));
  NAND2X1  g0955(.A(new_n1578_), .B(\in2[36] ), .Y(new_n1598_));
  NOR2X1   g0956(.A(new_n1598_), .B(new_n1597_), .Y(new_n1599_));
  AOI21X1  g0957(.A0(new_n1579_), .A1(\in2[37] ), .B0(new_n1599_), .Y(new_n1600_));
  INVX1    g0958(.A(\in3[39] ), .Y(new_n1601_));
  AND2X1   g0959(.A(\in3[39] ), .B(new_n1575_), .Y(new_n1602_));
  NOR3X1   g0960(.A(new_n1602_), .B(\in3[38] ), .C(new_n1574_), .Y(new_n1603_));
  AOI21X1  g0961(.A0(new_n1601_), .A1(\in2[39] ), .B0(new_n1603_), .Y(new_n1604_));
  OAI21X1  g0962(.A0(new_n1600_), .A1(new_n1577_), .B0(new_n1604_), .Y(new_n1605_));
  AOI21X1  g0963(.A0(new_n1596_), .A1(new_n1590_), .B0(new_n1605_), .Y(new_n1606_));
  OAI21X1  g0964(.A0(new_n1589_), .A1(new_n1573_), .B0(new_n1606_), .Y(new_n1607_));
  INVX1    g0965(.A(\in2[46] ), .Y(new_n1608_));
  INVX1    g0966(.A(\in2[47] ), .Y(new_n1609_));
  AOI22X1  g0967(.A0(\in3[47] ), .A1(new_n1609_), .B0(\in3[46] ), .B1(new_n1608_), .Y(new_n1610_));
  INVX1    g0968(.A(new_n1610_), .Y(new_n1611_));
  INVX1    g0969(.A(\in3[44] ), .Y(new_n1612_));
  INVX1    g0970(.A(\in3[45] ), .Y(new_n1613_));
  OAI22X1  g0971(.A0(new_n1613_), .A1(\in2[45] ), .B0(new_n1612_), .B1(\in2[44] ), .Y(new_n1614_));
  INVX1    g0972(.A(\in2[42] ), .Y(new_n1615_));
  INVX1    g0973(.A(\in2[43] ), .Y(new_n1616_));
  AOI22X1  g0974(.A0(\in3[43] ), .A1(new_n1616_), .B0(\in3[42] ), .B1(new_n1615_), .Y(new_n1617_));
  INVX1    g0975(.A(new_n1617_), .Y(new_n1618_));
  INVX1    g0976(.A(\in3[40] ), .Y(new_n1619_));
  INVX1    g0977(.A(\in3[41] ), .Y(new_n1620_));
  OAI22X1  g0978(.A0(new_n1620_), .A1(\in2[41] ), .B0(new_n1619_), .B1(\in2[40] ), .Y(new_n1621_));
  NOR4X1   g0979(.A(new_n1621_), .B(new_n1618_), .C(new_n1614_), .D(new_n1611_), .Y(new_n1622_));
  NOR2X1   g0980(.A(new_n1614_), .B(new_n1611_), .Y(new_n1623_));
  AND2X1   g0981(.A(new_n1619_), .B(\in2[40] ), .Y(new_n1624_));
  OAI21X1  g0982(.A0(new_n1620_), .A1(\in2[41] ), .B0(new_n1624_), .Y(new_n1625_));
  INVX1    g0983(.A(\in3[42] ), .Y(new_n1626_));
  AOI22X1  g0984(.A0(new_n1626_), .A1(\in2[42] ), .B0(new_n1620_), .B1(\in2[41] ), .Y(new_n1627_));
  AND2X1   g0985(.A(new_n1627_), .B(new_n1625_), .Y(new_n1628_));
  OAI22X1  g0986(.A0(new_n1628_), .A1(new_n1618_), .B0(\in3[43] ), .B1(new_n1616_), .Y(new_n1629_));
  NOR2X1   g0987(.A(new_n1613_), .B(\in2[45] ), .Y(new_n1630_));
  NAND2X1  g0988(.A(new_n1612_), .B(\in2[44] ), .Y(new_n1631_));
  NOR2X1   g0989(.A(new_n1631_), .B(new_n1630_), .Y(new_n1632_));
  AOI21X1  g0990(.A0(new_n1613_), .A1(\in2[45] ), .B0(new_n1632_), .Y(new_n1633_));
  INVX1    g0991(.A(\in3[47] ), .Y(new_n1634_));
  AND2X1   g0992(.A(\in3[47] ), .B(new_n1609_), .Y(new_n1635_));
  NOR3X1   g0993(.A(new_n1635_), .B(\in3[46] ), .C(new_n1608_), .Y(new_n1636_));
  AOI21X1  g0994(.A0(new_n1634_), .A1(\in2[47] ), .B0(new_n1636_), .Y(new_n1637_));
  OAI21X1  g0995(.A0(new_n1633_), .A1(new_n1611_), .B0(new_n1637_), .Y(new_n1638_));
  AOI21X1  g0996(.A0(new_n1629_), .A1(new_n1623_), .B0(new_n1638_), .Y(new_n1639_));
  INVX1    g0997(.A(new_n1639_), .Y(new_n1640_));
  AOI21X1  g0998(.A0(new_n1622_), .A1(new_n1607_), .B0(new_n1640_), .Y(new_n1641_));
  INVX1    g0999(.A(\in2[54] ), .Y(new_n1642_));
  INVX1    g1000(.A(\in2[55] ), .Y(new_n1643_));
  AOI22X1  g1001(.A0(\in3[55] ), .A1(new_n1643_), .B0(\in3[54] ), .B1(new_n1642_), .Y(new_n1644_));
  INVX1    g1002(.A(new_n1644_), .Y(new_n1645_));
  INVX1    g1003(.A(\in3[52] ), .Y(new_n1646_));
  INVX1    g1004(.A(\in3[53] ), .Y(new_n1647_));
  OAI22X1  g1005(.A0(new_n1647_), .A1(\in2[53] ), .B0(new_n1646_), .B1(\in2[52] ), .Y(new_n1648_));
  INVX1    g1006(.A(\in2[50] ), .Y(new_n1649_));
  INVX1    g1007(.A(\in2[51] ), .Y(new_n1650_));
  AOI22X1  g1008(.A0(\in3[51] ), .A1(new_n1650_), .B0(\in3[50] ), .B1(new_n1649_), .Y(new_n1651_));
  INVX1    g1009(.A(new_n1651_), .Y(new_n1652_));
  INVX1    g1010(.A(\in3[48] ), .Y(new_n1653_));
  INVX1    g1011(.A(\in3[49] ), .Y(new_n1654_));
  OAI22X1  g1012(.A0(new_n1654_), .A1(\in2[49] ), .B0(new_n1653_), .B1(\in2[48] ), .Y(new_n1655_));
  NOR4X1   g1013(.A(new_n1655_), .B(new_n1652_), .C(new_n1648_), .D(new_n1645_), .Y(new_n1656_));
  INVX1    g1014(.A(new_n1656_), .Y(new_n1657_));
  NOR2X1   g1015(.A(new_n1648_), .B(new_n1645_), .Y(new_n1658_));
  AND2X1   g1016(.A(new_n1653_), .B(\in2[48] ), .Y(new_n1659_));
  OAI21X1  g1017(.A0(new_n1654_), .A1(\in2[49] ), .B0(new_n1659_), .Y(new_n1660_));
  INVX1    g1018(.A(\in3[50] ), .Y(new_n1661_));
  AOI22X1  g1019(.A0(new_n1661_), .A1(\in2[50] ), .B0(new_n1654_), .B1(\in2[49] ), .Y(new_n1662_));
  AND2X1   g1020(.A(new_n1662_), .B(new_n1660_), .Y(new_n1663_));
  OAI22X1  g1021(.A0(new_n1663_), .A1(new_n1652_), .B0(\in3[51] ), .B1(new_n1650_), .Y(new_n1664_));
  AND2X1   g1022(.A(new_n1646_), .B(\in2[52] ), .Y(new_n1665_));
  OAI21X1  g1023(.A0(new_n1647_), .A1(\in2[53] ), .B0(new_n1665_), .Y(new_n1666_));
  INVX1    g1024(.A(\in3[54] ), .Y(new_n1667_));
  AOI22X1  g1025(.A0(new_n1667_), .A1(\in2[54] ), .B0(new_n1647_), .B1(\in2[53] ), .Y(new_n1668_));
  AND2X1   g1026(.A(new_n1668_), .B(new_n1666_), .Y(new_n1669_));
  OAI22X1  g1027(.A0(new_n1669_), .A1(new_n1645_), .B0(\in3[55] ), .B1(new_n1643_), .Y(new_n1670_));
  AOI21X1  g1028(.A0(new_n1664_), .A1(new_n1658_), .B0(new_n1670_), .Y(new_n1671_));
  OAI21X1  g1029(.A0(new_n1657_), .A1(new_n1641_), .B0(new_n1671_), .Y(new_n1672_));
  INVX1    g1030(.A(\in2[62] ), .Y(new_n1673_));
  INVX1    g1031(.A(\in2[63] ), .Y(new_n1674_));
  AOI22X1  g1032(.A0(\in3[63] ), .A1(new_n1674_), .B0(\in3[62] ), .B1(new_n1673_), .Y(new_n1675_));
  INVX1    g1033(.A(new_n1675_), .Y(new_n1676_));
  INVX1    g1034(.A(\in3[60] ), .Y(new_n1677_));
  INVX1    g1035(.A(\in3[61] ), .Y(new_n1678_));
  OAI22X1  g1036(.A0(new_n1678_), .A1(\in2[61] ), .B0(new_n1677_), .B1(\in2[60] ), .Y(new_n1679_));
  INVX1    g1037(.A(\in2[58] ), .Y(new_n1680_));
  INVX1    g1038(.A(\in2[59] ), .Y(new_n1681_));
  AOI22X1  g1039(.A0(\in3[59] ), .A1(new_n1681_), .B0(\in3[58] ), .B1(new_n1680_), .Y(new_n1682_));
  INVX1    g1040(.A(new_n1682_), .Y(new_n1683_));
  INVX1    g1041(.A(\in3[56] ), .Y(new_n1684_));
  INVX1    g1042(.A(\in3[57] ), .Y(new_n1685_));
  OAI22X1  g1043(.A0(new_n1685_), .A1(\in2[57] ), .B0(new_n1684_), .B1(\in2[56] ), .Y(new_n1686_));
  NOR4X1   g1044(.A(new_n1686_), .B(new_n1683_), .C(new_n1679_), .D(new_n1676_), .Y(new_n1687_));
  NOR2X1   g1045(.A(new_n1679_), .B(new_n1676_), .Y(new_n1688_));
  AND2X1   g1046(.A(new_n1684_), .B(\in2[56] ), .Y(new_n1689_));
  OAI21X1  g1047(.A0(new_n1685_), .A1(\in2[57] ), .B0(new_n1689_), .Y(new_n1690_));
  INVX1    g1048(.A(\in3[58] ), .Y(new_n1691_));
  AOI22X1  g1049(.A0(new_n1691_), .A1(\in2[58] ), .B0(new_n1685_), .B1(\in2[57] ), .Y(new_n1692_));
  AND2X1   g1050(.A(new_n1692_), .B(new_n1690_), .Y(new_n1693_));
  OAI22X1  g1051(.A0(new_n1693_), .A1(new_n1683_), .B0(\in3[59] ), .B1(new_n1681_), .Y(new_n1694_));
  NOR2X1   g1052(.A(new_n1678_), .B(\in2[61] ), .Y(new_n1695_));
  NAND2X1  g1053(.A(new_n1677_), .B(\in2[60] ), .Y(new_n1696_));
  NOR2X1   g1054(.A(new_n1696_), .B(new_n1695_), .Y(new_n1697_));
  AOI21X1  g1055(.A0(new_n1678_), .A1(\in2[61] ), .B0(new_n1697_), .Y(new_n1698_));
  INVX1    g1056(.A(\in3[63] ), .Y(new_n1699_));
  AND2X1   g1057(.A(\in3[63] ), .B(new_n1674_), .Y(new_n1700_));
  NOR3X1   g1058(.A(new_n1700_), .B(\in3[62] ), .C(new_n1673_), .Y(new_n1701_));
  AOI21X1  g1059(.A0(new_n1699_), .A1(\in2[63] ), .B0(new_n1701_), .Y(new_n1702_));
  OAI21X1  g1060(.A0(new_n1698_), .A1(new_n1676_), .B0(new_n1702_), .Y(new_n1703_));
  AOI21X1  g1061(.A0(new_n1694_), .A1(new_n1688_), .B0(new_n1703_), .Y(new_n1704_));
  INVX1    g1062(.A(new_n1704_), .Y(new_n1705_));
  AOI21X1  g1063(.A0(new_n1687_), .A1(new_n1672_), .B0(new_n1705_), .Y(new_n1706_));
  INVX1    g1064(.A(\in2[66] ), .Y(new_n1707_));
  INVX1    g1065(.A(\in2[67] ), .Y(new_n1708_));
  AOI22X1  g1066(.A0(\in3[67] ), .A1(new_n1708_), .B0(\in3[66] ), .B1(new_n1707_), .Y(new_n1709_));
  INVX1    g1067(.A(\in2[64] ), .Y(new_n1710_));
  INVX1    g1068(.A(\in2[65] ), .Y(new_n1711_));
  AOI22X1  g1069(.A0(\in3[65] ), .A1(new_n1711_), .B0(\in3[64] ), .B1(new_n1710_), .Y(new_n1712_));
  AND2X1   g1070(.A(new_n1712_), .B(new_n1709_), .Y(new_n1713_));
  INVX1    g1071(.A(new_n1713_), .Y(new_n1714_));
  OR2X1    g1072(.A(\in3[67] ), .B(new_n1708_), .Y(new_n1715_));
  AND2X1   g1073(.A(\in3[65] ), .B(new_n1711_), .Y(new_n1716_));
  NOR3X1   g1074(.A(new_n1716_), .B(\in3[64] ), .C(new_n1710_), .Y(new_n1717_));
  INVX1    g1075(.A(\in3[65] ), .Y(new_n1718_));
  INVX1    g1076(.A(\in3[66] ), .Y(new_n1719_));
  AOI22X1  g1077(.A0(new_n1719_), .A1(\in2[66] ), .B0(new_n1718_), .B1(\in2[65] ), .Y(new_n1720_));
  INVX1    g1078(.A(new_n1720_), .Y(new_n1721_));
  OAI21X1  g1079(.A0(new_n1721_), .A1(new_n1717_), .B0(new_n1709_), .Y(new_n1722_));
  AND2X1   g1080(.A(new_n1722_), .B(new_n1715_), .Y(new_n1723_));
  OAI21X1  g1081(.A0(new_n1714_), .A1(new_n1706_), .B0(new_n1723_), .Y(new_n1724_));
  INVX1    g1082(.A(\in2[70] ), .Y(new_n1725_));
  INVX1    g1083(.A(\in2[71] ), .Y(new_n1726_));
  AOI22X1  g1084(.A0(\in3[71] ), .A1(new_n1726_), .B0(\in3[70] ), .B1(new_n1725_), .Y(new_n1727_));
  INVX1    g1085(.A(\in2[68] ), .Y(new_n1728_));
  INVX1    g1086(.A(\in2[69] ), .Y(new_n1729_));
  AOI22X1  g1087(.A0(\in3[69] ), .A1(new_n1729_), .B0(\in3[68] ), .B1(new_n1728_), .Y(new_n1730_));
  AND2X1   g1088(.A(new_n1730_), .B(new_n1727_), .Y(new_n1731_));
  AND2X1   g1089(.A(\in3[69] ), .B(new_n1729_), .Y(new_n1732_));
  NOR3X1   g1090(.A(new_n1732_), .B(\in3[68] ), .C(new_n1728_), .Y(new_n1733_));
  INVX1    g1091(.A(\in3[69] ), .Y(new_n1734_));
  AND2X1   g1092(.A(new_n1734_), .B(\in2[69] ), .Y(new_n1735_));
  OAI21X1  g1093(.A0(new_n1735_), .A1(new_n1733_), .B0(new_n1727_), .Y(new_n1736_));
  INVX1    g1094(.A(\in3[71] ), .Y(new_n1737_));
  AND2X1   g1095(.A(\in3[71] ), .B(new_n1726_), .Y(new_n1738_));
  NOR3X1   g1096(.A(new_n1738_), .B(\in3[70] ), .C(new_n1725_), .Y(new_n1739_));
  AOI21X1  g1097(.A0(new_n1737_), .A1(\in2[71] ), .B0(new_n1739_), .Y(new_n1740_));
  AND2X1   g1098(.A(new_n1740_), .B(new_n1736_), .Y(new_n1741_));
  INVX1    g1099(.A(new_n1741_), .Y(new_n1742_));
  AOI21X1  g1100(.A0(new_n1731_), .A1(new_n1724_), .B0(new_n1742_), .Y(new_n1743_));
  INVX1    g1101(.A(\in2[74] ), .Y(new_n1744_));
  INVX1    g1102(.A(\in2[75] ), .Y(new_n1745_));
  AOI22X1  g1103(.A0(\in3[75] ), .A1(new_n1745_), .B0(\in3[74] ), .B1(new_n1744_), .Y(new_n1746_));
  INVX1    g1104(.A(\in2[72] ), .Y(new_n1747_));
  INVX1    g1105(.A(\in2[73] ), .Y(new_n1748_));
  AOI22X1  g1106(.A0(\in3[73] ), .A1(new_n1748_), .B0(\in3[72] ), .B1(new_n1747_), .Y(new_n1749_));
  AND2X1   g1107(.A(new_n1749_), .B(new_n1746_), .Y(new_n1750_));
  INVX1    g1108(.A(new_n1750_), .Y(new_n1751_));
  OR2X1    g1109(.A(\in3[75] ), .B(new_n1745_), .Y(new_n1752_));
  AND2X1   g1110(.A(\in3[73] ), .B(new_n1748_), .Y(new_n1753_));
  NOR3X1   g1111(.A(new_n1753_), .B(\in3[72] ), .C(new_n1747_), .Y(new_n1754_));
  INVX1    g1112(.A(\in3[73] ), .Y(new_n1755_));
  INVX1    g1113(.A(\in3[74] ), .Y(new_n1756_));
  AOI22X1  g1114(.A0(new_n1756_), .A1(\in2[74] ), .B0(new_n1755_), .B1(\in2[73] ), .Y(new_n1757_));
  INVX1    g1115(.A(new_n1757_), .Y(new_n1758_));
  OAI21X1  g1116(.A0(new_n1758_), .A1(new_n1754_), .B0(new_n1746_), .Y(new_n1759_));
  AND2X1   g1117(.A(new_n1759_), .B(new_n1752_), .Y(new_n1760_));
  OAI21X1  g1118(.A0(new_n1751_), .A1(new_n1743_), .B0(new_n1760_), .Y(new_n1761_));
  INVX1    g1119(.A(\in2[78] ), .Y(new_n1762_));
  INVX1    g1120(.A(\in2[79] ), .Y(new_n1763_));
  AOI22X1  g1121(.A0(\in3[79] ), .A1(new_n1763_), .B0(\in3[78] ), .B1(new_n1762_), .Y(new_n1764_));
  INVX1    g1122(.A(\in2[76] ), .Y(new_n1765_));
  INVX1    g1123(.A(\in2[77] ), .Y(new_n1766_));
  AOI22X1  g1124(.A0(\in3[77] ), .A1(new_n1766_), .B0(\in3[76] ), .B1(new_n1765_), .Y(new_n1767_));
  AND2X1   g1125(.A(new_n1767_), .B(new_n1764_), .Y(new_n1768_));
  AND2X1   g1126(.A(\in3[77] ), .B(new_n1766_), .Y(new_n1769_));
  NOR3X1   g1127(.A(new_n1769_), .B(\in3[76] ), .C(new_n1765_), .Y(new_n1770_));
  INVX1    g1128(.A(\in3[77] ), .Y(new_n1771_));
  AND2X1   g1129(.A(new_n1771_), .B(\in2[77] ), .Y(new_n1772_));
  OAI21X1  g1130(.A0(new_n1772_), .A1(new_n1770_), .B0(new_n1764_), .Y(new_n1773_));
  INVX1    g1131(.A(\in3[79] ), .Y(new_n1774_));
  AND2X1   g1132(.A(\in3[79] ), .B(new_n1763_), .Y(new_n1775_));
  NOR3X1   g1133(.A(new_n1775_), .B(\in3[78] ), .C(new_n1762_), .Y(new_n1776_));
  AOI21X1  g1134(.A0(new_n1774_), .A1(\in2[79] ), .B0(new_n1776_), .Y(new_n1777_));
  AND2X1   g1135(.A(new_n1777_), .B(new_n1773_), .Y(new_n1778_));
  INVX1    g1136(.A(new_n1778_), .Y(new_n1779_));
  AOI21X1  g1137(.A0(new_n1768_), .A1(new_n1761_), .B0(new_n1779_), .Y(new_n1780_));
  INVX1    g1138(.A(\in2[82] ), .Y(new_n1781_));
  INVX1    g1139(.A(\in2[83] ), .Y(new_n1782_));
  AOI22X1  g1140(.A0(\in3[83] ), .A1(new_n1782_), .B0(\in3[82] ), .B1(new_n1781_), .Y(new_n1783_));
  INVX1    g1141(.A(\in2[80] ), .Y(new_n1784_));
  INVX1    g1142(.A(\in2[81] ), .Y(new_n1785_));
  AOI22X1  g1143(.A0(\in3[81] ), .A1(new_n1785_), .B0(\in3[80] ), .B1(new_n1784_), .Y(new_n1786_));
  AND2X1   g1144(.A(new_n1786_), .B(new_n1783_), .Y(new_n1787_));
  INVX1    g1145(.A(new_n1787_), .Y(new_n1788_));
  OR2X1    g1146(.A(\in3[83] ), .B(new_n1782_), .Y(new_n1789_));
  AND2X1   g1147(.A(\in3[81] ), .B(new_n1785_), .Y(new_n1790_));
  NOR3X1   g1148(.A(new_n1790_), .B(\in3[80] ), .C(new_n1784_), .Y(new_n1791_));
  INVX1    g1149(.A(\in3[81] ), .Y(new_n1792_));
  INVX1    g1150(.A(\in3[82] ), .Y(new_n1793_));
  AOI22X1  g1151(.A0(new_n1793_), .A1(\in2[82] ), .B0(new_n1792_), .B1(\in2[81] ), .Y(new_n1794_));
  INVX1    g1152(.A(new_n1794_), .Y(new_n1795_));
  OAI21X1  g1153(.A0(new_n1795_), .A1(new_n1791_), .B0(new_n1783_), .Y(new_n1796_));
  AND2X1   g1154(.A(new_n1796_), .B(new_n1789_), .Y(new_n1797_));
  OAI21X1  g1155(.A0(new_n1788_), .A1(new_n1780_), .B0(new_n1797_), .Y(new_n1798_));
  INVX1    g1156(.A(\in2[86] ), .Y(new_n1799_));
  INVX1    g1157(.A(\in2[87] ), .Y(new_n1800_));
  AOI22X1  g1158(.A0(\in3[87] ), .A1(new_n1800_), .B0(\in3[86] ), .B1(new_n1799_), .Y(new_n1801_));
  INVX1    g1159(.A(\in2[84] ), .Y(new_n1802_));
  INVX1    g1160(.A(\in2[85] ), .Y(new_n1803_));
  AOI22X1  g1161(.A0(\in3[85] ), .A1(new_n1803_), .B0(\in3[84] ), .B1(new_n1802_), .Y(new_n1804_));
  AND2X1   g1162(.A(new_n1804_), .B(new_n1801_), .Y(new_n1805_));
  AND2X1   g1163(.A(\in3[85] ), .B(new_n1803_), .Y(new_n1806_));
  NOR3X1   g1164(.A(new_n1806_), .B(\in3[84] ), .C(new_n1802_), .Y(new_n1807_));
  INVX1    g1165(.A(\in3[85] ), .Y(new_n1808_));
  AND2X1   g1166(.A(new_n1808_), .B(\in2[85] ), .Y(new_n1809_));
  OAI21X1  g1167(.A0(new_n1809_), .A1(new_n1807_), .B0(new_n1801_), .Y(new_n1810_));
  INVX1    g1168(.A(\in3[87] ), .Y(new_n1811_));
  AND2X1   g1169(.A(\in3[87] ), .B(new_n1800_), .Y(new_n1812_));
  NOR3X1   g1170(.A(new_n1812_), .B(\in3[86] ), .C(new_n1799_), .Y(new_n1813_));
  AOI21X1  g1171(.A0(new_n1811_), .A1(\in2[87] ), .B0(new_n1813_), .Y(new_n1814_));
  AND2X1   g1172(.A(new_n1814_), .B(new_n1810_), .Y(new_n1815_));
  INVX1    g1173(.A(new_n1815_), .Y(new_n1816_));
  AOI21X1  g1174(.A0(new_n1805_), .A1(new_n1798_), .B0(new_n1816_), .Y(new_n1817_));
  INVX1    g1175(.A(\in2[90] ), .Y(new_n1818_));
  INVX1    g1176(.A(\in2[91] ), .Y(new_n1819_));
  AOI22X1  g1177(.A0(\in3[91] ), .A1(new_n1819_), .B0(\in3[90] ), .B1(new_n1818_), .Y(new_n1820_));
  INVX1    g1178(.A(\in2[88] ), .Y(new_n1821_));
  INVX1    g1179(.A(\in2[89] ), .Y(new_n1822_));
  AOI22X1  g1180(.A0(\in3[89] ), .A1(new_n1822_), .B0(\in3[88] ), .B1(new_n1821_), .Y(new_n1823_));
  AND2X1   g1181(.A(new_n1823_), .B(new_n1820_), .Y(new_n1824_));
  INVX1    g1182(.A(new_n1824_), .Y(new_n1825_));
  OR2X1    g1183(.A(\in3[91] ), .B(new_n1819_), .Y(new_n1826_));
  AND2X1   g1184(.A(\in3[89] ), .B(new_n1822_), .Y(new_n1827_));
  NOR3X1   g1185(.A(new_n1827_), .B(\in3[88] ), .C(new_n1821_), .Y(new_n1828_));
  INVX1    g1186(.A(\in3[89] ), .Y(new_n1829_));
  INVX1    g1187(.A(\in3[90] ), .Y(new_n1830_));
  AOI22X1  g1188(.A0(new_n1830_), .A1(\in2[90] ), .B0(new_n1829_), .B1(\in2[89] ), .Y(new_n1831_));
  INVX1    g1189(.A(new_n1831_), .Y(new_n1832_));
  OAI21X1  g1190(.A0(new_n1832_), .A1(new_n1828_), .B0(new_n1820_), .Y(new_n1833_));
  AND2X1   g1191(.A(new_n1833_), .B(new_n1826_), .Y(new_n1834_));
  OAI21X1  g1192(.A0(new_n1825_), .A1(new_n1817_), .B0(new_n1834_), .Y(new_n1835_));
  INVX1    g1193(.A(\in2[94] ), .Y(new_n1836_));
  INVX1    g1194(.A(\in2[95] ), .Y(new_n1837_));
  AOI22X1  g1195(.A0(\in3[95] ), .A1(new_n1837_), .B0(\in3[94] ), .B1(new_n1836_), .Y(new_n1838_));
  INVX1    g1196(.A(\in2[92] ), .Y(new_n1839_));
  INVX1    g1197(.A(\in2[93] ), .Y(new_n1840_));
  AOI22X1  g1198(.A0(\in3[93] ), .A1(new_n1840_), .B0(\in3[92] ), .B1(new_n1839_), .Y(new_n1841_));
  AND2X1   g1199(.A(new_n1841_), .B(new_n1838_), .Y(new_n1842_));
  AND2X1   g1200(.A(\in3[93] ), .B(new_n1840_), .Y(new_n1843_));
  NOR3X1   g1201(.A(new_n1843_), .B(\in3[92] ), .C(new_n1839_), .Y(new_n1844_));
  INVX1    g1202(.A(\in3[93] ), .Y(new_n1845_));
  AND2X1   g1203(.A(new_n1845_), .B(\in2[93] ), .Y(new_n1846_));
  OAI21X1  g1204(.A0(new_n1846_), .A1(new_n1844_), .B0(new_n1838_), .Y(new_n1847_));
  INVX1    g1205(.A(\in3[95] ), .Y(new_n1848_));
  AND2X1   g1206(.A(\in3[95] ), .B(new_n1837_), .Y(new_n1849_));
  NOR3X1   g1207(.A(new_n1849_), .B(\in3[94] ), .C(new_n1836_), .Y(new_n1850_));
  AOI21X1  g1208(.A0(new_n1848_), .A1(\in2[95] ), .B0(new_n1850_), .Y(new_n1851_));
  AND2X1   g1209(.A(new_n1851_), .B(new_n1847_), .Y(new_n1852_));
  INVX1    g1210(.A(new_n1852_), .Y(new_n1853_));
  AOI21X1  g1211(.A0(new_n1842_), .A1(new_n1835_), .B0(new_n1853_), .Y(new_n1854_));
  INVX1    g1212(.A(\in2[98] ), .Y(new_n1855_));
  INVX1    g1213(.A(\in2[99] ), .Y(new_n1856_));
  AOI22X1  g1214(.A0(\in3[99] ), .A1(new_n1856_), .B0(\in3[98] ), .B1(new_n1855_), .Y(new_n1857_));
  INVX1    g1215(.A(\in2[96] ), .Y(new_n1858_));
  INVX1    g1216(.A(\in2[97] ), .Y(new_n1859_));
  AOI22X1  g1217(.A0(\in3[97] ), .A1(new_n1859_), .B0(\in3[96] ), .B1(new_n1858_), .Y(new_n1860_));
  AND2X1   g1218(.A(new_n1860_), .B(new_n1857_), .Y(new_n1861_));
  INVX1    g1219(.A(new_n1861_), .Y(new_n1862_));
  OR2X1    g1220(.A(\in3[99] ), .B(new_n1856_), .Y(new_n1863_));
  AND2X1   g1221(.A(\in3[97] ), .B(new_n1859_), .Y(new_n1864_));
  NOR3X1   g1222(.A(new_n1864_), .B(\in3[96] ), .C(new_n1858_), .Y(new_n1865_));
  INVX1    g1223(.A(\in3[97] ), .Y(new_n1866_));
  INVX1    g1224(.A(\in3[98] ), .Y(new_n1867_));
  AOI22X1  g1225(.A0(new_n1867_), .A1(\in2[98] ), .B0(new_n1866_), .B1(\in2[97] ), .Y(new_n1868_));
  INVX1    g1226(.A(new_n1868_), .Y(new_n1869_));
  OAI21X1  g1227(.A0(new_n1869_), .A1(new_n1865_), .B0(new_n1857_), .Y(new_n1870_));
  AND2X1   g1228(.A(new_n1870_), .B(new_n1863_), .Y(new_n1871_));
  OAI21X1  g1229(.A0(new_n1862_), .A1(new_n1854_), .B0(new_n1871_), .Y(new_n1872_));
  INVX1    g1230(.A(\in2[102] ), .Y(new_n1873_));
  INVX1    g1231(.A(\in2[103] ), .Y(new_n1874_));
  AOI22X1  g1232(.A0(\in3[103] ), .A1(new_n1874_), .B0(\in3[102] ), .B1(new_n1873_), .Y(new_n1875_));
  INVX1    g1233(.A(\in2[100] ), .Y(new_n1876_));
  INVX1    g1234(.A(\in2[101] ), .Y(new_n1877_));
  AOI22X1  g1235(.A0(\in3[101] ), .A1(new_n1877_), .B0(\in3[100] ), .B1(new_n1876_), .Y(new_n1878_));
  AND2X1   g1236(.A(new_n1878_), .B(new_n1875_), .Y(new_n1879_));
  AND2X1   g1237(.A(\in3[101] ), .B(new_n1877_), .Y(new_n1880_));
  NOR3X1   g1238(.A(new_n1880_), .B(\in3[100] ), .C(new_n1876_), .Y(new_n1881_));
  INVX1    g1239(.A(\in3[101] ), .Y(new_n1882_));
  AND2X1   g1240(.A(new_n1882_), .B(\in2[101] ), .Y(new_n1883_));
  OAI21X1  g1241(.A0(new_n1883_), .A1(new_n1881_), .B0(new_n1875_), .Y(new_n1884_));
  INVX1    g1242(.A(\in3[103] ), .Y(new_n1885_));
  AND2X1   g1243(.A(\in3[103] ), .B(new_n1874_), .Y(new_n1886_));
  NOR3X1   g1244(.A(new_n1886_), .B(\in3[102] ), .C(new_n1873_), .Y(new_n1887_));
  AOI21X1  g1245(.A0(new_n1885_), .A1(\in2[103] ), .B0(new_n1887_), .Y(new_n1888_));
  AND2X1   g1246(.A(new_n1888_), .B(new_n1884_), .Y(new_n1889_));
  INVX1    g1247(.A(new_n1889_), .Y(new_n1890_));
  AOI21X1  g1248(.A0(new_n1879_), .A1(new_n1872_), .B0(new_n1890_), .Y(new_n1891_));
  INVX1    g1249(.A(\in2[106] ), .Y(new_n1892_));
  INVX1    g1250(.A(\in2[107] ), .Y(new_n1893_));
  AOI22X1  g1251(.A0(\in3[107] ), .A1(new_n1893_), .B0(\in3[106] ), .B1(new_n1892_), .Y(new_n1894_));
  INVX1    g1252(.A(\in2[104] ), .Y(new_n1895_));
  INVX1    g1253(.A(\in2[105] ), .Y(new_n1896_));
  AOI22X1  g1254(.A0(\in3[105] ), .A1(new_n1896_), .B0(\in3[104] ), .B1(new_n1895_), .Y(new_n1897_));
  AND2X1   g1255(.A(new_n1897_), .B(new_n1894_), .Y(new_n1898_));
  INVX1    g1256(.A(new_n1898_), .Y(new_n1899_));
  OR2X1    g1257(.A(\in3[107] ), .B(new_n1893_), .Y(new_n1900_));
  AND2X1   g1258(.A(\in3[105] ), .B(new_n1896_), .Y(new_n1901_));
  NOR3X1   g1259(.A(new_n1901_), .B(\in3[104] ), .C(new_n1895_), .Y(new_n1902_));
  INVX1    g1260(.A(\in3[105] ), .Y(new_n1903_));
  INVX1    g1261(.A(\in3[106] ), .Y(new_n1904_));
  AOI22X1  g1262(.A0(new_n1904_), .A1(\in2[106] ), .B0(new_n1903_), .B1(\in2[105] ), .Y(new_n1905_));
  INVX1    g1263(.A(new_n1905_), .Y(new_n1906_));
  OAI21X1  g1264(.A0(new_n1906_), .A1(new_n1902_), .B0(new_n1894_), .Y(new_n1907_));
  AND2X1   g1265(.A(new_n1907_), .B(new_n1900_), .Y(new_n1908_));
  OAI21X1  g1266(.A0(new_n1899_), .A1(new_n1891_), .B0(new_n1908_), .Y(new_n1909_));
  INVX1    g1267(.A(\in2[110] ), .Y(new_n1910_));
  INVX1    g1268(.A(\in2[111] ), .Y(new_n1911_));
  AOI22X1  g1269(.A0(\in3[111] ), .A1(new_n1911_), .B0(\in3[110] ), .B1(new_n1910_), .Y(new_n1912_));
  INVX1    g1270(.A(\in2[108] ), .Y(new_n1913_));
  INVX1    g1271(.A(\in2[109] ), .Y(new_n1914_));
  AOI22X1  g1272(.A0(\in3[109] ), .A1(new_n1914_), .B0(\in3[108] ), .B1(new_n1913_), .Y(new_n1915_));
  AND2X1   g1273(.A(new_n1915_), .B(new_n1912_), .Y(new_n1916_));
  AND2X1   g1274(.A(\in3[109] ), .B(new_n1914_), .Y(new_n1917_));
  NOR3X1   g1275(.A(new_n1917_), .B(\in3[108] ), .C(new_n1913_), .Y(new_n1918_));
  INVX1    g1276(.A(\in3[109] ), .Y(new_n1919_));
  AND2X1   g1277(.A(new_n1919_), .B(\in2[109] ), .Y(new_n1920_));
  OAI21X1  g1278(.A0(new_n1920_), .A1(new_n1918_), .B0(new_n1912_), .Y(new_n1921_));
  INVX1    g1279(.A(\in3[111] ), .Y(new_n1922_));
  AND2X1   g1280(.A(\in3[111] ), .B(new_n1911_), .Y(new_n1923_));
  NOR3X1   g1281(.A(new_n1923_), .B(\in3[110] ), .C(new_n1910_), .Y(new_n1924_));
  AOI21X1  g1282(.A0(new_n1922_), .A1(\in2[111] ), .B0(new_n1924_), .Y(new_n1925_));
  AND2X1   g1283(.A(new_n1925_), .B(new_n1921_), .Y(new_n1926_));
  INVX1    g1284(.A(new_n1926_), .Y(new_n1927_));
  AOI21X1  g1285(.A0(new_n1916_), .A1(new_n1909_), .B0(new_n1927_), .Y(new_n1928_));
  INVX1    g1286(.A(\in2[114] ), .Y(new_n1929_));
  INVX1    g1287(.A(\in2[115] ), .Y(new_n1930_));
  AOI22X1  g1288(.A0(\in3[115] ), .A1(new_n1930_), .B0(\in3[114] ), .B1(new_n1929_), .Y(new_n1931_));
  INVX1    g1289(.A(\in2[112] ), .Y(new_n1932_));
  INVX1    g1290(.A(\in2[113] ), .Y(new_n1933_));
  AOI22X1  g1291(.A0(\in3[113] ), .A1(new_n1933_), .B0(\in3[112] ), .B1(new_n1932_), .Y(new_n1934_));
  AND2X1   g1292(.A(new_n1934_), .B(new_n1931_), .Y(new_n1935_));
  INVX1    g1293(.A(new_n1935_), .Y(new_n1936_));
  OR2X1    g1294(.A(\in3[115] ), .B(new_n1930_), .Y(new_n1937_));
  AND2X1   g1295(.A(\in3[113] ), .B(new_n1933_), .Y(new_n1938_));
  NOR3X1   g1296(.A(new_n1938_), .B(\in3[112] ), .C(new_n1932_), .Y(new_n1939_));
  INVX1    g1297(.A(\in3[113] ), .Y(new_n1940_));
  INVX1    g1298(.A(\in3[114] ), .Y(new_n1941_));
  AOI22X1  g1299(.A0(new_n1941_), .A1(\in2[114] ), .B0(new_n1940_), .B1(\in2[113] ), .Y(new_n1942_));
  INVX1    g1300(.A(new_n1942_), .Y(new_n1943_));
  OAI21X1  g1301(.A0(new_n1943_), .A1(new_n1939_), .B0(new_n1931_), .Y(new_n1944_));
  AND2X1   g1302(.A(new_n1944_), .B(new_n1937_), .Y(new_n1945_));
  OAI21X1  g1303(.A0(new_n1936_), .A1(new_n1928_), .B0(new_n1945_), .Y(new_n1946_));
  INVX1    g1304(.A(\in2[118] ), .Y(new_n1947_));
  INVX1    g1305(.A(\in2[119] ), .Y(new_n1948_));
  AOI22X1  g1306(.A0(\in3[119] ), .A1(new_n1948_), .B0(\in3[118] ), .B1(new_n1947_), .Y(new_n1949_));
  INVX1    g1307(.A(\in2[116] ), .Y(new_n1950_));
  INVX1    g1308(.A(\in2[117] ), .Y(new_n1951_));
  AOI22X1  g1309(.A0(\in3[117] ), .A1(new_n1951_), .B0(\in3[116] ), .B1(new_n1950_), .Y(new_n1952_));
  AND2X1   g1310(.A(new_n1952_), .B(new_n1949_), .Y(new_n1953_));
  AND2X1   g1311(.A(\in3[117] ), .B(new_n1951_), .Y(new_n1954_));
  NOR3X1   g1312(.A(new_n1954_), .B(\in3[116] ), .C(new_n1950_), .Y(new_n1955_));
  INVX1    g1313(.A(\in3[117] ), .Y(new_n1956_));
  AND2X1   g1314(.A(new_n1956_), .B(\in2[117] ), .Y(new_n1957_));
  OAI21X1  g1315(.A0(new_n1957_), .A1(new_n1955_), .B0(new_n1949_), .Y(new_n1958_));
  INVX1    g1316(.A(\in3[119] ), .Y(new_n1959_));
  AND2X1   g1317(.A(\in3[119] ), .B(new_n1948_), .Y(new_n1960_));
  NOR3X1   g1318(.A(new_n1960_), .B(\in3[118] ), .C(new_n1947_), .Y(new_n1961_));
  AOI21X1  g1319(.A0(new_n1959_), .A1(\in2[119] ), .B0(new_n1961_), .Y(new_n1962_));
  AND2X1   g1320(.A(new_n1962_), .B(new_n1958_), .Y(new_n1963_));
  INVX1    g1321(.A(new_n1963_), .Y(new_n1964_));
  AOI21X1  g1322(.A0(new_n1953_), .A1(new_n1946_), .B0(new_n1964_), .Y(new_n1965_));
  INVX1    g1323(.A(\in2[122] ), .Y(new_n1966_));
  INVX1    g1324(.A(\in2[123] ), .Y(new_n1967_));
  AOI22X1  g1325(.A0(\in3[123] ), .A1(new_n1967_), .B0(\in3[122] ), .B1(new_n1966_), .Y(new_n1968_));
  INVX1    g1326(.A(\in2[120] ), .Y(new_n1969_));
  INVX1    g1327(.A(\in2[121] ), .Y(new_n1970_));
  AOI22X1  g1328(.A0(\in3[121] ), .A1(new_n1970_), .B0(\in3[120] ), .B1(new_n1969_), .Y(new_n1971_));
  AND2X1   g1329(.A(new_n1971_), .B(new_n1968_), .Y(new_n1972_));
  INVX1    g1330(.A(new_n1972_), .Y(new_n1973_));
  OR2X1    g1331(.A(\in3[123] ), .B(new_n1967_), .Y(new_n1974_));
  AND2X1   g1332(.A(\in3[121] ), .B(new_n1970_), .Y(new_n1975_));
  NOR3X1   g1333(.A(new_n1975_), .B(\in3[120] ), .C(new_n1969_), .Y(new_n1976_));
  INVX1    g1334(.A(\in3[121] ), .Y(new_n1977_));
  INVX1    g1335(.A(\in3[122] ), .Y(new_n1978_));
  AOI22X1  g1336(.A0(new_n1978_), .A1(\in2[122] ), .B0(new_n1977_), .B1(\in2[121] ), .Y(new_n1979_));
  INVX1    g1337(.A(new_n1979_), .Y(new_n1980_));
  OAI21X1  g1338(.A0(new_n1980_), .A1(new_n1976_), .B0(new_n1968_), .Y(new_n1981_));
  AND2X1   g1339(.A(new_n1981_), .B(new_n1974_), .Y(new_n1982_));
  OAI21X1  g1340(.A0(new_n1973_), .A1(new_n1965_), .B0(new_n1982_), .Y(new_n1983_));
  INVX1    g1341(.A(\in2[125] ), .Y(new_n1984_));
  INVX1    g1342(.A(\in2[126] ), .Y(new_n1985_));
  AOI22X1  g1343(.A0(\in3[126] ), .A1(new_n1985_), .B0(\in3[125] ), .B1(new_n1984_), .Y(new_n1986_));
  INVX1    g1344(.A(\in2[124] ), .Y(new_n1987_));
  AOI22X1  g1345(.A0(new_n1352_), .A1(\in2[127] ), .B0(\in3[124] ), .B1(new_n1987_), .Y(new_n1988_));
  AND2X1   g1346(.A(new_n1988_), .B(new_n1986_), .Y(new_n1989_));
  AND2X1   g1347(.A(new_n1352_), .B(\in2[127] ), .Y(new_n1990_));
  INVX1    g1348(.A(\in3[126] ), .Y(new_n1991_));
  INVX1    g1349(.A(\in3[124] ), .Y(new_n1992_));
  INVX1    g1350(.A(\in3[125] ), .Y(new_n1993_));
  AOI22X1  g1351(.A0(new_n1993_), .A1(\in2[125] ), .B0(new_n1992_), .B1(\in2[124] ), .Y(new_n1994_));
  INVX1    g1352(.A(new_n1994_), .Y(new_n1995_));
  AOI22X1  g1353(.A0(new_n1995_), .A1(new_n1986_), .B0(new_n1991_), .B1(\in2[126] ), .Y(new_n1996_));
  NOR2X1   g1354(.A(new_n1996_), .B(new_n1990_), .Y(new_n1997_));
  AOI21X1  g1355(.A0(new_n1989_), .A1(new_n1983_), .B0(new_n1997_), .Y(new_n1998_));
  AOI21X1  g1356(.A0(new_n1998_), .A1(new_n1352_), .B0(new_n1351_), .Y(new_n1999_));
  OAI21X1  g1357(.A0(new_n1284_), .A1(\in1[127] ), .B0(\in0[127] ), .Y(new_n2000_));
  AND2X1   g1358(.A(new_n2000_), .B(new_n1999_), .Y(new_n2001_));
  NOR3X1   g1359(.A(new_n1286_), .B(new_n1284_), .C(new_n855_), .Y(new_n2002_));
  AOI21X1  g1360(.A0(new_n1348_), .A1(new_n1347_), .B0(new_n644_), .Y(new_n2003_));
  INVX1    g1361(.A(new_n1357_), .Y(new_n2004_));
  INVX1    g1362(.A(new_n1362_), .Y(new_n2005_));
  INVX1    g1363(.A(new_n1367_), .Y(new_n2006_));
  AOI21X1  g1364(.A0(new_n1548_), .A1(new_n1528_), .B0(\in3[24] ), .Y(new_n2007_));
  AND2X1   g1365(.A(new_n1526_), .B(\in2[24] ), .Y(new_n2008_));
  NOR3X1   g1366(.A(new_n2008_), .B(new_n2007_), .C(\in2[25] ), .Y(new_n2009_));
  OAI21X1  g1367(.A0(new_n2008_), .A1(new_n2007_), .B0(\in2[25] ), .Y(new_n2010_));
  OAI21X1  g1368(.A0(new_n2009_), .A1(\in3[25] ), .B0(new_n2010_), .Y(new_n2011_));
  AOI21X1  g1369(.A0(new_n2011_), .A1(new_n2006_), .B0(new_n1554_), .Y(new_n2012_));
  INVX1    g1370(.A(new_n1558_), .Y(new_n2013_));
  OAI21X1  g1371(.A0(new_n2012_), .A1(new_n1364_), .B0(new_n2013_), .Y(new_n2014_));
  AOI21X1  g1372(.A0(new_n2014_), .A1(new_n2005_), .B0(new_n1561_), .Y(new_n2015_));
  INVX1    g1373(.A(new_n1565_), .Y(new_n2016_));
  OAI21X1  g1374(.A0(new_n2015_), .A1(new_n1359_), .B0(new_n2016_), .Y(new_n2017_));
  AOI21X1  g1375(.A0(new_n2017_), .A1(new_n2004_), .B0(new_n1568_), .Y(new_n2018_));
  INVX1    g1376(.A(new_n1572_), .Y(new_n2019_));
  OAI21X1  g1377(.A0(new_n2018_), .A1(new_n1354_), .B0(new_n2019_), .Y(new_n2020_));
  INVX1    g1378(.A(new_n1606_), .Y(new_n2021_));
  AOI21X1  g1379(.A0(new_n1588_), .A1(new_n2020_), .B0(new_n2021_), .Y(new_n2022_));
  INVX1    g1380(.A(new_n1622_), .Y(new_n2023_));
  OAI21X1  g1381(.A0(new_n2023_), .A1(new_n2022_), .B0(new_n1639_), .Y(new_n2024_));
  INVX1    g1382(.A(new_n1671_), .Y(new_n2025_));
  AOI21X1  g1383(.A0(new_n1656_), .A1(new_n2024_), .B0(new_n2025_), .Y(new_n2026_));
  INVX1    g1384(.A(new_n1687_), .Y(new_n2027_));
  OAI21X1  g1385(.A0(new_n2027_), .A1(new_n2026_), .B0(new_n1704_), .Y(new_n2028_));
  INVX1    g1386(.A(new_n1723_), .Y(new_n2029_));
  AOI21X1  g1387(.A0(new_n1713_), .A1(new_n2028_), .B0(new_n2029_), .Y(new_n2030_));
  INVX1    g1388(.A(new_n1731_), .Y(new_n2031_));
  OAI21X1  g1389(.A0(new_n2031_), .A1(new_n2030_), .B0(new_n1741_), .Y(new_n2032_));
  INVX1    g1390(.A(new_n1760_), .Y(new_n2033_));
  AOI21X1  g1391(.A0(new_n1750_), .A1(new_n2032_), .B0(new_n2033_), .Y(new_n2034_));
  INVX1    g1392(.A(new_n1768_), .Y(new_n2035_));
  OAI21X1  g1393(.A0(new_n2035_), .A1(new_n2034_), .B0(new_n1778_), .Y(new_n2036_));
  INVX1    g1394(.A(new_n1797_), .Y(new_n2037_));
  AOI21X1  g1395(.A0(new_n1787_), .A1(new_n2036_), .B0(new_n2037_), .Y(new_n2038_));
  INVX1    g1396(.A(new_n1805_), .Y(new_n2039_));
  OAI21X1  g1397(.A0(new_n2039_), .A1(new_n2038_), .B0(new_n1815_), .Y(new_n2040_));
  INVX1    g1398(.A(new_n1834_), .Y(new_n2041_));
  AOI21X1  g1399(.A0(new_n1824_), .A1(new_n2040_), .B0(new_n2041_), .Y(new_n2042_));
  INVX1    g1400(.A(new_n1842_), .Y(new_n2043_));
  OAI21X1  g1401(.A0(new_n2043_), .A1(new_n2042_), .B0(new_n1852_), .Y(new_n2044_));
  INVX1    g1402(.A(new_n1871_), .Y(new_n2045_));
  AOI21X1  g1403(.A0(new_n1861_), .A1(new_n2044_), .B0(new_n2045_), .Y(new_n2046_));
  INVX1    g1404(.A(new_n1879_), .Y(new_n2047_));
  OAI21X1  g1405(.A0(new_n2047_), .A1(new_n2046_), .B0(new_n1889_), .Y(new_n2048_));
  INVX1    g1406(.A(new_n1908_), .Y(new_n2049_));
  AOI21X1  g1407(.A0(new_n1898_), .A1(new_n2048_), .B0(new_n2049_), .Y(new_n2050_));
  INVX1    g1408(.A(new_n1916_), .Y(new_n2051_));
  OAI21X1  g1409(.A0(new_n2051_), .A1(new_n2050_), .B0(new_n1926_), .Y(new_n2052_));
  INVX1    g1410(.A(new_n1945_), .Y(new_n2053_));
  AOI21X1  g1411(.A0(new_n1935_), .A1(new_n2052_), .B0(new_n2053_), .Y(new_n2054_));
  INVX1    g1412(.A(new_n1953_), .Y(new_n2055_));
  OAI21X1  g1413(.A0(new_n2055_), .A1(new_n2054_), .B0(new_n1963_), .Y(new_n2056_));
  INVX1    g1414(.A(new_n1982_), .Y(new_n2057_));
  AOI21X1  g1415(.A0(new_n1972_), .A1(new_n2056_), .B0(new_n2057_), .Y(new_n2058_));
  INVX1    g1416(.A(new_n1989_), .Y(new_n2059_));
  OAI22X1  g1417(.A0(new_n1996_), .A1(new_n1990_), .B0(new_n2059_), .B1(new_n2058_), .Y(new_n2060_));
  AND2X1   g1418(.A(\in3[127] ), .B(new_n1351_), .Y(new_n2061_));
  NOR3X1   g1419(.A(new_n2061_), .B(new_n2060_), .C(new_n1571_), .Y(new_n2062_));
  INVX1    g1420(.A(new_n2061_), .Y(new_n2063_));
  AOI21X1  g1421(.A0(new_n2063_), .A1(new_n1998_), .B0(new_n1353_), .Y(new_n2064_));
  NOR2X1   g1422(.A(new_n2064_), .B(new_n2062_), .Y(new_n2065_));
  NOR3X1   g1423(.A(new_n2065_), .B(new_n2003_), .C(new_n2002_), .Y(new_n2066_));
  NOR3X1   g1424(.A(new_n1286_), .B(new_n1284_), .C(new_n852_), .Y(new_n2067_));
  AOI21X1  g1425(.A0(new_n1348_), .A1(new_n1347_), .B0(new_n646_), .Y(new_n2068_));
  NOR2X1   g1426(.A(new_n2068_), .B(new_n2067_), .Y(new_n2069_));
  INVX1    g1427(.A(new_n2069_), .Y(new_n2070_));
  OR2X1    g1428(.A(new_n2061_), .B(new_n2060_), .Y(new_n2071_));
  NOR3X1   g1429(.A(new_n2061_), .B(new_n2060_), .C(new_n1567_), .Y(new_n2072_));
  AOI21X1  g1430(.A0(new_n2071_), .A1(\in2[30] ), .B0(new_n2072_), .Y(new_n2073_));
  NOR3X1   g1431(.A(new_n1286_), .B(new_n1284_), .C(new_n848_), .Y(new_n2074_));
  AOI21X1  g1432(.A0(new_n1348_), .A1(new_n1347_), .B0(new_n649_), .Y(new_n2075_));
  NOR3X1   g1433(.A(new_n2061_), .B(new_n2060_), .C(new_n1564_), .Y(new_n2076_));
  AOI21X1  g1434(.A0(new_n2063_), .A1(new_n1998_), .B0(new_n1358_), .Y(new_n2077_));
  NOR2X1   g1435(.A(new_n2077_), .B(new_n2076_), .Y(new_n2078_));
  NOR3X1   g1436(.A(new_n2078_), .B(new_n2075_), .C(new_n2074_), .Y(new_n2079_));
  NOR3X1   g1437(.A(new_n1286_), .B(new_n1284_), .C(new_n845_), .Y(new_n2080_));
  AOI21X1  g1438(.A0(new_n1348_), .A1(new_n1347_), .B0(new_n651_), .Y(new_n2081_));
  NOR2X1   g1439(.A(new_n2081_), .B(new_n2080_), .Y(new_n2082_));
  INVX1    g1440(.A(new_n2082_), .Y(new_n2083_));
  NOR3X1   g1441(.A(new_n2061_), .B(new_n2060_), .C(new_n1560_), .Y(new_n2084_));
  AOI21X1  g1442(.A0(new_n2071_), .A1(\in2[28] ), .B0(new_n2084_), .Y(new_n2085_));
  NOR3X1   g1443(.A(new_n1286_), .B(new_n1284_), .C(new_n841_), .Y(new_n2086_));
  AOI21X1  g1444(.A0(new_n1348_), .A1(new_n1347_), .B0(new_n654_), .Y(new_n2087_));
  NOR3X1   g1445(.A(new_n2061_), .B(new_n2060_), .C(new_n1557_), .Y(new_n2088_));
  AOI21X1  g1446(.A0(new_n2063_), .A1(new_n1998_), .B0(new_n1363_), .Y(new_n2089_));
  NOR2X1   g1447(.A(new_n2089_), .B(new_n2088_), .Y(new_n2090_));
  NOR3X1   g1448(.A(new_n2090_), .B(new_n2087_), .C(new_n2086_), .Y(new_n2091_));
  NOR3X1   g1449(.A(new_n1286_), .B(new_n1284_), .C(new_n838_), .Y(new_n2092_));
  AOI21X1  g1450(.A0(new_n1348_), .A1(new_n1347_), .B0(new_n656_), .Y(new_n2093_));
  NOR2X1   g1451(.A(new_n2093_), .B(new_n2092_), .Y(new_n2094_));
  INVX1    g1452(.A(new_n2094_), .Y(new_n2095_));
  NOR3X1   g1453(.A(new_n2061_), .B(new_n2060_), .C(new_n1553_), .Y(new_n2096_));
  AOI21X1  g1454(.A0(new_n2071_), .A1(\in2[26] ), .B0(new_n2096_), .Y(new_n2097_));
  NOR3X1   g1455(.A(new_n2061_), .B(new_n2060_), .C(new_n1368_), .Y(new_n2098_));
  AOI21X1  g1456(.A0(new_n2063_), .A1(new_n1998_), .B0(new_n1369_), .Y(new_n2099_));
  NOR2X1   g1457(.A(new_n2099_), .B(new_n2098_), .Y(new_n2100_));
  INVX1    g1458(.A(new_n2100_), .Y(new_n2101_));
  NOR3X1   g1459(.A(new_n2061_), .B(new_n2060_), .C(new_n1370_), .Y(new_n2102_));
  AOI21X1  g1460(.A0(new_n2071_), .A1(\in2[24] ), .B0(new_n2102_), .Y(new_n2103_));
  NOR3X1   g1461(.A(new_n1286_), .B(new_n1284_), .C(new_n813_), .Y(new_n2104_));
  AOI21X1  g1462(.A0(new_n1348_), .A1(new_n1347_), .B0(new_n660_), .Y(new_n2105_));
  NOR2X1   g1463(.A(new_n2105_), .B(new_n2104_), .Y(new_n2106_));
  NOR3X1   g1464(.A(new_n2061_), .B(new_n2060_), .C(new_n1523_), .Y(new_n2107_));
  AOI21X1  g1465(.A0(new_n2063_), .A1(new_n1998_), .B0(new_n1371_), .Y(new_n2108_));
  OAI21X1  g1466(.A0(new_n2108_), .A1(new_n2107_), .B0(new_n2106_), .Y(new_n2109_));
  NOR3X1   g1467(.A(new_n1286_), .B(new_n1284_), .C(new_n809_), .Y(new_n2110_));
  AOI21X1  g1468(.A0(new_n1348_), .A1(new_n1347_), .B0(new_n663_), .Y(new_n2111_));
  NOR3X1   g1469(.A(new_n2061_), .B(new_n2060_), .C(new_n1520_), .Y(new_n2112_));
  AOI21X1  g1470(.A0(new_n2063_), .A1(new_n1998_), .B0(new_n1373_), .Y(new_n2113_));
  NOR2X1   g1471(.A(new_n2113_), .B(new_n2112_), .Y(new_n2114_));
  NOR3X1   g1472(.A(new_n2114_), .B(new_n2111_), .C(new_n2110_), .Y(new_n2115_));
  NOR3X1   g1473(.A(new_n1286_), .B(new_n1284_), .C(new_n806_), .Y(new_n2116_));
  AOI21X1  g1474(.A0(new_n1348_), .A1(new_n1347_), .B0(new_n665_), .Y(new_n2117_));
  NOR2X1   g1475(.A(new_n2117_), .B(new_n2116_), .Y(new_n2118_));
  NOR3X1   g1476(.A(new_n2061_), .B(new_n2060_), .C(new_n1516_), .Y(new_n2119_));
  AOI21X1  g1477(.A0(new_n2063_), .A1(new_n1998_), .B0(new_n1376_), .Y(new_n2120_));
  OAI21X1  g1478(.A0(new_n2120_), .A1(new_n2119_), .B0(new_n2118_), .Y(new_n2121_));
  NOR3X1   g1479(.A(new_n1286_), .B(new_n1284_), .C(new_n802_), .Y(new_n2122_));
  AOI21X1  g1480(.A0(new_n1348_), .A1(new_n1347_), .B0(new_n668_), .Y(new_n2123_));
  NOR3X1   g1481(.A(new_n2061_), .B(new_n2060_), .C(new_n1513_), .Y(new_n2124_));
  AOI21X1  g1482(.A0(new_n2063_), .A1(new_n1998_), .B0(new_n1378_), .Y(new_n2125_));
  NOR2X1   g1483(.A(new_n2125_), .B(new_n2124_), .Y(new_n2126_));
  NOR3X1   g1484(.A(new_n2126_), .B(new_n2123_), .C(new_n2122_), .Y(new_n2127_));
  NOR3X1   g1485(.A(new_n1286_), .B(new_n1284_), .C(new_n799_), .Y(new_n2128_));
  AOI21X1  g1486(.A0(new_n1348_), .A1(new_n1347_), .B0(new_n670_), .Y(new_n2129_));
  NOR2X1   g1487(.A(new_n2129_), .B(new_n2128_), .Y(new_n2130_));
  NOR3X1   g1488(.A(new_n2061_), .B(new_n2060_), .C(new_n1509_), .Y(new_n2131_));
  AOI21X1  g1489(.A0(new_n2063_), .A1(new_n1998_), .B0(new_n1381_), .Y(new_n2132_));
  OAI21X1  g1490(.A0(new_n2132_), .A1(new_n2131_), .B0(new_n2130_), .Y(new_n2133_));
  NOR3X1   g1491(.A(new_n1286_), .B(new_n1284_), .C(new_n795_), .Y(new_n2134_));
  AOI21X1  g1492(.A0(new_n1348_), .A1(new_n1347_), .B0(new_n673_), .Y(new_n2135_));
  NOR3X1   g1493(.A(new_n2061_), .B(new_n2060_), .C(new_n1506_), .Y(new_n2136_));
  AOI21X1  g1494(.A0(new_n2063_), .A1(new_n1998_), .B0(new_n1383_), .Y(new_n2137_));
  NOR2X1   g1495(.A(new_n2137_), .B(new_n2136_), .Y(new_n2138_));
  NOR3X1   g1496(.A(new_n2138_), .B(new_n2135_), .C(new_n2134_), .Y(new_n2139_));
  NOR3X1   g1497(.A(new_n2061_), .B(new_n2060_), .C(new_n1532_), .Y(new_n2140_));
  AOI21X1  g1498(.A0(new_n2071_), .A1(\in2[17] ), .B0(new_n2140_), .Y(new_n2141_));
  NOR3X1   g1499(.A(new_n2061_), .B(new_n2060_), .C(new_n1534_), .Y(new_n2142_));
  AOI21X1  g1500(.A0(new_n2063_), .A1(new_n1998_), .B0(new_n1386_), .Y(new_n2143_));
  NOR2X1   g1501(.A(new_n2143_), .B(new_n2142_), .Y(new_n2144_));
  INVX1    g1502(.A(new_n2144_), .Y(new_n2145_));
  NOR3X1   g1503(.A(new_n1286_), .B(new_n1284_), .C(new_n765_), .Y(new_n2146_));
  AOI21X1  g1504(.A0(new_n1348_), .A1(new_n1347_), .B0(new_n678_), .Y(new_n2147_));
  NOR2X1   g1505(.A(new_n2147_), .B(new_n2146_), .Y(new_n2148_));
  INVX1    g1506(.A(new_n2148_), .Y(new_n2149_));
  NOR3X1   g1507(.A(new_n2061_), .B(new_n2060_), .C(new_n1481_), .Y(new_n2150_));
  AOI21X1  g1508(.A0(new_n2063_), .A1(new_n1998_), .B0(new_n1387_), .Y(new_n2151_));
  NOR2X1   g1509(.A(new_n2151_), .B(new_n2150_), .Y(new_n2152_));
  NOR2X1   g1510(.A(new_n2152_), .B(new_n2149_), .Y(new_n2153_));
  NOR3X1   g1511(.A(new_n1286_), .B(new_n1284_), .C(new_n762_), .Y(new_n2154_));
  AOI21X1  g1512(.A0(new_n1348_), .A1(new_n1347_), .B0(new_n680_), .Y(new_n2155_));
  NOR2X1   g1513(.A(new_n2155_), .B(new_n2154_), .Y(new_n2156_));
  INVX1    g1514(.A(new_n2156_), .Y(new_n2157_));
  NOR3X1   g1515(.A(new_n2061_), .B(new_n2060_), .C(new_n1477_), .Y(new_n2158_));
  AOI21X1  g1516(.A0(new_n2063_), .A1(new_n1998_), .B0(new_n1390_), .Y(new_n2159_));
  NOR2X1   g1517(.A(new_n2159_), .B(new_n2158_), .Y(new_n2160_));
  NOR3X1   g1518(.A(new_n1286_), .B(new_n1284_), .C(new_n758_), .Y(new_n2161_));
  AOI21X1  g1519(.A0(new_n1348_), .A1(new_n1347_), .B0(new_n683_), .Y(new_n2162_));
  NOR2X1   g1520(.A(new_n2162_), .B(new_n2161_), .Y(new_n2163_));
  INVX1    g1521(.A(new_n2163_), .Y(new_n2164_));
  NOR3X1   g1522(.A(new_n2061_), .B(new_n2060_), .C(new_n1474_), .Y(new_n2165_));
  AOI21X1  g1523(.A0(new_n2063_), .A1(new_n1998_), .B0(new_n1392_), .Y(new_n2166_));
  NOR2X1   g1524(.A(new_n2166_), .B(new_n2165_), .Y(new_n2167_));
  NOR2X1   g1525(.A(new_n2167_), .B(new_n2164_), .Y(new_n2168_));
  NOR3X1   g1526(.A(new_n1286_), .B(new_n1284_), .C(new_n755_), .Y(new_n2169_));
  AOI21X1  g1527(.A0(new_n1348_), .A1(new_n1347_), .B0(new_n685_), .Y(new_n2170_));
  NOR2X1   g1528(.A(new_n2170_), .B(new_n2169_), .Y(new_n2171_));
  INVX1    g1529(.A(new_n2171_), .Y(new_n2172_));
  NOR3X1   g1530(.A(new_n2061_), .B(new_n2060_), .C(new_n1470_), .Y(new_n2173_));
  AOI21X1  g1531(.A0(new_n2063_), .A1(new_n1998_), .B0(new_n1395_), .Y(new_n2174_));
  NOR2X1   g1532(.A(new_n2174_), .B(new_n2173_), .Y(new_n2175_));
  NOR3X1   g1533(.A(new_n1286_), .B(new_n1284_), .C(new_n751_), .Y(new_n2176_));
  AOI21X1  g1534(.A0(new_n1348_), .A1(new_n1347_), .B0(new_n688_), .Y(new_n2177_));
  NOR2X1   g1535(.A(new_n2177_), .B(new_n2176_), .Y(new_n2178_));
  INVX1    g1536(.A(new_n2178_), .Y(new_n2179_));
  NOR3X1   g1537(.A(new_n2061_), .B(new_n2060_), .C(new_n1467_), .Y(new_n2180_));
  AOI21X1  g1538(.A0(new_n2063_), .A1(new_n1998_), .B0(new_n1397_), .Y(new_n2181_));
  NOR2X1   g1539(.A(new_n2181_), .B(new_n2180_), .Y(new_n2182_));
  NOR2X1   g1540(.A(new_n2182_), .B(new_n2179_), .Y(new_n2183_));
  NOR3X1   g1541(.A(new_n1286_), .B(new_n1284_), .C(new_n748_), .Y(new_n2184_));
  AOI21X1  g1542(.A0(new_n1348_), .A1(new_n1347_), .B0(new_n690_), .Y(new_n2185_));
  NOR2X1   g1543(.A(new_n2185_), .B(new_n2184_), .Y(new_n2186_));
  INVX1    g1544(.A(new_n2186_), .Y(new_n2187_));
  NOR3X1   g1545(.A(new_n2061_), .B(new_n2060_), .C(new_n1463_), .Y(new_n2188_));
  AOI21X1  g1546(.A0(new_n2063_), .A1(new_n1998_), .B0(new_n1400_), .Y(new_n2189_));
  NOR2X1   g1547(.A(new_n2189_), .B(new_n2188_), .Y(new_n2190_));
  NOR3X1   g1548(.A(new_n2061_), .B(new_n2060_), .C(new_n1402_), .Y(new_n2191_));
  AOI21X1  g1549(.A0(new_n2063_), .A1(new_n1998_), .B0(new_n1403_), .Y(new_n2192_));
  NOR2X1   g1550(.A(new_n2192_), .B(new_n2191_), .Y(new_n2193_));
  INVX1    g1551(.A(new_n2193_), .Y(new_n2194_));
  NOR3X1   g1552(.A(new_n2061_), .B(new_n2060_), .C(new_n1404_), .Y(new_n2195_));
  AOI21X1  g1553(.A0(new_n2063_), .A1(new_n1998_), .B0(new_n1446_), .Y(new_n2196_));
  NOR2X1   g1554(.A(new_n2196_), .B(new_n2195_), .Y(new_n2197_));
  NOR3X1   g1555(.A(new_n1286_), .B(new_n1284_), .C(new_n731_), .Y(new_n2198_));
  AOI21X1  g1556(.A0(new_n1348_), .A1(new_n1347_), .B0(new_n694_), .Y(new_n2199_));
  NOR2X1   g1557(.A(new_n2199_), .B(new_n2198_), .Y(new_n2200_));
  INVX1    g1558(.A(new_n2200_), .Y(new_n2201_));
  NOR3X1   g1559(.A(new_n2061_), .B(new_n2060_), .C(new_n1441_), .Y(new_n2202_));
  AOI21X1  g1560(.A0(new_n2063_), .A1(new_n1998_), .B0(new_n1405_), .Y(new_n2203_));
  NOR2X1   g1561(.A(new_n2203_), .B(new_n2202_), .Y(new_n2204_));
  NOR3X1   g1562(.A(new_n2061_), .B(new_n2060_), .C(new_n1438_), .Y(new_n2205_));
  AOI21X1  g1563(.A0(new_n2063_), .A1(new_n1998_), .B0(new_n1407_), .Y(new_n2206_));
  NOR2X1   g1564(.A(new_n2206_), .B(new_n2205_), .Y(new_n2207_));
  INVX1    g1565(.A(new_n2207_), .Y(new_n2208_));
  NOR3X1   g1566(.A(new_n1286_), .B(new_n1284_), .C(new_n727_), .Y(new_n2209_));
  AOI21X1  g1567(.A0(new_n1348_), .A1(new_n1347_), .B0(new_n697_), .Y(new_n2210_));
  NOR2X1   g1568(.A(new_n2210_), .B(new_n2209_), .Y(new_n2211_));
  NOR3X1   g1569(.A(new_n2061_), .B(new_n2060_), .C(new_n1448_), .Y(new_n2212_));
  AOI21X1  g1570(.A0(new_n2063_), .A1(new_n1998_), .B0(new_n1449_), .Y(new_n2213_));
  NOR2X1   g1571(.A(new_n2213_), .B(new_n2212_), .Y(new_n2214_));
  NOR3X1   g1572(.A(new_n1286_), .B(new_n1284_), .C(new_n699_), .Y(new_n2215_));
  AOI21X1  g1573(.A0(new_n1348_), .A1(new_n1347_), .B0(new_n700_), .Y(new_n2216_));
  NOR2X1   g1574(.A(new_n2216_), .B(new_n2215_), .Y(new_n2217_));
  NOR3X1   g1575(.A(new_n2061_), .B(new_n2060_), .C(new_n1450_), .Y(new_n2218_));
  AOI21X1  g1576(.A0(new_n2063_), .A1(new_n1998_), .B0(new_n1410_), .Y(new_n2219_));
  NOR2X1   g1577(.A(new_n2219_), .B(new_n2218_), .Y(new_n2220_));
  NOR3X1   g1578(.A(new_n1286_), .B(new_n1284_), .C(new_n701_), .Y(new_n2221_));
  AOI21X1  g1579(.A0(new_n1348_), .A1(new_n1347_), .B0(new_n714_), .Y(new_n2222_));
  NOR2X1   g1580(.A(new_n2222_), .B(new_n2221_), .Y(new_n2223_));
  INVX1    g1581(.A(new_n2223_), .Y(new_n2224_));
  AND2X1   g1582(.A(new_n1348_), .B(new_n1347_), .Y(new_n2225_));
  NAND3X1  g1583(.A(new_n1348_), .B(new_n1347_), .C(\in1[3] ), .Y(new_n2226_));
  OAI21X1  g1584(.A0(new_n2225_), .A1(new_n702_), .B0(new_n2226_), .Y(new_n2227_));
  NOR3X1   g1585(.A(new_n2061_), .B(new_n2060_), .C(new_n1422_), .Y(new_n2228_));
  AOI21X1  g1586(.A0(new_n2071_), .A1(\in2[3] ), .B0(new_n2228_), .Y(new_n2229_));
  NOR2X1   g1587(.A(new_n2229_), .B(new_n2227_), .Y(new_n2230_));
  NOR3X1   g1588(.A(new_n2061_), .B(new_n2060_), .C(new_n1415_), .Y(new_n2231_));
  AOI21X1  g1589(.A0(new_n2063_), .A1(new_n1998_), .B0(new_n1426_), .Y(new_n2232_));
  OR2X1    g1590(.A(new_n2232_), .B(new_n2231_), .Y(new_n2233_));
  NAND3X1  g1591(.A(new_n2063_), .B(new_n1998_), .C(\in3[0] ), .Y(new_n2234_));
  OAI21X1  g1592(.A0(new_n2061_), .A1(new_n2060_), .B0(\in2[0] ), .Y(new_n2235_));
  OR2X1    g1593(.A(new_n1349_), .B(new_n1287_), .Y(new_n2236_));
  NAND3X1  g1594(.A(new_n2236_), .B(new_n2235_), .C(new_n2234_), .Y(new_n2237_));
  NOR3X1   g1595(.A(new_n1286_), .B(new_n1284_), .C(new_n717_), .Y(new_n2238_));
  AOI21X1  g1596(.A0(new_n1348_), .A1(new_n1347_), .B0(new_n706_), .Y(new_n2239_));
  NOR2X1   g1597(.A(new_n2239_), .B(new_n2238_), .Y(new_n2240_));
  OAI21X1  g1598(.A0(new_n2237_), .A1(new_n2233_), .B0(new_n2240_), .Y(new_n2241_));
  NOR3X1   g1599(.A(new_n1286_), .B(new_n1284_), .C(new_n704_), .Y(new_n2242_));
  AOI21X1  g1600(.A0(new_n1348_), .A1(new_n1347_), .B0(new_n708_), .Y(new_n2243_));
  OR2X1    g1601(.A(new_n2243_), .B(new_n2242_), .Y(new_n2244_));
  NOR3X1   g1602(.A(new_n2061_), .B(new_n2060_), .C(new_n1419_), .Y(new_n2245_));
  AOI21X1  g1603(.A0(new_n2063_), .A1(new_n1998_), .B0(new_n1414_), .Y(new_n2246_));
  NOR2X1   g1604(.A(new_n2246_), .B(new_n2245_), .Y(new_n2247_));
  NOR2X1   g1605(.A(new_n2243_), .B(new_n2242_), .Y(new_n2248_));
  OR2X1    g1606(.A(new_n2246_), .B(new_n2245_), .Y(new_n2249_));
  AOI22X1  g1607(.A0(new_n2249_), .A1(new_n2248_), .B0(new_n2237_), .B1(new_n2233_), .Y(new_n2250_));
  AOI22X1  g1608(.A0(new_n2250_), .A1(new_n2241_), .B0(new_n2247_), .B1(new_n2244_), .Y(new_n2251_));
  NAND2X1  g1609(.A(new_n2229_), .B(new_n2227_), .Y(new_n2252_));
  OAI21X1  g1610(.A0(new_n2251_), .A1(new_n2230_), .B0(new_n2252_), .Y(new_n2253_));
  OAI21X1  g1611(.A0(new_n2253_), .A1(new_n2224_), .B0(new_n2220_), .Y(new_n2254_));
  OR2X1    g1612(.A(new_n2229_), .B(new_n2227_), .Y(new_n2255_));
  NOR2X1   g1613(.A(new_n2232_), .B(new_n2231_), .Y(new_n2256_));
  NOR3X1   g1614(.A(new_n2061_), .B(new_n2060_), .C(new_n1416_), .Y(new_n2257_));
  AOI21X1  g1615(.A0(new_n2063_), .A1(new_n1998_), .B0(new_n1427_), .Y(new_n2258_));
  NOR3X1   g1616(.A(new_n1350_), .B(new_n2258_), .C(new_n2257_), .Y(new_n2259_));
  OR2X1    g1617(.A(new_n2239_), .B(new_n2238_), .Y(new_n2260_));
  AOI21X1  g1618(.A0(new_n2259_), .A1(new_n2256_), .B0(new_n2260_), .Y(new_n2261_));
  OAI22X1  g1619(.A0(new_n2247_), .A1(new_n2244_), .B0(new_n2259_), .B1(new_n2256_), .Y(new_n2262_));
  OAI22X1  g1620(.A0(new_n2262_), .A1(new_n2261_), .B0(new_n2249_), .B1(new_n2248_), .Y(new_n2263_));
  AND2X1   g1621(.A(new_n2229_), .B(new_n2227_), .Y(new_n2264_));
  AOI21X1  g1622(.A0(new_n2263_), .A1(new_n2255_), .B0(new_n2264_), .Y(new_n2265_));
  OR2X1    g1623(.A(new_n2265_), .B(new_n2223_), .Y(new_n2266_));
  NAND3X1  g1624(.A(new_n2266_), .B(new_n2254_), .C(new_n2217_), .Y(new_n2267_));
  AOI21X1  g1625(.A0(new_n2266_), .A1(new_n2254_), .B0(new_n2217_), .Y(new_n2268_));
  AOI21X1  g1626(.A0(new_n2267_), .A1(new_n2214_), .B0(new_n2268_), .Y(new_n2269_));
  AOI21X1  g1627(.A0(new_n2269_), .A1(new_n2211_), .B0(new_n2208_), .Y(new_n2270_));
  INVX1    g1628(.A(new_n2211_), .Y(new_n2271_));
  INVX1    g1629(.A(new_n2214_), .Y(new_n2272_));
  INVX1    g1630(.A(new_n2217_), .Y(new_n2273_));
  INVX1    g1631(.A(new_n2220_), .Y(new_n2274_));
  AOI21X1  g1632(.A0(new_n2265_), .A1(new_n2223_), .B0(new_n2274_), .Y(new_n2275_));
  NOR2X1   g1633(.A(new_n2265_), .B(new_n2223_), .Y(new_n2276_));
  NOR3X1   g1634(.A(new_n2276_), .B(new_n2275_), .C(new_n2273_), .Y(new_n2277_));
  OAI21X1  g1635(.A0(new_n2276_), .A1(new_n2275_), .B0(new_n2273_), .Y(new_n2278_));
  OAI21X1  g1636(.A0(new_n2277_), .A1(new_n2272_), .B0(new_n2278_), .Y(new_n2279_));
  AND2X1   g1637(.A(new_n2279_), .B(new_n2271_), .Y(new_n2280_));
  OAI22X1  g1638(.A0(new_n2280_), .A1(new_n2270_), .B0(new_n2204_), .B1(new_n2201_), .Y(new_n2281_));
  NOR3X1   g1639(.A(new_n2203_), .B(new_n2202_), .C(new_n2200_), .Y(new_n2282_));
  INVX1    g1640(.A(new_n2282_), .Y(new_n2283_));
  NOR3X1   g1641(.A(new_n1286_), .B(new_n1284_), .C(new_n776_), .Y(new_n2284_));
  AOI21X1  g1642(.A0(new_n1348_), .A1(new_n1347_), .B0(new_n693_), .Y(new_n2285_));
  NOR2X1   g1643(.A(new_n2285_), .B(new_n2284_), .Y(new_n2286_));
  NAND3X1  g1644(.A(new_n2286_), .B(new_n2283_), .C(new_n2281_), .Y(new_n2287_));
  AOI21X1  g1645(.A0(new_n2283_), .A1(new_n2281_), .B0(new_n2286_), .Y(new_n2288_));
  AOI21X1  g1646(.A0(new_n2287_), .A1(new_n2197_), .B0(new_n2288_), .Y(new_n2289_));
  NOR3X1   g1647(.A(new_n1286_), .B(new_n1284_), .C(new_n774_), .Y(new_n2290_));
  AOI21X1  g1648(.A0(new_n1348_), .A1(new_n1347_), .B0(new_n775_), .Y(new_n2291_));
  NOR2X1   g1649(.A(new_n2291_), .B(new_n2290_), .Y(new_n2292_));
  AOI21X1  g1650(.A0(new_n2292_), .A1(new_n2289_), .B0(new_n2194_), .Y(new_n2293_));
  INVX1    g1651(.A(new_n2197_), .Y(new_n2294_));
  NOR2X1   g1652(.A(new_n2204_), .B(new_n2201_), .Y(new_n2295_));
  OAI21X1  g1653(.A0(new_n2279_), .A1(new_n2271_), .B0(new_n2207_), .Y(new_n2296_));
  NAND2X1  g1654(.A(new_n2279_), .B(new_n2271_), .Y(new_n2297_));
  AOI21X1  g1655(.A0(new_n2297_), .A1(new_n2296_), .B0(new_n2295_), .Y(new_n2298_));
  INVX1    g1656(.A(new_n2286_), .Y(new_n2299_));
  NOR3X1   g1657(.A(new_n2299_), .B(new_n2282_), .C(new_n2298_), .Y(new_n2300_));
  OAI21X1  g1658(.A0(new_n2282_), .A1(new_n2298_), .B0(new_n2299_), .Y(new_n2301_));
  OAI21X1  g1659(.A0(new_n2300_), .A1(new_n2294_), .B0(new_n2301_), .Y(new_n2302_));
  INVX1    g1660(.A(new_n2292_), .Y(new_n2303_));
  AND2X1   g1661(.A(new_n2303_), .B(new_n2302_), .Y(new_n2304_));
  OAI22X1  g1662(.A0(new_n2304_), .A1(new_n2293_), .B0(new_n2190_), .B1(new_n2187_), .Y(new_n2305_));
  NOR3X1   g1663(.A(new_n2189_), .B(new_n2188_), .C(new_n2186_), .Y(new_n2306_));
  INVX1    g1664(.A(new_n2306_), .Y(new_n2307_));
  AOI21X1  g1665(.A0(new_n2307_), .A1(new_n2305_), .B0(new_n2183_), .Y(new_n2308_));
  NOR3X1   g1666(.A(new_n2181_), .B(new_n2180_), .C(new_n2178_), .Y(new_n2309_));
  OAI22X1  g1667(.A0(new_n2309_), .A1(new_n2308_), .B0(new_n2175_), .B1(new_n2172_), .Y(new_n2310_));
  NOR3X1   g1668(.A(new_n2174_), .B(new_n2173_), .C(new_n2171_), .Y(new_n2311_));
  INVX1    g1669(.A(new_n2311_), .Y(new_n2312_));
  AOI21X1  g1670(.A0(new_n2312_), .A1(new_n2310_), .B0(new_n2168_), .Y(new_n2313_));
  NOR3X1   g1671(.A(new_n2166_), .B(new_n2165_), .C(new_n2163_), .Y(new_n2314_));
  OAI22X1  g1672(.A0(new_n2314_), .A1(new_n2313_), .B0(new_n2160_), .B1(new_n2157_), .Y(new_n2315_));
  NOR3X1   g1673(.A(new_n2159_), .B(new_n2158_), .C(new_n2156_), .Y(new_n2316_));
  INVX1    g1674(.A(new_n2316_), .Y(new_n2317_));
  AOI21X1  g1675(.A0(new_n2317_), .A1(new_n2315_), .B0(new_n2153_), .Y(new_n2318_));
  NOR3X1   g1676(.A(new_n2151_), .B(new_n2150_), .C(new_n2148_), .Y(new_n2319_));
  NOR3X1   g1677(.A(new_n1286_), .B(new_n1284_), .C(new_n677_), .Y(new_n2320_));
  AOI21X1  g1678(.A0(new_n1348_), .A1(new_n1347_), .B0(new_n770_), .Y(new_n2321_));
  NOR2X1   g1679(.A(new_n2321_), .B(new_n2320_), .Y(new_n2322_));
  INVX1    g1680(.A(new_n2322_), .Y(new_n2323_));
  NOR3X1   g1681(.A(new_n2323_), .B(new_n2319_), .C(new_n2318_), .Y(new_n2324_));
  OAI21X1  g1682(.A0(new_n2319_), .A1(new_n2318_), .B0(new_n2323_), .Y(new_n2325_));
  OAI21X1  g1683(.A0(new_n2324_), .A1(new_n2145_), .B0(new_n2325_), .Y(new_n2326_));
  NOR3X1   g1684(.A(new_n1286_), .B(new_n1284_), .C(new_n675_), .Y(new_n2327_));
  AOI21X1  g1685(.A0(new_n1348_), .A1(new_n1347_), .B0(new_n676_), .Y(new_n2328_));
  NOR2X1   g1686(.A(new_n2328_), .B(new_n2327_), .Y(new_n2329_));
  INVX1    g1687(.A(new_n2329_), .Y(new_n2330_));
  OAI21X1  g1688(.A0(new_n2330_), .A1(new_n2326_), .B0(new_n2141_), .Y(new_n2331_));
  NAND2X1  g1689(.A(new_n2330_), .B(new_n2326_), .Y(new_n2332_));
  AOI21X1  g1690(.A0(new_n2332_), .A1(new_n2331_), .B0(new_n2139_), .Y(new_n2333_));
  NOR2X1   g1691(.A(new_n2135_), .B(new_n2134_), .Y(new_n2334_));
  NOR3X1   g1692(.A(new_n2137_), .B(new_n2136_), .C(new_n2334_), .Y(new_n2335_));
  OAI21X1  g1693(.A0(new_n2335_), .A1(new_n2333_), .B0(new_n2133_), .Y(new_n2336_));
  NOR3X1   g1694(.A(new_n2132_), .B(new_n2131_), .C(new_n2130_), .Y(new_n2337_));
  INVX1    g1695(.A(new_n2337_), .Y(new_n2338_));
  AOI21X1  g1696(.A0(new_n2338_), .A1(new_n2336_), .B0(new_n2127_), .Y(new_n2339_));
  NOR2X1   g1697(.A(new_n2123_), .B(new_n2122_), .Y(new_n2340_));
  NOR3X1   g1698(.A(new_n2125_), .B(new_n2124_), .C(new_n2340_), .Y(new_n2341_));
  OAI21X1  g1699(.A0(new_n2341_), .A1(new_n2339_), .B0(new_n2121_), .Y(new_n2342_));
  NOR3X1   g1700(.A(new_n2120_), .B(new_n2119_), .C(new_n2118_), .Y(new_n2343_));
  INVX1    g1701(.A(new_n2343_), .Y(new_n2344_));
  AOI21X1  g1702(.A0(new_n2344_), .A1(new_n2342_), .B0(new_n2115_), .Y(new_n2345_));
  NOR2X1   g1703(.A(new_n2111_), .B(new_n2110_), .Y(new_n2346_));
  NOR3X1   g1704(.A(new_n2113_), .B(new_n2112_), .C(new_n2346_), .Y(new_n2347_));
  OAI21X1  g1705(.A0(new_n2347_), .A1(new_n2345_), .B0(new_n2109_), .Y(new_n2348_));
  NOR3X1   g1706(.A(new_n2108_), .B(new_n2107_), .C(new_n2106_), .Y(new_n2349_));
  INVX1    g1707(.A(new_n2349_), .Y(new_n2350_));
  AOI21X1  g1708(.A0(new_n1348_), .A1(new_n1347_), .B0(new_n659_), .Y(new_n2351_));
  AOI21X1  g1709(.A0(new_n2225_), .A1(\in1[24] ), .B0(new_n2351_), .Y(new_n2352_));
  NAND3X1  g1710(.A(new_n2352_), .B(new_n2350_), .C(new_n2348_), .Y(new_n2353_));
  AOI21X1  g1711(.A0(new_n2350_), .A1(new_n2348_), .B0(new_n2352_), .Y(new_n2354_));
  AOI21X1  g1712(.A0(new_n2353_), .A1(new_n2103_), .B0(new_n2354_), .Y(new_n2355_));
  AOI21X1  g1713(.A0(new_n1348_), .A1(new_n1347_), .B0(new_n1292_), .Y(new_n2356_));
  AOI21X1  g1714(.A0(new_n2225_), .A1(\in1[25] ), .B0(new_n2356_), .Y(new_n2357_));
  AOI21X1  g1715(.A0(new_n2357_), .A1(new_n2355_), .B0(new_n2101_), .Y(new_n2358_));
  NOR2X1   g1716(.A(new_n2357_), .B(new_n2355_), .Y(new_n2359_));
  OAI22X1  g1717(.A0(new_n2359_), .A1(new_n2358_), .B0(new_n2097_), .B1(new_n2095_), .Y(new_n2360_));
  NAND2X1  g1718(.A(new_n2097_), .B(new_n2095_), .Y(new_n2361_));
  AOI21X1  g1719(.A0(new_n2361_), .A1(new_n2360_), .B0(new_n2091_), .Y(new_n2362_));
  NOR2X1   g1720(.A(new_n2087_), .B(new_n2086_), .Y(new_n2363_));
  NOR3X1   g1721(.A(new_n2089_), .B(new_n2088_), .C(new_n2363_), .Y(new_n2364_));
  OAI22X1  g1722(.A0(new_n2364_), .A1(new_n2362_), .B0(new_n2085_), .B1(new_n2083_), .Y(new_n2365_));
  NAND2X1  g1723(.A(new_n2085_), .B(new_n2083_), .Y(new_n2366_));
  AOI21X1  g1724(.A0(new_n2366_), .A1(new_n2365_), .B0(new_n2079_), .Y(new_n2367_));
  NOR2X1   g1725(.A(new_n2075_), .B(new_n2074_), .Y(new_n2368_));
  NOR3X1   g1726(.A(new_n2077_), .B(new_n2076_), .C(new_n2368_), .Y(new_n2369_));
  OAI22X1  g1727(.A0(new_n2369_), .A1(new_n2367_), .B0(new_n2073_), .B1(new_n2070_), .Y(new_n2370_));
  NAND2X1  g1728(.A(new_n2073_), .B(new_n2070_), .Y(new_n2371_));
  AOI21X1  g1729(.A0(new_n2371_), .A1(new_n2370_), .B0(new_n2066_), .Y(new_n2372_));
  NOR2X1   g1730(.A(new_n2003_), .B(new_n2002_), .Y(new_n2373_));
  NOR3X1   g1731(.A(new_n2064_), .B(new_n2062_), .C(new_n2373_), .Y(new_n2374_));
  NOR3X1   g1732(.A(new_n2061_), .B(new_n2060_), .C(new_n1593_), .Y(new_n2375_));
  AOI21X1  g1733(.A0(new_n2071_), .A1(\in2[34] ), .B0(new_n2375_), .Y(new_n2376_));
  NOR3X1   g1734(.A(new_n1286_), .B(new_n1284_), .C(new_n877_), .Y(new_n2377_));
  AOI21X1  g1735(.A0(new_n1348_), .A1(new_n1347_), .B0(new_n866_), .Y(new_n2378_));
  NOR2X1   g1736(.A(new_n2378_), .B(new_n2377_), .Y(new_n2379_));
  INVX1    g1737(.A(new_n2379_), .Y(new_n2380_));
  NOR2X1   g1738(.A(new_n2380_), .B(new_n2376_), .Y(new_n2381_));
  INVX1    g1739(.A(new_n2225_), .Y(new_n2382_));
  NOR3X1   g1740(.A(new_n1286_), .B(new_n1284_), .C(new_n871_), .Y(new_n2383_));
  AOI21X1  g1741(.A0(new_n2382_), .A1(\in0[33] ), .B0(new_n2383_), .Y(new_n2384_));
  INVX1    g1742(.A(new_n2384_), .Y(new_n2385_));
  NOR3X1   g1743(.A(new_n2061_), .B(new_n2060_), .C(new_n1586_), .Y(new_n2386_));
  AOI21X1  g1744(.A0(new_n2071_), .A1(\in2[33] ), .B0(new_n2386_), .Y(new_n2387_));
  AOI21X1  g1745(.A0(new_n1348_), .A1(new_n1347_), .B0(new_n867_), .Y(new_n2388_));
  AOI21X1  g1746(.A0(new_n2225_), .A1(\in1[35] ), .B0(new_n2388_), .Y(new_n2389_));
  INVX1    g1747(.A(new_n2389_), .Y(new_n2390_));
  INVX1    g1748(.A(new_n2071_), .Y(new_n2391_));
  AOI21X1  g1749(.A0(new_n2063_), .A1(new_n1998_), .B0(new_n1582_), .Y(new_n2392_));
  AOI21X1  g1750(.A0(new_n2391_), .A1(\in3[35] ), .B0(new_n2392_), .Y(new_n2393_));
  OAI22X1  g1751(.A0(new_n2393_), .A1(new_n2390_), .B0(new_n2387_), .B1(new_n2385_), .Y(new_n2394_));
  OR2X1    g1752(.A(new_n2394_), .B(new_n2381_), .Y(new_n2395_));
  NOR3X1   g1753(.A(new_n2061_), .B(new_n2060_), .C(new_n1585_), .Y(new_n2396_));
  AOI21X1  g1754(.A0(new_n2071_), .A1(\in2[32] ), .B0(new_n2396_), .Y(new_n2397_));
  NOR3X1   g1755(.A(new_n1286_), .B(new_n1284_), .C(new_n870_), .Y(new_n2398_));
  AND2X1   g1756(.A(new_n2382_), .B(\in0[32] ), .Y(new_n2399_));
  NOR3X1   g1757(.A(new_n2399_), .B(new_n2398_), .C(new_n2397_), .Y(new_n2400_));
  NOR3X1   g1758(.A(new_n1286_), .B(new_n1284_), .C(new_n886_), .Y(new_n2401_));
  AOI21X1  g1759(.A0(new_n1348_), .A1(new_n1347_), .B0(new_n860_), .Y(new_n2402_));
  NOR2X1   g1760(.A(new_n2402_), .B(new_n2401_), .Y(new_n2403_));
  INVX1    g1761(.A(new_n2403_), .Y(new_n2404_));
  NOR3X1   g1762(.A(new_n2061_), .B(new_n2060_), .C(new_n1601_), .Y(new_n2405_));
  AOI21X1  g1763(.A0(new_n2071_), .A1(\in2[39] ), .B0(new_n2405_), .Y(new_n2406_));
  AOI21X1  g1764(.A0(new_n2063_), .A1(new_n1998_), .B0(new_n1574_), .Y(new_n2407_));
  AOI21X1  g1765(.A0(new_n2391_), .A1(\in3[38] ), .B0(new_n2407_), .Y(new_n2408_));
  AOI21X1  g1766(.A0(new_n1348_), .A1(new_n1347_), .B0(new_n859_), .Y(new_n2409_));
  AOI21X1  g1767(.A0(new_n2225_), .A1(\in1[38] ), .B0(new_n2409_), .Y(new_n2410_));
  INVX1    g1768(.A(new_n2410_), .Y(new_n2411_));
  OAI22X1  g1769(.A0(new_n2411_), .A1(new_n2408_), .B0(new_n2406_), .B1(new_n2404_), .Y(new_n2412_));
  NOR3X1   g1770(.A(new_n1286_), .B(new_n1284_), .C(new_n863_), .Y(new_n2413_));
  AOI21X1  g1771(.A0(new_n1348_), .A1(new_n1347_), .B0(new_n881_), .Y(new_n2414_));
  NOR2X1   g1772(.A(new_n2414_), .B(new_n2413_), .Y(new_n2415_));
  INVX1    g1773(.A(new_n2415_), .Y(new_n2416_));
  NOR3X1   g1774(.A(new_n2061_), .B(new_n2060_), .C(new_n1578_), .Y(new_n2417_));
  AOI21X1  g1775(.A0(new_n2071_), .A1(\in2[36] ), .B0(new_n2417_), .Y(new_n2418_));
  NOR3X1   g1776(.A(new_n1286_), .B(new_n1284_), .C(new_n864_), .Y(new_n2419_));
  AOI21X1  g1777(.A0(new_n1348_), .A1(new_n1347_), .B0(new_n882_), .Y(new_n2420_));
  NOR2X1   g1778(.A(new_n2420_), .B(new_n2419_), .Y(new_n2421_));
  INVX1    g1779(.A(new_n2421_), .Y(new_n2422_));
  NOR3X1   g1780(.A(new_n2061_), .B(new_n2060_), .C(new_n1579_), .Y(new_n2423_));
  AOI21X1  g1781(.A0(new_n2071_), .A1(\in2[37] ), .B0(new_n2423_), .Y(new_n2424_));
  OAI22X1  g1782(.A0(new_n2424_), .A1(new_n2422_), .B0(new_n2418_), .B1(new_n2416_), .Y(new_n2425_));
  NOR4X1   g1783(.A(new_n2425_), .B(new_n2412_), .C(new_n2400_), .D(new_n2395_), .Y(new_n2426_));
  OAI21X1  g1784(.A0(new_n2374_), .A1(new_n2372_), .B0(new_n2426_), .Y(new_n2427_));
  NOR2X1   g1785(.A(new_n2425_), .B(new_n2412_), .Y(new_n2428_));
  AOI21X1  g1786(.A0(new_n2382_), .A1(\in0[32] ), .B0(new_n2398_), .Y(new_n2429_));
  INVX1    g1787(.A(new_n2429_), .Y(new_n2430_));
  AOI22X1  g1788(.A0(new_n2430_), .A1(new_n2397_), .B0(new_n2387_), .B1(new_n2385_), .Y(new_n2431_));
  NAND2X1  g1789(.A(new_n2393_), .B(new_n2390_), .Y(new_n2432_));
  AND2X1   g1790(.A(new_n2380_), .B(new_n2376_), .Y(new_n2433_));
  OAI21X1  g1791(.A0(new_n2393_), .A1(new_n2390_), .B0(new_n2433_), .Y(new_n2434_));
  AND2X1   g1792(.A(new_n2434_), .B(new_n2432_), .Y(new_n2435_));
  OAI21X1  g1793(.A0(new_n2431_), .A1(new_n2395_), .B0(new_n2435_), .Y(new_n2436_));
  AND2X1   g1794(.A(new_n2418_), .B(new_n2416_), .Y(new_n2437_));
  OAI21X1  g1795(.A0(new_n2424_), .A1(new_n2422_), .B0(new_n2437_), .Y(new_n2438_));
  NAND2X1  g1796(.A(new_n2424_), .B(new_n2422_), .Y(new_n2439_));
  AOI21X1  g1797(.A0(new_n2439_), .A1(new_n2438_), .B0(new_n2412_), .Y(new_n2440_));
  NOR2X1   g1798(.A(new_n2406_), .B(new_n2404_), .Y(new_n2441_));
  NAND2X1  g1799(.A(new_n2406_), .B(new_n2404_), .Y(new_n2442_));
  NAND2X1  g1800(.A(new_n2411_), .B(new_n2408_), .Y(new_n2443_));
  OAI21X1  g1801(.A0(new_n2443_), .A1(new_n2441_), .B0(new_n2442_), .Y(new_n2444_));
  OR2X1    g1802(.A(new_n2444_), .B(new_n2440_), .Y(new_n2445_));
  AOI21X1  g1803(.A0(new_n2436_), .A1(new_n2428_), .B0(new_n2445_), .Y(new_n2446_));
  NOR3X1   g1804(.A(new_n1286_), .B(new_n1284_), .C(new_n922_), .Y(new_n2447_));
  AOI21X1  g1805(.A0(new_n1348_), .A1(new_n1347_), .B0(new_n895_), .Y(new_n2448_));
  NOR2X1   g1806(.A(new_n2448_), .B(new_n2447_), .Y(new_n2449_));
  INVX1    g1807(.A(new_n2449_), .Y(new_n2450_));
  NOR3X1   g1808(.A(new_n2061_), .B(new_n2060_), .C(new_n1634_), .Y(new_n2451_));
  AOI21X1  g1809(.A0(new_n2071_), .A1(\in2[47] ), .B0(new_n2451_), .Y(new_n2452_));
  OR2X1    g1810(.A(new_n2452_), .B(new_n2450_), .Y(new_n2453_));
  AOI21X1  g1811(.A0(new_n2063_), .A1(new_n1998_), .B0(new_n1608_), .Y(new_n2454_));
  AOI21X1  g1812(.A0(new_n2391_), .A1(\in3[46] ), .B0(new_n2454_), .Y(new_n2455_));
  AOI21X1  g1813(.A0(new_n1348_), .A1(new_n1347_), .B0(new_n894_), .Y(new_n2456_));
  AOI21X1  g1814(.A0(new_n2225_), .A1(\in1[46] ), .B0(new_n2456_), .Y(new_n2457_));
  INVX1    g1815(.A(new_n2457_), .Y(new_n2458_));
  OAI21X1  g1816(.A0(new_n2458_), .A1(new_n2455_), .B0(new_n2453_), .Y(new_n2459_));
  NOR3X1   g1817(.A(new_n1286_), .B(new_n1284_), .C(new_n898_), .Y(new_n2460_));
  AOI21X1  g1818(.A0(new_n1348_), .A1(new_n1347_), .B0(new_n917_), .Y(new_n2461_));
  NOR2X1   g1819(.A(new_n2461_), .B(new_n2460_), .Y(new_n2462_));
  INVX1    g1820(.A(new_n2462_), .Y(new_n2463_));
  NOR3X1   g1821(.A(new_n2061_), .B(new_n2060_), .C(new_n1612_), .Y(new_n2464_));
  AOI21X1  g1822(.A0(new_n2071_), .A1(\in2[44] ), .B0(new_n2464_), .Y(new_n2465_));
  NOR3X1   g1823(.A(new_n1286_), .B(new_n1284_), .C(new_n899_), .Y(new_n2466_));
  AOI21X1  g1824(.A0(new_n1348_), .A1(new_n1347_), .B0(new_n918_), .Y(new_n2467_));
  NOR2X1   g1825(.A(new_n2467_), .B(new_n2466_), .Y(new_n2468_));
  INVX1    g1826(.A(new_n2468_), .Y(new_n2469_));
  NOR3X1   g1827(.A(new_n2061_), .B(new_n2060_), .C(new_n1613_), .Y(new_n2470_));
  AOI21X1  g1828(.A0(new_n2071_), .A1(\in2[45] ), .B0(new_n2470_), .Y(new_n2471_));
  OAI22X1  g1829(.A0(new_n2471_), .A1(new_n2469_), .B0(new_n2465_), .B1(new_n2463_), .Y(new_n2472_));
  NOR2X1   g1830(.A(new_n2472_), .B(new_n2459_), .Y(new_n2473_));
  AOI21X1  g1831(.A0(new_n1348_), .A1(new_n1347_), .B0(new_n902_), .Y(new_n2474_));
  AOI21X1  g1832(.A0(new_n2225_), .A1(\in1[43] ), .B0(new_n2474_), .Y(new_n2475_));
  AOI21X1  g1833(.A0(new_n2063_), .A1(new_n1998_), .B0(new_n1616_), .Y(new_n2476_));
  AOI21X1  g1834(.A0(new_n2391_), .A1(\in3[43] ), .B0(new_n2476_), .Y(new_n2477_));
  INVX1    g1835(.A(new_n2477_), .Y(new_n2478_));
  AOI21X1  g1836(.A0(new_n1348_), .A1(new_n1347_), .B0(new_n901_), .Y(new_n2479_));
  AOI21X1  g1837(.A0(new_n2225_), .A1(\in1[42] ), .B0(new_n2479_), .Y(new_n2480_));
  NOR3X1   g1838(.A(new_n2061_), .B(new_n2060_), .C(new_n1626_), .Y(new_n2481_));
  AOI21X1  g1839(.A0(new_n2063_), .A1(new_n1998_), .B0(new_n1615_), .Y(new_n2482_));
  NOR2X1   g1840(.A(new_n2482_), .B(new_n2481_), .Y(new_n2483_));
  INVX1    g1841(.A(new_n2483_), .Y(new_n2484_));
  AOI22X1  g1842(.A0(new_n2484_), .A1(new_n2480_), .B0(new_n2478_), .B1(new_n2475_), .Y(new_n2485_));
  NOR3X1   g1843(.A(new_n1286_), .B(new_n1284_), .C(new_n906_), .Y(new_n2486_));
  AND2X1   g1844(.A(new_n2382_), .B(\in0[41] ), .Y(new_n2487_));
  NOR3X1   g1845(.A(new_n2061_), .B(new_n2060_), .C(new_n1620_), .Y(new_n2488_));
  AOI21X1  g1846(.A0(new_n2071_), .A1(\in2[41] ), .B0(new_n2488_), .Y(new_n2489_));
  NOR3X1   g1847(.A(new_n2489_), .B(new_n2487_), .C(new_n2486_), .Y(new_n2490_));
  NOR3X1   g1848(.A(new_n1286_), .B(new_n1284_), .C(new_n905_), .Y(new_n2491_));
  AOI21X1  g1849(.A0(new_n2382_), .A1(\in0[40] ), .B0(new_n2491_), .Y(new_n2492_));
  NOR3X1   g1850(.A(new_n2061_), .B(new_n2060_), .C(new_n1619_), .Y(new_n2493_));
  AOI21X1  g1851(.A0(new_n2071_), .A1(\in2[40] ), .B0(new_n2493_), .Y(new_n2494_));
  INVX1    g1852(.A(new_n2494_), .Y(new_n2495_));
  AOI21X1  g1853(.A0(new_n2495_), .A1(new_n2492_), .B0(new_n2490_), .Y(new_n2496_));
  NAND3X1  g1854(.A(new_n2496_), .B(new_n2485_), .C(new_n2473_), .Y(new_n2497_));
  AOI21X1  g1855(.A0(new_n2446_), .A1(new_n2427_), .B0(new_n2497_), .Y(new_n2498_));
  INVX1    g1856(.A(new_n2473_), .Y(new_n2499_));
  OR2X1    g1857(.A(new_n2478_), .B(new_n2475_), .Y(new_n2500_));
  NOR3X1   g1858(.A(new_n2495_), .B(new_n2492_), .C(new_n2490_), .Y(new_n2501_));
  OAI21X1  g1859(.A0(new_n2487_), .A1(new_n2486_), .B0(new_n2489_), .Y(new_n2502_));
  OAI21X1  g1860(.A0(new_n2484_), .A1(new_n2480_), .B0(new_n2502_), .Y(new_n2503_));
  OAI21X1  g1861(.A0(new_n2503_), .A1(new_n2501_), .B0(new_n2485_), .Y(new_n2504_));
  AOI21X1  g1862(.A0(new_n2504_), .A1(new_n2500_), .B0(new_n2499_), .Y(new_n2505_));
  OR2X1    g1863(.A(new_n2471_), .B(new_n2469_), .Y(new_n2506_));
  NAND3X1  g1864(.A(new_n2506_), .B(new_n2465_), .C(new_n2463_), .Y(new_n2507_));
  NAND2X1  g1865(.A(new_n2471_), .B(new_n2469_), .Y(new_n2508_));
  AOI21X1  g1866(.A0(new_n2508_), .A1(new_n2507_), .B0(new_n2459_), .Y(new_n2509_));
  AND2X1   g1867(.A(new_n2452_), .B(new_n2450_), .Y(new_n2510_));
  AND2X1   g1868(.A(new_n2458_), .B(new_n2455_), .Y(new_n2511_));
  AND2X1   g1869(.A(new_n2511_), .B(new_n2453_), .Y(new_n2512_));
  OR4X1    g1870(.A(new_n2512_), .B(new_n2510_), .C(new_n2509_), .D(new_n2505_), .Y(new_n2513_));
  NOR3X1   g1871(.A(new_n2061_), .B(new_n2060_), .C(new_n1661_), .Y(new_n2514_));
  AOI21X1  g1872(.A0(new_n2071_), .A1(\in2[50] ), .B0(new_n2514_), .Y(new_n2515_));
  NOR3X1   g1873(.A(new_n1286_), .B(new_n1284_), .C(new_n947_), .Y(new_n2516_));
  AOI21X1  g1874(.A0(new_n1348_), .A1(new_n1347_), .B0(new_n936_), .Y(new_n2517_));
  NOR2X1   g1875(.A(new_n2517_), .B(new_n2516_), .Y(new_n2518_));
  INVX1    g1876(.A(new_n2518_), .Y(new_n2519_));
  NOR2X1   g1877(.A(new_n2519_), .B(new_n2515_), .Y(new_n2520_));
  NOR3X1   g1878(.A(new_n1286_), .B(new_n1284_), .C(new_n941_), .Y(new_n2521_));
  AOI21X1  g1879(.A0(new_n2382_), .A1(\in0[49] ), .B0(new_n2521_), .Y(new_n2522_));
  INVX1    g1880(.A(new_n2522_), .Y(new_n2523_));
  NOR3X1   g1881(.A(new_n2061_), .B(new_n2060_), .C(new_n1654_), .Y(new_n2524_));
  AOI21X1  g1882(.A0(new_n2071_), .A1(\in2[49] ), .B0(new_n2524_), .Y(new_n2525_));
  AOI21X1  g1883(.A0(new_n1348_), .A1(new_n1347_), .B0(new_n937_), .Y(new_n2526_));
  AOI21X1  g1884(.A0(new_n2225_), .A1(\in1[51] ), .B0(new_n2526_), .Y(new_n2527_));
  INVX1    g1885(.A(new_n2527_), .Y(new_n2528_));
  AOI21X1  g1886(.A0(new_n2063_), .A1(new_n1998_), .B0(new_n1650_), .Y(new_n2529_));
  AOI21X1  g1887(.A0(new_n2391_), .A1(\in3[51] ), .B0(new_n2529_), .Y(new_n2530_));
  OAI22X1  g1888(.A0(new_n2530_), .A1(new_n2528_), .B0(new_n2525_), .B1(new_n2523_), .Y(new_n2531_));
  OR2X1    g1889(.A(new_n2531_), .B(new_n2520_), .Y(new_n2532_));
  NOR3X1   g1890(.A(new_n2061_), .B(new_n2060_), .C(new_n1653_), .Y(new_n2533_));
  AOI21X1  g1891(.A0(new_n2071_), .A1(\in2[48] ), .B0(new_n2533_), .Y(new_n2534_));
  NOR3X1   g1892(.A(new_n1286_), .B(new_n1284_), .C(new_n940_), .Y(new_n2535_));
  AND2X1   g1893(.A(new_n2382_), .B(\in0[48] ), .Y(new_n2536_));
  NOR3X1   g1894(.A(new_n2536_), .B(new_n2535_), .C(new_n2534_), .Y(new_n2537_));
  AOI21X1  g1895(.A0(new_n1348_), .A1(new_n1347_), .B0(new_n930_), .Y(new_n2538_));
  AOI21X1  g1896(.A0(new_n2225_), .A1(\in1[55] ), .B0(new_n2538_), .Y(new_n2539_));
  AOI21X1  g1897(.A0(new_n2063_), .A1(new_n1998_), .B0(new_n1643_), .Y(new_n2540_));
  AOI21X1  g1898(.A0(new_n2391_), .A1(\in3[55] ), .B0(new_n2540_), .Y(new_n2541_));
  INVX1    g1899(.A(new_n2541_), .Y(new_n2542_));
  NOR3X1   g1900(.A(new_n2061_), .B(new_n2060_), .C(new_n1667_), .Y(new_n2543_));
  AOI21X1  g1901(.A0(new_n2063_), .A1(new_n1998_), .B0(new_n1642_), .Y(new_n2544_));
  NOR2X1   g1902(.A(new_n2544_), .B(new_n2543_), .Y(new_n2545_));
  INVX1    g1903(.A(new_n2545_), .Y(new_n2546_));
  AOI21X1  g1904(.A0(new_n1348_), .A1(new_n1347_), .B0(new_n929_), .Y(new_n2547_));
  AOI21X1  g1905(.A0(new_n2225_), .A1(\in1[54] ), .B0(new_n2547_), .Y(new_n2548_));
  AOI22X1  g1906(.A0(new_n2548_), .A1(new_n2546_), .B0(new_n2542_), .B1(new_n2539_), .Y(new_n2549_));
  INVX1    g1907(.A(new_n2549_), .Y(new_n2550_));
  NOR3X1   g1908(.A(new_n1286_), .B(new_n1284_), .C(new_n934_), .Y(new_n2551_));
  AOI21X1  g1909(.A0(new_n2382_), .A1(\in0[53] ), .B0(new_n2551_), .Y(new_n2552_));
  NOR3X1   g1910(.A(new_n2061_), .B(new_n2060_), .C(new_n1647_), .Y(new_n2553_));
  AND2X1   g1911(.A(new_n2071_), .B(\in2[53] ), .Y(new_n2554_));
  OAI21X1  g1912(.A0(new_n2554_), .A1(new_n2553_), .B0(new_n2552_), .Y(new_n2555_));
  NOR3X1   g1913(.A(new_n2061_), .B(new_n2060_), .C(new_n1646_), .Y(new_n2556_));
  AOI21X1  g1914(.A0(new_n2071_), .A1(\in2[52] ), .B0(new_n2556_), .Y(new_n2557_));
  NOR3X1   g1915(.A(new_n1286_), .B(new_n1284_), .C(new_n933_), .Y(new_n2558_));
  AOI21X1  g1916(.A0(new_n2382_), .A1(\in0[52] ), .B0(new_n2558_), .Y(new_n2559_));
  INVX1    g1917(.A(new_n2559_), .Y(new_n2560_));
  OAI21X1  g1918(.A0(new_n2560_), .A1(new_n2557_), .B0(new_n2555_), .Y(new_n2561_));
  NOR4X1   g1919(.A(new_n2561_), .B(new_n2550_), .C(new_n2537_), .D(new_n2532_), .Y(new_n2562_));
  OAI21X1  g1920(.A0(new_n2513_), .A1(new_n2498_), .B0(new_n2562_), .Y(new_n2563_));
  NOR2X1   g1921(.A(new_n2561_), .B(new_n2550_), .Y(new_n2564_));
  AOI21X1  g1922(.A0(new_n2382_), .A1(\in0[48] ), .B0(new_n2535_), .Y(new_n2565_));
  INVX1    g1923(.A(new_n2565_), .Y(new_n2566_));
  AOI22X1  g1924(.A0(new_n2566_), .A1(new_n2534_), .B0(new_n2525_), .B1(new_n2523_), .Y(new_n2567_));
  NAND2X1  g1925(.A(new_n2530_), .B(new_n2528_), .Y(new_n2568_));
  AND2X1   g1926(.A(new_n2519_), .B(new_n2515_), .Y(new_n2569_));
  OAI21X1  g1927(.A0(new_n2530_), .A1(new_n2528_), .B0(new_n2569_), .Y(new_n2570_));
  AND2X1   g1928(.A(new_n2570_), .B(new_n2568_), .Y(new_n2571_));
  OAI21X1  g1929(.A0(new_n2567_), .A1(new_n2532_), .B0(new_n2571_), .Y(new_n2572_));
  AND2X1   g1930(.A(new_n2071_), .B(\in2[52] ), .Y(new_n2573_));
  NOR3X1   g1931(.A(new_n2559_), .B(new_n2573_), .C(new_n2556_), .Y(new_n2574_));
  AND2X1   g1932(.A(new_n2574_), .B(new_n2555_), .Y(new_n2575_));
  AND2X1   g1933(.A(new_n2382_), .B(\in0[53] ), .Y(new_n2576_));
  AOI21X1  g1934(.A0(new_n2071_), .A1(\in2[53] ), .B0(new_n2553_), .Y(new_n2577_));
  OAI21X1  g1935(.A0(new_n2576_), .A1(new_n2551_), .B0(new_n2577_), .Y(new_n2578_));
  OAI21X1  g1936(.A0(new_n2548_), .A1(new_n2546_), .B0(new_n2578_), .Y(new_n2579_));
  OAI21X1  g1937(.A0(new_n2579_), .A1(new_n2575_), .B0(new_n2549_), .Y(new_n2580_));
  OAI21X1  g1938(.A0(new_n2542_), .A1(new_n2539_), .B0(new_n2580_), .Y(new_n2581_));
  AOI21X1  g1939(.A0(new_n2572_), .A1(new_n2564_), .B0(new_n2581_), .Y(new_n2582_));
  NOR3X1   g1940(.A(new_n1286_), .B(new_n1284_), .C(new_n988_), .Y(new_n2583_));
  AOI21X1  g1941(.A0(new_n1348_), .A1(new_n1347_), .B0(new_n961_), .Y(new_n2584_));
  NOR2X1   g1942(.A(new_n2584_), .B(new_n2583_), .Y(new_n2585_));
  INVX1    g1943(.A(new_n2585_), .Y(new_n2586_));
  NOR3X1   g1944(.A(new_n2061_), .B(new_n2060_), .C(new_n1699_), .Y(new_n2587_));
  AOI21X1  g1945(.A0(new_n2071_), .A1(\in2[63] ), .B0(new_n2587_), .Y(new_n2588_));
  OR2X1    g1946(.A(new_n2588_), .B(new_n2586_), .Y(new_n2589_));
  AOI21X1  g1947(.A0(new_n2063_), .A1(new_n1998_), .B0(new_n1673_), .Y(new_n2590_));
  AOI21X1  g1948(.A0(new_n2391_), .A1(\in3[62] ), .B0(new_n2590_), .Y(new_n2591_));
  AOI21X1  g1949(.A0(new_n1348_), .A1(new_n1347_), .B0(new_n960_), .Y(new_n2592_));
  AOI21X1  g1950(.A0(new_n2225_), .A1(\in1[62] ), .B0(new_n2592_), .Y(new_n2593_));
  INVX1    g1951(.A(new_n2593_), .Y(new_n2594_));
  OAI21X1  g1952(.A0(new_n2594_), .A1(new_n2591_), .B0(new_n2589_), .Y(new_n2595_));
  NOR3X1   g1953(.A(new_n1286_), .B(new_n1284_), .C(new_n964_), .Y(new_n2596_));
  AOI21X1  g1954(.A0(new_n1348_), .A1(new_n1347_), .B0(new_n983_), .Y(new_n2597_));
  NOR2X1   g1955(.A(new_n2597_), .B(new_n2596_), .Y(new_n2598_));
  INVX1    g1956(.A(new_n2598_), .Y(new_n2599_));
  NOR3X1   g1957(.A(new_n2061_), .B(new_n2060_), .C(new_n1677_), .Y(new_n2600_));
  AOI21X1  g1958(.A0(new_n2071_), .A1(\in2[60] ), .B0(new_n2600_), .Y(new_n2601_));
  NOR3X1   g1959(.A(new_n1286_), .B(new_n1284_), .C(new_n965_), .Y(new_n2602_));
  AOI21X1  g1960(.A0(new_n1348_), .A1(new_n1347_), .B0(new_n984_), .Y(new_n2603_));
  NOR2X1   g1961(.A(new_n2603_), .B(new_n2602_), .Y(new_n2604_));
  INVX1    g1962(.A(new_n2604_), .Y(new_n2605_));
  NOR3X1   g1963(.A(new_n2061_), .B(new_n2060_), .C(new_n1678_), .Y(new_n2606_));
  AOI21X1  g1964(.A0(new_n2071_), .A1(\in2[61] ), .B0(new_n2606_), .Y(new_n2607_));
  OAI22X1  g1965(.A0(new_n2607_), .A1(new_n2605_), .B0(new_n2601_), .B1(new_n2599_), .Y(new_n2608_));
  NOR2X1   g1966(.A(new_n2608_), .B(new_n2595_), .Y(new_n2609_));
  AOI21X1  g1967(.A0(new_n1348_), .A1(new_n1347_), .B0(new_n968_), .Y(new_n2610_));
  AOI21X1  g1968(.A0(new_n2225_), .A1(\in1[59] ), .B0(new_n2610_), .Y(new_n2611_));
  AOI21X1  g1969(.A0(new_n2063_), .A1(new_n1998_), .B0(new_n1681_), .Y(new_n2612_));
  AOI21X1  g1970(.A0(new_n2391_), .A1(\in3[59] ), .B0(new_n2612_), .Y(new_n2613_));
  INVX1    g1971(.A(new_n2613_), .Y(new_n2614_));
  AOI21X1  g1972(.A0(new_n1348_), .A1(new_n1347_), .B0(new_n967_), .Y(new_n2615_));
  AOI21X1  g1973(.A0(new_n2225_), .A1(\in1[58] ), .B0(new_n2615_), .Y(new_n2616_));
  NOR3X1   g1974(.A(new_n2061_), .B(new_n2060_), .C(new_n1691_), .Y(new_n2617_));
  AOI21X1  g1975(.A0(new_n2063_), .A1(new_n1998_), .B0(new_n1680_), .Y(new_n2618_));
  NOR2X1   g1976(.A(new_n2618_), .B(new_n2617_), .Y(new_n2619_));
  INVX1    g1977(.A(new_n2619_), .Y(new_n2620_));
  AOI22X1  g1978(.A0(new_n2620_), .A1(new_n2616_), .B0(new_n2614_), .B1(new_n2611_), .Y(new_n2621_));
  NOR3X1   g1979(.A(new_n1286_), .B(new_n1284_), .C(new_n972_), .Y(new_n2622_));
  AND2X1   g1980(.A(new_n2382_), .B(\in0[57] ), .Y(new_n2623_));
  NOR3X1   g1981(.A(new_n2061_), .B(new_n2060_), .C(new_n1685_), .Y(new_n2624_));
  AOI21X1  g1982(.A0(new_n2071_), .A1(\in2[57] ), .B0(new_n2624_), .Y(new_n2625_));
  NOR3X1   g1983(.A(new_n2625_), .B(new_n2623_), .C(new_n2622_), .Y(new_n2626_));
  NOR3X1   g1984(.A(new_n1286_), .B(new_n1284_), .C(new_n971_), .Y(new_n2627_));
  AOI21X1  g1985(.A0(new_n2382_), .A1(\in0[56] ), .B0(new_n2627_), .Y(new_n2628_));
  NOR3X1   g1986(.A(new_n2061_), .B(new_n2060_), .C(new_n1684_), .Y(new_n2629_));
  AOI21X1  g1987(.A0(new_n2071_), .A1(\in2[56] ), .B0(new_n2629_), .Y(new_n2630_));
  INVX1    g1988(.A(new_n2630_), .Y(new_n2631_));
  AOI21X1  g1989(.A0(new_n2631_), .A1(new_n2628_), .B0(new_n2626_), .Y(new_n2632_));
  NAND3X1  g1990(.A(new_n2632_), .B(new_n2621_), .C(new_n2609_), .Y(new_n2633_));
  AOI21X1  g1991(.A0(new_n2582_), .A1(new_n2563_), .B0(new_n2633_), .Y(new_n2634_));
  INVX1    g1992(.A(new_n2609_), .Y(new_n2635_));
  OR2X1    g1993(.A(new_n2614_), .B(new_n2611_), .Y(new_n2636_));
  NOR3X1   g1994(.A(new_n2631_), .B(new_n2628_), .C(new_n2626_), .Y(new_n2637_));
  OAI21X1  g1995(.A0(new_n2623_), .A1(new_n2622_), .B0(new_n2625_), .Y(new_n2638_));
  OAI21X1  g1996(.A0(new_n2620_), .A1(new_n2616_), .B0(new_n2638_), .Y(new_n2639_));
  OAI21X1  g1997(.A0(new_n2639_), .A1(new_n2637_), .B0(new_n2621_), .Y(new_n2640_));
  AOI21X1  g1998(.A0(new_n2640_), .A1(new_n2636_), .B0(new_n2635_), .Y(new_n2641_));
  OR2X1    g1999(.A(new_n2607_), .B(new_n2605_), .Y(new_n2642_));
  NAND3X1  g2000(.A(new_n2642_), .B(new_n2601_), .C(new_n2599_), .Y(new_n2643_));
  NAND2X1  g2001(.A(new_n2607_), .B(new_n2605_), .Y(new_n2644_));
  AOI21X1  g2002(.A0(new_n2644_), .A1(new_n2643_), .B0(new_n2595_), .Y(new_n2645_));
  AND2X1   g2003(.A(new_n2588_), .B(new_n2586_), .Y(new_n2646_));
  AND2X1   g2004(.A(new_n2594_), .B(new_n2591_), .Y(new_n2647_));
  AND2X1   g2005(.A(new_n2647_), .B(new_n2589_), .Y(new_n2648_));
  OR4X1    g2006(.A(new_n2648_), .B(new_n2646_), .C(new_n2645_), .D(new_n2641_), .Y(new_n2649_));
  AOI21X1  g2007(.A0(new_n1348_), .A1(new_n1347_), .B0(new_n996_), .Y(new_n2650_));
  AOI21X1  g2008(.A0(new_n2225_), .A1(\in1[67] ), .B0(new_n2650_), .Y(new_n2651_));
  INVX1    g2009(.A(new_n2651_), .Y(new_n2652_));
  AOI21X1  g2010(.A0(new_n2063_), .A1(new_n1998_), .B0(new_n1708_), .Y(new_n2653_));
  AOI21X1  g2011(.A0(new_n2391_), .A1(\in3[67] ), .B0(new_n2653_), .Y(new_n2654_));
  NOR3X1   g2012(.A(new_n2061_), .B(new_n2060_), .C(new_n1719_), .Y(new_n2655_));
  AOI21X1  g2013(.A0(new_n2071_), .A1(\in2[66] ), .B0(new_n2655_), .Y(new_n2656_));
  NOR3X1   g2014(.A(new_n1286_), .B(new_n1284_), .C(new_n1006_), .Y(new_n2657_));
  AOI21X1  g2015(.A0(new_n1348_), .A1(new_n1347_), .B0(new_n995_), .Y(new_n2658_));
  NOR2X1   g2016(.A(new_n2658_), .B(new_n2657_), .Y(new_n2659_));
  INVX1    g2017(.A(new_n2659_), .Y(new_n2660_));
  OAI22X1  g2018(.A0(new_n2660_), .A1(new_n2656_), .B0(new_n2654_), .B1(new_n2652_), .Y(new_n2661_));
  AOI21X1  g2019(.A0(new_n2063_), .A1(new_n1998_), .B0(new_n1710_), .Y(new_n2662_));
  AOI21X1  g2020(.A0(new_n2391_), .A1(\in3[64] ), .B0(new_n2662_), .Y(new_n2663_));
  AOI21X1  g2021(.A0(new_n1348_), .A1(new_n1347_), .B0(new_n998_), .Y(new_n2664_));
  AOI21X1  g2022(.A0(new_n2225_), .A1(\in1[64] ), .B0(new_n2664_), .Y(new_n2665_));
  INVX1    g2023(.A(new_n2665_), .Y(new_n2666_));
  NOR3X1   g2024(.A(new_n1286_), .B(new_n1284_), .C(new_n1005_), .Y(new_n2667_));
  AOI21X1  g2025(.A0(new_n1348_), .A1(new_n1347_), .B0(new_n999_), .Y(new_n2668_));
  NOR2X1   g2026(.A(new_n2668_), .B(new_n2667_), .Y(new_n2669_));
  INVX1    g2027(.A(new_n2669_), .Y(new_n2670_));
  NOR3X1   g2028(.A(new_n2061_), .B(new_n2060_), .C(new_n1718_), .Y(new_n2671_));
  AOI21X1  g2029(.A0(new_n2071_), .A1(\in2[65] ), .B0(new_n2671_), .Y(new_n2672_));
  OAI22X1  g2030(.A0(new_n2672_), .A1(new_n2670_), .B0(new_n2666_), .B1(new_n2663_), .Y(new_n2673_));
  NOR2X1   g2031(.A(new_n2673_), .B(new_n2661_), .Y(new_n2674_));
  OAI21X1  g2032(.A0(new_n2649_), .A1(new_n2634_), .B0(new_n2674_), .Y(new_n2675_));
  AND2X1   g2033(.A(new_n2666_), .B(new_n2663_), .Y(new_n2676_));
  OAI21X1  g2034(.A0(new_n2672_), .A1(new_n2670_), .B0(new_n2676_), .Y(new_n2677_));
  AOI22X1  g2035(.A0(new_n2672_), .A1(new_n2670_), .B0(new_n2660_), .B1(new_n2656_), .Y(new_n2678_));
  AOI21X1  g2036(.A0(new_n2678_), .A1(new_n2677_), .B0(new_n2661_), .Y(new_n2679_));
  AOI21X1  g2037(.A0(new_n2654_), .A1(new_n2652_), .B0(new_n2679_), .Y(new_n2680_));
  NOR3X1   g2038(.A(new_n1286_), .B(new_n1284_), .C(new_n1026_), .Y(new_n2681_));
  AOI21X1  g2039(.A0(new_n1348_), .A1(new_n1347_), .B0(new_n1014_), .Y(new_n2682_));
  NOR2X1   g2040(.A(new_n2682_), .B(new_n2681_), .Y(new_n2683_));
  INVX1    g2041(.A(new_n2683_), .Y(new_n2684_));
  NOR3X1   g2042(.A(new_n2061_), .B(new_n2060_), .C(new_n1737_), .Y(new_n2685_));
  AOI21X1  g2043(.A0(new_n2071_), .A1(\in2[71] ), .B0(new_n2685_), .Y(new_n2686_));
  AOI21X1  g2044(.A0(new_n2063_), .A1(new_n1998_), .B0(new_n1725_), .Y(new_n2687_));
  AOI21X1  g2045(.A0(new_n2391_), .A1(\in3[70] ), .B0(new_n2687_), .Y(new_n2688_));
  AOI21X1  g2046(.A0(new_n1348_), .A1(new_n1347_), .B0(new_n1013_), .Y(new_n2689_));
  AOI21X1  g2047(.A0(new_n2225_), .A1(\in1[70] ), .B0(new_n2689_), .Y(new_n2690_));
  INVX1    g2048(.A(new_n2690_), .Y(new_n2691_));
  OAI22X1  g2049(.A0(new_n2691_), .A1(new_n2688_), .B0(new_n2686_), .B1(new_n2684_), .Y(new_n2692_));
  NOR3X1   g2050(.A(new_n1286_), .B(new_n1284_), .C(new_n1023_), .Y(new_n2693_));
  AOI21X1  g2051(.A0(new_n1348_), .A1(new_n1347_), .B0(new_n1017_), .Y(new_n2694_));
  NOR2X1   g2052(.A(new_n2694_), .B(new_n2693_), .Y(new_n2695_));
  INVX1    g2053(.A(new_n2695_), .Y(new_n2696_));
  NOR3X1   g2054(.A(new_n2061_), .B(new_n2060_), .C(new_n1734_), .Y(new_n2697_));
  AOI21X1  g2055(.A0(new_n2071_), .A1(\in2[69] ), .B0(new_n2697_), .Y(new_n2698_));
  AOI21X1  g2056(.A0(new_n1348_), .A1(new_n1347_), .B0(new_n1016_), .Y(new_n2699_));
  AOI21X1  g2057(.A0(new_n2225_), .A1(\in1[68] ), .B0(new_n2699_), .Y(new_n2700_));
  INVX1    g2058(.A(new_n2700_), .Y(new_n2701_));
  AOI21X1  g2059(.A0(new_n2063_), .A1(new_n1998_), .B0(new_n1728_), .Y(new_n2702_));
  AOI21X1  g2060(.A0(new_n2391_), .A1(\in3[68] ), .B0(new_n2702_), .Y(new_n2703_));
  OAI22X1  g2061(.A0(new_n2703_), .A1(new_n2701_), .B0(new_n2698_), .B1(new_n2696_), .Y(new_n2704_));
  OR2X1    g2062(.A(new_n2704_), .B(new_n2692_), .Y(new_n2705_));
  AOI21X1  g2063(.A0(new_n2680_), .A1(new_n2675_), .B0(new_n2705_), .Y(new_n2706_));
  AND2X1   g2064(.A(new_n2703_), .B(new_n2701_), .Y(new_n2707_));
  OAI21X1  g2065(.A0(new_n2698_), .A1(new_n2696_), .B0(new_n2707_), .Y(new_n2708_));
  NAND2X1  g2066(.A(new_n2698_), .B(new_n2696_), .Y(new_n2709_));
  AOI21X1  g2067(.A0(new_n2709_), .A1(new_n2708_), .B0(new_n2692_), .Y(new_n2710_));
  NOR2X1   g2068(.A(new_n2686_), .B(new_n2684_), .Y(new_n2711_));
  NAND2X1  g2069(.A(new_n2686_), .B(new_n2684_), .Y(new_n2712_));
  NAND2X1  g2070(.A(new_n2691_), .B(new_n2688_), .Y(new_n2713_));
  OAI21X1  g2071(.A0(new_n2713_), .A1(new_n2711_), .B0(new_n2712_), .Y(new_n2714_));
  OR2X1    g2072(.A(new_n2714_), .B(new_n2710_), .Y(new_n2715_));
  AOI21X1  g2073(.A0(new_n1348_), .A1(new_n1347_), .B0(new_n1033_), .Y(new_n2716_));
  AOI21X1  g2074(.A0(new_n2225_), .A1(\in1[75] ), .B0(new_n2716_), .Y(new_n2717_));
  INVX1    g2075(.A(new_n2717_), .Y(new_n2718_));
  AOI21X1  g2076(.A0(new_n2063_), .A1(new_n1998_), .B0(new_n1745_), .Y(new_n2719_));
  AOI21X1  g2077(.A0(new_n2391_), .A1(\in3[75] ), .B0(new_n2719_), .Y(new_n2720_));
  NOR3X1   g2078(.A(new_n2061_), .B(new_n2060_), .C(new_n1756_), .Y(new_n2721_));
  AOI21X1  g2079(.A0(new_n2071_), .A1(\in2[74] ), .B0(new_n2721_), .Y(new_n2722_));
  NOR3X1   g2080(.A(new_n1286_), .B(new_n1284_), .C(new_n1043_), .Y(new_n2723_));
  AOI21X1  g2081(.A0(new_n1348_), .A1(new_n1347_), .B0(new_n1032_), .Y(new_n2724_));
  NOR2X1   g2082(.A(new_n2724_), .B(new_n2723_), .Y(new_n2725_));
  INVX1    g2083(.A(new_n2725_), .Y(new_n2726_));
  OAI22X1  g2084(.A0(new_n2726_), .A1(new_n2722_), .B0(new_n2720_), .B1(new_n2718_), .Y(new_n2727_));
  NOR3X1   g2085(.A(new_n1286_), .B(new_n1284_), .C(new_n1042_), .Y(new_n2728_));
  AOI21X1  g2086(.A0(new_n1348_), .A1(new_n1347_), .B0(new_n1036_), .Y(new_n2729_));
  NOR2X1   g2087(.A(new_n2729_), .B(new_n2728_), .Y(new_n2730_));
  INVX1    g2088(.A(new_n2730_), .Y(new_n2731_));
  NOR3X1   g2089(.A(new_n2061_), .B(new_n2060_), .C(new_n1755_), .Y(new_n2732_));
  AOI21X1  g2090(.A0(new_n2071_), .A1(\in2[73] ), .B0(new_n2732_), .Y(new_n2733_));
  AOI21X1  g2091(.A0(new_n2063_), .A1(new_n1998_), .B0(new_n1747_), .Y(new_n2734_));
  AOI21X1  g2092(.A0(new_n2391_), .A1(\in3[72] ), .B0(new_n2734_), .Y(new_n2735_));
  AOI21X1  g2093(.A0(new_n1348_), .A1(new_n1347_), .B0(new_n1035_), .Y(new_n2736_));
  AOI21X1  g2094(.A0(new_n2225_), .A1(\in1[72] ), .B0(new_n2736_), .Y(new_n2737_));
  INVX1    g2095(.A(new_n2737_), .Y(new_n2738_));
  OAI22X1  g2096(.A0(new_n2738_), .A1(new_n2735_), .B0(new_n2733_), .B1(new_n2731_), .Y(new_n2739_));
  NOR2X1   g2097(.A(new_n2739_), .B(new_n2727_), .Y(new_n2740_));
  OAI21X1  g2098(.A0(new_n2715_), .A1(new_n2706_), .B0(new_n2740_), .Y(new_n2741_));
  AND2X1   g2099(.A(new_n2738_), .B(new_n2735_), .Y(new_n2742_));
  OAI21X1  g2100(.A0(new_n2733_), .A1(new_n2731_), .B0(new_n2742_), .Y(new_n2743_));
  AOI22X1  g2101(.A0(new_n2733_), .A1(new_n2731_), .B0(new_n2726_), .B1(new_n2722_), .Y(new_n2744_));
  AOI21X1  g2102(.A0(new_n2744_), .A1(new_n2743_), .B0(new_n2727_), .Y(new_n2745_));
  AOI21X1  g2103(.A0(new_n2720_), .A1(new_n2718_), .B0(new_n2745_), .Y(new_n2746_));
  NOR3X1   g2104(.A(new_n1286_), .B(new_n1284_), .C(new_n1063_), .Y(new_n2747_));
  AOI21X1  g2105(.A0(new_n1348_), .A1(new_n1347_), .B0(new_n1051_), .Y(new_n2748_));
  NOR2X1   g2106(.A(new_n2748_), .B(new_n2747_), .Y(new_n2749_));
  INVX1    g2107(.A(new_n2749_), .Y(new_n2750_));
  NOR3X1   g2108(.A(new_n2061_), .B(new_n2060_), .C(new_n1774_), .Y(new_n2751_));
  AOI21X1  g2109(.A0(new_n2071_), .A1(\in2[79] ), .B0(new_n2751_), .Y(new_n2752_));
  AOI21X1  g2110(.A0(new_n2063_), .A1(new_n1998_), .B0(new_n1762_), .Y(new_n2753_));
  AOI21X1  g2111(.A0(new_n2391_), .A1(\in3[78] ), .B0(new_n2753_), .Y(new_n2754_));
  AOI21X1  g2112(.A0(new_n1348_), .A1(new_n1347_), .B0(new_n1050_), .Y(new_n2755_));
  AOI21X1  g2113(.A0(new_n2225_), .A1(\in1[78] ), .B0(new_n2755_), .Y(new_n2756_));
  INVX1    g2114(.A(new_n2756_), .Y(new_n2757_));
  OAI22X1  g2115(.A0(new_n2757_), .A1(new_n2754_), .B0(new_n2752_), .B1(new_n2750_), .Y(new_n2758_));
  NOR3X1   g2116(.A(new_n1286_), .B(new_n1284_), .C(new_n1060_), .Y(new_n2759_));
  AOI21X1  g2117(.A0(new_n1348_), .A1(new_n1347_), .B0(new_n1054_), .Y(new_n2760_));
  NOR2X1   g2118(.A(new_n2760_), .B(new_n2759_), .Y(new_n2761_));
  INVX1    g2119(.A(new_n2761_), .Y(new_n2762_));
  NOR3X1   g2120(.A(new_n2061_), .B(new_n2060_), .C(new_n1771_), .Y(new_n2763_));
  AOI21X1  g2121(.A0(new_n2071_), .A1(\in2[77] ), .B0(new_n2763_), .Y(new_n2764_));
  AOI21X1  g2122(.A0(new_n1348_), .A1(new_n1347_), .B0(new_n1053_), .Y(new_n2765_));
  AOI21X1  g2123(.A0(new_n2225_), .A1(\in1[76] ), .B0(new_n2765_), .Y(new_n2766_));
  INVX1    g2124(.A(new_n2766_), .Y(new_n2767_));
  AOI21X1  g2125(.A0(new_n2063_), .A1(new_n1998_), .B0(new_n1765_), .Y(new_n2768_));
  AOI21X1  g2126(.A0(new_n2391_), .A1(\in3[76] ), .B0(new_n2768_), .Y(new_n2769_));
  OAI22X1  g2127(.A0(new_n2769_), .A1(new_n2767_), .B0(new_n2764_), .B1(new_n2762_), .Y(new_n2770_));
  OR2X1    g2128(.A(new_n2770_), .B(new_n2758_), .Y(new_n2771_));
  AOI21X1  g2129(.A0(new_n2746_), .A1(new_n2741_), .B0(new_n2771_), .Y(new_n2772_));
  AND2X1   g2130(.A(new_n2769_), .B(new_n2767_), .Y(new_n2773_));
  OAI21X1  g2131(.A0(new_n2764_), .A1(new_n2762_), .B0(new_n2773_), .Y(new_n2774_));
  NAND2X1  g2132(.A(new_n2764_), .B(new_n2762_), .Y(new_n2775_));
  AOI21X1  g2133(.A0(new_n2775_), .A1(new_n2774_), .B0(new_n2758_), .Y(new_n2776_));
  NOR2X1   g2134(.A(new_n2752_), .B(new_n2750_), .Y(new_n2777_));
  NAND2X1  g2135(.A(new_n2752_), .B(new_n2750_), .Y(new_n2778_));
  NAND2X1  g2136(.A(new_n2757_), .B(new_n2754_), .Y(new_n2779_));
  OAI21X1  g2137(.A0(new_n2779_), .A1(new_n2777_), .B0(new_n2778_), .Y(new_n2780_));
  OR2X1    g2138(.A(new_n2780_), .B(new_n2776_), .Y(new_n2781_));
  AOI21X1  g2139(.A0(new_n1348_), .A1(new_n1347_), .B0(new_n1070_), .Y(new_n2782_));
  AOI21X1  g2140(.A0(new_n2225_), .A1(\in1[83] ), .B0(new_n2782_), .Y(new_n2783_));
  INVX1    g2141(.A(new_n2783_), .Y(new_n2784_));
  AOI21X1  g2142(.A0(new_n2063_), .A1(new_n1998_), .B0(new_n1782_), .Y(new_n2785_));
  AOI21X1  g2143(.A0(new_n2391_), .A1(\in3[83] ), .B0(new_n2785_), .Y(new_n2786_));
  NOR3X1   g2144(.A(new_n2061_), .B(new_n2060_), .C(new_n1793_), .Y(new_n2787_));
  AOI21X1  g2145(.A0(new_n2071_), .A1(\in2[82] ), .B0(new_n2787_), .Y(new_n2788_));
  NOR3X1   g2146(.A(new_n1286_), .B(new_n1284_), .C(new_n1080_), .Y(new_n2789_));
  AOI21X1  g2147(.A0(new_n1348_), .A1(new_n1347_), .B0(new_n1069_), .Y(new_n2790_));
  NOR2X1   g2148(.A(new_n2790_), .B(new_n2789_), .Y(new_n2791_));
  INVX1    g2149(.A(new_n2791_), .Y(new_n2792_));
  OAI22X1  g2150(.A0(new_n2792_), .A1(new_n2788_), .B0(new_n2786_), .B1(new_n2784_), .Y(new_n2793_));
  AOI21X1  g2151(.A0(new_n2063_), .A1(new_n1998_), .B0(new_n1784_), .Y(new_n2794_));
  AOI21X1  g2152(.A0(new_n2391_), .A1(\in3[80] ), .B0(new_n2794_), .Y(new_n2795_));
  AOI21X1  g2153(.A0(new_n1348_), .A1(new_n1347_), .B0(new_n1072_), .Y(new_n2796_));
  AOI21X1  g2154(.A0(new_n2225_), .A1(\in1[80] ), .B0(new_n2796_), .Y(new_n2797_));
  INVX1    g2155(.A(new_n2797_), .Y(new_n2798_));
  NOR3X1   g2156(.A(new_n1286_), .B(new_n1284_), .C(new_n1079_), .Y(new_n2799_));
  AOI21X1  g2157(.A0(new_n1348_), .A1(new_n1347_), .B0(new_n1073_), .Y(new_n2800_));
  NOR2X1   g2158(.A(new_n2800_), .B(new_n2799_), .Y(new_n2801_));
  INVX1    g2159(.A(new_n2801_), .Y(new_n2802_));
  NOR3X1   g2160(.A(new_n2061_), .B(new_n2060_), .C(new_n1792_), .Y(new_n2803_));
  AOI21X1  g2161(.A0(new_n2071_), .A1(\in2[81] ), .B0(new_n2803_), .Y(new_n2804_));
  OAI22X1  g2162(.A0(new_n2804_), .A1(new_n2802_), .B0(new_n2798_), .B1(new_n2795_), .Y(new_n2805_));
  NOR2X1   g2163(.A(new_n2805_), .B(new_n2793_), .Y(new_n2806_));
  OAI21X1  g2164(.A0(new_n2781_), .A1(new_n2772_), .B0(new_n2806_), .Y(new_n2807_));
  AND2X1   g2165(.A(new_n2798_), .B(new_n2795_), .Y(new_n2808_));
  OAI21X1  g2166(.A0(new_n2804_), .A1(new_n2802_), .B0(new_n2808_), .Y(new_n2809_));
  AOI22X1  g2167(.A0(new_n2804_), .A1(new_n2802_), .B0(new_n2792_), .B1(new_n2788_), .Y(new_n2810_));
  AOI21X1  g2168(.A0(new_n2810_), .A1(new_n2809_), .B0(new_n2793_), .Y(new_n2811_));
  AOI21X1  g2169(.A0(new_n2786_), .A1(new_n2784_), .B0(new_n2811_), .Y(new_n2812_));
  NOR3X1   g2170(.A(new_n1286_), .B(new_n1284_), .C(new_n1100_), .Y(new_n2813_));
  AOI21X1  g2171(.A0(new_n1348_), .A1(new_n1347_), .B0(new_n1088_), .Y(new_n2814_));
  NOR2X1   g2172(.A(new_n2814_), .B(new_n2813_), .Y(new_n2815_));
  INVX1    g2173(.A(new_n2815_), .Y(new_n2816_));
  NOR3X1   g2174(.A(new_n2061_), .B(new_n2060_), .C(new_n1811_), .Y(new_n2817_));
  AOI21X1  g2175(.A0(new_n2071_), .A1(\in2[87] ), .B0(new_n2817_), .Y(new_n2818_));
  AOI21X1  g2176(.A0(new_n2063_), .A1(new_n1998_), .B0(new_n1799_), .Y(new_n2819_));
  AOI21X1  g2177(.A0(new_n2391_), .A1(\in3[86] ), .B0(new_n2819_), .Y(new_n2820_));
  AOI21X1  g2178(.A0(new_n1348_), .A1(new_n1347_), .B0(new_n1087_), .Y(new_n2821_));
  AOI21X1  g2179(.A0(new_n2225_), .A1(\in1[86] ), .B0(new_n2821_), .Y(new_n2822_));
  INVX1    g2180(.A(new_n2822_), .Y(new_n2823_));
  OAI22X1  g2181(.A0(new_n2823_), .A1(new_n2820_), .B0(new_n2818_), .B1(new_n2816_), .Y(new_n2824_));
  NOR3X1   g2182(.A(new_n1286_), .B(new_n1284_), .C(new_n1097_), .Y(new_n2825_));
  AOI21X1  g2183(.A0(new_n1348_), .A1(new_n1347_), .B0(new_n1091_), .Y(new_n2826_));
  NOR2X1   g2184(.A(new_n2826_), .B(new_n2825_), .Y(new_n2827_));
  INVX1    g2185(.A(new_n2827_), .Y(new_n2828_));
  NOR3X1   g2186(.A(new_n2061_), .B(new_n2060_), .C(new_n1808_), .Y(new_n2829_));
  AOI21X1  g2187(.A0(new_n2071_), .A1(\in2[85] ), .B0(new_n2829_), .Y(new_n2830_));
  AOI21X1  g2188(.A0(new_n1348_), .A1(new_n1347_), .B0(new_n1090_), .Y(new_n2831_));
  AOI21X1  g2189(.A0(new_n2225_), .A1(\in1[84] ), .B0(new_n2831_), .Y(new_n2832_));
  INVX1    g2190(.A(new_n2832_), .Y(new_n2833_));
  AOI21X1  g2191(.A0(new_n2063_), .A1(new_n1998_), .B0(new_n1802_), .Y(new_n2834_));
  AOI21X1  g2192(.A0(new_n2391_), .A1(\in3[84] ), .B0(new_n2834_), .Y(new_n2835_));
  OAI22X1  g2193(.A0(new_n2835_), .A1(new_n2833_), .B0(new_n2830_), .B1(new_n2828_), .Y(new_n2836_));
  OR2X1    g2194(.A(new_n2836_), .B(new_n2824_), .Y(new_n2837_));
  AOI21X1  g2195(.A0(new_n2812_), .A1(new_n2807_), .B0(new_n2837_), .Y(new_n2838_));
  AND2X1   g2196(.A(new_n2835_), .B(new_n2833_), .Y(new_n2839_));
  OAI21X1  g2197(.A0(new_n2830_), .A1(new_n2828_), .B0(new_n2839_), .Y(new_n2840_));
  NAND2X1  g2198(.A(new_n2830_), .B(new_n2828_), .Y(new_n2841_));
  AOI21X1  g2199(.A0(new_n2841_), .A1(new_n2840_), .B0(new_n2824_), .Y(new_n2842_));
  NOR2X1   g2200(.A(new_n2818_), .B(new_n2816_), .Y(new_n2843_));
  NAND2X1  g2201(.A(new_n2818_), .B(new_n2816_), .Y(new_n2844_));
  NAND2X1  g2202(.A(new_n2823_), .B(new_n2820_), .Y(new_n2845_));
  OAI21X1  g2203(.A0(new_n2845_), .A1(new_n2843_), .B0(new_n2844_), .Y(new_n2846_));
  OR2X1    g2204(.A(new_n2846_), .B(new_n2842_), .Y(new_n2847_));
  AOI21X1  g2205(.A0(new_n1348_), .A1(new_n1347_), .B0(new_n1107_), .Y(new_n2848_));
  AOI21X1  g2206(.A0(new_n2225_), .A1(\in1[91] ), .B0(new_n2848_), .Y(new_n2849_));
  INVX1    g2207(.A(new_n2849_), .Y(new_n2850_));
  AOI21X1  g2208(.A0(new_n2063_), .A1(new_n1998_), .B0(new_n1819_), .Y(new_n2851_));
  AOI21X1  g2209(.A0(new_n2391_), .A1(\in3[91] ), .B0(new_n2851_), .Y(new_n2852_));
  NOR3X1   g2210(.A(new_n2061_), .B(new_n2060_), .C(new_n1830_), .Y(new_n2853_));
  AOI21X1  g2211(.A0(new_n2071_), .A1(\in2[90] ), .B0(new_n2853_), .Y(new_n2854_));
  NOR3X1   g2212(.A(new_n1286_), .B(new_n1284_), .C(new_n1117_), .Y(new_n2855_));
  AOI21X1  g2213(.A0(new_n1348_), .A1(new_n1347_), .B0(new_n1106_), .Y(new_n2856_));
  NOR2X1   g2214(.A(new_n2856_), .B(new_n2855_), .Y(new_n2857_));
  INVX1    g2215(.A(new_n2857_), .Y(new_n2858_));
  OAI22X1  g2216(.A0(new_n2858_), .A1(new_n2854_), .B0(new_n2852_), .B1(new_n2850_), .Y(new_n2859_));
  NOR3X1   g2217(.A(new_n1286_), .B(new_n1284_), .C(new_n1116_), .Y(new_n2860_));
  AOI21X1  g2218(.A0(new_n1348_), .A1(new_n1347_), .B0(new_n1110_), .Y(new_n2861_));
  NOR2X1   g2219(.A(new_n2861_), .B(new_n2860_), .Y(new_n2862_));
  INVX1    g2220(.A(new_n2862_), .Y(new_n2863_));
  NOR3X1   g2221(.A(new_n2061_), .B(new_n2060_), .C(new_n1829_), .Y(new_n2864_));
  AOI21X1  g2222(.A0(new_n2071_), .A1(\in2[89] ), .B0(new_n2864_), .Y(new_n2865_));
  AOI21X1  g2223(.A0(new_n2063_), .A1(new_n1998_), .B0(new_n1821_), .Y(new_n2866_));
  AOI21X1  g2224(.A0(new_n2391_), .A1(\in3[88] ), .B0(new_n2866_), .Y(new_n2867_));
  AOI21X1  g2225(.A0(new_n1348_), .A1(new_n1347_), .B0(new_n1109_), .Y(new_n2868_));
  AOI21X1  g2226(.A0(new_n2225_), .A1(\in1[88] ), .B0(new_n2868_), .Y(new_n2869_));
  INVX1    g2227(.A(new_n2869_), .Y(new_n2870_));
  OAI22X1  g2228(.A0(new_n2870_), .A1(new_n2867_), .B0(new_n2865_), .B1(new_n2863_), .Y(new_n2871_));
  NOR2X1   g2229(.A(new_n2871_), .B(new_n2859_), .Y(new_n2872_));
  OAI21X1  g2230(.A0(new_n2847_), .A1(new_n2838_), .B0(new_n2872_), .Y(new_n2873_));
  AND2X1   g2231(.A(new_n2870_), .B(new_n2867_), .Y(new_n2874_));
  OAI21X1  g2232(.A0(new_n2865_), .A1(new_n2863_), .B0(new_n2874_), .Y(new_n2875_));
  AOI22X1  g2233(.A0(new_n2865_), .A1(new_n2863_), .B0(new_n2858_), .B1(new_n2854_), .Y(new_n2876_));
  AOI21X1  g2234(.A0(new_n2876_), .A1(new_n2875_), .B0(new_n2859_), .Y(new_n2877_));
  AOI21X1  g2235(.A0(new_n2852_), .A1(new_n2850_), .B0(new_n2877_), .Y(new_n2878_));
  NOR3X1   g2236(.A(new_n1286_), .B(new_n1284_), .C(new_n1137_), .Y(new_n2879_));
  AOI21X1  g2237(.A0(new_n1348_), .A1(new_n1347_), .B0(new_n1125_), .Y(new_n2880_));
  NOR2X1   g2238(.A(new_n2880_), .B(new_n2879_), .Y(new_n2881_));
  INVX1    g2239(.A(new_n2881_), .Y(new_n2882_));
  NOR3X1   g2240(.A(new_n2061_), .B(new_n2060_), .C(new_n1848_), .Y(new_n2883_));
  AOI21X1  g2241(.A0(new_n2071_), .A1(\in2[95] ), .B0(new_n2883_), .Y(new_n2884_));
  AOI21X1  g2242(.A0(new_n2063_), .A1(new_n1998_), .B0(new_n1836_), .Y(new_n2885_));
  AOI21X1  g2243(.A0(new_n2391_), .A1(\in3[94] ), .B0(new_n2885_), .Y(new_n2886_));
  AOI21X1  g2244(.A0(new_n1348_), .A1(new_n1347_), .B0(new_n1124_), .Y(new_n2887_));
  AOI21X1  g2245(.A0(new_n2225_), .A1(\in1[94] ), .B0(new_n2887_), .Y(new_n2888_));
  INVX1    g2246(.A(new_n2888_), .Y(new_n2889_));
  OAI22X1  g2247(.A0(new_n2889_), .A1(new_n2886_), .B0(new_n2884_), .B1(new_n2882_), .Y(new_n2890_));
  NOR3X1   g2248(.A(new_n1286_), .B(new_n1284_), .C(new_n1134_), .Y(new_n2891_));
  AOI21X1  g2249(.A0(new_n1348_), .A1(new_n1347_), .B0(new_n1128_), .Y(new_n2892_));
  NOR2X1   g2250(.A(new_n2892_), .B(new_n2891_), .Y(new_n2893_));
  INVX1    g2251(.A(new_n2893_), .Y(new_n2894_));
  NOR3X1   g2252(.A(new_n2061_), .B(new_n2060_), .C(new_n1845_), .Y(new_n2895_));
  AOI21X1  g2253(.A0(new_n2071_), .A1(\in2[93] ), .B0(new_n2895_), .Y(new_n2896_));
  AOI21X1  g2254(.A0(new_n1348_), .A1(new_n1347_), .B0(new_n1127_), .Y(new_n2897_));
  AOI21X1  g2255(.A0(new_n2225_), .A1(\in1[92] ), .B0(new_n2897_), .Y(new_n2898_));
  INVX1    g2256(.A(new_n2898_), .Y(new_n2899_));
  AOI21X1  g2257(.A0(new_n2063_), .A1(new_n1998_), .B0(new_n1839_), .Y(new_n2900_));
  AOI21X1  g2258(.A0(new_n2391_), .A1(\in3[92] ), .B0(new_n2900_), .Y(new_n2901_));
  OAI22X1  g2259(.A0(new_n2901_), .A1(new_n2899_), .B0(new_n2896_), .B1(new_n2894_), .Y(new_n2902_));
  OR2X1    g2260(.A(new_n2902_), .B(new_n2890_), .Y(new_n2903_));
  AOI21X1  g2261(.A0(new_n2878_), .A1(new_n2873_), .B0(new_n2903_), .Y(new_n2904_));
  AND2X1   g2262(.A(new_n2901_), .B(new_n2899_), .Y(new_n2905_));
  OAI21X1  g2263(.A0(new_n2896_), .A1(new_n2894_), .B0(new_n2905_), .Y(new_n2906_));
  NAND2X1  g2264(.A(new_n2896_), .B(new_n2894_), .Y(new_n2907_));
  AOI21X1  g2265(.A0(new_n2907_), .A1(new_n2906_), .B0(new_n2890_), .Y(new_n2908_));
  NOR2X1   g2266(.A(new_n2884_), .B(new_n2882_), .Y(new_n2909_));
  NAND2X1  g2267(.A(new_n2884_), .B(new_n2882_), .Y(new_n2910_));
  NAND2X1  g2268(.A(new_n2889_), .B(new_n2886_), .Y(new_n2911_));
  OAI21X1  g2269(.A0(new_n2911_), .A1(new_n2909_), .B0(new_n2910_), .Y(new_n2912_));
  OR2X1    g2270(.A(new_n2912_), .B(new_n2908_), .Y(new_n2913_));
  AOI21X1  g2271(.A0(new_n1348_), .A1(new_n1347_), .B0(new_n1144_), .Y(new_n2914_));
  AOI21X1  g2272(.A0(new_n2225_), .A1(\in1[99] ), .B0(new_n2914_), .Y(new_n2915_));
  INVX1    g2273(.A(new_n2915_), .Y(new_n2916_));
  AOI21X1  g2274(.A0(new_n2063_), .A1(new_n1998_), .B0(new_n1856_), .Y(new_n2917_));
  AOI21X1  g2275(.A0(new_n2391_), .A1(\in3[99] ), .B0(new_n2917_), .Y(new_n2918_));
  NOR3X1   g2276(.A(new_n2061_), .B(new_n2060_), .C(new_n1867_), .Y(new_n2919_));
  AOI21X1  g2277(.A0(new_n2071_), .A1(\in2[98] ), .B0(new_n2919_), .Y(new_n2920_));
  NOR3X1   g2278(.A(new_n1286_), .B(new_n1284_), .C(new_n1154_), .Y(new_n2921_));
  AOI21X1  g2279(.A0(new_n1348_), .A1(new_n1347_), .B0(new_n1143_), .Y(new_n2922_));
  NOR2X1   g2280(.A(new_n2922_), .B(new_n2921_), .Y(new_n2923_));
  INVX1    g2281(.A(new_n2923_), .Y(new_n2924_));
  OAI22X1  g2282(.A0(new_n2924_), .A1(new_n2920_), .B0(new_n2918_), .B1(new_n2916_), .Y(new_n2925_));
  AOI21X1  g2283(.A0(new_n2063_), .A1(new_n1998_), .B0(new_n1858_), .Y(new_n2926_));
  AOI21X1  g2284(.A0(new_n2391_), .A1(\in3[96] ), .B0(new_n2926_), .Y(new_n2927_));
  AOI21X1  g2285(.A0(new_n1348_), .A1(new_n1347_), .B0(new_n1146_), .Y(new_n2928_));
  AOI21X1  g2286(.A0(new_n2225_), .A1(\in1[96] ), .B0(new_n2928_), .Y(new_n2929_));
  INVX1    g2287(.A(new_n2929_), .Y(new_n2930_));
  NOR3X1   g2288(.A(new_n1286_), .B(new_n1284_), .C(new_n1153_), .Y(new_n2931_));
  AOI21X1  g2289(.A0(new_n1348_), .A1(new_n1347_), .B0(new_n1147_), .Y(new_n2932_));
  NOR2X1   g2290(.A(new_n2932_), .B(new_n2931_), .Y(new_n2933_));
  INVX1    g2291(.A(new_n2933_), .Y(new_n2934_));
  NOR3X1   g2292(.A(new_n2061_), .B(new_n2060_), .C(new_n1866_), .Y(new_n2935_));
  AOI21X1  g2293(.A0(new_n2071_), .A1(\in2[97] ), .B0(new_n2935_), .Y(new_n2936_));
  OAI22X1  g2294(.A0(new_n2936_), .A1(new_n2934_), .B0(new_n2930_), .B1(new_n2927_), .Y(new_n2937_));
  NOR2X1   g2295(.A(new_n2937_), .B(new_n2925_), .Y(new_n2938_));
  OAI21X1  g2296(.A0(new_n2913_), .A1(new_n2904_), .B0(new_n2938_), .Y(new_n2939_));
  AND2X1   g2297(.A(new_n2930_), .B(new_n2927_), .Y(new_n2940_));
  OAI21X1  g2298(.A0(new_n2936_), .A1(new_n2934_), .B0(new_n2940_), .Y(new_n2941_));
  AOI22X1  g2299(.A0(new_n2936_), .A1(new_n2934_), .B0(new_n2924_), .B1(new_n2920_), .Y(new_n2942_));
  AOI21X1  g2300(.A0(new_n2942_), .A1(new_n2941_), .B0(new_n2925_), .Y(new_n2943_));
  AOI21X1  g2301(.A0(new_n2918_), .A1(new_n2916_), .B0(new_n2943_), .Y(new_n2944_));
  NOR3X1   g2302(.A(new_n1286_), .B(new_n1284_), .C(new_n1174_), .Y(new_n2945_));
  AOI21X1  g2303(.A0(new_n1348_), .A1(new_n1347_), .B0(new_n1162_), .Y(new_n2946_));
  NOR2X1   g2304(.A(new_n2946_), .B(new_n2945_), .Y(new_n2947_));
  INVX1    g2305(.A(new_n2947_), .Y(new_n2948_));
  NOR3X1   g2306(.A(new_n2061_), .B(new_n2060_), .C(new_n1885_), .Y(new_n2949_));
  AOI21X1  g2307(.A0(new_n2071_), .A1(\in2[103] ), .B0(new_n2949_), .Y(new_n2950_));
  AOI21X1  g2308(.A0(new_n2063_), .A1(new_n1998_), .B0(new_n1873_), .Y(new_n2951_));
  AOI21X1  g2309(.A0(new_n2391_), .A1(\in3[102] ), .B0(new_n2951_), .Y(new_n2952_));
  AOI21X1  g2310(.A0(new_n1348_), .A1(new_n1347_), .B0(new_n1161_), .Y(new_n2953_));
  AOI21X1  g2311(.A0(new_n2225_), .A1(\in1[102] ), .B0(new_n2953_), .Y(new_n2954_));
  INVX1    g2312(.A(new_n2954_), .Y(new_n2955_));
  OAI22X1  g2313(.A0(new_n2955_), .A1(new_n2952_), .B0(new_n2950_), .B1(new_n2948_), .Y(new_n2956_));
  NOR3X1   g2314(.A(new_n1286_), .B(new_n1284_), .C(new_n1171_), .Y(new_n2957_));
  AOI21X1  g2315(.A0(new_n1348_), .A1(new_n1347_), .B0(new_n1165_), .Y(new_n2958_));
  NOR2X1   g2316(.A(new_n2958_), .B(new_n2957_), .Y(new_n2959_));
  INVX1    g2317(.A(new_n2959_), .Y(new_n2960_));
  NOR3X1   g2318(.A(new_n2061_), .B(new_n2060_), .C(new_n1882_), .Y(new_n2961_));
  AOI21X1  g2319(.A0(new_n2071_), .A1(\in2[101] ), .B0(new_n2961_), .Y(new_n2962_));
  AOI21X1  g2320(.A0(new_n1348_), .A1(new_n1347_), .B0(new_n1164_), .Y(new_n2963_));
  AOI21X1  g2321(.A0(new_n2225_), .A1(\in1[100] ), .B0(new_n2963_), .Y(new_n2964_));
  INVX1    g2322(.A(new_n2964_), .Y(new_n2965_));
  AOI21X1  g2323(.A0(new_n2063_), .A1(new_n1998_), .B0(new_n1876_), .Y(new_n2966_));
  AOI21X1  g2324(.A0(new_n2391_), .A1(\in3[100] ), .B0(new_n2966_), .Y(new_n2967_));
  OAI22X1  g2325(.A0(new_n2967_), .A1(new_n2965_), .B0(new_n2962_), .B1(new_n2960_), .Y(new_n2968_));
  OR2X1    g2326(.A(new_n2968_), .B(new_n2956_), .Y(new_n2969_));
  AOI21X1  g2327(.A0(new_n2944_), .A1(new_n2939_), .B0(new_n2969_), .Y(new_n2970_));
  AND2X1   g2328(.A(new_n2967_), .B(new_n2965_), .Y(new_n2971_));
  OAI21X1  g2329(.A0(new_n2962_), .A1(new_n2960_), .B0(new_n2971_), .Y(new_n2972_));
  NAND2X1  g2330(.A(new_n2962_), .B(new_n2960_), .Y(new_n2973_));
  AOI21X1  g2331(.A0(new_n2973_), .A1(new_n2972_), .B0(new_n2956_), .Y(new_n2974_));
  NOR2X1   g2332(.A(new_n2950_), .B(new_n2948_), .Y(new_n2975_));
  NAND2X1  g2333(.A(new_n2950_), .B(new_n2948_), .Y(new_n2976_));
  NAND2X1  g2334(.A(new_n2955_), .B(new_n2952_), .Y(new_n2977_));
  OAI21X1  g2335(.A0(new_n2977_), .A1(new_n2975_), .B0(new_n2976_), .Y(new_n2978_));
  OR2X1    g2336(.A(new_n2978_), .B(new_n2974_), .Y(new_n2979_));
  AOI21X1  g2337(.A0(new_n1348_), .A1(new_n1347_), .B0(new_n1181_), .Y(new_n2980_));
  AOI21X1  g2338(.A0(new_n2225_), .A1(\in1[107] ), .B0(new_n2980_), .Y(new_n2981_));
  INVX1    g2339(.A(new_n2981_), .Y(new_n2982_));
  AOI21X1  g2340(.A0(new_n2063_), .A1(new_n1998_), .B0(new_n1893_), .Y(new_n2983_));
  AOI21X1  g2341(.A0(new_n2391_), .A1(\in3[107] ), .B0(new_n2983_), .Y(new_n2984_));
  NOR3X1   g2342(.A(new_n2061_), .B(new_n2060_), .C(new_n1904_), .Y(new_n2985_));
  AOI21X1  g2343(.A0(new_n2071_), .A1(\in2[106] ), .B0(new_n2985_), .Y(new_n2986_));
  NOR3X1   g2344(.A(new_n1286_), .B(new_n1284_), .C(new_n1191_), .Y(new_n2987_));
  AOI21X1  g2345(.A0(new_n1348_), .A1(new_n1347_), .B0(new_n1180_), .Y(new_n2988_));
  NOR2X1   g2346(.A(new_n2988_), .B(new_n2987_), .Y(new_n2989_));
  INVX1    g2347(.A(new_n2989_), .Y(new_n2990_));
  OAI22X1  g2348(.A0(new_n2990_), .A1(new_n2986_), .B0(new_n2984_), .B1(new_n2982_), .Y(new_n2991_));
  NOR3X1   g2349(.A(new_n1286_), .B(new_n1284_), .C(new_n1190_), .Y(new_n2992_));
  AOI21X1  g2350(.A0(new_n1348_), .A1(new_n1347_), .B0(new_n1184_), .Y(new_n2993_));
  NOR2X1   g2351(.A(new_n2993_), .B(new_n2992_), .Y(new_n2994_));
  INVX1    g2352(.A(new_n2994_), .Y(new_n2995_));
  NOR3X1   g2353(.A(new_n2061_), .B(new_n2060_), .C(new_n1903_), .Y(new_n2996_));
  AOI21X1  g2354(.A0(new_n2071_), .A1(\in2[105] ), .B0(new_n2996_), .Y(new_n2997_));
  AOI21X1  g2355(.A0(new_n2063_), .A1(new_n1998_), .B0(new_n1895_), .Y(new_n2998_));
  AOI21X1  g2356(.A0(new_n2391_), .A1(\in3[104] ), .B0(new_n2998_), .Y(new_n2999_));
  AOI21X1  g2357(.A0(new_n1348_), .A1(new_n1347_), .B0(new_n1183_), .Y(new_n3000_));
  AOI21X1  g2358(.A0(new_n2225_), .A1(\in1[104] ), .B0(new_n3000_), .Y(new_n3001_));
  INVX1    g2359(.A(new_n3001_), .Y(new_n3002_));
  OAI22X1  g2360(.A0(new_n3002_), .A1(new_n2999_), .B0(new_n2997_), .B1(new_n2995_), .Y(new_n3003_));
  NOR2X1   g2361(.A(new_n3003_), .B(new_n2991_), .Y(new_n3004_));
  OAI21X1  g2362(.A0(new_n2979_), .A1(new_n2970_), .B0(new_n3004_), .Y(new_n3005_));
  AND2X1   g2363(.A(new_n3002_), .B(new_n2999_), .Y(new_n3006_));
  OAI21X1  g2364(.A0(new_n2997_), .A1(new_n2995_), .B0(new_n3006_), .Y(new_n3007_));
  AOI22X1  g2365(.A0(new_n2997_), .A1(new_n2995_), .B0(new_n2990_), .B1(new_n2986_), .Y(new_n3008_));
  AOI21X1  g2366(.A0(new_n3008_), .A1(new_n3007_), .B0(new_n2991_), .Y(new_n3009_));
  AOI21X1  g2367(.A0(new_n2984_), .A1(new_n2982_), .B0(new_n3009_), .Y(new_n3010_));
  NOR3X1   g2368(.A(new_n1286_), .B(new_n1284_), .C(new_n1211_), .Y(new_n3011_));
  AOI21X1  g2369(.A0(new_n1348_), .A1(new_n1347_), .B0(new_n1199_), .Y(new_n3012_));
  NOR2X1   g2370(.A(new_n3012_), .B(new_n3011_), .Y(new_n3013_));
  INVX1    g2371(.A(new_n3013_), .Y(new_n3014_));
  NOR3X1   g2372(.A(new_n2061_), .B(new_n2060_), .C(new_n1922_), .Y(new_n3015_));
  AOI21X1  g2373(.A0(new_n2071_), .A1(\in2[111] ), .B0(new_n3015_), .Y(new_n3016_));
  AOI21X1  g2374(.A0(new_n2063_), .A1(new_n1998_), .B0(new_n1910_), .Y(new_n3017_));
  AOI21X1  g2375(.A0(new_n2391_), .A1(\in3[110] ), .B0(new_n3017_), .Y(new_n3018_));
  AOI21X1  g2376(.A0(new_n1348_), .A1(new_n1347_), .B0(new_n1198_), .Y(new_n3019_));
  AOI21X1  g2377(.A0(new_n2225_), .A1(\in1[110] ), .B0(new_n3019_), .Y(new_n3020_));
  INVX1    g2378(.A(new_n3020_), .Y(new_n3021_));
  OAI22X1  g2379(.A0(new_n3021_), .A1(new_n3018_), .B0(new_n3016_), .B1(new_n3014_), .Y(new_n3022_));
  NOR3X1   g2380(.A(new_n1286_), .B(new_n1284_), .C(new_n1208_), .Y(new_n3023_));
  AOI21X1  g2381(.A0(new_n1348_), .A1(new_n1347_), .B0(new_n1202_), .Y(new_n3024_));
  NOR2X1   g2382(.A(new_n3024_), .B(new_n3023_), .Y(new_n3025_));
  INVX1    g2383(.A(new_n3025_), .Y(new_n3026_));
  NOR3X1   g2384(.A(new_n2061_), .B(new_n2060_), .C(new_n1919_), .Y(new_n3027_));
  AOI21X1  g2385(.A0(new_n2071_), .A1(\in2[109] ), .B0(new_n3027_), .Y(new_n3028_));
  AOI21X1  g2386(.A0(new_n1348_), .A1(new_n1347_), .B0(new_n1201_), .Y(new_n3029_));
  AOI21X1  g2387(.A0(new_n2225_), .A1(\in1[108] ), .B0(new_n3029_), .Y(new_n3030_));
  INVX1    g2388(.A(new_n3030_), .Y(new_n3031_));
  AOI21X1  g2389(.A0(new_n2063_), .A1(new_n1998_), .B0(new_n1913_), .Y(new_n3032_));
  AOI21X1  g2390(.A0(new_n2391_), .A1(\in3[108] ), .B0(new_n3032_), .Y(new_n3033_));
  OAI22X1  g2391(.A0(new_n3033_), .A1(new_n3031_), .B0(new_n3028_), .B1(new_n3026_), .Y(new_n3034_));
  OR2X1    g2392(.A(new_n3034_), .B(new_n3022_), .Y(new_n3035_));
  AOI21X1  g2393(.A0(new_n3010_), .A1(new_n3005_), .B0(new_n3035_), .Y(new_n3036_));
  AND2X1   g2394(.A(new_n3033_), .B(new_n3031_), .Y(new_n3037_));
  OAI21X1  g2395(.A0(new_n3028_), .A1(new_n3026_), .B0(new_n3037_), .Y(new_n3038_));
  NAND2X1  g2396(.A(new_n3028_), .B(new_n3026_), .Y(new_n3039_));
  AOI21X1  g2397(.A0(new_n3039_), .A1(new_n3038_), .B0(new_n3022_), .Y(new_n3040_));
  NOR2X1   g2398(.A(new_n3016_), .B(new_n3014_), .Y(new_n3041_));
  NAND2X1  g2399(.A(new_n3016_), .B(new_n3014_), .Y(new_n3042_));
  NAND2X1  g2400(.A(new_n3021_), .B(new_n3018_), .Y(new_n3043_));
  OAI21X1  g2401(.A0(new_n3043_), .A1(new_n3041_), .B0(new_n3042_), .Y(new_n3044_));
  OR2X1    g2402(.A(new_n3044_), .B(new_n3040_), .Y(new_n3045_));
  AOI21X1  g2403(.A0(new_n1348_), .A1(new_n1347_), .B0(new_n1218_), .Y(new_n3046_));
  AOI21X1  g2404(.A0(new_n2225_), .A1(\in1[115] ), .B0(new_n3046_), .Y(new_n3047_));
  INVX1    g2405(.A(new_n3047_), .Y(new_n3048_));
  AOI21X1  g2406(.A0(new_n2063_), .A1(new_n1998_), .B0(new_n1930_), .Y(new_n3049_));
  AOI21X1  g2407(.A0(new_n2391_), .A1(\in3[115] ), .B0(new_n3049_), .Y(new_n3050_));
  NOR3X1   g2408(.A(new_n2061_), .B(new_n2060_), .C(new_n1941_), .Y(new_n3051_));
  AOI21X1  g2409(.A0(new_n2071_), .A1(\in2[114] ), .B0(new_n3051_), .Y(new_n3052_));
  NOR3X1   g2410(.A(new_n1286_), .B(new_n1284_), .C(new_n1228_), .Y(new_n3053_));
  AOI21X1  g2411(.A0(new_n1348_), .A1(new_n1347_), .B0(new_n1217_), .Y(new_n3054_));
  NOR2X1   g2412(.A(new_n3054_), .B(new_n3053_), .Y(new_n3055_));
  INVX1    g2413(.A(new_n3055_), .Y(new_n3056_));
  OAI22X1  g2414(.A0(new_n3056_), .A1(new_n3052_), .B0(new_n3050_), .B1(new_n3048_), .Y(new_n3057_));
  AOI21X1  g2415(.A0(new_n2063_), .A1(new_n1998_), .B0(new_n1932_), .Y(new_n3058_));
  AOI21X1  g2416(.A0(new_n2391_), .A1(\in3[112] ), .B0(new_n3058_), .Y(new_n3059_));
  AOI21X1  g2417(.A0(new_n1348_), .A1(new_n1347_), .B0(new_n1220_), .Y(new_n3060_));
  AOI21X1  g2418(.A0(new_n2225_), .A1(\in1[112] ), .B0(new_n3060_), .Y(new_n3061_));
  INVX1    g2419(.A(new_n3061_), .Y(new_n3062_));
  NOR3X1   g2420(.A(new_n1286_), .B(new_n1284_), .C(new_n1227_), .Y(new_n3063_));
  AOI21X1  g2421(.A0(new_n1348_), .A1(new_n1347_), .B0(new_n1221_), .Y(new_n3064_));
  NOR2X1   g2422(.A(new_n3064_), .B(new_n3063_), .Y(new_n3065_));
  INVX1    g2423(.A(new_n3065_), .Y(new_n3066_));
  NOR3X1   g2424(.A(new_n2061_), .B(new_n2060_), .C(new_n1940_), .Y(new_n3067_));
  AOI21X1  g2425(.A0(new_n2071_), .A1(\in2[113] ), .B0(new_n3067_), .Y(new_n3068_));
  OAI22X1  g2426(.A0(new_n3068_), .A1(new_n3066_), .B0(new_n3062_), .B1(new_n3059_), .Y(new_n3069_));
  NOR2X1   g2427(.A(new_n3069_), .B(new_n3057_), .Y(new_n3070_));
  OAI21X1  g2428(.A0(new_n3045_), .A1(new_n3036_), .B0(new_n3070_), .Y(new_n3071_));
  AND2X1   g2429(.A(new_n3062_), .B(new_n3059_), .Y(new_n3072_));
  OAI21X1  g2430(.A0(new_n3068_), .A1(new_n3066_), .B0(new_n3072_), .Y(new_n3073_));
  AOI22X1  g2431(.A0(new_n3068_), .A1(new_n3066_), .B0(new_n3056_), .B1(new_n3052_), .Y(new_n3074_));
  AOI21X1  g2432(.A0(new_n3074_), .A1(new_n3073_), .B0(new_n3057_), .Y(new_n3075_));
  AOI21X1  g2433(.A0(new_n3050_), .A1(new_n3048_), .B0(new_n3075_), .Y(new_n3076_));
  NOR3X1   g2434(.A(new_n1286_), .B(new_n1284_), .C(new_n1248_), .Y(new_n3077_));
  AOI21X1  g2435(.A0(new_n1348_), .A1(new_n1347_), .B0(new_n1236_), .Y(new_n3078_));
  NOR2X1   g2436(.A(new_n3078_), .B(new_n3077_), .Y(new_n3079_));
  INVX1    g2437(.A(new_n3079_), .Y(new_n3080_));
  NOR3X1   g2438(.A(new_n2061_), .B(new_n2060_), .C(new_n1959_), .Y(new_n3081_));
  AOI21X1  g2439(.A0(new_n2071_), .A1(\in2[119] ), .B0(new_n3081_), .Y(new_n3082_));
  AOI21X1  g2440(.A0(new_n2063_), .A1(new_n1998_), .B0(new_n1947_), .Y(new_n3083_));
  AOI21X1  g2441(.A0(new_n2391_), .A1(\in3[118] ), .B0(new_n3083_), .Y(new_n3084_));
  AOI21X1  g2442(.A0(new_n1348_), .A1(new_n1347_), .B0(new_n1235_), .Y(new_n3085_));
  AOI21X1  g2443(.A0(new_n2225_), .A1(\in1[118] ), .B0(new_n3085_), .Y(new_n3086_));
  INVX1    g2444(.A(new_n3086_), .Y(new_n3087_));
  OAI22X1  g2445(.A0(new_n3087_), .A1(new_n3084_), .B0(new_n3082_), .B1(new_n3080_), .Y(new_n3088_));
  NOR3X1   g2446(.A(new_n1286_), .B(new_n1284_), .C(new_n1245_), .Y(new_n3089_));
  AOI21X1  g2447(.A0(new_n1348_), .A1(new_n1347_), .B0(new_n1239_), .Y(new_n3090_));
  NOR2X1   g2448(.A(new_n3090_), .B(new_n3089_), .Y(new_n3091_));
  INVX1    g2449(.A(new_n3091_), .Y(new_n3092_));
  NOR3X1   g2450(.A(new_n2061_), .B(new_n2060_), .C(new_n1956_), .Y(new_n3093_));
  AOI21X1  g2451(.A0(new_n2071_), .A1(\in2[117] ), .B0(new_n3093_), .Y(new_n3094_));
  AOI21X1  g2452(.A0(new_n1348_), .A1(new_n1347_), .B0(new_n1238_), .Y(new_n3095_));
  AOI21X1  g2453(.A0(new_n2225_), .A1(\in1[116] ), .B0(new_n3095_), .Y(new_n3096_));
  INVX1    g2454(.A(new_n3096_), .Y(new_n3097_));
  AOI21X1  g2455(.A0(new_n2063_), .A1(new_n1998_), .B0(new_n1950_), .Y(new_n3098_));
  AOI21X1  g2456(.A0(new_n2391_), .A1(\in3[116] ), .B0(new_n3098_), .Y(new_n3099_));
  OAI22X1  g2457(.A0(new_n3099_), .A1(new_n3097_), .B0(new_n3094_), .B1(new_n3092_), .Y(new_n3100_));
  OR2X1    g2458(.A(new_n3100_), .B(new_n3088_), .Y(new_n3101_));
  AOI21X1  g2459(.A0(new_n3076_), .A1(new_n3071_), .B0(new_n3101_), .Y(new_n3102_));
  AND2X1   g2460(.A(new_n3099_), .B(new_n3097_), .Y(new_n3103_));
  OAI21X1  g2461(.A0(new_n3094_), .A1(new_n3092_), .B0(new_n3103_), .Y(new_n3104_));
  NAND2X1  g2462(.A(new_n3094_), .B(new_n3092_), .Y(new_n3105_));
  AOI21X1  g2463(.A0(new_n3105_), .A1(new_n3104_), .B0(new_n3088_), .Y(new_n3106_));
  NOR2X1   g2464(.A(new_n3082_), .B(new_n3080_), .Y(new_n3107_));
  NAND2X1  g2465(.A(new_n3082_), .B(new_n3080_), .Y(new_n3108_));
  NAND2X1  g2466(.A(new_n3087_), .B(new_n3084_), .Y(new_n3109_));
  OAI21X1  g2467(.A0(new_n3109_), .A1(new_n3107_), .B0(new_n3108_), .Y(new_n3110_));
  OR2X1    g2468(.A(new_n3110_), .B(new_n3106_), .Y(new_n3111_));
  AOI21X1  g2469(.A0(new_n1348_), .A1(new_n1347_), .B0(new_n1255_), .Y(new_n3112_));
  AOI21X1  g2470(.A0(new_n2225_), .A1(\in1[123] ), .B0(new_n3112_), .Y(new_n3113_));
  INVX1    g2471(.A(new_n3113_), .Y(new_n3114_));
  AOI21X1  g2472(.A0(new_n2063_), .A1(new_n1998_), .B0(new_n1967_), .Y(new_n3115_));
  AOI21X1  g2473(.A0(new_n2391_), .A1(\in3[123] ), .B0(new_n3115_), .Y(new_n3116_));
  NOR3X1   g2474(.A(new_n2061_), .B(new_n2060_), .C(new_n1978_), .Y(new_n3117_));
  AOI21X1  g2475(.A0(new_n2071_), .A1(\in2[122] ), .B0(new_n3117_), .Y(new_n3118_));
  NOR3X1   g2476(.A(new_n1286_), .B(new_n1284_), .C(new_n1265_), .Y(new_n3119_));
  AOI21X1  g2477(.A0(new_n1348_), .A1(new_n1347_), .B0(new_n1254_), .Y(new_n3120_));
  NOR2X1   g2478(.A(new_n3120_), .B(new_n3119_), .Y(new_n3121_));
  INVX1    g2479(.A(new_n3121_), .Y(new_n3122_));
  OAI22X1  g2480(.A0(new_n3122_), .A1(new_n3118_), .B0(new_n3116_), .B1(new_n3114_), .Y(new_n3123_));
  NOR3X1   g2481(.A(new_n1286_), .B(new_n1284_), .C(new_n1264_), .Y(new_n3124_));
  AOI21X1  g2482(.A0(new_n1348_), .A1(new_n1347_), .B0(new_n1258_), .Y(new_n3125_));
  NOR2X1   g2483(.A(new_n3125_), .B(new_n3124_), .Y(new_n3126_));
  INVX1    g2484(.A(new_n3126_), .Y(new_n3127_));
  NOR3X1   g2485(.A(new_n2061_), .B(new_n2060_), .C(new_n1977_), .Y(new_n3128_));
  AOI21X1  g2486(.A0(new_n2071_), .A1(\in2[121] ), .B0(new_n3128_), .Y(new_n3129_));
  AOI21X1  g2487(.A0(new_n2063_), .A1(new_n1998_), .B0(new_n1969_), .Y(new_n3130_));
  AOI21X1  g2488(.A0(new_n2391_), .A1(\in3[120] ), .B0(new_n3130_), .Y(new_n3131_));
  AOI21X1  g2489(.A0(new_n1348_), .A1(new_n1347_), .B0(new_n1257_), .Y(new_n3132_));
  AOI21X1  g2490(.A0(new_n2225_), .A1(\in1[120] ), .B0(new_n3132_), .Y(new_n3133_));
  INVX1    g2491(.A(new_n3133_), .Y(new_n3134_));
  OAI22X1  g2492(.A0(new_n3134_), .A1(new_n3131_), .B0(new_n3129_), .B1(new_n3127_), .Y(new_n3135_));
  NOR2X1   g2493(.A(new_n3135_), .B(new_n3123_), .Y(new_n3136_));
  OAI21X1  g2494(.A0(new_n3111_), .A1(new_n3102_), .B0(new_n3136_), .Y(new_n3137_));
  AND2X1   g2495(.A(new_n3134_), .B(new_n3131_), .Y(new_n3138_));
  OAI21X1  g2496(.A0(new_n3129_), .A1(new_n3127_), .B0(new_n3138_), .Y(new_n3139_));
  AOI22X1  g2497(.A0(new_n3129_), .A1(new_n3127_), .B0(new_n3122_), .B1(new_n3118_), .Y(new_n3140_));
  AOI21X1  g2498(.A0(new_n3140_), .A1(new_n3139_), .B0(new_n3123_), .Y(new_n3141_));
  AOI21X1  g2499(.A0(new_n3116_), .A1(new_n3114_), .B0(new_n3141_), .Y(new_n3142_));
  NOR3X1   g2500(.A(new_n1286_), .B(new_n1284_), .C(new_n1281_), .Y(new_n3143_));
  AOI21X1  g2501(.A0(new_n1348_), .A1(new_n1347_), .B0(new_n1275_), .Y(new_n3144_));
  NOR2X1   g2502(.A(new_n3144_), .B(new_n3143_), .Y(new_n3145_));
  INVX1    g2503(.A(new_n3145_), .Y(new_n3146_));
  NOR3X1   g2504(.A(new_n2061_), .B(new_n2060_), .C(new_n1991_), .Y(new_n3147_));
  AOI21X1  g2505(.A0(new_n2071_), .A1(\in2[126] ), .B0(new_n3147_), .Y(new_n3148_));
  NOR2X1   g2506(.A(new_n3148_), .B(new_n3146_), .Y(new_n3149_));
  AOI21X1  g2507(.A0(new_n1348_), .A1(new_n1347_), .B0(new_n1274_), .Y(new_n3150_));
  AOI21X1  g2508(.A0(new_n2225_), .A1(\in1[125] ), .B0(new_n3150_), .Y(new_n3151_));
  NOR3X1   g2509(.A(new_n2061_), .B(new_n2060_), .C(new_n1993_), .Y(new_n3152_));
  AOI21X1  g2510(.A0(new_n2063_), .A1(new_n1998_), .B0(new_n1984_), .Y(new_n3153_));
  NOR2X1   g2511(.A(new_n3153_), .B(new_n3152_), .Y(new_n3154_));
  INVX1    g2512(.A(new_n3154_), .Y(new_n3155_));
  AOI21X1  g2513(.A0(new_n3155_), .A1(new_n3151_), .B0(new_n3149_), .Y(new_n3156_));
  AOI21X1  g2514(.A0(new_n1348_), .A1(new_n1347_), .B0(new_n1277_), .Y(new_n3157_));
  AOI21X1  g2515(.A0(new_n2225_), .A1(\in1[124] ), .B0(new_n3157_), .Y(new_n3158_));
  NOR3X1   g2516(.A(new_n2061_), .B(new_n2060_), .C(new_n1992_), .Y(new_n3159_));
  AOI21X1  g2517(.A0(new_n2063_), .A1(new_n1998_), .B0(new_n1987_), .Y(new_n3160_));
  NOR2X1   g2518(.A(new_n3160_), .B(new_n3159_), .Y(new_n3161_));
  INVX1    g2519(.A(new_n3161_), .Y(new_n3162_));
  NOR2X1   g2520(.A(new_n2000_), .B(new_n1999_), .Y(new_n3163_));
  AOI21X1  g2521(.A0(new_n3162_), .A1(new_n3158_), .B0(new_n3163_), .Y(new_n3164_));
  NAND2X1  g2522(.A(new_n3164_), .B(new_n3156_), .Y(new_n3165_));
  AOI21X1  g2523(.A0(new_n3142_), .A1(new_n3137_), .B0(new_n3165_), .Y(new_n3166_));
  OAI22X1  g2524(.A0(new_n3162_), .A1(new_n3158_), .B0(new_n3155_), .B1(new_n3151_), .Y(new_n3167_));
  AOI22X1  g2525(.A0(new_n3167_), .A1(new_n3156_), .B0(new_n3148_), .B1(new_n3146_), .Y(new_n3168_));
  NOR2X1   g2526(.A(new_n3168_), .B(new_n3163_), .Y(new_n3169_));
  NOR3X1   g2527(.A(new_n3169_), .B(new_n3166_), .C(new_n2001_), .Y(\address[1] ));
  AND2X1   g2528(.A(new_n2235_), .B(new_n2234_), .Y(new_n3171_));
  OR4X1    g2529(.A(new_n3169_), .B(new_n3166_), .C(new_n2001_), .D(new_n3171_), .Y(new_n3172_));
  OAI21X1  g2530(.A0(\address[1] ), .A1(new_n1350_), .B0(new_n3172_), .Y(\result[0] ));
  OR4X1    g2531(.A(new_n3169_), .B(new_n3166_), .C(new_n2256_), .D(new_n2001_), .Y(new_n3174_));
  OAI21X1  g2532(.A0(\address[1] ), .A1(new_n2240_), .B0(new_n3174_), .Y(\result[1] ));
  OR4X1    g2533(.A(new_n3169_), .B(new_n3166_), .C(new_n2247_), .D(new_n2001_), .Y(new_n3176_));
  OAI21X1  g2534(.A0(\address[1] ), .A1(new_n2248_), .B0(new_n3176_), .Y(\result[2] ));
  INVX1    g2535(.A(new_n2227_), .Y(new_n3178_));
  OR4X1    g2536(.A(new_n3169_), .B(new_n3166_), .C(new_n2229_), .D(new_n2001_), .Y(new_n3179_));
  OAI21X1  g2537(.A0(\address[1] ), .A1(new_n3178_), .B0(new_n3179_), .Y(\result[3] ));
  OR4X1    g2538(.A(new_n3169_), .B(new_n3166_), .C(new_n2220_), .D(new_n2001_), .Y(new_n3181_));
  OAI21X1  g2539(.A0(\address[1] ), .A1(new_n2223_), .B0(new_n3181_), .Y(\result[4] ));
  OR4X1    g2540(.A(new_n3169_), .B(new_n3166_), .C(new_n2214_), .D(new_n2001_), .Y(new_n3183_));
  OAI21X1  g2541(.A0(\address[1] ), .A1(new_n2217_), .B0(new_n3183_), .Y(\result[5] ));
  OR4X1    g2542(.A(new_n3169_), .B(new_n3166_), .C(new_n2207_), .D(new_n2001_), .Y(new_n3185_));
  OAI21X1  g2543(.A0(\address[1] ), .A1(new_n2211_), .B0(new_n3185_), .Y(\result[6] ));
  OR4X1    g2544(.A(new_n3169_), .B(new_n3166_), .C(new_n2204_), .D(new_n2001_), .Y(new_n3187_));
  OAI21X1  g2545(.A0(\address[1] ), .A1(new_n2200_), .B0(new_n3187_), .Y(\result[7] ));
  OR4X1    g2546(.A(new_n3169_), .B(new_n3166_), .C(new_n2197_), .D(new_n2001_), .Y(new_n3189_));
  OAI21X1  g2547(.A0(\address[1] ), .A1(new_n2286_), .B0(new_n3189_), .Y(\result[8] ));
  OR4X1    g2548(.A(new_n3169_), .B(new_n3166_), .C(new_n2193_), .D(new_n2001_), .Y(new_n3191_));
  OAI21X1  g2549(.A0(\address[1] ), .A1(new_n2292_), .B0(new_n3191_), .Y(\result[9] ));
  OR4X1    g2550(.A(new_n3169_), .B(new_n3166_), .C(new_n2190_), .D(new_n2001_), .Y(new_n3193_));
  OAI21X1  g2551(.A0(\address[1] ), .A1(new_n2186_), .B0(new_n3193_), .Y(\result[10] ));
  OR4X1    g2552(.A(new_n3169_), .B(new_n3166_), .C(new_n2182_), .D(new_n2001_), .Y(new_n3195_));
  OAI21X1  g2553(.A0(\address[1] ), .A1(new_n2178_), .B0(new_n3195_), .Y(\result[11] ));
  OR4X1    g2554(.A(new_n3169_), .B(new_n3166_), .C(new_n2175_), .D(new_n2001_), .Y(new_n3197_));
  OAI21X1  g2555(.A0(\address[1] ), .A1(new_n2171_), .B0(new_n3197_), .Y(\result[12] ));
  OR4X1    g2556(.A(new_n3169_), .B(new_n3166_), .C(new_n2167_), .D(new_n2001_), .Y(new_n3199_));
  OAI21X1  g2557(.A0(\address[1] ), .A1(new_n2163_), .B0(new_n3199_), .Y(\result[13] ));
  OR4X1    g2558(.A(new_n3169_), .B(new_n3166_), .C(new_n2160_), .D(new_n2001_), .Y(new_n3201_));
  OAI21X1  g2559(.A0(\address[1] ), .A1(new_n2156_), .B0(new_n3201_), .Y(\result[14] ));
  OR4X1    g2560(.A(new_n3169_), .B(new_n3166_), .C(new_n2152_), .D(new_n2001_), .Y(new_n3203_));
  OAI21X1  g2561(.A0(\address[1] ), .A1(new_n2148_), .B0(new_n3203_), .Y(\result[15] ));
  OR4X1    g2562(.A(new_n3169_), .B(new_n3166_), .C(new_n2144_), .D(new_n2001_), .Y(new_n3205_));
  OAI21X1  g2563(.A0(\address[1] ), .A1(new_n2322_), .B0(new_n3205_), .Y(\result[16] ));
  OR4X1    g2564(.A(new_n3169_), .B(new_n3166_), .C(new_n2141_), .D(new_n2001_), .Y(new_n3207_));
  OAI21X1  g2565(.A0(\address[1] ), .A1(new_n2329_), .B0(new_n3207_), .Y(\result[17] ));
  OR4X1    g2566(.A(new_n3169_), .B(new_n3166_), .C(new_n2138_), .D(new_n2001_), .Y(new_n3209_));
  OAI21X1  g2567(.A0(\address[1] ), .A1(new_n2334_), .B0(new_n3209_), .Y(\result[18] ));
  NOR2X1   g2568(.A(new_n2132_), .B(new_n2131_), .Y(new_n3211_));
  OR4X1    g2569(.A(new_n3169_), .B(new_n3166_), .C(new_n3211_), .D(new_n2001_), .Y(new_n3212_));
  OAI21X1  g2570(.A0(\address[1] ), .A1(new_n2130_), .B0(new_n3212_), .Y(\result[19] ));
  OR4X1    g2571(.A(new_n3169_), .B(new_n3166_), .C(new_n2126_), .D(new_n2001_), .Y(new_n3214_));
  OAI21X1  g2572(.A0(\address[1] ), .A1(new_n2340_), .B0(new_n3214_), .Y(\result[20] ));
  NOR2X1   g2573(.A(new_n2120_), .B(new_n2119_), .Y(new_n3216_));
  OR4X1    g2574(.A(new_n3169_), .B(new_n3166_), .C(new_n3216_), .D(new_n2001_), .Y(new_n3217_));
  OAI21X1  g2575(.A0(\address[1] ), .A1(new_n2118_), .B0(new_n3217_), .Y(\result[21] ));
  OR4X1    g2576(.A(new_n3169_), .B(new_n3166_), .C(new_n2114_), .D(new_n2001_), .Y(new_n3219_));
  OAI21X1  g2577(.A0(\address[1] ), .A1(new_n2346_), .B0(new_n3219_), .Y(\result[22] ));
  NOR2X1   g2578(.A(new_n2108_), .B(new_n2107_), .Y(new_n3221_));
  OR4X1    g2579(.A(new_n3169_), .B(new_n3166_), .C(new_n3221_), .D(new_n2001_), .Y(new_n3222_));
  OAI21X1  g2580(.A0(\address[1] ), .A1(new_n2106_), .B0(new_n3222_), .Y(\result[23] ));
  OR4X1    g2581(.A(new_n3169_), .B(new_n3166_), .C(new_n2103_), .D(new_n2001_), .Y(new_n3224_));
  OAI21X1  g2582(.A0(\address[1] ), .A1(new_n2352_), .B0(new_n3224_), .Y(\result[24] ));
  OR4X1    g2583(.A(new_n3169_), .B(new_n3166_), .C(new_n2100_), .D(new_n2001_), .Y(new_n3226_));
  OAI21X1  g2584(.A0(\address[1] ), .A1(new_n2357_), .B0(new_n3226_), .Y(\result[25] ));
  OR4X1    g2585(.A(new_n3169_), .B(new_n3166_), .C(new_n2097_), .D(new_n2001_), .Y(new_n3228_));
  OAI21X1  g2586(.A0(\address[1] ), .A1(new_n2094_), .B0(new_n3228_), .Y(\result[26] ));
  OR4X1    g2587(.A(new_n3169_), .B(new_n3166_), .C(new_n2090_), .D(new_n2001_), .Y(new_n3230_));
  OAI21X1  g2588(.A0(\address[1] ), .A1(new_n2363_), .B0(new_n3230_), .Y(\result[27] ));
  OR4X1    g2589(.A(new_n3169_), .B(new_n3166_), .C(new_n2085_), .D(new_n2001_), .Y(new_n3232_));
  OAI21X1  g2590(.A0(\address[1] ), .A1(new_n2082_), .B0(new_n3232_), .Y(\result[28] ));
  OR4X1    g2591(.A(new_n3169_), .B(new_n3166_), .C(new_n2078_), .D(new_n2001_), .Y(new_n3234_));
  OAI21X1  g2592(.A0(\address[1] ), .A1(new_n2368_), .B0(new_n3234_), .Y(\result[29] ));
  OR4X1    g2593(.A(new_n3169_), .B(new_n3166_), .C(new_n2073_), .D(new_n2001_), .Y(new_n3236_));
  OAI21X1  g2594(.A0(\address[1] ), .A1(new_n2069_), .B0(new_n3236_), .Y(\result[30] ));
  OR4X1    g2595(.A(new_n3169_), .B(new_n3166_), .C(new_n2065_), .D(new_n2001_), .Y(new_n3238_));
  OAI21X1  g2596(.A0(\address[1] ), .A1(new_n2373_), .B0(new_n3238_), .Y(\result[31] ));
  OR4X1    g2597(.A(new_n3169_), .B(new_n3166_), .C(new_n2397_), .D(new_n2001_), .Y(new_n3240_));
  OAI21X1  g2598(.A0(\address[1] ), .A1(new_n2429_), .B0(new_n3240_), .Y(\result[32] ));
  OR4X1    g2599(.A(new_n3169_), .B(new_n3166_), .C(new_n2387_), .D(new_n2001_), .Y(new_n3242_));
  OAI21X1  g2600(.A0(\address[1] ), .A1(new_n2384_), .B0(new_n3242_), .Y(\result[33] ));
  OR4X1    g2601(.A(new_n3169_), .B(new_n3166_), .C(new_n2376_), .D(new_n2001_), .Y(new_n3244_));
  OAI21X1  g2602(.A0(\address[1] ), .A1(new_n2379_), .B0(new_n3244_), .Y(\result[34] ));
  OR4X1    g2603(.A(new_n3169_), .B(new_n3166_), .C(new_n2393_), .D(new_n2001_), .Y(new_n3246_));
  OAI21X1  g2604(.A0(\address[1] ), .A1(new_n2389_), .B0(new_n3246_), .Y(\result[35] ));
  OR4X1    g2605(.A(new_n3169_), .B(new_n3166_), .C(new_n2418_), .D(new_n2001_), .Y(new_n3248_));
  OAI21X1  g2606(.A0(\address[1] ), .A1(new_n2415_), .B0(new_n3248_), .Y(\result[36] ));
  OR4X1    g2607(.A(new_n3169_), .B(new_n3166_), .C(new_n2424_), .D(new_n2001_), .Y(new_n3250_));
  OAI21X1  g2608(.A0(\address[1] ), .A1(new_n2421_), .B0(new_n3250_), .Y(\result[37] ));
  OR4X1    g2609(.A(new_n3169_), .B(new_n3166_), .C(new_n2408_), .D(new_n2001_), .Y(new_n3252_));
  OAI21X1  g2610(.A0(\address[1] ), .A1(new_n2410_), .B0(new_n3252_), .Y(\result[38] ));
  OR4X1    g2611(.A(new_n3169_), .B(new_n3166_), .C(new_n2406_), .D(new_n2001_), .Y(new_n3254_));
  OAI21X1  g2612(.A0(\address[1] ), .A1(new_n2403_), .B0(new_n3254_), .Y(\result[39] ));
  OR4X1    g2613(.A(new_n3169_), .B(new_n3166_), .C(new_n2494_), .D(new_n2001_), .Y(new_n3256_));
  OAI21X1  g2614(.A0(\address[1] ), .A1(new_n2492_), .B0(new_n3256_), .Y(\result[40] ));
  AOI21X1  g2615(.A0(new_n2382_), .A1(\in0[41] ), .B0(new_n2486_), .Y(new_n3258_));
  OR4X1    g2616(.A(new_n3169_), .B(new_n3166_), .C(new_n2489_), .D(new_n2001_), .Y(new_n3259_));
  OAI21X1  g2617(.A0(\address[1] ), .A1(new_n3258_), .B0(new_n3259_), .Y(\result[41] ));
  OR4X1    g2618(.A(new_n3169_), .B(new_n3166_), .C(new_n2483_), .D(new_n2001_), .Y(new_n3261_));
  OAI21X1  g2619(.A0(\address[1] ), .A1(new_n2480_), .B0(new_n3261_), .Y(\result[42] ));
  OR4X1    g2620(.A(new_n3169_), .B(new_n3166_), .C(new_n2477_), .D(new_n2001_), .Y(new_n3263_));
  OAI21X1  g2621(.A0(\address[1] ), .A1(new_n2475_), .B0(new_n3263_), .Y(\result[43] ));
  OR4X1    g2622(.A(new_n3169_), .B(new_n3166_), .C(new_n2465_), .D(new_n2001_), .Y(new_n3265_));
  OAI21X1  g2623(.A0(\address[1] ), .A1(new_n2462_), .B0(new_n3265_), .Y(\result[44] ));
  OR4X1    g2624(.A(new_n3169_), .B(new_n3166_), .C(new_n2471_), .D(new_n2001_), .Y(new_n3267_));
  OAI21X1  g2625(.A0(\address[1] ), .A1(new_n2468_), .B0(new_n3267_), .Y(\result[45] ));
  OR4X1    g2626(.A(new_n3169_), .B(new_n3166_), .C(new_n2455_), .D(new_n2001_), .Y(new_n3269_));
  OAI21X1  g2627(.A0(\address[1] ), .A1(new_n2457_), .B0(new_n3269_), .Y(\result[46] ));
  OR4X1    g2628(.A(new_n3169_), .B(new_n3166_), .C(new_n2452_), .D(new_n2001_), .Y(new_n3271_));
  OAI21X1  g2629(.A0(\address[1] ), .A1(new_n2449_), .B0(new_n3271_), .Y(\result[47] ));
  OR4X1    g2630(.A(new_n3169_), .B(new_n3166_), .C(new_n2534_), .D(new_n2001_), .Y(new_n3273_));
  OAI21X1  g2631(.A0(\address[1] ), .A1(new_n2565_), .B0(new_n3273_), .Y(\result[48] ));
  OR4X1    g2632(.A(new_n3169_), .B(new_n3166_), .C(new_n2525_), .D(new_n2001_), .Y(new_n3275_));
  OAI21X1  g2633(.A0(\address[1] ), .A1(new_n2522_), .B0(new_n3275_), .Y(\result[49] ));
  OR4X1    g2634(.A(new_n3169_), .B(new_n3166_), .C(new_n2515_), .D(new_n2001_), .Y(new_n3277_));
  OAI21X1  g2635(.A0(\address[1] ), .A1(new_n2518_), .B0(new_n3277_), .Y(\result[50] ));
  OR4X1    g2636(.A(new_n3169_), .B(new_n3166_), .C(new_n2530_), .D(new_n2001_), .Y(new_n3279_));
  OAI21X1  g2637(.A0(\address[1] ), .A1(new_n2527_), .B0(new_n3279_), .Y(\result[51] ));
  OR4X1    g2638(.A(new_n3169_), .B(new_n3166_), .C(new_n2557_), .D(new_n2001_), .Y(new_n3281_));
  OAI21X1  g2639(.A0(\address[1] ), .A1(new_n2559_), .B0(new_n3281_), .Y(\result[52] ));
  OR4X1    g2640(.A(new_n3169_), .B(new_n3166_), .C(new_n2577_), .D(new_n2001_), .Y(new_n3283_));
  OAI21X1  g2641(.A0(\address[1] ), .A1(new_n2552_), .B0(new_n3283_), .Y(\result[53] ));
  OR4X1    g2642(.A(new_n3169_), .B(new_n3166_), .C(new_n2545_), .D(new_n2001_), .Y(new_n3285_));
  OAI21X1  g2643(.A0(\address[1] ), .A1(new_n2548_), .B0(new_n3285_), .Y(\result[54] ));
  OR4X1    g2644(.A(new_n3169_), .B(new_n3166_), .C(new_n2541_), .D(new_n2001_), .Y(new_n3287_));
  OAI21X1  g2645(.A0(\address[1] ), .A1(new_n2539_), .B0(new_n3287_), .Y(\result[55] ));
  OR4X1    g2646(.A(new_n3169_), .B(new_n3166_), .C(new_n2630_), .D(new_n2001_), .Y(new_n3289_));
  OAI21X1  g2647(.A0(\address[1] ), .A1(new_n2628_), .B0(new_n3289_), .Y(\result[56] ));
  AOI21X1  g2648(.A0(new_n2382_), .A1(\in0[57] ), .B0(new_n2622_), .Y(new_n3291_));
  OR4X1    g2649(.A(new_n3169_), .B(new_n3166_), .C(new_n2625_), .D(new_n2001_), .Y(new_n3292_));
  OAI21X1  g2650(.A0(\address[1] ), .A1(new_n3291_), .B0(new_n3292_), .Y(\result[57] ));
  OR4X1    g2651(.A(new_n3169_), .B(new_n3166_), .C(new_n2619_), .D(new_n2001_), .Y(new_n3294_));
  OAI21X1  g2652(.A0(\address[1] ), .A1(new_n2616_), .B0(new_n3294_), .Y(\result[58] ));
  OR4X1    g2653(.A(new_n3169_), .B(new_n3166_), .C(new_n2613_), .D(new_n2001_), .Y(new_n3296_));
  OAI21X1  g2654(.A0(\address[1] ), .A1(new_n2611_), .B0(new_n3296_), .Y(\result[59] ));
  OR4X1    g2655(.A(new_n3169_), .B(new_n3166_), .C(new_n2601_), .D(new_n2001_), .Y(new_n3298_));
  OAI21X1  g2656(.A0(\address[1] ), .A1(new_n2598_), .B0(new_n3298_), .Y(\result[60] ));
  OR4X1    g2657(.A(new_n3169_), .B(new_n3166_), .C(new_n2607_), .D(new_n2001_), .Y(new_n3300_));
  OAI21X1  g2658(.A0(\address[1] ), .A1(new_n2604_), .B0(new_n3300_), .Y(\result[61] ));
  OR4X1    g2659(.A(new_n3169_), .B(new_n3166_), .C(new_n2591_), .D(new_n2001_), .Y(new_n3302_));
  OAI21X1  g2660(.A0(\address[1] ), .A1(new_n2593_), .B0(new_n3302_), .Y(\result[62] ));
  OR4X1    g2661(.A(new_n3169_), .B(new_n3166_), .C(new_n2588_), .D(new_n2001_), .Y(new_n3304_));
  OAI21X1  g2662(.A0(\address[1] ), .A1(new_n2585_), .B0(new_n3304_), .Y(\result[63] ));
  OR4X1    g2663(.A(new_n3169_), .B(new_n3166_), .C(new_n2663_), .D(new_n2001_), .Y(new_n3306_));
  OAI21X1  g2664(.A0(\address[1] ), .A1(new_n2665_), .B0(new_n3306_), .Y(\result[64] ));
  OR4X1    g2665(.A(new_n3169_), .B(new_n3166_), .C(new_n2672_), .D(new_n2001_), .Y(new_n3308_));
  OAI21X1  g2666(.A0(\address[1] ), .A1(new_n2669_), .B0(new_n3308_), .Y(\result[65] ));
  OR4X1    g2667(.A(new_n3169_), .B(new_n3166_), .C(new_n2656_), .D(new_n2001_), .Y(new_n3310_));
  OAI21X1  g2668(.A0(\address[1] ), .A1(new_n2659_), .B0(new_n3310_), .Y(\result[66] ));
  OR4X1    g2669(.A(new_n3169_), .B(new_n3166_), .C(new_n2654_), .D(new_n2001_), .Y(new_n3312_));
  OAI21X1  g2670(.A0(\address[1] ), .A1(new_n2651_), .B0(new_n3312_), .Y(\result[67] ));
  OR4X1    g2671(.A(new_n3169_), .B(new_n3166_), .C(new_n2703_), .D(new_n2001_), .Y(new_n3314_));
  OAI21X1  g2672(.A0(\address[1] ), .A1(new_n2700_), .B0(new_n3314_), .Y(\result[68] ));
  OR4X1    g2673(.A(new_n3169_), .B(new_n3166_), .C(new_n2698_), .D(new_n2001_), .Y(new_n3316_));
  OAI21X1  g2674(.A0(\address[1] ), .A1(new_n2695_), .B0(new_n3316_), .Y(\result[69] ));
  OR4X1    g2675(.A(new_n3169_), .B(new_n3166_), .C(new_n2688_), .D(new_n2001_), .Y(new_n3318_));
  OAI21X1  g2676(.A0(\address[1] ), .A1(new_n2690_), .B0(new_n3318_), .Y(\result[70] ));
  OR4X1    g2677(.A(new_n3169_), .B(new_n3166_), .C(new_n2686_), .D(new_n2001_), .Y(new_n3320_));
  OAI21X1  g2678(.A0(\address[1] ), .A1(new_n2683_), .B0(new_n3320_), .Y(\result[71] ));
  OR4X1    g2679(.A(new_n3169_), .B(new_n3166_), .C(new_n2735_), .D(new_n2001_), .Y(new_n3322_));
  OAI21X1  g2680(.A0(\address[1] ), .A1(new_n2737_), .B0(new_n3322_), .Y(\result[72] ));
  OR4X1    g2681(.A(new_n3169_), .B(new_n3166_), .C(new_n2733_), .D(new_n2001_), .Y(new_n3324_));
  OAI21X1  g2682(.A0(\address[1] ), .A1(new_n2730_), .B0(new_n3324_), .Y(\result[73] ));
  OR4X1    g2683(.A(new_n3169_), .B(new_n3166_), .C(new_n2722_), .D(new_n2001_), .Y(new_n3326_));
  OAI21X1  g2684(.A0(\address[1] ), .A1(new_n2725_), .B0(new_n3326_), .Y(\result[74] ));
  OR4X1    g2685(.A(new_n3169_), .B(new_n3166_), .C(new_n2720_), .D(new_n2001_), .Y(new_n3328_));
  OAI21X1  g2686(.A0(\address[1] ), .A1(new_n2717_), .B0(new_n3328_), .Y(\result[75] ));
  OR4X1    g2687(.A(new_n3169_), .B(new_n3166_), .C(new_n2769_), .D(new_n2001_), .Y(new_n3330_));
  OAI21X1  g2688(.A0(\address[1] ), .A1(new_n2766_), .B0(new_n3330_), .Y(\result[76] ));
  OR4X1    g2689(.A(new_n3169_), .B(new_n3166_), .C(new_n2764_), .D(new_n2001_), .Y(new_n3332_));
  OAI21X1  g2690(.A0(\address[1] ), .A1(new_n2761_), .B0(new_n3332_), .Y(\result[77] ));
  OR4X1    g2691(.A(new_n3169_), .B(new_n3166_), .C(new_n2754_), .D(new_n2001_), .Y(new_n3334_));
  OAI21X1  g2692(.A0(\address[1] ), .A1(new_n2756_), .B0(new_n3334_), .Y(\result[78] ));
  OR4X1    g2693(.A(new_n3169_), .B(new_n3166_), .C(new_n2752_), .D(new_n2001_), .Y(new_n3336_));
  OAI21X1  g2694(.A0(\address[1] ), .A1(new_n2749_), .B0(new_n3336_), .Y(\result[79] ));
  OR4X1    g2695(.A(new_n3169_), .B(new_n3166_), .C(new_n2795_), .D(new_n2001_), .Y(new_n3338_));
  OAI21X1  g2696(.A0(\address[1] ), .A1(new_n2797_), .B0(new_n3338_), .Y(\result[80] ));
  OR4X1    g2697(.A(new_n3169_), .B(new_n3166_), .C(new_n2804_), .D(new_n2001_), .Y(new_n3340_));
  OAI21X1  g2698(.A0(\address[1] ), .A1(new_n2801_), .B0(new_n3340_), .Y(\result[81] ));
  OR4X1    g2699(.A(new_n3169_), .B(new_n3166_), .C(new_n2788_), .D(new_n2001_), .Y(new_n3342_));
  OAI21X1  g2700(.A0(\address[1] ), .A1(new_n2791_), .B0(new_n3342_), .Y(\result[82] ));
  OR4X1    g2701(.A(new_n3169_), .B(new_n3166_), .C(new_n2786_), .D(new_n2001_), .Y(new_n3344_));
  OAI21X1  g2702(.A0(\address[1] ), .A1(new_n2783_), .B0(new_n3344_), .Y(\result[83] ));
  OR4X1    g2703(.A(new_n3169_), .B(new_n3166_), .C(new_n2835_), .D(new_n2001_), .Y(new_n3346_));
  OAI21X1  g2704(.A0(\address[1] ), .A1(new_n2832_), .B0(new_n3346_), .Y(\result[84] ));
  OR4X1    g2705(.A(new_n3169_), .B(new_n3166_), .C(new_n2830_), .D(new_n2001_), .Y(new_n3348_));
  OAI21X1  g2706(.A0(\address[1] ), .A1(new_n2827_), .B0(new_n3348_), .Y(\result[85] ));
  OR4X1    g2707(.A(new_n3169_), .B(new_n3166_), .C(new_n2820_), .D(new_n2001_), .Y(new_n3350_));
  OAI21X1  g2708(.A0(\address[1] ), .A1(new_n2822_), .B0(new_n3350_), .Y(\result[86] ));
  OR4X1    g2709(.A(new_n3169_), .B(new_n3166_), .C(new_n2818_), .D(new_n2001_), .Y(new_n3352_));
  OAI21X1  g2710(.A0(\address[1] ), .A1(new_n2815_), .B0(new_n3352_), .Y(\result[87] ));
  OR4X1    g2711(.A(new_n3169_), .B(new_n3166_), .C(new_n2867_), .D(new_n2001_), .Y(new_n3354_));
  OAI21X1  g2712(.A0(\address[1] ), .A1(new_n2869_), .B0(new_n3354_), .Y(\result[88] ));
  OR4X1    g2713(.A(new_n3169_), .B(new_n3166_), .C(new_n2865_), .D(new_n2001_), .Y(new_n3356_));
  OAI21X1  g2714(.A0(\address[1] ), .A1(new_n2862_), .B0(new_n3356_), .Y(\result[89] ));
  OR4X1    g2715(.A(new_n3169_), .B(new_n3166_), .C(new_n2854_), .D(new_n2001_), .Y(new_n3358_));
  OAI21X1  g2716(.A0(\address[1] ), .A1(new_n2857_), .B0(new_n3358_), .Y(\result[90] ));
  OR4X1    g2717(.A(new_n3169_), .B(new_n3166_), .C(new_n2852_), .D(new_n2001_), .Y(new_n3360_));
  OAI21X1  g2718(.A0(\address[1] ), .A1(new_n2849_), .B0(new_n3360_), .Y(\result[91] ));
  OR4X1    g2719(.A(new_n3169_), .B(new_n3166_), .C(new_n2901_), .D(new_n2001_), .Y(new_n3362_));
  OAI21X1  g2720(.A0(\address[1] ), .A1(new_n2898_), .B0(new_n3362_), .Y(\result[92] ));
  OR4X1    g2721(.A(new_n3169_), .B(new_n3166_), .C(new_n2896_), .D(new_n2001_), .Y(new_n3364_));
  OAI21X1  g2722(.A0(\address[1] ), .A1(new_n2893_), .B0(new_n3364_), .Y(\result[93] ));
  OR4X1    g2723(.A(new_n3169_), .B(new_n3166_), .C(new_n2886_), .D(new_n2001_), .Y(new_n3366_));
  OAI21X1  g2724(.A0(\address[1] ), .A1(new_n2888_), .B0(new_n3366_), .Y(\result[94] ));
  OR4X1    g2725(.A(new_n3169_), .B(new_n3166_), .C(new_n2884_), .D(new_n2001_), .Y(new_n3368_));
  OAI21X1  g2726(.A0(\address[1] ), .A1(new_n2881_), .B0(new_n3368_), .Y(\result[95] ));
  OR4X1    g2727(.A(new_n3169_), .B(new_n3166_), .C(new_n2927_), .D(new_n2001_), .Y(new_n3370_));
  OAI21X1  g2728(.A0(\address[1] ), .A1(new_n2929_), .B0(new_n3370_), .Y(\result[96] ));
  OR4X1    g2729(.A(new_n3169_), .B(new_n3166_), .C(new_n2936_), .D(new_n2001_), .Y(new_n3372_));
  OAI21X1  g2730(.A0(\address[1] ), .A1(new_n2933_), .B0(new_n3372_), .Y(\result[97] ));
  OR4X1    g2731(.A(new_n3169_), .B(new_n3166_), .C(new_n2920_), .D(new_n2001_), .Y(new_n3374_));
  OAI21X1  g2732(.A0(\address[1] ), .A1(new_n2923_), .B0(new_n3374_), .Y(\result[98] ));
  OR4X1    g2733(.A(new_n3169_), .B(new_n3166_), .C(new_n2918_), .D(new_n2001_), .Y(new_n3376_));
  OAI21X1  g2734(.A0(\address[1] ), .A1(new_n2915_), .B0(new_n3376_), .Y(\result[99] ));
  OR4X1    g2735(.A(new_n3169_), .B(new_n3166_), .C(new_n2967_), .D(new_n2001_), .Y(new_n3378_));
  OAI21X1  g2736(.A0(\address[1] ), .A1(new_n2964_), .B0(new_n3378_), .Y(\result[100] ));
  OR4X1    g2737(.A(new_n3169_), .B(new_n3166_), .C(new_n2962_), .D(new_n2001_), .Y(new_n3380_));
  OAI21X1  g2738(.A0(\address[1] ), .A1(new_n2959_), .B0(new_n3380_), .Y(\result[101] ));
  OR4X1    g2739(.A(new_n3169_), .B(new_n3166_), .C(new_n2952_), .D(new_n2001_), .Y(new_n3382_));
  OAI21X1  g2740(.A0(\address[1] ), .A1(new_n2954_), .B0(new_n3382_), .Y(\result[102] ));
  OR4X1    g2741(.A(new_n3169_), .B(new_n3166_), .C(new_n2950_), .D(new_n2001_), .Y(new_n3384_));
  OAI21X1  g2742(.A0(\address[1] ), .A1(new_n2947_), .B0(new_n3384_), .Y(\result[103] ));
  OR4X1    g2743(.A(new_n3169_), .B(new_n3166_), .C(new_n2999_), .D(new_n2001_), .Y(new_n3386_));
  OAI21X1  g2744(.A0(\address[1] ), .A1(new_n3001_), .B0(new_n3386_), .Y(\result[104] ));
  OR4X1    g2745(.A(new_n3169_), .B(new_n3166_), .C(new_n2997_), .D(new_n2001_), .Y(new_n3388_));
  OAI21X1  g2746(.A0(\address[1] ), .A1(new_n2994_), .B0(new_n3388_), .Y(\result[105] ));
  OR4X1    g2747(.A(new_n3169_), .B(new_n3166_), .C(new_n2986_), .D(new_n2001_), .Y(new_n3390_));
  OAI21X1  g2748(.A0(\address[1] ), .A1(new_n2989_), .B0(new_n3390_), .Y(\result[106] ));
  OR4X1    g2749(.A(new_n3169_), .B(new_n3166_), .C(new_n2984_), .D(new_n2001_), .Y(new_n3392_));
  OAI21X1  g2750(.A0(\address[1] ), .A1(new_n2981_), .B0(new_n3392_), .Y(\result[107] ));
  OR4X1    g2751(.A(new_n3169_), .B(new_n3166_), .C(new_n3033_), .D(new_n2001_), .Y(new_n3394_));
  OAI21X1  g2752(.A0(\address[1] ), .A1(new_n3030_), .B0(new_n3394_), .Y(\result[108] ));
  OR4X1    g2753(.A(new_n3169_), .B(new_n3166_), .C(new_n3028_), .D(new_n2001_), .Y(new_n3396_));
  OAI21X1  g2754(.A0(\address[1] ), .A1(new_n3025_), .B0(new_n3396_), .Y(\result[109] ));
  OR4X1    g2755(.A(new_n3169_), .B(new_n3166_), .C(new_n3018_), .D(new_n2001_), .Y(new_n3398_));
  OAI21X1  g2756(.A0(\address[1] ), .A1(new_n3020_), .B0(new_n3398_), .Y(\result[110] ));
  OR4X1    g2757(.A(new_n3169_), .B(new_n3166_), .C(new_n3016_), .D(new_n2001_), .Y(new_n3400_));
  OAI21X1  g2758(.A0(\address[1] ), .A1(new_n3013_), .B0(new_n3400_), .Y(\result[111] ));
  OR4X1    g2759(.A(new_n3169_), .B(new_n3166_), .C(new_n3059_), .D(new_n2001_), .Y(new_n3402_));
  OAI21X1  g2760(.A0(\address[1] ), .A1(new_n3061_), .B0(new_n3402_), .Y(\result[112] ));
  OR4X1    g2761(.A(new_n3169_), .B(new_n3166_), .C(new_n3068_), .D(new_n2001_), .Y(new_n3404_));
  OAI21X1  g2762(.A0(\address[1] ), .A1(new_n3065_), .B0(new_n3404_), .Y(\result[113] ));
  OR4X1    g2763(.A(new_n3169_), .B(new_n3166_), .C(new_n3052_), .D(new_n2001_), .Y(new_n3406_));
  OAI21X1  g2764(.A0(\address[1] ), .A1(new_n3055_), .B0(new_n3406_), .Y(\result[114] ));
  OR4X1    g2765(.A(new_n3169_), .B(new_n3166_), .C(new_n3050_), .D(new_n2001_), .Y(new_n3408_));
  OAI21X1  g2766(.A0(\address[1] ), .A1(new_n3047_), .B0(new_n3408_), .Y(\result[115] ));
  OR4X1    g2767(.A(new_n3169_), .B(new_n3166_), .C(new_n3099_), .D(new_n2001_), .Y(new_n3410_));
  OAI21X1  g2768(.A0(\address[1] ), .A1(new_n3096_), .B0(new_n3410_), .Y(\result[116] ));
  OR4X1    g2769(.A(new_n3169_), .B(new_n3166_), .C(new_n3094_), .D(new_n2001_), .Y(new_n3412_));
  OAI21X1  g2770(.A0(\address[1] ), .A1(new_n3091_), .B0(new_n3412_), .Y(\result[117] ));
  OR4X1    g2771(.A(new_n3169_), .B(new_n3166_), .C(new_n3084_), .D(new_n2001_), .Y(new_n3414_));
  OAI21X1  g2772(.A0(\address[1] ), .A1(new_n3086_), .B0(new_n3414_), .Y(\result[118] ));
  OR4X1    g2773(.A(new_n3169_), .B(new_n3166_), .C(new_n3082_), .D(new_n2001_), .Y(new_n3416_));
  OAI21X1  g2774(.A0(\address[1] ), .A1(new_n3079_), .B0(new_n3416_), .Y(\result[119] ));
  OR4X1    g2775(.A(new_n3169_), .B(new_n3166_), .C(new_n3131_), .D(new_n2001_), .Y(new_n3418_));
  OAI21X1  g2776(.A0(\address[1] ), .A1(new_n3133_), .B0(new_n3418_), .Y(\result[120] ));
  OR4X1    g2777(.A(new_n3169_), .B(new_n3166_), .C(new_n3129_), .D(new_n2001_), .Y(new_n3420_));
  OAI21X1  g2778(.A0(\address[1] ), .A1(new_n3126_), .B0(new_n3420_), .Y(\result[121] ));
  OR4X1    g2779(.A(new_n3169_), .B(new_n3166_), .C(new_n3118_), .D(new_n2001_), .Y(new_n3422_));
  OAI21X1  g2780(.A0(\address[1] ), .A1(new_n3121_), .B0(new_n3422_), .Y(\result[122] ));
  OR4X1    g2781(.A(new_n3169_), .B(new_n3166_), .C(new_n3116_), .D(new_n2001_), .Y(new_n3424_));
  OAI21X1  g2782(.A0(\address[1] ), .A1(new_n3113_), .B0(new_n3424_), .Y(\result[123] ));
  OR4X1    g2783(.A(new_n3169_), .B(new_n3166_), .C(new_n3161_), .D(new_n2001_), .Y(new_n3426_));
  OAI21X1  g2784(.A0(\address[1] ), .A1(new_n3158_), .B0(new_n3426_), .Y(\result[124] ));
  OR4X1    g2785(.A(new_n3169_), .B(new_n3166_), .C(new_n3154_), .D(new_n2001_), .Y(new_n3428_));
  OAI21X1  g2786(.A0(\address[1] ), .A1(new_n3151_), .B0(new_n3428_), .Y(\result[125] ));
  OR4X1    g2787(.A(new_n3169_), .B(new_n3166_), .C(new_n3148_), .D(new_n2001_), .Y(new_n3430_));
  OAI21X1  g2788(.A0(\address[1] ), .A1(new_n3145_), .B0(new_n3430_), .Y(\result[126] ));
  NOR3X1   g2789(.A(new_n3169_), .B(new_n3166_), .C(new_n1999_), .Y(new_n3432_));
  NOR2X1   g2790(.A(new_n3432_), .B(new_n2000_), .Y(\result[127] ));
  OR4X1    g2791(.A(new_n3169_), .B(new_n3166_), .C(new_n2001_), .D(new_n2071_), .Y(new_n3434_));
  OAI21X1  g2792(.A0(\address[1] ), .A1(new_n2382_), .B0(new_n3434_), .Y(\address[0] ));
endmodule


