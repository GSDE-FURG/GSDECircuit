//Converted to Combinational (Partial output: n2564) , Module name: s38584_n2564 , Timestamp: 2018-12-03T15:51:16.442941 
module s38584_n2564 ( g113, g134, g99, g37, g2741, g2610, g2476, g2342, g2051, g2208, g1917, g1783, g2748, g2756, g2619, g2485, g1657, g2351, g2060, g2217, g1926, g1792, g72, g2759, g73, g2763, g1648, n2564 );
input g113, g134, g99, g37, g2741, g2610, g2476, g2342, g2051, g2208, g1917, g1783, g2748, g2756, g2619, g2485, g1657, g2351, g2060, g2217, g1926, g1792, g72, g2759, g73, g2763, g1648;
output n2564;
wire n7528, n4928, n4947, n4946, n4908, n4920_1, n4927, n4936, n4945, n4824, n4809, n4919, n4914, n4917, n4918, n4926, n4922, n4924, n4925_1, n4935, n4930_1, n4931, n4933, n4944_1, n4938, n4940, n4942, n4916, n4909, n4913, n4923, n4921, n4934_1, n4929, g25167, n4932, n4943, n4937, n4939_1, n4941, n4912, n4910_1, n4915_1, n4911, n4629;
OAI21X1  g2884(.A0(n4947), .A1(n4928), .B0(n7528), .Y(n2564));
NAND2X1  g2883(.A(n4946), .B(n4928), .Y(n7528));
OAI21X1  g0308(.A0(n4927), .A1(n4920_1), .B0(n4908), .Y(n4928));
NOR2X1   g0327(.A(n4946), .B(n4928), .Y(n4947));
OR2X1    g0326(.A(n4945), .B(n4936), .Y(n4946));
NOR2X1   g0288(.A(n4809), .B(n4824), .Y(n4908));
NAND4X1  g0300(.A(n4918), .B(n4917), .C(n4914), .D(n4919), .Y(n4920_1));
NAND4X1  g0307(.A(n4925_1), .B(n4924), .C(n4922), .D(n4926), .Y(n4927));
NAND4X1  g0316(.A(n4933), .B(n4931), .C(n4930_1), .D(n4935), .Y(n4936));
NAND4X1  g0325(.A(n4942), .B(n4940), .C(n4938), .D(n4944_1), .Y(n4945));
INVX1    g0204(.A(g113), .Y(n4824));
AOI21X1  g0189(.A0(g37), .A1(g99), .B0(g134), .Y(n4809));
NAND2X1  g0299(.A(n4916), .B(g2741), .Y(n4919));
NAND2X1  g0294(.A(n4913), .B(n4909), .Y(n4914));
NAND2X1  g0297(.A(n4916), .B(n4909), .Y(n4917));
NAND2X1  g0298(.A(n4913), .B(g2741), .Y(n4918));
NAND2X1  g0306(.A(n4923), .B(g2741), .Y(n4926));
NAND2X1  g0302(.A(n4921), .B(n4909), .Y(n4922));
NAND2X1  g0304(.A(n4923), .B(n4909), .Y(n4924));
NAND2X1  g0305(.A(n4921), .B(g2741), .Y(n4925_1));
NAND4X1  g0315(.A(g2741), .B(n4934_1), .C(g2610), .D(n4916), .Y(n4935));
NAND4X1  g0310(.A(n4909), .B(g2476), .C(n4929), .D(n4916), .Y(n4930_1));
NAND3X1  g0311(.A(n4921), .B(g25167), .C(n4909), .Y(n4931));
NAND4X1  g0313(.A(g2741), .B(n4932), .C(g2342), .D(n4913), .Y(n4933));
NAND4X1  g0324(.A(n4943), .B(g2051), .C(g2741), .D(n4923), .Y(n4944_1));
NAND4X1  g0318(.A(n4937), .B(n4909), .C(g2208), .D(n4913), .Y(n4938));
NAND4X1  g0320(.A(n4909), .B(g1917), .C(n4939_1), .D(n4923), .Y(n4940));
NAND4X1  g0322(.A(n4941), .B(g2741), .C(g1783), .D(n4921), .Y(n4942));
NOR4X1   g0296(.A(n4911), .B(n4915_1), .C(n4910_1), .D(n4912), .Y(n4916));
INVX1    g0289(.A(g2741), .Y(n4909));
NOR4X1   g0293(.A(n4911), .B(g2748), .C(n4910_1), .D(n4912), .Y(n4913));
NOR4X1   g0303(.A(n4911), .B(n4915_1), .C(g2756), .D(n4912), .Y(n4923));
NOR4X1   g0301(.A(n4911), .B(g2748), .C(g2756), .D(n4912), .Y(n4921));
INVX1    g0314(.A(g2619), .Y(n4934_1));
INVX1    g0309(.A(g2485), .Y(n4929));
NOR2X1   g0010(.A(n4629), .B(g1657), .Y(g25167));
INVX1    g0312(.A(g2351), .Y(n4932));
INVX1    g0323(.A(g2060), .Y(n4943));
INVX1    g0317(.A(g2217), .Y(n4937));
INVX1    g0319(.A(g1926), .Y(n4939_1));
INVX1    g0321(.A(g1792), .Y(n4941));
XOR2X1   g0292(.A(g2759), .B(g72), .Y(n4912));
INVX1    g0290(.A(g2756), .Y(n4910_1));
INVX1    g0295(.A(g2748), .Y(n4915_1));
XOR2X1   g0291(.A(g2763), .B(g73), .Y(n4911));
INVX1    g0009(.A(g1648), .Y(n4629));

endmodule
