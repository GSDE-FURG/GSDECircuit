//Converted to Combinational (Partial output: n3574) , Module name: s38417_n3574 , Timestamp: 2018-12-03T15:51:13.656565 
module s38417_n3574 ( g2896, g2903, g2908, g1001, g1000, g999, g2892, g2900, g1004, g1003, g1005, g1007, g1006, g1002, g767, g1088, g1092, g963, g762, g749, g758, g744, g740, g776, g753, g771, g780, g897, g853, g823, g894, g826, g900, g906, g903, g891, g873, g879, g876, g945, g951, g948, g936, g942, g939, g888, g885, g909, g915, g912, g882, g954, g960, g957, g918, g924, g921, g927, g933, g930, n3574 );
input g2896, g2903, g2908, g1001, g1000, g999, g2892, g2900, g1004, g1003, g1005, g1007, g1006, g1002, g767, g1088, g1092, g963, g762, g749, g758, g744, g740, g776, g753, g771, g780, g897, g853, g823, g894, g826, g900, g906, g903, g891, g873, g879, g876, g945, g951, g948, g936, g942, g939, g888, g885, g909, g915, g912, g882, g954, g960, g957, g918, g924, g921, g927, g933, g930;
output n3574;
wire n3569, n6965, n6980, n6752, n5399, n6590, n6588, n6571, n6599, n6969, n6974, n6979, n6569_1, n6564_1, n6567, n6568, n5398, n6589, n6566, n6560, n6563, n6565, n6570, n6596_1, n6598, n6966_1, n6967, n6968, n6973, n6970, n6971_1, n6972, n6978, n6975, n6562, n6561, n6559_1, n6595, n6501, n6533, n6546, n6597, n6529_1, n6538, n6542, n6711, n6509_1, n6719, n6715_1, n6724, n6492, n6728, n6696, n6720_1, n6496, n6976_1, n6977, n6508, n6494_1, n6495, n6507, n6499_1, n6500, n6531, n6532, n6544_1, n6545, n6504_1, n6484_1, n6485, n6503, n6521, n6522, n6536, n6537, n6540, n6541, n6505;
OAI21X1  g1937(.A0(n6980), .A1(n6965), .B0(n3569), .Y(n3574));
AOI21X1  g1710(.A0(n6590), .A1(n5399), .B0(n6752), .Y(n3569));
NOR3X1   g1921(.A(n6599), .B(n6571), .C(n6588), .Y(n6965));
NOR3X1   g1936(.A(n6979), .B(n6974), .C(n6969), .Y(n6980));
NOR4X1   g1709(.A(n6568), .B(n6567), .C(n6564_1), .D(n6569_1), .Y(n6752));
NOR4X1   g0357(.A(g2908), .B(g2903), .C(g2896), .D(n5398), .Y(n5399));
INVX1    g1547(.A(n6589), .Y(n6590));
OR4X1    g1545(.A(n6565), .B(n6563), .C(n6560), .D(n6566), .Y(n6588));
INVX1    g1528(.A(n6570), .Y(n6571));
OR2X1    g1556(.A(n6598), .B(n6596_1), .Y(n6599));
NAND3X1  g1925(.A(n6968), .B(n6967), .C(n6966_1), .Y(n6969));
NAND4X1  g1930(.A(n6972), .B(n6971_1), .C(n6970), .D(n6973), .Y(n6974));
OR4X1    g1935(.A(n6975), .B(n6752), .C(n5399), .D(n6978), .Y(n6979));
OAI22X1  g1526(.A0(g1000), .A1(n6561), .B0(n6562), .B1(g1001), .Y(n6569_1));
NOR2X1   g1521(.A(n6563), .B(n6560), .Y(n6564_1));
NOR2X1   g1524(.A(n6566), .B(n6565), .Y(n6567));
NOR2X1   g1525(.A(g999), .B(n6559_1), .Y(n6568));
OR2X1    g0356(.A(g2900), .B(g2892), .Y(n5398));
NOR3X1   g1546(.A(n6569_1), .B(n6568), .C(n6588), .Y(n6589));
OAI22X1  g1523(.A0(g1003), .A1(n6561), .B0(n6562), .B1(g1004), .Y(n6566));
NOR2X1   g1517(.A(g1005), .B(n6559_1), .Y(n6560));
OAI22X1  g1520(.A0(g1006), .A1(n6561), .B0(n6562), .B1(g1007), .Y(n6563));
NOR2X1   g1522(.A(g1002), .B(n6559_1), .Y(n6565));
NOR2X1   g1527(.A(n6569_1), .B(n6568), .Y(n6570));
OR4X1    g1553(.A(n6546), .B(n6533), .C(n6501), .D(n6595), .Y(n6596_1));
OR4X1    g1555(.A(n6542), .B(n6538), .C(n6529_1), .D(n6597), .Y(n6598));
XOR2X1   g1922(.A(n6509_1), .B(n6711), .Y(n6966_1));
XOR2X1   g1923(.A(n6533), .B(n6719), .Y(n6967));
XOR2X1   g1924(.A(n6546), .B(n6715_1), .Y(n6968));
XOR2X1   g1929(.A(n6492), .B(n6724), .Y(n6973));
XOR2X1   g1926(.A(n6529_1), .B(n6728), .Y(n6970));
XOR2X1   g1927(.A(n6538), .B(n6696), .Y(n6971_1));
XOR2X1   g1928(.A(n6496), .B(n6720_1), .Y(n6972));
OR2X1    g1934(.A(n6977), .B(n6976_1), .Y(n6978));
XOR2X1   g1931(.A(n6542), .B(g767), .Y(n6975));
INVX1    g1519(.A(g1088), .Y(n6562));
INVX1    g1518(.A(g1092), .Y(n6561));
INVX1    g1516(.A(g963), .Y(n6559_1));
NAND4X1  g1552(.A(n6507), .B(n6495), .C(n6494_1), .D(n6508), .Y(n6595));
NAND2X1  g1458(.A(n6500), .B(n6499_1), .Y(n6501));
NAND2X1  g1490(.A(n6532), .B(n6531), .Y(n6533));
NAND2X1  g1503(.A(n6545), .B(n6544_1), .Y(n6546));
NAND4X1  g1554(.A(n6503), .B(n6485), .C(n6484_1), .D(n6504_1), .Y(n6597));
NAND2X1  g1486(.A(n6522), .B(n6521), .Y(n6529_1));
NAND2X1  g1495(.A(n6537), .B(n6536), .Y(n6538));
NAND2X1  g1499(.A(n6541), .B(n6540), .Y(n6542));
INVX1    g1668(.A(g762), .Y(n6711));
NAND2X1  g1466(.A(n6508), .B(n6507), .Y(n6509_1));
INVX1    g1676(.A(g749), .Y(n6719));
INVX1    g1672(.A(g758), .Y(n6715_1));
INVX1    g1681(.A(g744), .Y(n6724));
NAND2X1  g1449(.A(n6485), .B(n6484_1), .Y(n6492));
INVX1    g1685(.A(g740), .Y(n6728));
INVX1    g1653(.A(g776), .Y(n6696));
INVX1    g1677(.A(g753), .Y(n6720_1));
NAND2X1  g1453(.A(n6495), .B(n6494_1), .Y(n6496));
XOR2X1   g1932(.A(n6505), .B(g771), .Y(n6976_1));
XOR2X1   g1933(.A(n6501), .B(g780), .Y(n6977));
AOI22X1  g1465(.A0(g894), .A1(g823), .B0(g853), .B1(g897), .Y(n6508));
NAND2X1  g1451(.A(g900), .B(g826), .Y(n6494_1));
AOI22X1  g1452(.A0(g903), .A1(g823), .B0(g853), .B1(g906), .Y(n6495));
NAND2X1  g1464(.A(g891), .B(g826), .Y(n6507));
NAND2X1  g1456(.A(g873), .B(g826), .Y(n6499_1));
AOI22X1  g1457(.A0(g876), .A1(g823), .B0(g853), .B1(g879), .Y(n6500));
NAND2X1  g1488(.A(g945), .B(g826), .Y(n6531));
AOI22X1  g1489(.A0(g948), .A1(g823), .B0(g853), .B1(g951), .Y(n6532));
NAND2X1  g1501(.A(g936), .B(g826), .Y(n6544_1));
AOI22X1  g1502(.A0(g939), .A1(g823), .B0(g853), .B1(g942), .Y(n6545));
AOI22X1  g1461(.A0(g885), .A1(g823), .B0(g853), .B1(g888), .Y(n6504_1));
NAND2X1  g1441(.A(g909), .B(g826), .Y(n6484_1));
AOI22X1  g1442(.A0(g912), .A1(g823), .B0(g853), .B1(g915), .Y(n6485));
NAND2X1  g1460(.A(g882), .B(g826), .Y(n6503));
NAND2X1  g1478(.A(g954), .B(g826), .Y(n6521));
AOI22X1  g1479(.A0(g957), .A1(g823), .B0(g853), .B1(g960), .Y(n6522));
NAND2X1  g1493(.A(g918), .B(g826), .Y(n6536));
AOI22X1  g1494(.A0(g921), .A1(g823), .B0(g853), .B1(g924), .Y(n6537));
NAND2X1  g1497(.A(g927), .B(g826), .Y(n6540));
AOI22X1  g1498(.A0(g930), .A1(g823), .B0(g853), .B1(g933), .Y(n6541));
NAND2X1  g1462(.A(n6504_1), .B(n6503), .Y(n6505));

endmodule
